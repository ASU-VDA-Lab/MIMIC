module fake_netlist_5_2147_n_1201 (n_137, n_210, n_168, n_260, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_248, n_124, n_86, n_136, n_146, n_268, n_182, n_143, n_83, n_132, n_61, n_237, n_90, n_241, n_127, n_75, n_101, n_180, n_184, n_226, n_235, n_65, n_78, n_74, n_144, n_207, n_240, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_229, n_108, n_231, n_257, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_236, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_249, n_271, n_46, n_233, n_21, n_94, n_203, n_245, n_205, n_113, n_38, n_123, n_139, n_105, n_246, n_80, n_4, n_179, n_125, n_35, n_269, n_167, n_128, n_73, n_234, n_17, n_92, n_19, n_267, n_149, n_120, n_232, n_135, n_30, n_156, n_5, n_33, n_126, n_254, n_14, n_225, n_84, n_23, n_202, n_130, n_266, n_272, n_219, n_157, n_258, n_265, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_244, n_251, n_25, n_53, n_160, n_198, n_223, n_247, n_188, n_190, n_8, n_201, n_158, n_263, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_264, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_243, n_239, n_175, n_252, n_169, n_59, n_262, n_26, n_255, n_133, n_238, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_242, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_259, n_270, n_222, n_230, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_253, n_261, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_256, n_48, n_204, n_50, n_250, n_52, n_88, n_110, n_216, n_1201);

input n_137;
input n_210;
input n_168;
input n_260;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_268;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_237;
input n_90;
input n_241;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_235;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_240;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_257;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_236;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_249;
input n_271;
input n_46;
input n_233;
input n_21;
input n_94;
input n_203;
input n_245;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_246;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_269;
input n_167;
input n_128;
input n_73;
input n_234;
input n_17;
input n_92;
input n_19;
input n_267;
input n_149;
input n_120;
input n_232;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_254;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_266;
input n_272;
input n_219;
input n_157;
input n_258;
input n_265;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_244;
input n_251;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_247;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_264;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_243;
input n_239;
input n_175;
input n_252;
input n_169;
input n_59;
input n_262;
input n_26;
input n_255;
input n_133;
input n_238;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_242;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_259;
input n_270;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_253;
input n_261;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_256;
input n_48;
input n_204;
input n_50;
input n_250;
input n_52;
input n_88;
input n_110;
input n_216;

output n_1201;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_380;
wire n_419;
wire n_318;
wire n_977;
wire n_653;
wire n_1194;
wire n_611;
wire n_444;
wire n_1126;
wire n_642;
wire n_1166;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_1141;
wire n_316;
wire n_785;
wire n_389;
wire n_855;
wire n_843;
wire n_1178;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_912;
wire n_315;
wire n_523;
wire n_913;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_1161;
wire n_678;
wire n_664;
wire n_697;
wire n_376;
wire n_503;
wire n_967;
wire n_1150;
wire n_605;
wire n_776;
wire n_928;
wire n_1139;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_620;
wire n_643;
wire n_367;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_525;
wire n_493;
wire n_397;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_1191;
wire n_1198;
wire n_721;
wire n_998;
wire n_1157;
wire n_1099;
wire n_841;
wire n_1050;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_1128;
wire n_280;
wire n_744;
wire n_1021;
wire n_629;
wire n_590;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_690;
wire n_1013;
wire n_583;
wire n_718;
wire n_671;
wire n_819;
wire n_302;
wire n_1022;
wire n_526;
wire n_915;
wire n_1120;
wire n_719;
wire n_443;
wire n_293;
wire n_372;
wire n_677;
wire n_859;
wire n_864;
wire n_1110;
wire n_951;
wire n_1121;
wire n_821;
wire n_714;
wire n_447;
wire n_314;
wire n_368;
wire n_604;
wire n_433;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_1179;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_946;
wire n_417;
wire n_932;
wire n_1048;
wire n_612;
wire n_1001;
wire n_498;
wire n_516;
wire n_385;
wire n_933;
wire n_788;
wire n_507;
wire n_1152;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_1195;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_947;
wire n_373;
wire n_820;
wire n_1090;
wire n_757;
wire n_936;
wire n_1200;
wire n_307;
wire n_633;
wire n_1192;
wire n_439;
wire n_530;
wire n_1024;
wire n_1063;
wire n_556;
wire n_1107;
wire n_448;
wire n_758;
wire n_999;
wire n_1185;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1032;
wire n_1143;
wire n_804;
wire n_867;
wire n_1124;
wire n_537;
wire n_1158;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_1104;
wire n_563;
wire n_1182;
wire n_756;
wire n_1145;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_394;
wire n_579;
wire n_992;
wire n_1049;
wire n_1153;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_1154;
wire n_286;
wire n_883;
wire n_1135;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_1163;
wire n_406;
wire n_519;
wire n_470;
wire n_919;
wire n_782;
wire n_908;
wire n_1108;
wire n_325;
wire n_449;
wire n_1073;
wire n_1100;
wire n_862;
wire n_900;
wire n_1016;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_942;
wire n_381;
wire n_291;
wire n_1147;
wire n_731;
wire n_390;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_592;
wire n_1169;
wire n_920;
wire n_894;
wire n_1046;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_1172;
wire n_1096;
wire n_976;
wire n_1095;
wire n_343;
wire n_308;
wire n_379;
wire n_833;
wire n_428;
wire n_514;
wire n_570;
wire n_457;
wire n_1045;
wire n_297;
wire n_1079;
wire n_853;
wire n_603;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_1168;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_1142;
wire n_660;
wire n_1114;
wire n_1129;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_1148;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_995;
wire n_961;
wire n_955;
wire n_387;
wire n_771;
wire n_1176;
wire n_374;
wire n_276;
wire n_339;
wire n_1149;
wire n_882;
wire n_398;
wire n_1146;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_522;
wire n_550;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_1020;
wire n_662;
wire n_459;
wire n_1062;
wire n_646;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_622;
wire n_1171;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1188;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_1165;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_584;
wire n_681;
wire n_336;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_1177;
wire n_680;
wire n_974;
wire n_432;
wire n_553;
wire n_727;
wire n_395;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_1159;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_1167;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_829;
wire n_749;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_1151;
wire n_1134;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_482;
wire n_342;
wire n_517;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_1173;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_796;
wire n_573;
wire n_1069;
wire n_969;
wire n_866;
wire n_1075;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_571;
wire n_461;
wire n_693;
wire n_333;
wire n_338;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_1193;
wire n_567;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_1122;
wire n_1197;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_1031;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_1028;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1187;
wire n_1015;
wire n_1000;
wire n_891;
wire n_1140;
wire n_466;
wire n_1164;
wire n_630;
wire n_420;
wire n_489;
wire n_632;
wire n_699;
wire n_1174;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_1101;
wire n_273;
wire n_585;
wire n_349;
wire n_1106;
wire n_1190;
wire n_616;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_289;
wire n_745;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1116;
wire n_767;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_1175;
wire n_861;
wire n_534;
wire n_948;
wire n_1183;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1131;
wire n_1059;
wire n_1084;
wire n_1133;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_607;
wire n_575;
wire n_647;
wire n_480;
wire n_354;
wire n_425;
wire n_513;
wire n_710;
wire n_795;
wire n_527;
wire n_707;
wire n_407;
wire n_679;
wire n_832;
wire n_695;
wire n_857;
wire n_1072;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_495;
wire n_487;
wire n_665;
wire n_602;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1130;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_1156;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_404;
wire n_686;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_1136;
wire n_815;
wire n_596;
wire n_1125;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_327;
wire n_1109;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_1160;
wire n_1080;
wire n_1162;
wire n_491;
wire n_1074;
wire n_427;
wire n_1199;
wire n_791;
wire n_732;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_1181;
wire n_1196;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_952;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_870;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_803;
wire n_868;
wire n_1092;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_1138;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_1186;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_1155;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_1123;
wire n_1184;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_1189;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_1180;
wire n_424;
wire n_1003;
wire n_1144;
wire n_1137;
wire n_706;
wire n_746;
wire n_305;
wire n_533;
wire n_950;
wire n_1170;
wire n_747;
wire n_278;
wire n_784;

INVx1_ASAP7_75t_L g273 ( 
.A(n_120),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_50),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_200),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_55),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_141),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_58),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_54),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_201),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_89),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_224),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_66),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_29),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_179),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_163),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_194),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_156),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_35),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_245),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_198),
.B(n_181),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_170),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_138),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_180),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_9),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_155),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_205),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_139),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_251),
.Y(n_299)
);

INVxp33_ASAP7_75t_L g300 ( 
.A(n_136),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_211),
.B(n_85),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_42),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_215),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_253),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_159),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_221),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_206),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_209),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_117),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_7),
.Y(n_310)
);

INVxp33_ASAP7_75t_L g311 ( 
.A(n_258),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_243),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_199),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_80),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_190),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_153),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_39),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_234),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_254),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_266),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_124),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_225),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_204),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_2),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_152),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_236),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_164),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_213),
.Y(n_328)
);

NOR2xp67_ASAP7_75t_L g329 ( 
.A(n_150),
.B(n_178),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_52),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_207),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_270),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_263),
.Y(n_333)
);

NOR2xp67_ASAP7_75t_L g334 ( 
.A(n_100),
.B(n_31),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_121),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_262),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_86),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_143),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_113),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_37),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_36),
.Y(n_341)
);

NOR2xp67_ASAP7_75t_L g342 ( 
.A(n_46),
.B(n_203),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_59),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_84),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_165),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_174),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_184),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_269),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_31),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_149),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_191),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_144),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_264),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_219),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_14),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_94),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_134),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_145),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_137),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_212),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_19),
.Y(n_361)
);

NOR2xp67_ASAP7_75t_L g362 ( 
.A(n_72),
.B(n_247),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_271),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_0),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_193),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_105),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_112),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_202),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_241),
.Y(n_369)
);

INVxp33_ASAP7_75t_L g370 ( 
.A(n_95),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_38),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_185),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_157),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_23),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_12),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_229),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_104),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_250),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_214),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_192),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_21),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_33),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_102),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_230),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_176),
.Y(n_385)
);

NOR2xp67_ASAP7_75t_L g386 ( 
.A(n_11),
.B(n_256),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_40),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_15),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_242),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_130),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_96),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_2),
.Y(n_392)
);

BUFx8_ASAP7_75t_SL g393 ( 
.A(n_27),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_25),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_63),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_103),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_183),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_76),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_30),
.Y(n_399)
);

INVx4_ASAP7_75t_R g400 ( 
.A(n_33),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_173),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_182),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_210),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_98),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_172),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_69),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_126),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_56),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_189),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_14),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_252),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_135),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_99),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_208),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_146),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_223),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_240),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_132),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_160),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_45),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_26),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_17),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_74),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_7),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_265),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_114),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_61),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_217),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_110),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_81),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_197),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_257),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_244),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_106),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_49),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_44),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_73),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_13),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_232),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_88),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_168),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_83),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_24),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_122),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_10),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_169),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_119),
.B(n_195),
.Y(n_447)
);

CKINVDCx14_ASAP7_75t_R g448 ( 
.A(n_259),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_188),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_255),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_111),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_71),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_148),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_231),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_6),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_20),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_261),
.Y(n_457)
);

NOR2xp67_ASAP7_75t_L g458 ( 
.A(n_218),
.B(n_70),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_260),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_62),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_65),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_388),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_393),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_402),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_388),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_445),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_402),
.Y(n_467)
);

INVx6_ASAP7_75t_L g468 ( 
.A(n_402),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_388),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_388),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_421),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_373),
.B(n_1),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_421),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_421),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_448),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_402),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_403),
.Y(n_477)
);

INVx5_ASAP7_75t_L g478 ( 
.A(n_403),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_421),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_361),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_403),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_324),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_341),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_374),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_423),
.B(n_8),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_375),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_381),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_306),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_284),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_394),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_422),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_456),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_295),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_349),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_273),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_403),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_274),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_355),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_392),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_409),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_300),
.B(n_8),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_409),
.Y(n_502)
);

OA21x2_ASAP7_75t_L g503 ( 
.A1(n_276),
.A2(n_9),
.B(n_10),
.Y(n_503)
);

INVx5_ASAP7_75t_L g504 ( 
.A(n_409),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_278),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_280),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_282),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_409),
.Y(n_508)
);

OA21x2_ASAP7_75t_L g509 ( 
.A1(n_283),
.A2(n_11),
.B(n_12),
.Y(n_509)
);

OA21x2_ASAP7_75t_L g510 ( 
.A1(n_285),
.A2(n_287),
.B(n_286),
.Y(n_510)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_415),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_364),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_423),
.B(n_16),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_288),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_290),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_294),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_399),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_415),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_415),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_353),
.B(n_17),
.Y(n_520)
);

OA21x2_ASAP7_75t_L g521 ( 
.A1(n_296),
.A2(n_18),
.B(n_19),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_404),
.B(n_18),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_382),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_415),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_460),
.B(n_22),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_410),
.Y(n_526)
);

OA21x2_ASAP7_75t_L g527 ( 
.A1(n_298),
.A2(n_23),
.B(n_24),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_304),
.Y(n_528)
);

OAI22x1_ASAP7_75t_SL g529 ( 
.A1(n_424),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_438),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_419),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_365),
.B(n_28),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_310),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_307),
.Y(n_534)
);

INVx1_ASAP7_75t_SL g535 ( 
.A(n_443),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_313),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_315),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_277),
.B(n_32),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_316),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_319),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_320),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_419),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_419),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_419),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_293),
.B(n_32),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_436),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_281),
.B(n_34),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_322),
.B(n_34),
.Y(n_548)
);

AND2x2_ASAP7_75t_SL g549 ( 
.A(n_291),
.B(n_41),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_455),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_321),
.Y(n_551)
);

INVx4_ASAP7_75t_L g552 ( 
.A(n_436),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_281),
.B(n_272),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_436),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_436),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_301),
.B(n_43),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_325),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_334),
.Y(n_558)
);

BUFx8_ASAP7_75t_L g559 ( 
.A(n_461),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_335),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_337),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_461),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_340),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_292),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_461),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_461),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_314),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_347),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_348),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_386),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_469),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_474),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_474),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_510),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_508),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_473),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_462),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_464),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_465),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_532),
.B(n_311),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_464),
.Y(n_581)
);

NAND2xp33_ASAP7_75t_L g582 ( 
.A(n_520),
.B(n_370),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_508),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_463),
.Y(n_584)
);

NAND2xp33_ASAP7_75t_L g585 ( 
.A(n_525),
.B(n_275),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_470),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_464),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_531),
.Y(n_588)
);

AND3x2_ASAP7_75t_L g589 ( 
.A(n_501),
.B(n_398),
.C(n_328),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_531),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_546),
.Y(n_591)
);

BUFx4f_ASAP7_75t_L g592 ( 
.A(n_510),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_546),
.Y(n_593)
);

OR2x6_ASAP7_75t_L g594 ( 
.A(n_532),
.B(n_328),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_565),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_489),
.Y(n_596)
);

OAI22xp33_ASAP7_75t_L g597 ( 
.A1(n_466),
.A2(n_439),
.B1(n_398),
.B2(n_317),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_SL g598 ( 
.A(n_549),
.B(n_434),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_471),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_565),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_559),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_479),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_569),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_502),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_569),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_564),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_493),
.B(n_498),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_493),
.B(n_326),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_468),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_482),
.A2(n_439),
.B1(n_302),
.B2(n_351),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_518),
.Y(n_611)
);

INVx5_ASAP7_75t_L g612 ( 
.A(n_478),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_489),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_468),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_524),
.Y(n_615)
);

NAND2xp33_ASAP7_75t_SL g616 ( 
.A(n_485),
.B(n_435),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_535),
.B(n_368),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_498),
.B(n_344),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_468),
.Y(n_619)
);

OR2x6_ASAP7_75t_L g620 ( 
.A(n_512),
.B(n_329),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_495),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_535),
.B(n_396),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_542),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_497),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_505),
.Y(n_625)
);

AO21x2_ASAP7_75t_L g626 ( 
.A1(n_485),
.A2(n_362),
.B(n_342),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_558),
.B(n_408),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_558),
.B(n_417),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_506),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_522),
.B(n_458),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_522),
.B(n_501),
.Y(n_631)
);

BUFx10_ASAP7_75t_L g632 ( 
.A(n_463),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_543),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_507),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_513),
.B(n_279),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_544),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_514),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_467),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_467),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_513),
.B(n_289),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_515),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_467),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_476),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_476),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_476),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_477),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_472),
.B(n_297),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_477),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_477),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_517),
.Y(n_650)
);

BUFx4f_ASAP7_75t_L g651 ( 
.A(n_549),
.Y(n_651)
);

OAI22xp33_ASAP7_75t_SL g652 ( 
.A1(n_545),
.A2(n_459),
.B1(n_454),
.B2(n_450),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_481),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_516),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_481),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_SL g656 ( 
.A1(n_620),
.A2(n_512),
.B1(n_523),
.B2(n_556),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_617),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_622),
.B(n_494),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_638),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_621),
.Y(n_660)
);

OR2x2_ASAP7_75t_SL g661 ( 
.A(n_597),
.B(n_545),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_581),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_624),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_594),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_638),
.Y(n_665)
);

INVxp67_ASAP7_75t_L g666 ( 
.A(n_627),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_574),
.B(n_555),
.Y(n_667)
);

NAND2xp33_ASAP7_75t_L g668 ( 
.A(n_580),
.B(n_553),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_581),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_574),
.B(n_555),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_639),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_580),
.B(n_517),
.Y(n_672)
);

AO221x1_ASAP7_75t_L g673 ( 
.A1(n_597),
.A2(n_533),
.B1(n_372),
.B2(n_380),
.C(n_383),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_625),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_626),
.B(n_631),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_589),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_626),
.B(n_528),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_627),
.B(n_628),
.Y(n_678)
);

INVx4_ASAP7_75t_L g679 ( 
.A(n_612),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_631),
.B(n_575),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_607),
.B(n_499),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_629),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_589),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_639),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_642),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_635),
.B(n_640),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_628),
.B(n_530),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_651),
.A2(n_538),
.B1(n_548),
.B2(n_472),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_575),
.B(n_534),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_598),
.A2(n_530),
.B1(n_475),
.B2(n_488),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_583),
.B(n_536),
.Y(n_691)
);

AO221x1_ASAP7_75t_L g692 ( 
.A1(n_610),
.A2(n_533),
.B1(n_357),
.B2(n_366),
.C(n_369),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_642),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_596),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_635),
.B(n_488),
.Y(n_695)
);

NAND2x1p5_ASAP7_75t_L g696 ( 
.A(n_651),
.B(n_503),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_594),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_581),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_644),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_594),
.A2(n_548),
.B1(n_538),
.B2(n_509),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_583),
.B(n_588),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_609),
.B(n_484),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_644),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_581),
.Y(n_704)
);

INVxp67_ASAP7_75t_L g705 ( 
.A(n_613),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_630),
.A2(n_503),
.B1(n_527),
.B2(n_509),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_630),
.A2(n_521),
.B1(n_527),
.B2(n_570),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_650),
.B(n_553),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_650),
.B(n_526),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_634),
.B(n_526),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_652),
.B(n_550),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_646),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_637),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_614),
.B(n_491),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_608),
.B(n_550),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_588),
.B(n_537),
.Y(n_716)
);

OAI221xp5_ASAP7_75t_L g717 ( 
.A1(n_582),
.A2(n_547),
.B1(n_570),
.B2(n_483),
.C(n_561),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_590),
.B(n_539),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_590),
.B(n_541),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_645),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_591),
.B(n_551),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_640),
.B(n_567),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_619),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_601),
.B(n_547),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_641),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_654),
.B(n_540),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_645),
.Y(n_727)
);

NAND2xp33_ASAP7_75t_L g728 ( 
.A(n_616),
.B(n_299),
.Y(n_728)
);

NOR3xp33_ASAP7_75t_L g729 ( 
.A(n_616),
.B(n_563),
.C(n_560),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_601),
.B(n_303),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_L g731 ( 
.A1(n_620),
.A2(n_492),
.B1(n_486),
.B2(n_490),
.Y(n_731)
);

INVxp67_ASAP7_75t_L g732 ( 
.A(n_620),
.Y(n_732)
);

NOR2xp67_ASAP7_75t_L g733 ( 
.A(n_584),
.B(n_478),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_L g734 ( 
.A(n_618),
.B(n_305),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_648),
.Y(n_735)
);

NOR2x1p5_ASAP7_75t_L g736 ( 
.A(n_577),
.B(n_480),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_702),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_675),
.B(n_592),
.Y(n_738)
);

A2O1A1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_686),
.A2(n_592),
.B(n_647),
.C(n_585),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_675),
.B(n_647),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_658),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_657),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_681),
.Y(n_743)
);

AOI21x1_ASAP7_75t_L g744 ( 
.A1(n_667),
.A2(n_593),
.B(n_591),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_702),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_667),
.A2(n_670),
.B(n_680),
.Y(n_746)
);

NOR2x1_ASAP7_75t_L g747 ( 
.A(n_708),
.B(n_447),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_666),
.B(n_606),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_723),
.Y(n_749)
);

BUFx2_ASAP7_75t_SL g750 ( 
.A(n_733),
.Y(n_750)
);

O2A1O1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_668),
.A2(n_557),
.B(n_568),
.C(n_540),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_670),
.A2(n_680),
.B(n_677),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_678),
.B(n_648),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_714),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_661),
.A2(n_521),
.B1(n_486),
.B2(n_492),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_687),
.B(n_649),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_714),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_688),
.B(n_649),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_672),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_677),
.A2(n_612),
.B(n_504),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_660),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_700),
.B(n_604),
.Y(n_762)
);

A2O1A1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_695),
.A2(n_425),
.B(n_426),
.C(n_416),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_710),
.B(n_632),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_706),
.B(n_604),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_663),
.Y(n_766)
);

NAND3xp33_ASAP7_75t_L g767 ( 
.A(n_729),
.B(n_568),
.C(n_557),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_701),
.A2(n_691),
.B(n_689),
.Y(n_768)
);

A2O1A1Ixp33_ASAP7_75t_L g769 ( 
.A1(n_722),
.A2(n_413),
.B(n_429),
.C(n_430),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_707),
.B(n_611),
.Y(n_770)
);

BUFx2_ASAP7_75t_L g771 ( 
.A(n_732),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_701),
.A2(n_612),
.B(n_504),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_674),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_689),
.A2(n_612),
.B(n_504),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_691),
.A2(n_504),
.B(n_478),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_716),
.A2(n_478),
.B(n_593),
.Y(n_776)
);

OAI22xp33_ASAP7_75t_SL g777 ( 
.A1(n_717),
.A2(n_411),
.B1(n_350),
.B2(n_385),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_682),
.B(n_611),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_715),
.B(n_308),
.Y(n_779)
);

NOR2xp67_ASAP7_75t_L g780 ( 
.A(n_694),
.B(n_579),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_713),
.B(n_725),
.Y(n_781)
);

O2A1O1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_731),
.A2(n_490),
.B(n_339),
.C(n_603),
.Y(n_782)
);

INVxp67_ASAP7_75t_L g783 ( 
.A(n_726),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_659),
.B(n_615),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_R g785 ( 
.A(n_728),
.B(n_606),
.Y(n_785)
);

O2A1O1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_731),
.A2(n_605),
.B(n_433),
.C(n_444),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_727),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_696),
.B(n_595),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_716),
.A2(n_600),
.B(n_595),
.Y(n_789)
);

CKINVDCx8_ASAP7_75t_R g790 ( 
.A(n_692),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_705),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_718),
.A2(n_600),
.B(n_615),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_718),
.A2(n_633),
.B(n_623),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_696),
.B(n_623),
.Y(n_794)
);

NAND3xp33_ASAP7_75t_L g795 ( 
.A(n_690),
.B(n_599),
.C(n_586),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_719),
.A2(n_636),
.B(n_633),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_719),
.A2(n_636),
.B(n_573),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_665),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_671),
.B(n_572),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_721),
.A2(n_573),
.B(n_572),
.Y(n_800)
);

OAI21xp5_ASAP7_75t_L g801 ( 
.A1(n_711),
.A2(n_391),
.B(n_389),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_684),
.B(n_578),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_697),
.A2(n_318),
.B1(n_309),
.B2(n_312),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_SL g804 ( 
.A(n_664),
.B(n_632),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_709),
.B(n_480),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_721),
.A2(n_602),
.B(n_646),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_676),
.B(n_323),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_685),
.B(n_578),
.Y(n_808)
);

BUFx12f_ASAP7_75t_L g809 ( 
.A(n_683),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_693),
.B(n_587),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_734),
.A2(n_327),
.B1(n_330),
.B2(n_331),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_699),
.B(n_587),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_703),
.B(n_643),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_662),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_720),
.A2(n_653),
.B(n_646),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_735),
.A2(n_653),
.B(n_646),
.Y(n_816)
);

OAI21x1_ASAP7_75t_L g817 ( 
.A1(n_744),
.A2(n_704),
.B(n_669),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_740),
.B(n_724),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_740),
.B(n_669),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_752),
.A2(n_698),
.B(n_662),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_759),
.B(n_704),
.Y(n_821)
);

NOR2xp67_ASAP7_75t_L g822 ( 
.A(n_795),
.B(n_571),
.Y(n_822)
);

OAI21x1_ASAP7_75t_L g823 ( 
.A1(n_746),
.A2(n_736),
.B(n_730),
.Y(n_823)
);

AOI221x1_ASAP7_75t_L g824 ( 
.A1(n_755),
.A2(n_414),
.B1(n_432),
.B2(n_446),
.C(n_427),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_742),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_738),
.A2(n_371),
.B(n_358),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_738),
.A2(n_418),
.B(n_576),
.Y(n_827)
);

NAND3xp33_ASAP7_75t_L g828 ( 
.A(n_739),
.B(n_333),
.C(n_332),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_761),
.Y(n_829)
);

NAND2x1_ASAP7_75t_L g830 ( 
.A(n_814),
.B(n_662),
.Y(n_830)
);

OR2x2_ASAP7_75t_L g831 ( 
.A(n_741),
.B(n_656),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_766),
.Y(n_832)
);

INVxp67_ASAP7_75t_SL g833 ( 
.A(n_814),
.Y(n_833)
);

AOI22xp5_ASAP7_75t_L g834 ( 
.A1(n_755),
.A2(n_673),
.B1(n_336),
.B2(n_420),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_801),
.A2(n_407),
.B(n_343),
.C(n_345),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_768),
.A2(n_751),
.B(n_747),
.C(n_758),
.Y(n_836)
);

NOR2x1_ASAP7_75t_R g837 ( 
.A(n_743),
.B(n_791),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_777),
.A2(n_437),
.B1(n_346),
.B2(n_352),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_753),
.B(n_698),
.Y(n_839)
);

OAI21x1_ASAP7_75t_L g840 ( 
.A1(n_788),
.A2(n_655),
.B(n_643),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_765),
.A2(n_770),
.B(n_788),
.Y(n_841)
);

OAI21x1_ASAP7_75t_L g842 ( 
.A1(n_794),
.A2(n_655),
.B(n_487),
.Y(n_842)
);

OAI21xp5_ASAP7_75t_L g843 ( 
.A1(n_794),
.A2(n_440),
.B(n_354),
.Y(n_843)
);

OAI21x1_ASAP7_75t_L g844 ( 
.A1(n_789),
.A2(n_487),
.B(n_712),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_773),
.Y(n_845)
);

OAI21x1_ASAP7_75t_L g846 ( 
.A1(n_800),
.A2(n_698),
.B(n_712),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_756),
.B(n_712),
.Y(n_847)
);

OAI21x1_ASAP7_75t_L g848 ( 
.A1(n_797),
.A2(n_47),
.B(n_48),
.Y(n_848)
);

BUFx2_ASAP7_75t_L g849 ( 
.A(n_764),
.Y(n_849)
);

INVxp67_ASAP7_75t_SL g850 ( 
.A(n_814),
.Y(n_850)
);

OAI21xp33_ASAP7_75t_L g851 ( 
.A1(n_769),
.A2(n_406),
.B(n_356),
.Y(n_851)
);

BUFx10_ASAP7_75t_L g852 ( 
.A(n_748),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_778),
.Y(n_853)
);

NAND3xp33_ASAP7_75t_SL g854 ( 
.A(n_785),
.B(n_405),
.C(n_359),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_783),
.B(n_338),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_805),
.B(n_360),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_781),
.B(n_363),
.Y(n_857)
);

AO31x2_ASAP7_75t_L g858 ( 
.A1(n_763),
.A2(n_511),
.A3(n_519),
.B(n_552),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_790),
.B(n_367),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_762),
.B(n_376),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_760),
.A2(n_679),
.B(n_653),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_749),
.B(n_51),
.Y(n_862)
);

AND2x2_ASAP7_75t_SL g863 ( 
.A(n_804),
.B(n_529),
.Y(n_863)
);

BUFx2_ASAP7_75t_L g864 ( 
.A(n_809),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_787),
.Y(n_865)
);

NAND2x1p5_ASAP7_75t_L g866 ( 
.A(n_737),
.B(n_653),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_798),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_807),
.A2(n_442),
.B1(n_378),
.B2(n_379),
.Y(n_868)
);

BUFx4_ASAP7_75t_SL g869 ( 
.A(n_771),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_799),
.A2(n_679),
.B(n_566),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_745),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_750),
.B(n_377),
.Y(n_872)
);

INVxp67_ASAP7_75t_SL g873 ( 
.A(n_754),
.Y(n_873)
);

AOI211x1_ASAP7_75t_L g874 ( 
.A1(n_767),
.A2(n_793),
.B(n_796),
.C(n_792),
.Y(n_874)
);

OAI21x1_ASAP7_75t_L g875 ( 
.A1(n_806),
.A2(n_810),
.B(n_802),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_818),
.B(n_779),
.Y(n_876)
);

OAI21x1_ASAP7_75t_L g877 ( 
.A1(n_840),
.A2(n_816),
.B(n_808),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_829),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_832),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_834),
.A2(n_757),
.B1(n_784),
.B2(n_803),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_856),
.A2(n_780),
.B1(n_811),
.B2(n_812),
.Y(n_881)
);

OAI21x1_ASAP7_75t_L g882 ( 
.A1(n_842),
.A2(n_813),
.B(n_815),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_849),
.B(n_782),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_834),
.A2(n_559),
.B1(n_384),
.B2(n_453),
.Y(n_884)
);

OAI21x1_ASAP7_75t_L g885 ( 
.A1(n_817),
.A2(n_776),
.B(n_786),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_853),
.B(n_387),
.Y(n_886)
);

OAI21x1_ASAP7_75t_L g887 ( 
.A1(n_875),
.A2(n_772),
.B(n_774),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_871),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_841),
.A2(n_775),
.B(n_566),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_844),
.Y(n_890)
);

AOI21x1_ASAP7_75t_L g891 ( 
.A1(n_820),
.A2(n_566),
.B(n_562),
.Y(n_891)
);

OAI21xp5_ASAP7_75t_L g892 ( 
.A1(n_836),
.A2(n_431),
.B(n_395),
.Y(n_892)
);

AOI221xp5_ASAP7_75t_L g893 ( 
.A1(n_831),
.A2(n_452),
.B1(n_397),
.B2(n_401),
.C(n_412),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_871),
.B(n_53),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_845),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_865),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_852),
.B(n_390),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_867),
.Y(n_898)
);

OAI21x1_ASAP7_75t_L g899 ( 
.A1(n_846),
.A2(n_57),
.B(n_60),
.Y(n_899)
);

INVxp67_ASAP7_75t_SL g900 ( 
.A(n_833),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_871),
.B(n_64),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_857),
.B(n_428),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_830),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_869),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_828),
.A2(n_441),
.B1(n_449),
.B2(n_451),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_828),
.A2(n_457),
.B(n_519),
.Y(n_906)
);

OAI222xp33_ASAP7_75t_L g907 ( 
.A1(n_838),
.A2(n_400),
.B1(n_552),
.B2(n_511),
.C1(n_77),
.C2(n_78),
.Y(n_907)
);

AOI21xp33_ASAP7_75t_SL g908 ( 
.A1(n_863),
.A2(n_825),
.B(n_859),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_819),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_873),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_874),
.Y(n_911)
);

A2O1A1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_826),
.A2(n_562),
.B(n_554),
.C(n_500),
.Y(n_912)
);

OR2x2_ASAP7_75t_L g913 ( 
.A(n_855),
.B(n_67),
.Y(n_913)
);

AOI221xp5_ASAP7_75t_L g914 ( 
.A1(n_868),
.A2(n_562),
.B1(n_554),
.B2(n_500),
.C(n_496),
.Y(n_914)
);

OAI21x1_ASAP7_75t_L g915 ( 
.A1(n_823),
.A2(n_68),
.B(n_75),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_874),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_827),
.A2(n_79),
.B(n_82),
.Y(n_917)
);

OA21x2_ASAP7_75t_L g918 ( 
.A1(n_824),
.A2(n_554),
.B(n_500),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_862),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_909),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_878),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_900),
.Y(n_922)
);

OA21x2_ASAP7_75t_L g923 ( 
.A1(n_911),
.A2(n_916),
.B(n_890),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_909),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_879),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_876),
.B(n_862),
.Y(n_926)
);

AOI222xp33_ASAP7_75t_L g927 ( 
.A1(n_884),
.A2(n_837),
.B1(n_852),
.B2(n_854),
.C1(n_843),
.C2(n_851),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_888),
.Y(n_928)
);

INVx5_ASAP7_75t_L g929 ( 
.A(n_888),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_895),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_896),
.Y(n_931)
);

OAI21x1_ASAP7_75t_L g932 ( 
.A1(n_899),
.A2(n_915),
.B(n_887),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_888),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_898),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_910),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_919),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_900),
.Y(n_937)
);

NOR2x1_ASAP7_75t_L g938 ( 
.A(n_913),
.B(n_872),
.Y(n_938)
);

BUFx5_ASAP7_75t_L g939 ( 
.A(n_894),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_917),
.A2(n_847),
.B(n_839),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_919),
.B(n_894),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_919),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_894),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_888),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_911),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_904),
.Y(n_946)
);

OA21x2_ASAP7_75t_L g947 ( 
.A1(n_916),
.A2(n_848),
.B(n_860),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_876),
.A2(n_835),
.B(n_822),
.Y(n_948)
);

NAND2x1p5_ASAP7_75t_L g949 ( 
.A(n_901),
.B(n_822),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_919),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_901),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_890),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_901),
.B(n_850),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_891),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_883),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_903),
.B(n_821),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_886),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_955),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_923),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_926),
.B(n_884),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_946),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_957),
.B(n_908),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_923),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_929),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_926),
.B(n_837),
.Y(n_965)
);

INVxp67_ASAP7_75t_SL g966 ( 
.A(n_922),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_923),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_920),
.B(n_897),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_945),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_952),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_920),
.B(n_897),
.Y(n_971)
);

NAND2x1p5_ASAP7_75t_L g972 ( 
.A(n_922),
.B(n_885),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_924),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_941),
.B(n_903),
.Y(n_974)
);

OR2x2_ASAP7_75t_L g975 ( 
.A(n_937),
.B(n_892),
.Y(n_975)
);

INVx4_ASAP7_75t_R g976 ( 
.A(n_951),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_924),
.B(n_880),
.Y(n_977)
);

BUFx2_ASAP7_75t_L g978 ( 
.A(n_951),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_945),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_943),
.B(n_921),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_921),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_931),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_952),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_931),
.B(n_880),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_939),
.B(n_858),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_939),
.B(n_858),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_932),
.Y(n_987)
);

HB1xp67_ASAP7_75t_L g988 ( 
.A(n_928),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_939),
.B(n_858),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_939),
.B(n_906),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_925),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_939),
.B(n_902),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_929),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_933),
.Y(n_994)
);

AOI22xp33_ASAP7_75t_SL g995 ( 
.A1(n_939),
.A2(n_907),
.B1(n_864),
.B2(n_918),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_939),
.B(n_949),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_991),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_959),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_991),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_977),
.B(n_925),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_959),
.Y(n_1001)
);

BUFx2_ASAP7_75t_SL g1002 ( 
.A(n_958),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_969),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_969),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_980),
.B(n_930),
.Y(n_1005)
);

OR2x2_ASAP7_75t_L g1006 ( 
.A(n_968),
.B(n_930),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_980),
.B(n_948),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_978),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_984),
.B(n_934),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_984),
.B(n_941),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_979),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_988),
.Y(n_1012)
);

INVx4_ASAP7_75t_R g1013 ( 
.A(n_993),
.Y(n_1013)
);

INVxp67_ASAP7_75t_SL g1014 ( 
.A(n_966),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_971),
.B(n_935),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_960),
.B(n_938),
.Y(n_1016)
);

OR2x2_ASAP7_75t_L g1017 ( 
.A(n_977),
.B(n_947),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_979),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_960),
.B(n_941),
.Y(n_1019)
);

INVx5_ASAP7_75t_L g1020 ( 
.A(n_963),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_981),
.B(n_949),
.Y(n_1021)
);

OR2x2_ASAP7_75t_L g1022 ( 
.A(n_967),
.B(n_947),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_981),
.B(n_949),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_983),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_959),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_983),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_973),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_982),
.B(n_944),
.Y(n_1028)
);

INVx4_ASAP7_75t_L g1029 ( 
.A(n_993),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_982),
.B(n_947),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_962),
.B(n_994),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_996),
.B(n_953),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_996),
.B(n_953),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_992),
.B(n_927),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_963),
.Y(n_1035)
);

OR2x2_ASAP7_75t_L g1036 ( 
.A(n_967),
.B(n_940),
.Y(n_1036)
);

OR2x2_ASAP7_75t_L g1037 ( 
.A(n_975),
.B(n_954),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1034),
.B(n_973),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_997),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_1007),
.B(n_963),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_1007),
.B(n_963),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_1019),
.B(n_985),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1016),
.B(n_990),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_1031),
.B(n_990),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_1037),
.B(n_975),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_1019),
.B(n_985),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_1015),
.A2(n_965),
.B1(n_995),
.B2(n_905),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1009),
.B(n_978),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_1008),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_1006),
.B(n_974),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_999),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_1010),
.B(n_1033),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1003),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_1037),
.B(n_972),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_998),
.Y(n_1055)
);

NAND2x1_ASAP7_75t_L g1056 ( 
.A(n_1013),
.B(n_976),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_1032),
.B(n_986),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_1010),
.B(n_986),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1004),
.Y(n_1059)
);

NOR3xp33_ASAP7_75t_L g1060 ( 
.A(n_1012),
.B(n_893),
.C(n_851),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1011),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_1033),
.B(n_989),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_1009),
.B(n_989),
.Y(n_1063)
);

OR2x2_ASAP7_75t_L g1064 ( 
.A(n_1000),
.B(n_972),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1018),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1024),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_1017),
.B(n_972),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_1017),
.B(n_987),
.Y(n_1068)
);

INVx2_ASAP7_75t_SL g1069 ( 
.A(n_1008),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1026),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1039),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1051),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_1040),
.B(n_1035),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1053),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_1049),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_1040),
.B(n_1035),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_SL g1077 ( 
.A(n_1047),
.B(n_961),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_1041),
.B(n_998),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1044),
.B(n_1014),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1059),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_1041),
.B(n_1001),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1061),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1043),
.B(n_1002),
.Y(n_1083)
);

INVxp67_ASAP7_75t_SL g1084 ( 
.A(n_1045),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1067),
.B(n_1001),
.Y(n_1085)
);

INVx2_ASAP7_75t_SL g1086 ( 
.A(n_1049),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_1055),
.Y(n_1087)
);

NAND2x1p5_ASAP7_75t_L g1088 ( 
.A(n_1056),
.B(n_1020),
.Y(n_1088)
);

OR2x2_ASAP7_75t_L g1089 ( 
.A(n_1068),
.B(n_1036),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1055),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1065),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1038),
.B(n_1000),
.Y(n_1092)
);

AOI332xp33_ASAP7_75t_L g1093 ( 
.A1(n_1071),
.A2(n_1070),
.A3(n_1066),
.B1(n_1048),
.B2(n_1005),
.B3(n_1068),
.C1(n_1063),
.C2(n_1067),
.Y(n_1093)
);

OAI211xp5_ASAP7_75t_L g1094 ( 
.A1(n_1077),
.A2(n_1060),
.B(n_905),
.C(n_1050),
.Y(n_1094)
);

INVx1_ASAP7_75t_SL g1095 ( 
.A(n_1083),
.Y(n_1095)
);

AOI21xp33_ASAP7_75t_L g1096 ( 
.A1(n_1079),
.A2(n_1050),
.B(n_1036),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_1084),
.B(n_1085),
.Y(n_1097)
);

OR2x2_ASAP7_75t_L g1098 ( 
.A(n_1089),
.B(n_1064),
.Y(n_1098)
);

OAI32xp33_ASAP7_75t_L g1099 ( 
.A1(n_1092),
.A2(n_1054),
.A3(n_1069),
.B1(n_1063),
.B2(n_1062),
.Y(n_1099)
);

AOI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1088),
.A2(n_1032),
.B1(n_1057),
.B2(n_974),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1089),
.B(n_1069),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_1085),
.B(n_1062),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_1075),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_1086),
.B(n_1075),
.Y(n_1104)
);

NAND2xp33_ASAP7_75t_L g1105 ( 
.A(n_1088),
.B(n_946),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1072),
.Y(n_1106)
);

OR2x2_ASAP7_75t_L g1107 ( 
.A(n_1073),
.B(n_1042),
.Y(n_1107)
);

AOI22xp33_ASAP7_75t_SL g1108 ( 
.A1(n_1088),
.A2(n_1057),
.B1(n_1032),
.B2(n_1029),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1074),
.B(n_1058),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1073),
.B(n_1057),
.Y(n_1110)
);

OR2x2_ASAP7_75t_L g1111 ( 
.A(n_1076),
.B(n_1042),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1080),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1076),
.B(n_1046),
.Y(n_1113)
);

INVxp67_ASAP7_75t_L g1114 ( 
.A(n_1101),
.Y(n_1114)
);

OAI21xp33_ASAP7_75t_SL g1115 ( 
.A1(n_1100),
.A2(n_1086),
.B(n_1091),
.Y(n_1115)
);

OAI21xp33_ASAP7_75t_L g1116 ( 
.A1(n_1094),
.A2(n_1082),
.B(n_1046),
.Y(n_1116)
);

INVx2_ASAP7_75t_SL g1117 ( 
.A(n_1104),
.Y(n_1117)
);

O2A1O1Ixp5_ASAP7_75t_L g1118 ( 
.A1(n_1094),
.A2(n_1087),
.B(n_1090),
.C(n_1081),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1106),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_1104),
.Y(n_1120)
);

NAND3xp33_ASAP7_75t_L g1121 ( 
.A(n_1096),
.B(n_1021),
.C(n_1023),
.Y(n_1121)
);

NAND3xp33_ASAP7_75t_L g1122 ( 
.A(n_1096),
.B(n_1021),
.C(n_1023),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_1095),
.B(n_1052),
.Y(n_1123)
);

NAND2xp33_ASAP7_75t_SL g1124 ( 
.A(n_1105),
.B(n_1052),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1112),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_1093),
.A2(n_1058),
.B(n_1081),
.C(n_1078),
.Y(n_1126)
);

AOI222xp33_ASAP7_75t_L g1127 ( 
.A1(n_1099),
.A2(n_1005),
.B1(n_1078),
.B2(n_914),
.C1(n_1027),
.C2(n_1090),
.Y(n_1127)
);

OAI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_1109),
.A2(n_1029),
.B1(n_1020),
.B2(n_1028),
.Y(n_1128)
);

INVx1_ASAP7_75t_SL g1129 ( 
.A(n_1101),
.Y(n_1129)
);

OAI211xp5_ASAP7_75t_L g1130 ( 
.A1(n_1108),
.A2(n_1087),
.B(n_881),
.C(n_1029),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1098),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_1110),
.B(n_1020),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1116),
.A2(n_1109),
.B1(n_1111),
.B2(n_1107),
.Y(n_1133)
);

AO22x1_ASAP7_75t_L g1134 ( 
.A1(n_1120),
.A2(n_1103),
.B1(n_1097),
.B2(n_1102),
.Y(n_1134)
);

AOI21xp33_ASAP7_75t_L g1135 ( 
.A1(n_1130),
.A2(n_974),
.B(n_1113),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_1114),
.B(n_936),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_1118),
.A2(n_993),
.B(n_974),
.C(n_953),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_1115),
.A2(n_912),
.B(n_936),
.C(n_942),
.Y(n_1138)
);

AOI21xp33_ASAP7_75t_L g1139 ( 
.A1(n_1128),
.A2(n_964),
.B(n_1020),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1119),
.Y(n_1140)
);

NOR4xp25_ASAP7_75t_L g1141 ( 
.A(n_1126),
.B(n_912),
.C(n_1025),
.D(n_1030),
.Y(n_1141)
);

AOI211xp5_ASAP7_75t_L g1142 ( 
.A1(n_1124),
.A2(n_950),
.B(n_942),
.C(n_956),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1121),
.A2(n_1122),
.B(n_1129),
.Y(n_1143)
);

OAI221xp5_ASAP7_75t_L g1144 ( 
.A1(n_1117),
.A2(n_964),
.B1(n_1020),
.B2(n_866),
.C(n_1025),
.Y(n_1144)
);

NAND3xp33_ASAP7_75t_L g1145 ( 
.A(n_1127),
.B(n_956),
.C(n_889),
.Y(n_1145)
);

NAND3xp33_ASAP7_75t_L g1146 ( 
.A(n_1125),
.B(n_956),
.C(n_1030),
.Y(n_1146)
);

O2A1O1Ixp5_ASAP7_75t_L g1147 ( 
.A1(n_1131),
.A2(n_970),
.B(n_1022),
.C(n_987),
.Y(n_1147)
);

OAI21xp33_ASAP7_75t_L g1148 ( 
.A1(n_1123),
.A2(n_1132),
.B(n_1022),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_1132),
.B(n_970),
.Y(n_1149)
);

NOR3xp33_ASAP7_75t_L g1150 ( 
.A(n_1116),
.B(n_970),
.C(n_932),
.Y(n_1150)
);

AOI222xp33_ASAP7_75t_L g1151 ( 
.A1(n_1116),
.A2(n_496),
.B1(n_481),
.B2(n_954),
.C1(n_987),
.C2(n_929),
.Y(n_1151)
);

NAND4xp25_ASAP7_75t_SL g1152 ( 
.A(n_1115),
.B(n_976),
.C(n_861),
.D(n_91),
.Y(n_1152)
);

NOR3xp33_ASAP7_75t_L g1153 ( 
.A(n_1116),
.B(n_882),
.C(n_877),
.Y(n_1153)
);

OAI221xp5_ASAP7_75t_L g1154 ( 
.A1(n_1141),
.A2(n_496),
.B1(n_929),
.B2(n_870),
.C(n_918),
.Y(n_1154)
);

AOI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1134),
.A2(n_918),
.B(n_929),
.Y(n_1155)
);

NOR3xp33_ASAP7_75t_L g1156 ( 
.A(n_1145),
.B(n_1152),
.C(n_1139),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_1133),
.B(n_87),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1140),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1142),
.B(n_268),
.Y(n_1159)
);

NOR3xp33_ASAP7_75t_L g1160 ( 
.A(n_1150),
.B(n_90),
.C(n_92),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1143),
.B(n_93),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1138),
.A2(n_97),
.B(n_101),
.Y(n_1162)
);

NOR2x1_ASAP7_75t_L g1163 ( 
.A(n_1136),
.B(n_107),
.Y(n_1163)
);

NAND3xp33_ASAP7_75t_L g1164 ( 
.A(n_1156),
.B(n_1151),
.C(n_1153),
.Y(n_1164)
);

NOR3xp33_ASAP7_75t_L g1165 ( 
.A(n_1161),
.B(n_1144),
.C(n_1135),
.Y(n_1165)
);

NAND4xp75_ASAP7_75t_L g1166 ( 
.A(n_1162),
.B(n_1147),
.C(n_1149),
.D(n_1137),
.Y(n_1166)
);

NAND4xp75_ASAP7_75t_L g1167 ( 
.A(n_1163),
.B(n_1148),
.C(n_1146),
.D(n_115),
.Y(n_1167)
);

NAND3xp33_ASAP7_75t_L g1168 ( 
.A(n_1160),
.B(n_108),
.C(n_109),
.Y(n_1168)
);

NOR3xp33_ASAP7_75t_L g1169 ( 
.A(n_1157),
.B(n_1159),
.C(n_1158),
.Y(n_1169)
);

NAND4xp75_ASAP7_75t_L g1170 ( 
.A(n_1154),
.B(n_116),
.C(n_118),
.D(n_123),
.Y(n_1170)
);

AOI211xp5_ASAP7_75t_SL g1171 ( 
.A1(n_1155),
.A2(n_125),
.B(n_127),
.C(n_128),
.Y(n_1171)
);

NOR2x1_ASAP7_75t_L g1172 ( 
.A(n_1161),
.B(n_129),
.Y(n_1172)
);

OAI211xp5_ASAP7_75t_L g1173 ( 
.A1(n_1156),
.A2(n_131),
.B(n_133),
.C(n_140),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_1172),
.B(n_142),
.Y(n_1174)
);

INVxp67_ASAP7_75t_L g1175 ( 
.A(n_1169),
.Y(n_1175)
);

NOR2x1_ASAP7_75t_L g1176 ( 
.A(n_1173),
.B(n_147),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1164),
.A2(n_151),
.B1(n_154),
.B2(n_158),
.Y(n_1177)
);

OAI21xp33_ASAP7_75t_L g1178 ( 
.A1(n_1165),
.A2(n_161),
.B(n_162),
.Y(n_1178)
);

NAND4xp75_ASAP7_75t_L g1179 ( 
.A(n_1171),
.B(n_166),
.C(n_167),
.D(n_171),
.Y(n_1179)
);

NOR2xp67_ASAP7_75t_L g1180 ( 
.A(n_1168),
.B(n_175),
.Y(n_1180)
);

XOR2xp5_ASAP7_75t_L g1181 ( 
.A(n_1177),
.B(n_1179),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1174),
.Y(n_1182)
);

NAND4xp75_ASAP7_75t_L g1183 ( 
.A(n_1176),
.B(n_1166),
.C(n_1167),
.D(n_1170),
.Y(n_1183)
);

NAND4xp75_ASAP7_75t_L g1184 ( 
.A(n_1180),
.B(n_177),
.C(n_186),
.D(n_187),
.Y(n_1184)
);

XOR2xp5_ASAP7_75t_L g1185 ( 
.A(n_1175),
.B(n_196),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1178),
.Y(n_1186)
);

NOR2x1_ASAP7_75t_L g1187 ( 
.A(n_1174),
.B(n_216),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1187),
.Y(n_1188)
);

XNOR2xp5_ASAP7_75t_L g1189 ( 
.A(n_1185),
.B(n_267),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1182),
.Y(n_1190)
);

AOI21xp33_ASAP7_75t_SL g1191 ( 
.A1(n_1188),
.A2(n_1181),
.B(n_1186),
.Y(n_1191)
);

INVx1_ASAP7_75t_SL g1192 ( 
.A(n_1190),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1192),
.Y(n_1193)
);

INVxp67_ASAP7_75t_L g1194 ( 
.A(n_1191),
.Y(n_1194)
);

OA21x2_ASAP7_75t_L g1195 ( 
.A1(n_1194),
.A2(n_1183),
.B(n_1189),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1193),
.A2(n_1184),
.B1(n_222),
.B2(n_226),
.Y(n_1196)
);

OR2x6_ASAP7_75t_L g1197 ( 
.A(n_1195),
.B(n_220),
.Y(n_1197)
);

AOI221xp5_ASAP7_75t_L g1198 ( 
.A1(n_1196),
.A2(n_227),
.B1(n_228),
.B2(n_233),
.C(n_235),
.Y(n_1198)
);

OR2x6_ASAP7_75t_L g1199 ( 
.A(n_1197),
.B(n_237),
.Y(n_1199)
);

AO21x1_ASAP7_75t_L g1200 ( 
.A1(n_1199),
.A2(n_1198),
.B(n_239),
.Y(n_1200)
);

AOI221xp5_ASAP7_75t_L g1201 ( 
.A1(n_1200),
.A2(n_238),
.B1(n_246),
.B2(n_248),
.C(n_249),
.Y(n_1201)
);


endmodule