module real_aes_3_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_519;
wire n_92;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_119;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_0), .B(n_226), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_1), .A2(n_221), .B(n_268), .Y(n_267) );
AO22x2_ASAP7_75t_L g102 ( .A1(n_2), .A2(n_50), .B1(n_90), .B2(n_103), .Y(n_102) );
OAI22xp5_ASAP7_75t_L g79 ( .A1(n_3), .A2(n_80), .B1(n_81), .B2(n_180), .Y(n_79) );
INVx1_ASAP7_75t_L g180 ( .A(n_3), .Y(n_180) );
AOI22xp5_ASAP7_75t_L g163 ( .A1(n_4), .A2(n_21), .B1(n_164), .B2(n_167), .Y(n_163) );
INVx1_ASAP7_75t_L g201 ( .A(n_5), .Y(n_201) );
INVx1_ASAP7_75t_L g119 ( .A(n_6), .Y(n_119) );
INVx1_ASAP7_75t_L g156 ( .A(n_7), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_8), .B(n_237), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_9), .B(n_237), .Y(n_276) );
INVx1_ASAP7_75t_L g105 ( .A(n_10), .Y(n_105) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_11), .A2(n_25), .B1(n_90), .B2(n_100), .Y(n_99) );
NAND2xp33_ASAP7_75t_L g288 ( .A(n_12), .B(n_235), .Y(n_288) );
INVx2_ASAP7_75t_L g218 ( .A(n_13), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_14), .A2(n_184), .B1(n_185), .B2(n_186), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_14), .Y(n_184) );
AOI221x1_ASAP7_75t_L g220 ( .A1(n_14), .A2(n_22), .B1(n_221), .B2(n_226), .C(n_233), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_15), .B(n_226), .Y(n_284) );
AO21x2_ASAP7_75t_L g281 ( .A1(n_16), .A2(n_282), .B(n_283), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_17), .B(n_216), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_18), .B(n_237), .Y(n_296) );
AO21x1_ASAP7_75t_L g307 ( .A1(n_19), .A2(n_226), .B(n_308), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g186 ( .A1(n_20), .A2(n_38), .B1(n_187), .B2(n_188), .Y(n_186) );
INVx1_ASAP7_75t_L g188 ( .A(n_20), .Y(n_188) );
NAND2x1_ASAP7_75t_L g245 ( .A(n_23), .B(n_237), .Y(n_245) );
NAND2x1_ASAP7_75t_L g275 ( .A(n_24), .B(n_235), .Y(n_275) );
OAI221xp5_ASAP7_75t_L g193 ( .A1(n_25), .A2(n_50), .B1(n_57), .B2(n_194), .C(n_196), .Y(n_193) );
OR2x2_ASAP7_75t_L g219 ( .A(n_26), .B(n_66), .Y(n_219) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_26), .A2(n_66), .B(n_218), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_27), .B(n_235), .Y(n_270) );
INVx3_ASAP7_75t_L g90 ( .A(n_28), .Y(n_90) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_29), .B(n_237), .Y(n_287) );
INVx1_ASAP7_75t_L g139 ( .A(n_30), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_31), .B(n_235), .Y(n_311) );
INVx1_ASAP7_75t_L g536 ( .A(n_31), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_32), .A2(n_221), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_SL g95 ( .A(n_33), .Y(n_95) );
INVx1_ASAP7_75t_L g203 ( .A(n_34), .Y(n_203) );
AND2x2_ASAP7_75t_L g222 ( .A(n_34), .B(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g232 ( .A(n_34), .B(n_201), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_35), .B(n_226), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g300 ( .A(n_36), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_37), .B(n_235), .Y(n_257) );
INVx1_ASAP7_75t_L g187 ( .A(n_38), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_39), .A2(n_221), .B(n_274), .Y(n_273) );
AO22x2_ASAP7_75t_L g89 ( .A1(n_40), .A2(n_57), .B1(n_90), .B2(n_91), .Y(n_89) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_41), .B(n_235), .Y(n_246) );
INVx1_ASAP7_75t_L g225 ( .A(n_42), .Y(n_225) );
INVx1_ASAP7_75t_L g229 ( .A(n_42), .Y(n_229) );
INVx1_ASAP7_75t_L g96 ( .A(n_43), .Y(n_96) );
INVx1_ASAP7_75t_L g161 ( .A(n_44), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_45), .B(n_237), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_46), .A2(n_221), .B(n_244), .Y(n_243) );
AO21x1_ASAP7_75t_L g309 ( .A1(n_47), .A2(n_221), .B(n_310), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_47), .A2(n_80), .B1(n_81), .B2(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_47), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_48), .B(n_226), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_49), .B(n_226), .Y(n_277) );
INVxp33_ASAP7_75t_L g198 ( .A(n_50), .Y(n_198) );
AND2x2_ASAP7_75t_L g260 ( .A(n_51), .B(n_217), .Y(n_260) );
INVx1_ASAP7_75t_L g223 ( .A(n_52), .Y(n_223) );
INVx1_ASAP7_75t_L g231 ( .A(n_52), .Y(n_231) );
AND2x2_ASAP7_75t_L g279 ( .A(n_53), .B(n_249), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g172 ( .A1(n_54), .A2(n_56), .B1(n_173), .B2(n_176), .Y(n_172) );
AOI221x1_ASAP7_75t_L g125 ( .A1(n_55), .A2(n_59), .B1(n_126), .B2(n_129), .C(n_132), .Y(n_125) );
INVxp67_ASAP7_75t_L g197 ( .A(n_57), .Y(n_197) );
INVx1_ASAP7_75t_L g104 ( .A(n_58), .Y(n_104) );
AND2x2_ASAP7_75t_L g264 ( .A(n_60), .B(n_249), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_61), .B(n_226), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_62), .A2(n_80), .B1(n_81), .B2(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_62), .Y(n_529) );
AND2x2_ASAP7_75t_L g308 ( .A(n_63), .B(n_289), .Y(n_308) );
INVx1_ASAP7_75t_L g138 ( .A(n_64), .Y(n_138) );
INVx1_ASAP7_75t_L g115 ( .A(n_65), .Y(n_115) );
AND2x2_ASAP7_75t_L g252 ( .A(n_67), .B(n_249), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_68), .B(n_235), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_69), .B(n_237), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_70), .B(n_235), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_71), .A2(n_221), .B(n_295), .Y(n_294) );
OAI22xp5_ASAP7_75t_SL g181 ( .A1(n_72), .A2(n_182), .B1(n_183), .B2(n_189), .Y(n_181) );
INVx1_ASAP7_75t_L g189 ( .A(n_72), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_73), .B(n_237), .Y(n_269) );
INVx1_ASAP7_75t_L g145 ( .A(n_74), .Y(n_145) );
BUFx2_ASAP7_75t_SL g195 ( .A(n_75), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_76), .A2(n_221), .B(n_286), .Y(n_285) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_190), .B1(n_204), .B2(n_512), .C(n_519), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_181), .Y(n_78) );
INVx1_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
INVxp33_ASAP7_75t_SL g81 ( .A(n_82), .Y(n_81) );
NAND3xp33_ASAP7_75t_L g82 ( .A(n_83), .B(n_125), .C(n_143), .Y(n_82) );
NOR2xp33_ASAP7_75t_L g83 ( .A(n_84), .B(n_114), .Y(n_83) );
OAI22xp33_ASAP7_75t_L g84 ( .A1(n_85), .A2(n_104), .B1(n_105), .B2(n_106), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
BUFx2_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_97), .Y(n_87) );
AND2x2_ASAP7_75t_L g137 ( .A(n_88), .B(n_112), .Y(n_137) );
AND2x4_ASAP7_75t_L g175 ( .A(n_88), .B(n_124), .Y(n_175) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_92), .Y(n_88) );
INVx2_ASAP7_75t_L g111 ( .A(n_89), .Y(n_111) );
BUFx2_ASAP7_75t_L g142 ( .A(n_89), .Y(n_142) );
AND2x2_ASAP7_75t_L g151 ( .A(n_89), .B(n_93), .Y(n_151) );
INVx1_ASAP7_75t_L g91 ( .A(n_90), .Y(n_91) );
OAI22x1_ASAP7_75t_L g93 ( .A1(n_90), .A2(n_94), .B1(n_95), .B2(n_96), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_90), .Y(n_94) );
INVx2_ASAP7_75t_L g100 ( .A(n_90), .Y(n_100) );
INVx1_ASAP7_75t_L g103 ( .A(n_90), .Y(n_103) );
AND2x4_ASAP7_75t_L g110 ( .A(n_92), .B(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
AND2x2_ASAP7_75t_L g118 ( .A(n_93), .B(n_111), .Y(n_118) );
HB1xp67_ASAP7_75t_L g155 ( .A(n_93), .Y(n_155) );
AND2x4_ASAP7_75t_L g117 ( .A(n_97), .B(n_118), .Y(n_117) );
AND2x4_ASAP7_75t_L g128 ( .A(n_97), .B(n_110), .Y(n_128) );
AND2x2_ASAP7_75t_L g150 ( .A(n_97), .B(n_151), .Y(n_150) );
AND2x4_ASAP7_75t_L g97 ( .A(n_98), .B(n_101), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
INVx1_ASAP7_75t_L g113 ( .A(n_99), .Y(n_113) );
AND2x4_ASAP7_75t_L g124 ( .A(n_99), .B(n_101), .Y(n_124) );
AND2x2_ASAP7_75t_L g131 ( .A(n_99), .B(n_102), .Y(n_131) );
INVxp67_ASAP7_75t_L g179 ( .A(n_101), .Y(n_179) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_L g112 ( .A(n_102), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx8_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x4_ASAP7_75t_L g109 ( .A(n_110), .B(n_112), .Y(n_109) );
AND2x4_ASAP7_75t_L g123 ( .A(n_110), .B(n_124), .Y(n_123) );
AND2x4_ASAP7_75t_L g130 ( .A(n_110), .B(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g166 ( .A(n_112), .B(n_118), .Y(n_166) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_113), .Y(n_171) );
OAI22xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_116), .B1(n_119), .B2(n_120), .Y(n_114) );
INVx6_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AND2x2_ASAP7_75t_L g160 ( .A(n_118), .B(n_124), .Y(n_160) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx3_ASAP7_75t_SL g126 ( .A(n_127), .Y(n_126) );
INVx8_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx2_ASAP7_75t_SL g129 ( .A(n_130), .Y(n_129) );
AND2x4_ASAP7_75t_L g141 ( .A(n_131), .B(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_L g154 ( .A(n_131), .B(n_155), .Y(n_154) );
OAI22xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_138), .B1(n_139), .B2(n_140), .Y(n_132) );
HB1xp67_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx5_ASAP7_75t_SL g140 ( .A(n_141), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_144), .B(n_162), .Y(n_143) );
OAI222xp33_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_146), .B1(n_152), .B2(n_156), .C1(n_157), .C2(n_161), .Y(n_144) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx3_ASAP7_75t_SL g148 ( .A(n_149), .Y(n_148) );
INVx6_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x4_ASAP7_75t_L g169 ( .A(n_151), .B(n_170), .Y(n_169) );
AND2x4_ASAP7_75t_L g178 ( .A(n_151), .B(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx12f_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_163), .B(n_172), .Y(n_162) );
BUFx6f_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_SL g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
BUFx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx6_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_183), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_186), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_191), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_192), .Y(n_191) );
AND3x1_ASAP7_75t_SL g192 ( .A(n_193), .B(n_199), .C(n_202), .Y(n_192) );
INVxp67_ASAP7_75t_L g527 ( .A(n_193), .Y(n_527) );
CKINVDCx8_ASAP7_75t_R g194 ( .A(n_195), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
CKINVDCx16_ASAP7_75t_R g525 ( .A(n_199), .Y(n_525) );
AOI21xp33_ASAP7_75t_L g532 ( .A1(n_199), .A2(n_533), .B(n_534), .Y(n_532) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g516 ( .A(n_200), .B(n_517), .Y(n_516) );
OR2x2_ASAP7_75t_SL g530 ( .A(n_200), .B(n_202), .Y(n_530) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g224 ( .A(n_201), .B(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_202), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x4_ASAP7_75t_L g207 ( .A(n_208), .B(n_424), .Y(n_207) );
AND4x1_ASAP7_75t_L g208 ( .A(n_209), .B(n_336), .C(n_363), .D(n_398), .Y(n_208) );
AOI221xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_261), .B1(n_301), .B2(n_316), .C(n_320), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_212), .B(n_240), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_212), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
OR2x2_ASAP7_75t_L g377 ( .A(n_213), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g432 ( .A(n_213), .B(n_387), .Y(n_432) );
BUFx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g335 ( .A(n_214), .B(n_253), .Y(n_335) );
AND2x4_ASAP7_75t_L g371 ( .A(n_214), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g385 ( .A(n_214), .B(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g302 ( .A(n_215), .Y(n_302) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_215), .Y(n_474) );
OA21x2_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_220), .B(n_239), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_216), .A2(n_266), .B(n_267), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_216), .Y(n_278) );
OA21x2_ASAP7_75t_L g348 ( .A1(n_216), .A2(n_220), .B(n_239), .Y(n_348) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_SL g217 ( .A(n_218), .B(n_219), .Y(n_217) );
AND2x4_ASAP7_75t_L g289 ( .A(n_218), .B(n_219), .Y(n_289) );
AND2x6_ASAP7_75t_L g221 ( .A(n_222), .B(n_224), .Y(n_221) );
BUFx3_ASAP7_75t_L g518 ( .A(n_222), .Y(n_518) );
AND2x6_ASAP7_75t_L g235 ( .A(n_223), .B(n_228), .Y(n_235) );
AND2x4_ASAP7_75t_L g237 ( .A(n_225), .B(n_230), .Y(n_237) );
INVx2_ASAP7_75t_L g517 ( .A(n_225), .Y(n_517) );
AND2x4_ASAP7_75t_L g226 ( .A(n_227), .B(n_232), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_228), .B(n_230), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx5_ASAP7_75t_L g238 ( .A(n_232), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_236), .B(n_238), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_238), .A2(n_245), .B(n_246), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_238), .A2(n_257), .B(n_258), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_238), .A2(n_269), .B(n_270), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_238), .A2(n_275), .B(n_276), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_238), .A2(n_287), .B(n_288), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_238), .A2(n_296), .B(n_297), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_238), .A2(n_311), .B(n_312), .Y(n_310) );
A2O1A1Ixp33_ASAP7_75t_SL g329 ( .A1(n_240), .A2(n_302), .B(n_330), .C(n_334), .Y(n_329) );
AND2x2_ASAP7_75t_L g350 ( .A(n_240), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_240), .B(n_302), .Y(n_490) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_253), .Y(n_240) );
INVx2_ASAP7_75t_L g370 ( .A(n_241), .Y(n_370) );
BUFx3_ASAP7_75t_L g386 ( .A(n_241), .Y(n_386) );
INVxp67_ASAP7_75t_L g390 ( .A(n_241), .Y(n_390) );
AO21x2_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_248), .B(n_252), .Y(n_241) );
AO21x2_ASAP7_75t_L g340 ( .A1(n_242), .A2(n_248), .B(n_252), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_247), .Y(n_242) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_248), .A2(n_254), .B(n_260), .Y(n_253) );
AO21x2_ASAP7_75t_L g315 ( .A1(n_248), .A2(n_254), .B(n_260), .Y(n_315) );
INVx3_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx4_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
BUFx4f_ASAP7_75t_L g282 ( .A(n_251), .Y(n_282) );
INVx2_ASAP7_75t_L g369 ( .A(n_253), .Y(n_369) );
AND2x2_ASAP7_75t_L g375 ( .A(n_253), .B(n_348), .Y(n_375) );
AND2x2_ASAP7_75t_L g401 ( .A(n_253), .B(n_370), .Y(n_401) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_255), .B(n_259), .Y(n_254) );
AOI211xp5_ASAP7_75t_L g398 ( .A1(n_261), .A2(n_399), .B(n_402), .C(n_412), .Y(n_398) );
AND2x2_ASAP7_75t_SL g261 ( .A(n_262), .B(n_280), .Y(n_261) );
OAI321xp33_ASAP7_75t_L g373 ( .A1(n_262), .A2(n_321), .A3(n_374), .B1(n_376), .B2(n_377), .C(n_379), .Y(n_373) );
AND2x2_ASAP7_75t_L g494 ( .A(n_262), .B(n_469), .Y(n_494) );
INVx1_ASAP7_75t_L g497 ( .A(n_262), .Y(n_497) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_271), .Y(n_262) );
INVx5_ASAP7_75t_L g319 ( .A(n_263), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_263), .B(n_333), .Y(n_332) );
NOR2x1_ASAP7_75t_SL g364 ( .A(n_263), .B(n_365), .Y(n_364) );
BUFx2_ASAP7_75t_L g409 ( .A(n_263), .Y(n_409) );
AND2x2_ASAP7_75t_L g511 ( .A(n_263), .B(n_281), .Y(n_511) );
OR2x6_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
AND2x2_ASAP7_75t_L g318 ( .A(n_271), .B(n_319), .Y(n_318) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_271), .Y(n_328) );
INVx4_ASAP7_75t_L g333 ( .A(n_271), .Y(n_333) );
AO21x2_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_278), .B(n_279), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_277), .Y(n_272) );
INVx1_ASAP7_75t_L g376 ( .A(n_280), .Y(n_376) );
A2O1A1Ixp33_ASAP7_75t_R g479 ( .A1(n_280), .A2(n_318), .B(n_350), .C(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g499 ( .A(n_280), .B(n_324), .Y(n_499) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_290), .Y(n_280) );
INVx1_ASAP7_75t_L g317 ( .A(n_281), .Y(n_317) );
INVx2_ASAP7_75t_L g323 ( .A(n_281), .Y(n_323) );
OR2x2_ASAP7_75t_L g342 ( .A(n_281), .B(n_333), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_281), .B(n_365), .Y(n_411) );
BUFx3_ASAP7_75t_L g418 ( .A(n_281), .Y(n_418) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_285), .B(n_289), .Y(n_283) );
INVx1_ASAP7_75t_SL g292 ( .A(n_289), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_289), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g381 ( .A(n_290), .Y(n_381) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_290), .Y(n_394) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g327 ( .A(n_291), .Y(n_327) );
INVx1_ASAP7_75t_L g436 ( .A(n_291), .Y(n_436) );
AO21x2_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_293), .B(n_299), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_292), .B(n_300), .Y(n_299) );
AO21x2_ASAP7_75t_L g365 ( .A1(n_292), .A2(n_293), .B(n_299), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_298), .Y(n_293) );
AND2x2_ASAP7_75t_L g337 ( .A(n_301), .B(n_338), .Y(n_337) );
OAI31xp33_ASAP7_75t_L g488 ( .A1(n_301), .A2(n_489), .A3(n_491), .B(n_494), .Y(n_488) );
INVx1_ASAP7_75t_SL g506 ( .A(n_301), .Y(n_506) );
AND2x4_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
AOI21xp33_ASAP7_75t_L g320 ( .A1(n_302), .A2(n_321), .B(n_329), .Y(n_320) );
NAND2x1_ASAP7_75t_L g400 ( .A(n_302), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g429 ( .A(n_302), .Y(n_429) );
INVx2_ASAP7_75t_L g378 ( .A(n_303), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_303), .B(n_361), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_303), .B(n_360), .Y(n_470) );
NOR2xp33_ASAP7_75t_SL g478 ( .A(n_303), .B(n_429), .Y(n_478) );
AND2x4_ASAP7_75t_L g303 ( .A(n_304), .B(n_315), .Y(n_303) );
AND2x2_ASAP7_75t_SL g347 ( .A(n_304), .B(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g358 ( .A(n_304), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g387 ( .A(n_304), .B(n_369), .Y(n_387) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx2_ASAP7_75t_L g351 ( .A(n_305), .Y(n_351) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g372 ( .A(n_306), .Y(n_372) );
OAI21x1_ASAP7_75t_SL g306 ( .A1(n_307), .A2(n_309), .B(n_313), .Y(n_306) );
INVx1_ASAP7_75t_L g314 ( .A(n_308), .Y(n_314) );
INVx2_ASAP7_75t_L g359 ( .A(n_315), .Y(n_359) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_315), .Y(n_419) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_L g355 ( .A(n_317), .Y(n_355) );
AND2x2_ASAP7_75t_L g434 ( .A(n_317), .B(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g345 ( .A(n_318), .B(n_339), .Y(n_345) );
INVx2_ASAP7_75t_SL g393 ( .A(n_318), .Y(n_393) );
INVx4_ASAP7_75t_L g324 ( .A(n_319), .Y(n_324) );
AND2x2_ASAP7_75t_L g422 ( .A(n_319), .B(n_365), .Y(n_422) );
AND2x2_ASAP7_75t_SL g440 ( .A(n_319), .B(n_435), .Y(n_440) );
NAND2x1p5_ASAP7_75t_L g457 ( .A(n_319), .B(n_333), .Y(n_457) );
INVx1_ASAP7_75t_L g463 ( .A(n_321), .Y(n_463) );
OR2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_325), .Y(n_321) );
INVx1_ASAP7_75t_L g382 ( .A(n_322), .Y(n_382) );
OR2x2_ASAP7_75t_L g395 ( .A(n_322), .B(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
OR2x2_ASAP7_75t_L g447 ( .A(n_323), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g477 ( .A(n_323), .B(n_365), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_324), .B(n_327), .Y(n_353) );
AND2x2_ASAP7_75t_L g445 ( .A(n_324), .B(n_435), .Y(n_445) );
AND2x4_ASAP7_75t_L g507 ( .A(n_324), .B(n_386), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
INVx2_ASAP7_75t_L g331 ( .A(n_326), .Y(n_331) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NOR2xp67_ASAP7_75t_SL g330 ( .A(n_331), .B(n_332), .Y(n_330) );
OAI322xp33_ASAP7_75t_SL g343 ( .A1(n_331), .A2(n_344), .A3(n_346), .B1(n_349), .B2(n_352), .C1(n_354), .C2(n_356), .Y(n_343) );
INVx1_ASAP7_75t_L g501 ( .A(n_331), .Y(n_501) );
OR2x2_ASAP7_75t_L g354 ( .A(n_332), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g380 ( .A(n_333), .B(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_333), .B(n_381), .Y(n_396) );
INVx2_ASAP7_75t_L g423 ( .A(n_333), .Y(n_423) );
AND2x4_ASAP7_75t_L g435 ( .A(n_333), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_SL g438 ( .A(n_335), .B(n_351), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_341), .B(n_343), .Y(n_336) );
AND2x2_ASAP7_75t_L g404 ( .A(n_338), .B(n_371), .Y(n_404) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_339), .B(n_493), .Y(n_492) );
BUFx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g362 ( .A(n_340), .Y(n_362) );
AND2x4_ASAP7_75t_SL g444 ( .A(n_340), .B(n_359), .Y(n_444) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g352 ( .A(n_342), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_345), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g480 ( .A(n_347), .B(n_444), .Y(n_480) );
NOR4xp25_ASAP7_75t_L g484 ( .A(n_347), .B(n_361), .C(n_401), .D(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g361 ( .A(n_348), .B(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g397 ( .A(n_348), .B(n_372), .Y(n_397) );
AND2x4_ASAP7_75t_L g461 ( .A(n_348), .B(n_372), .Y(n_461) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_351), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_358), .B(n_360), .Y(n_357) );
OR2x2_ASAP7_75t_L g450 ( .A(n_358), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g504 ( .A(n_358), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_359), .B(n_371), .Y(n_405) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
AOI211xp5_ASAP7_75t_SL g363 ( .A1(n_364), .A2(n_366), .B(n_373), .C(n_388), .Y(n_363) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_371), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_369), .B(n_372), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_370), .B(n_375), .Y(n_374) );
BUFx2_ASAP7_75t_L g452 ( .A(n_370), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_371), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g467 ( .A(n_371), .Y(n_467) );
OAI21xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_382), .B(n_383), .Y(n_379) );
AND2x4_ASAP7_75t_L g416 ( .A(n_380), .B(n_417), .Y(n_416) );
AND2x4_ASAP7_75t_L g510 ( .A(n_380), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
INVx1_ASAP7_75t_SL g414 ( .A(n_386), .Y(n_414) );
AND2x2_ASAP7_75t_L g473 ( .A(n_387), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g487 ( .A(n_387), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_SL g388 ( .A1(n_389), .A2(n_391), .B(n_395), .C(n_397), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_389), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g465 ( .A(n_390), .B(n_466), .Y(n_465) );
OR2x2_ASAP7_75t_L g486 ( .A(n_390), .B(n_487), .Y(n_486) );
INVxp67_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
OR2x2_ASAP7_75t_L g475 ( .A(n_393), .B(n_417), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_396), .A2(n_403), .B1(n_405), .B2(n_406), .Y(n_402) );
INVx1_ASAP7_75t_SL g493 ( .A(n_397), .Y(n_493) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_410), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_408), .B(n_417), .Y(n_459) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVxp67_ASAP7_75t_SL g469 ( .A(n_411), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_415), .B1(n_419), .B2(n_420), .Y(n_412) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AOI21xp5_ASAP7_75t_SL g426 ( .A1(n_417), .A2(n_427), .B(n_430), .Y(n_426) );
AND2x2_ASAP7_75t_L g455 ( .A(n_417), .B(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AND3x2_ASAP7_75t_L g421 ( .A(n_418), .B(n_422), .C(n_423), .Y(n_421) );
AND2x2_ASAP7_75t_L g483 ( .A(n_418), .B(n_440), .Y(n_483) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g468 ( .A(n_423), .B(n_469), .Y(n_468) );
NOR2xp67_ASAP7_75t_L g424 ( .A(n_425), .B(n_481), .Y(n_424) );
NAND4xp25_ASAP7_75t_L g425 ( .A(n_426), .B(n_441), .C(n_462), .D(n_479), .Y(n_425) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_433), .B1(n_437), .B2(n_439), .Y(n_430) );
INVx1_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_433), .A2(n_447), .B1(n_467), .B2(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g448 ( .A(n_435), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_437), .A2(n_460), .B(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx3_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
AOI221xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_445), .B1(n_446), .B2(n_449), .C(n_453), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_458), .B1(n_459), .B2(n_460), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_456), .B(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_456), .B(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AOI221xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_464), .B1(n_468), .B2(n_470), .C(n_471), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_465), .B(n_467), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_475), .B1(n_476), .B2(n_478), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OAI211xp5_ASAP7_75t_SL g496 ( .A1(n_477), .A2(n_497), .B(n_498), .C(n_500), .Y(n_496) );
OAI211xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_484), .B(n_488), .C(n_495), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
AOI221xp5_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_502), .B1(n_505), .B2(n_507), .C(n_508), .Y(n_495) );
INVx1_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_SL g509 ( .A(n_510), .Y(n_509) );
CKINVDCx16_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x4_ASAP7_75t_L g515 ( .A(n_516), .B(n_518), .Y(n_515) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_517), .Y(n_533) );
INVx1_ASAP7_75t_L g535 ( .A(n_518), .Y(n_535) );
OAI222xp33_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_522), .B1(n_528), .B2(n_530), .C1(n_531), .C2(n_536), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_523), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_524), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
INVx1_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
INVxp67_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
endmodule