module real_jpeg_29417_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_340, n_11, n_14, n_7, n_3, n_5, n_4, n_339, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_340;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_339;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_0),
.A2(n_30),
.B1(n_31),
.B2(n_218),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_0),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_0),
.A2(n_35),
.B1(n_37),
.B2(n_218),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_0),
.A2(n_101),
.B1(n_102),
.B2(n_218),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_0),
.A2(n_160),
.B1(n_166),
.B2(n_218),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_1),
.A2(n_30),
.B1(n_31),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_1),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_1),
.A2(n_35),
.B1(n_37),
.B2(n_156),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_1),
.A2(n_101),
.B1(n_102),
.B2(n_156),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_1),
.A2(n_156),
.B1(n_160),
.B2(n_166),
.Y(n_300)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_2),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_3),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_3),
.A2(n_35),
.B1(n_37),
.B2(n_139),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_3),
.A2(n_101),
.B1(n_102),
.B2(n_139),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_3),
.A2(n_139),
.B1(n_160),
.B2(n_166),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_4),
.B(n_37),
.Y(n_36)
);

A2O1A1O1Ixp25_ASAP7_75t_L g39 ( 
.A1(n_4),
.A2(n_36),
.B(n_37),
.C(n_40),
.D(n_44),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_4),
.B(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_4),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_L g88 ( 
.A1(n_4),
.A2(n_61),
.B(n_65),
.Y(n_88)
);

A2O1A1O1Ixp25_ASAP7_75t_L g100 ( 
.A1(n_4),
.A2(n_101),
.B(n_103),
.C(n_104),
.D(n_108),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_4),
.B(n_101),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_4),
.A2(n_102),
.B(n_136),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_4),
.A2(n_83),
.B1(n_160),
.B2(n_166),
.Y(n_167)
);

BUFx12_ASAP7_75t_L g136 ( 
.A(n_5),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_6),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_6),
.A2(n_35),
.B1(n_37),
.B2(n_200),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_6),
.A2(n_101),
.B1(n_102),
.B2(n_200),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_6),
.A2(n_160),
.B1(n_166),
.B2(n_200),
.Y(n_322)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_8),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_9),
.A2(n_35),
.B1(n_37),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_46),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_9),
.A2(n_46),
.B1(n_101),
.B2(n_102),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_9),
.A2(n_46),
.B1(n_160),
.B2(n_166),
.Y(n_170)
);

BUFx24_ASAP7_75t_L g102 ( 
.A(n_10),
.Y(n_102)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_11),
.B(n_31),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_11),
.B(n_37),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_12),
.A2(n_35),
.B1(n_37),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_12),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_12),
.A2(n_30),
.B1(n_31),
.B2(n_57),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_12),
.A2(n_57),
.B1(n_101),
.B2(n_102),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_12),
.A2(n_57),
.B1(n_160),
.B2(n_166),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_13),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_13),
.A2(n_35),
.B1(n_37),
.B2(n_118),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_13),
.A2(n_101),
.B1(n_102),
.B2(n_118),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_13),
.A2(n_118),
.B1(n_160),
.B2(n_166),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_64),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_14),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_14),
.A2(n_35),
.B1(n_37),
.B2(n_64),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_14),
.A2(n_64),
.B1(n_101),
.B2(n_102),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_14),
.A2(n_64),
.B1(n_160),
.B2(n_166),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_15),
.A2(n_35),
.B1(n_37),
.B2(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_15),
.Y(n_107)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_16),
.Y(n_33)
);

AO21x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_332),
.B(n_335),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_327),
.B(n_331),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_314),
.B(n_326),
.Y(n_19)
);

OAI321xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_278),
.A3(n_307),
.B1(n_312),
.B2(n_313),
.C(n_339),
.Y(n_20)
);

AOI321xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_228),
.A3(n_267),
.B1(n_272),
.B2(n_277),
.C(n_340),
.Y(n_21)
);

NOR3xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_180),
.C(n_224),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_147),
.B(n_179),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_123),
.B(n_146),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_96),
.B(n_122),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_70),
.B(n_95),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_48),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_28),
.B(n_48),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_39),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_29),
.B(n_39),
.Y(n_79)
);

AOI32xp33_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_34),
.A3(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_30),
.B(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_31),
.B(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_35),
.Y(n_37)
);

NAND2xp33_ASAP7_75t_SL g121 ( 
.A(n_35),
.B(n_106),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_41),
.B(n_42),
.C(n_43),
.Y(n_40)
);

AOI32xp33_ASAP7_75t_L g119 ( 
.A1(n_37),
.A2(n_102),
.A3(n_103),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_40),
.B(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_40),
.A2(n_43),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_40),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_40),
.A2(n_43),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_40),
.A2(n_43),
.B1(n_244),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_44),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_47),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_45),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_56),
.B(n_58),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_47),
.B(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_47),
.A2(n_58),
.B(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_47),
.A2(n_143),
.B1(n_178),
.B2(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_47),
.A2(n_143),
.B1(n_202),
.B2(n_220),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_47),
.A2(n_143),
.B(n_253),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_60),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_55),
.C(n_60),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_52),
.B(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_52),
.A2(n_104),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_52),
.A2(n_104),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_52),
.A2(n_104),
.B1(n_256),
.B2(n_285),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_52),
.A2(n_104),
.B(n_319),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_53),
.A2(n_101),
.B1(n_102),
.B2(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_56),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_63),
.B(n_65),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_67),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_61),
.A2(n_78),
.B1(n_117),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_61),
.A2(n_69),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_61),
.A2(n_78),
.B1(n_199),
.B2(n_217),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_61),
.A2(n_78),
.B(n_217),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_68),
.A2(n_86),
.B(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_68),
.A2(n_75),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_80),
.B(n_94),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_79),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_72),
.B(n_79),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_74),
.A2(n_78),
.B(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_87),
.B(n_93),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_84),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_82),
.B(n_84),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_83),
.B(n_133),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_83),
.A2(n_135),
.B(n_159),
.C(n_160),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_97),
.B(n_98),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_114),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_111),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_111),
.C(n_114),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_101),
.A2(n_102),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_104),
.B(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_104),
.Y(n_188)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_108),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_128),
.B(n_129),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_110),
.A2(n_129),
.B(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_110),
.A2(n_188),
.B1(n_214),
.B2(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_110),
.A2(n_188),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_113),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_119),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_119),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_124),
.B(n_125),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_140),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_141),
.C(n_142),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_131),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_132),
.C(n_137),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_128),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_137),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_133),
.A2(n_192),
.B(n_194),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_133),
.A2(n_194),
.B(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_133),
.A2(n_235),
.B1(n_263),
.B2(n_290),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_133),
.A2(n_235),
.B1(n_290),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_134),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_134),
.B(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_134),
.A2(n_164),
.B1(n_193),
.B2(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_134),
.A2(n_164),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_134),
.A2(n_164),
.B1(n_322),
.B2(n_329),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_134),
.A2(n_164),
.B(n_329),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_136),
.B1(n_160),
.B2(n_166),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_138),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_144),
.B(n_145),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_148),
.B(n_149),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_162),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_151),
.B(n_152),
.C(n_162),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_157),
.B1(n_158),
.B2(n_161),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_155),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_161),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_160),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_171),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_173),
.C(n_176),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_167),
.B(n_168),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_164),
.B(n_170),
.Y(n_194)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_164),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_169),
.A2(n_235),
.B(n_236),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_176),
.B2(n_177),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_175),
.Y(n_189)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_181),
.A2(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_204),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_182),
.B(n_204),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_196),
.C(n_203),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_183),
.B(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_186),
.C(n_195),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_191),
.B2(n_195),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B(n_190),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_191),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_203),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_201),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_201),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_204)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_215),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_206),
.B(n_215),
.C(n_223),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_207),
.B(n_210),
.C(n_212),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_212),
.B2(n_213),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_211),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_219),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_220),
.Y(n_243)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_221),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_225),
.B(n_226),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_248),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_229),
.B(n_248),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_240),
.C(n_247),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_230),
.B(n_240),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_239),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_231),
.Y(n_239)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_237),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_237),
.C(n_239),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_238),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_245),
.B2(n_246),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_246),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_245),
.A2(n_246),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

AOI21xp33_ASAP7_75t_L g294 ( 
.A1(n_246),
.A2(n_261),
.B(n_264),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_266),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_258),
.B1(n_259),
.B2(n_265),
.Y(n_249)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

OAI21xp33_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_254),
.B(n_257),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_254),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_257),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_257),
.A2(n_280),
.B1(n_281),
.B2(n_292),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_258),
.B(n_265),
.C(n_266),
.Y(n_308)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_264),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_268),
.A2(n_273),
.B(n_276),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_269),
.B(n_270),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_295),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_279),
.B(n_295),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_292),
.C(n_293),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_289),
.B2(n_291),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_284),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_288),
.C(n_289),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_285),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_286),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_286),
.A2(n_288),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_288),
.B(n_299),
.C(n_303),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_289),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_289),
.A2(n_291),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_298),
.C(n_306),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_293),
.A2(n_294),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_306),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_300),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_303),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_305),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_308),
.B(n_309),
.Y(n_312)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_316),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_325),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_320),
.B1(n_323),
.B2(n_324),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_318),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_320),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_324),
.C(n_325),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_330),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_328),
.B(n_330),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_333),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_328),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_337),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_336),
.Y(n_335)
);


endmodule