module fake_jpeg_17480_n_45 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_45);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_45;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_0),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_30),
.B(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_29),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_19),
.B1(n_12),
.B2(n_3),
.Y(n_28)
);

AO21x2_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_2),
.B(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_35),
.B1(n_8),
.B2(n_9),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_5),
.B(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_33),
.Y(n_36)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_32),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_39),
.B(n_38),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_40),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_42),
.A2(n_36),
.B(n_13),
.Y(n_43)
);

AO21x1_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_11),
.B(n_14),
.Y(n_44)
);

OAI21x1_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_15),
.B(n_17),
.Y(n_45)
);


endmodule