module fake_netlist_5_101_n_1777 (n_137, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1777);

input n_137;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1777;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_604;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1155;
wire n_1418;
wire n_1689;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_130),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_124),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_136),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_138),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_137),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_146),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_64),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_159),
.Y(n_174)
);

BUFx10_ASAP7_75t_L g175 ( 
.A(n_104),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_23),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_42),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_20),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_156),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_1),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_15),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_86),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_73),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_118),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_102),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_48),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_74),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_78),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_105),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_0),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_81),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_38),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_75),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_114),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_153),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_113),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_63),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_127),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_47),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_76),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_143),
.Y(n_201)
);

INVxp67_ASAP7_75t_SL g202 ( 
.A(n_147),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_103),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_24),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_24),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_5),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_77),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_23),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_25),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_101),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_45),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_97),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_90),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_164),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_5),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_72),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_69),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_25),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_4),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_84),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_149),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_120),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_65),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_51),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_0),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_13),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_35),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_6),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_155),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_112),
.Y(n_230)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_133),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_88),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_35),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_49),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_39),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_121),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_135),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_128),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_12),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_117),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_36),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_142),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_57),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_49),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_34),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_61),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_56),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_96),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_6),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_123),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_157),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_33),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_134),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_8),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_39),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_13),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_19),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_21),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_126),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_87),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_83),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_55),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_48),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_7),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_71),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_144),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_107),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_7),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_34),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_158),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_115),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_9),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_47),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_10),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_11),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_141),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_1),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_99),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_151),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_44),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_59),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_10),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_28),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_14),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_89),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_110),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_145),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_82),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_152),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_66),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_106),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_36),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_132),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_27),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_93),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_139),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_53),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_148),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_154),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_56),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_44),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_162),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_21),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_62),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_38),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_161),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_62),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_14),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_37),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_2),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_33),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_32),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_28),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_108),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_27),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_91),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_15),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_57),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_8),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_51),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_61),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_116),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_58),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_31),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_29),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_160),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_46),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_297),
.Y(n_328)
);

INVxp33_ASAP7_75t_L g329 ( 
.A(n_176),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_231),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_165),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_236),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_167),
.Y(n_333)
);

INVxp33_ASAP7_75t_SL g334 ( 
.A(n_173),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_168),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_184),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_200),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_287),
.B(n_2),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_176),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_248),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_297),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_177),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_169),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_297),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_170),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_231),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_177),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_169),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_261),
.B(n_3),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_180),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_180),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_181),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_297),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_179),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_182),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_236),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_183),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_277),
.Y(n_358)
);

INVxp33_ASAP7_75t_SL g359 ( 
.A(n_178),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_185),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_297),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_297),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_187),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_303),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_188),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_189),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_181),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_172),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_191),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_193),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_194),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_261),
.B(n_3),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_303),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_195),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_303),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_231),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_186),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_303),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_166),
.B(n_4),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_303),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_186),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_203),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_303),
.B(n_9),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_213),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_325),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_214),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_217),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_325),
.B(n_11),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_325),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_220),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_222),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_325),
.B(n_12),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_230),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_231),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_325),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_325),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_237),
.Y(n_397)
);

NOR2xp67_ASAP7_75t_L g398 ( 
.A(n_279),
.B(n_16),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_233),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_233),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_238),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_282),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_204),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_282),
.B(n_294),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_240),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_328),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_328),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_404),
.B(n_172),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_368),
.B(n_242),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_341),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_398),
.B(n_172),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_330),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_341),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_344),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_330),
.Y(n_415)
);

INVx5_ASAP7_75t_L g416 ( 
.A(n_330),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_344),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_353),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_353),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_343),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_346),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_361),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_368),
.B(n_250),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_346),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_361),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_362),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_362),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_332),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_364),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_364),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_373),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_373),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_375),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_375),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_378),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_378),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_380),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_380),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_385),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_385),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_404),
.B(n_295),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_389),
.Y(n_442)
);

NOR2x1_ASAP7_75t_L g443 ( 
.A(n_398),
.B(n_279),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_346),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_389),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_376),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_376),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_376),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_395),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_368),
.Y(n_450)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_394),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_395),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_396),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_396),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_394),
.Y(n_455)
);

NAND2xp33_ASAP7_75t_SL g456 ( 
.A(n_329),
.B(n_190),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_404),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_394),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_399),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_383),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_399),
.Y(n_461)
);

INVx6_ASAP7_75t_L g462 ( 
.A(n_332),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_400),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_400),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_349),
.B(n_251),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_402),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_402),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_383),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_336),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_372),
.B(n_260),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_338),
.B(n_334),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_359),
.B(n_332),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_337),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_356),
.B(n_174),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_342),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_356),
.B(n_265),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_356),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_342),
.B(n_266),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_352),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_450),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_410),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_471),
.A2(n_300),
.B1(n_226),
.B2(n_379),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_451),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_471),
.B(n_331),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_469),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_451),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_410),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_451),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_450),
.Y(n_489)
);

NAND3xp33_ASAP7_75t_L g490 ( 
.A(n_460),
.B(n_392),
.C(n_388),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_451),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_473),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_456),
.A2(n_292),
.B1(n_348),
.B2(n_197),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_475),
.B(n_333),
.Y(n_494)
);

INVx4_ASAP7_75t_L g495 ( 
.A(n_460),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_474),
.B(n_335),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_450),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_412),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_474),
.B(n_345),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_475),
.B(n_354),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_477),
.B(n_295),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_460),
.B(n_355),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_451),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_477),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_410),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g506 ( 
.A(n_456),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_477),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_457),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_413),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_462),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_462),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_412),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_457),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_412),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_412),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_413),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_413),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_414),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_412),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_460),
.Y(n_520)
);

AND3x2_ASAP7_75t_L g521 ( 
.A(n_428),
.B(n_392),
.C(n_388),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_414),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_406),
.Y(n_523)
);

AND2x2_ASAP7_75t_SL g524 ( 
.A(n_460),
.B(n_279),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_460),
.B(n_365),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_479),
.B(n_366),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_472),
.B(n_371),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_472),
.B(n_384),
.Y(n_528)
);

BUFx8_ASAP7_75t_SL g529 ( 
.A(n_420),
.Y(n_529)
);

INVx5_ASAP7_75t_L g530 ( 
.A(n_412),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_478),
.B(n_386),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_406),
.Y(n_532)
);

NAND3xp33_ASAP7_75t_L g533 ( 
.A(n_460),
.B(n_352),
.C(n_279),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_407),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_462),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_407),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_417),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_417),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_478),
.B(n_387),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_414),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_479),
.B(n_390),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_428),
.B(n_391),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_418),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_408),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_412),
.Y(n_545)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_468),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_408),
.B(n_351),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_418),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_462),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_419),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_462),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_420),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_465),
.B(n_393),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_419),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_415),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_425),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_SL g557 ( 
.A(n_465),
.B(n_357),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_425),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_L g559 ( 
.A(n_468),
.B(n_397),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_422),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_470),
.B(n_405),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_470),
.A2(n_370),
.B1(n_401),
.B2(n_382),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_427),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_468),
.B(n_295),
.Y(n_564)
);

OR2x2_ASAP7_75t_L g565 ( 
.A(n_476),
.B(n_358),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_422),
.Y(n_566)
);

AO21x2_ASAP7_75t_L g567 ( 
.A1(n_409),
.A2(n_171),
.B(n_166),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_427),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_468),
.B(n_299),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_408),
.B(n_441),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_431),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_476),
.B(n_358),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_422),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_468),
.A2(n_360),
.B1(n_374),
.B2(n_369),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_426),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_426),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_409),
.B(n_363),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_431),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_415),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_426),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_441),
.B(n_171),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_433),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_423),
.B(n_340),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_468),
.A2(n_294),
.B1(n_257),
.B2(n_206),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_468),
.B(n_267),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_429),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_423),
.B(n_271),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_441),
.B(n_403),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_411),
.A2(n_257),
.B1(n_206),
.B2(n_268),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_415),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_429),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_411),
.B(n_175),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_411),
.B(n_278),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_415),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_415),
.Y(n_595)
);

XOR2x2_ASAP7_75t_L g596 ( 
.A(n_443),
.B(n_339),
.Y(n_596)
);

INVx5_ASAP7_75t_L g597 ( 
.A(n_415),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_415),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_421),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_411),
.B(n_462),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_429),
.Y(n_601)
);

INVx5_ASAP7_75t_L g602 ( 
.A(n_421),
.Y(n_602)
);

INVxp67_ASAP7_75t_SL g603 ( 
.A(n_421),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_433),
.Y(n_604)
);

AND2x6_ASAP7_75t_L g605 ( 
.A(n_411),
.B(n_196),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_443),
.B(n_175),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_430),
.Y(n_607)
);

AND3x2_ASAP7_75t_L g608 ( 
.A(n_459),
.B(n_276),
.C(n_196),
.Y(n_608)
);

NAND2xp33_ASAP7_75t_R g609 ( 
.A(n_459),
.B(n_192),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_467),
.B(n_175),
.Y(n_610)
);

BUFx4f_ASAP7_75t_L g611 ( 
.A(n_421),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_434),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_434),
.Y(n_613)
);

INVx4_ASAP7_75t_L g614 ( 
.A(n_421),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_435),
.Y(n_615)
);

AND2x2_ASAP7_75t_SL g616 ( 
.A(n_421),
.B(n_276),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_461),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_461),
.B(n_351),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_435),
.B(n_285),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_430),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_463),
.A2(n_280),
.B1(n_244),
.B2(n_243),
.Y(n_621)
);

BUFx10_ASAP7_75t_L g622 ( 
.A(n_463),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_421),
.Y(n_623)
);

INVx8_ASAP7_75t_L g624 ( 
.A(n_424),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_464),
.B(n_175),
.Y(n_625)
);

NAND3xp33_ASAP7_75t_L g626 ( 
.A(n_464),
.B(n_201),
.C(n_198),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_437),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_424),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_467),
.B(n_377),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_430),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_553),
.B(n_424),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_521),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_544),
.Y(n_633)
);

NAND3xp33_ASAP7_75t_L g634 ( 
.A(n_494),
.B(n_347),
.C(n_339),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_524),
.B(n_495),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_569),
.B(n_424),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_570),
.B(n_424),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_508),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_570),
.B(n_424),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_570),
.B(n_424),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_524),
.B(n_444),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_570),
.B(n_508),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_513),
.B(n_444),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_500),
.B(n_199),
.Y(n_644)
);

OAI22xp5_ASAP7_75t_SL g645 ( 
.A1(n_482),
.A2(n_269),
.B1(n_273),
.B2(n_283),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_489),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_513),
.B(n_444),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_489),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_524),
.B(n_444),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_617),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_495),
.B(n_444),
.Y(n_651)
);

NOR2xp67_ASAP7_75t_L g652 ( 
.A(n_574),
.B(n_377),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_617),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_481),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_526),
.B(n_205),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_547),
.B(n_347),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_523),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_523),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_547),
.B(n_350),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_497),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_588),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_495),
.B(n_444),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_502),
.B(n_525),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_541),
.B(n_444),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_483),
.B(n_446),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_484),
.B(n_209),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_483),
.B(n_446),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_532),
.Y(n_668)
);

AO221x1_ASAP7_75t_L g669 ( 
.A1(n_506),
.A2(n_252),
.B1(n_249),
.B2(n_327),
.C(n_256),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_486),
.B(n_446),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_532),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g672 ( 
.A(n_609),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_481),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_565),
.B(n_211),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_534),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_534),
.Y(n_676)
);

BUFx5_ASAP7_75t_L g677 ( 
.A(n_605),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_520),
.B(n_446),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_486),
.B(n_446),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_520),
.B(n_446),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_488),
.B(n_446),
.Y(n_681)
);

NOR2xp67_ASAP7_75t_SL g682 ( 
.A(n_520),
.B(n_198),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_488),
.B(n_447),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_565),
.B(n_215),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_496),
.B(n_218),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_491),
.B(n_447),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_491),
.B(n_447),
.Y(n_687)
);

INVx1_ASAP7_75t_SL g688 ( 
.A(n_552),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_588),
.B(n_350),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_499),
.B(n_224),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_546),
.B(n_447),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_561),
.B(n_227),
.Y(n_692)
);

NOR2x1p5_ASAP7_75t_L g693 ( 
.A(n_552),
.B(n_228),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_501),
.Y(n_694)
);

INVxp67_ASAP7_75t_SL g695 ( 
.A(n_546),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_536),
.Y(n_696)
);

AND2x4_ASAP7_75t_L g697 ( 
.A(n_497),
.B(n_201),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_510),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_546),
.B(n_447),
.Y(n_699)
);

BUFx6f_ASAP7_75t_SL g700 ( 
.A(n_581),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_616),
.B(n_447),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_480),
.B(n_207),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_616),
.B(n_447),
.Y(n_703)
);

OR2x6_ASAP7_75t_L g704 ( 
.A(n_506),
.B(n_367),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_503),
.B(n_455),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_531),
.B(n_234),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_539),
.B(n_235),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_616),
.B(n_455),
.Y(n_708)
);

INVx4_ASAP7_75t_L g709 ( 
.A(n_498),
.Y(n_709)
);

INVxp67_ASAP7_75t_SL g710 ( 
.A(n_498),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_503),
.B(n_587),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_557),
.B(n_239),
.Y(n_712)
);

INVx4_ASAP7_75t_L g713 ( 
.A(n_498),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_536),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_487),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_537),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_618),
.B(n_367),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_581),
.B(n_455),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_487),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_505),
.Y(n_720)
);

INVxp33_ASAP7_75t_L g721 ( 
.A(n_529),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_581),
.B(n_455),
.Y(n_722)
);

AND2x6_ASAP7_75t_L g723 ( 
.A(n_581),
.B(n_207),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_583),
.A2(n_202),
.B1(n_298),
.B2(n_302),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_537),
.B(n_455),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_559),
.A2(n_306),
.B1(n_286),
.B2(n_289),
.Y(n_726)
);

BUFx6f_ASAP7_75t_SL g727 ( 
.A(n_501),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_501),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_501),
.B(n_210),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_538),
.B(n_455),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_629),
.B(n_596),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_538),
.B(n_543),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_596),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_490),
.B(n_458),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_505),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_482),
.B(n_381),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_600),
.A2(n_416),
.B(n_448),
.Y(n_737)
);

OAI21xp33_ASAP7_75t_L g738 ( 
.A1(n_621),
.A2(n_493),
.B(n_589),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_490),
.B(n_458),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_543),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_L g741 ( 
.A1(n_593),
.A2(n_316),
.B1(n_221),
.B2(n_212),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_527),
.B(n_245),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_548),
.B(n_458),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_548),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_550),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_509),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_550),
.B(n_554),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_554),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_622),
.B(n_458),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_533),
.B(n_210),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_528),
.B(n_246),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_567),
.A2(n_275),
.B1(n_225),
.B2(n_219),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_509),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_556),
.B(n_458),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_542),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_622),
.B(n_458),
.Y(n_756)
);

NOR2x1p5_ASAP7_75t_L g757 ( 
.A(n_485),
.B(n_247),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_567),
.A2(n_225),
.B1(n_275),
.B2(n_268),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_567),
.A2(n_281),
.B1(n_208),
.B2(n_204),
.Y(n_759)
);

A2O1A1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_533),
.A2(n_281),
.B(n_219),
.C(n_241),
.Y(n_760)
);

NOR2xp67_ASAP7_75t_L g761 ( 
.A(n_562),
.B(n_381),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_622),
.B(n_403),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_510),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_516),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_556),
.B(n_458),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_558),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_558),
.B(n_448),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_622),
.B(n_231),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_585),
.B(n_231),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_563),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_563),
.B(n_448),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_568),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_568),
.B(n_448),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_511),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_571),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_564),
.B(n_231),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_571),
.B(n_448),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_578),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_572),
.A2(n_293),
.B1(n_291),
.B2(n_290),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_578),
.B(n_437),
.Y(n_780)
);

NOR2xp67_ASAP7_75t_SL g781 ( 
.A(n_626),
.B(n_212),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_582),
.B(n_438),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_582),
.Y(n_783)
);

INVxp67_ASAP7_75t_L g784 ( 
.A(n_493),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_604),
.B(n_438),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_577),
.B(n_254),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_604),
.B(n_612),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_612),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_613),
.B(n_439),
.Y(n_789)
);

INVxp33_ASAP7_75t_L g790 ( 
.A(n_621),
.Y(n_790)
);

BUFx8_ASAP7_75t_L g791 ( 
.A(n_492),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_613),
.B(n_439),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_615),
.B(n_440),
.Y(n_793)
);

NOR2xp67_ASAP7_75t_L g794 ( 
.A(n_626),
.B(n_314),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_615),
.B(n_440),
.Y(n_795)
);

NOR3xp33_ASAP7_75t_L g796 ( 
.A(n_610),
.B(n_307),
.C(n_301),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_619),
.B(n_255),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_504),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_627),
.B(n_603),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_627),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_660),
.B(n_592),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_635),
.A2(n_535),
.B1(n_551),
.B2(n_549),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_717),
.B(n_625),
.Y(n_803)
);

BUFx4f_ASAP7_75t_L g804 ( 
.A(n_632),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_663),
.A2(n_624),
.B(n_631),
.Y(n_805)
);

AO21x1_ASAP7_75t_L g806 ( 
.A1(n_644),
.A2(n_221),
.B(n_216),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_791),
.Y(n_807)
);

A2O1A1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_738),
.A2(n_208),
.B(n_274),
.C(n_264),
.Y(n_808)
);

NOR3xp33_ASAP7_75t_L g809 ( 
.A(n_666),
.B(n_606),
.C(n_223),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_SL g810 ( 
.A(n_688),
.B(n_270),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_636),
.A2(n_624),
.B(n_611),
.Y(n_811)
);

OAI21xp5_ASAP7_75t_L g812 ( 
.A1(n_734),
.A2(n_611),
.B(n_535),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_644),
.B(n_504),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_655),
.B(n_507),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_637),
.A2(n_624),
.B(n_611),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_728),
.Y(n_816)
);

NOR2x1_ASAP7_75t_L g817 ( 
.A(n_634),
.B(n_511),
.Y(n_817)
);

INVx3_ASAP7_75t_L g818 ( 
.A(n_728),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_677),
.B(n_498),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_787),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_787),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_639),
.A2(n_624),
.B(n_623),
.Y(n_822)
);

OR2x2_ASAP7_75t_L g823 ( 
.A(n_633),
.B(n_584),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_640),
.A2(n_624),
.B(n_623),
.Y(n_824)
);

NOR2x1_ASAP7_75t_L g825 ( 
.A(n_757),
.B(n_549),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_798),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_664),
.A2(n_623),
.B(n_614),
.Y(n_827)
);

INVxp67_ASAP7_75t_L g828 ( 
.A(n_656),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_666),
.B(n_507),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_638),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_655),
.B(n_605),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_791),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_677),
.B(n_498),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_762),
.B(n_605),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_797),
.B(n_605),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_797),
.B(n_605),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_677),
.B(n_515),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_649),
.A2(n_614),
.B(n_551),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_651),
.A2(n_614),
.B(n_519),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_711),
.B(n_605),
.Y(n_840)
);

BUFx2_ASAP7_75t_L g841 ( 
.A(n_704),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_651),
.A2(n_519),
.B(n_515),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_677),
.B(n_642),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_677),
.B(n_515),
.Y(n_844)
);

AOI21x1_ASAP7_75t_L g845 ( 
.A1(n_749),
.A2(n_517),
.B(n_516),
.Y(n_845)
);

INVx4_ASAP7_75t_L g846 ( 
.A(n_660),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_646),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_657),
.Y(n_848)
);

BUFx4f_ASAP7_75t_L g849 ( 
.A(n_704),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_658),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_662),
.A2(n_519),
.B(n_515),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_662),
.A2(n_519),
.B(n_515),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_668),
.Y(n_853)
);

O2A1O1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_661),
.A2(n_232),
.B(n_296),
.C(n_253),
.Y(n_854)
);

AOI21xp33_ASAP7_75t_L g855 ( 
.A1(n_790),
.A2(n_223),
.B(n_216),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_650),
.B(n_605),
.Y(n_856)
);

O2A1O1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_661),
.A2(n_253),
.B(n_232),
.C(n_229),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_653),
.B(n_671),
.Y(n_858)
);

NAND2xp33_ASAP7_75t_L g859 ( 
.A(n_677),
.B(n_519),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_675),
.B(n_512),
.Y(n_860)
);

NAND2x1_ASAP7_75t_L g861 ( 
.A(n_709),
.B(n_512),
.Y(n_861)
);

BUFx12f_ASAP7_75t_L g862 ( 
.A(n_704),
.Y(n_862)
);

INVx4_ASAP7_75t_L g863 ( 
.A(n_660),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_798),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_676),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_696),
.B(n_512),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_672),
.B(n_784),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_714),
.B(n_514),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_633),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_L g870 ( 
.A1(n_734),
.A2(n_590),
.B(n_514),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_678),
.A2(n_691),
.B(n_680),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_716),
.B(n_514),
.Y(n_872)
);

OAI21xp33_ASAP7_75t_L g873 ( 
.A1(n_736),
.A2(n_284),
.B(n_258),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_739),
.A2(n_545),
.B(n_555),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_740),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_635),
.B(n_579),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_678),
.A2(n_691),
.B(n_680),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_699),
.A2(n_579),
.B(n_628),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_755),
.B(n_579),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_744),
.B(n_745),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_748),
.Y(n_881)
);

OAI21xp33_ASAP7_75t_L g882 ( 
.A1(n_712),
.A2(n_313),
.B(n_309),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_766),
.Y(n_883)
);

O2A1O1Ixp5_ASAP7_75t_L g884 ( 
.A1(n_768),
.A2(n_739),
.B(n_769),
.C(n_682),
.Y(n_884)
);

OAI21xp33_ASAP7_75t_L g885 ( 
.A1(n_712),
.A2(n_305),
.B(n_320),
.Y(n_885)
);

O2A1O1Ixp5_ASAP7_75t_L g886 ( 
.A1(n_768),
.A2(n_545),
.B(n_555),
.C(n_590),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_685),
.A2(n_598),
.B1(n_555),
.B2(n_590),
.Y(n_887)
);

AOI21x1_ASAP7_75t_L g888 ( 
.A1(n_749),
.A2(n_630),
.B(n_517),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_641),
.A2(n_545),
.B(n_594),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_674),
.B(n_594),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_699),
.A2(n_628),
.B(n_579),
.Y(n_891)
);

O2A1O1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_760),
.A2(n_229),
.B(n_259),
.C(n_288),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_770),
.B(n_594),
.Y(n_893)
);

AOI21xp33_ASAP7_75t_L g894 ( 
.A1(n_786),
.A2(n_296),
.B(n_259),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_674),
.B(n_598),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_700),
.Y(n_896)
);

OAI21xp5_ASAP7_75t_L g897 ( 
.A1(n_641),
.A2(n_598),
.B(n_599),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_695),
.A2(n_316),
.B1(n_599),
.B2(n_288),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_660),
.B(n_608),
.Y(n_899)
);

A2O1A1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_731),
.A2(n_241),
.B(n_249),
.C(n_327),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_718),
.A2(n_628),
.B(n_579),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_659),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_722),
.A2(n_628),
.B(n_595),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_772),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_701),
.A2(n_628),
.B(n_595),
.Y(n_905)
);

OAI21xp33_ASAP7_75t_L g906 ( 
.A1(n_786),
.A2(n_318),
.B(n_263),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_646),
.A2(n_599),
.B1(n_595),
.B2(n_322),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_775),
.B(n_778),
.Y(n_908)
);

BUFx12f_ASAP7_75t_L g909 ( 
.A(n_693),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_783),
.B(n_595),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_788),
.B(n_595),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_701),
.A2(n_416),
.B(n_530),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_703),
.A2(n_416),
.B(n_530),
.Y(n_913)
);

OAI21xp5_ASAP7_75t_L g914 ( 
.A1(n_703),
.A2(n_630),
.B(n_620),
.Y(n_914)
);

INVx1_ASAP7_75t_SL g915 ( 
.A(n_689),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_750),
.B(n_652),
.Y(n_916)
);

AO21x1_ASAP7_75t_L g917 ( 
.A1(n_769),
.A2(n_252),
.B(n_256),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_800),
.B(n_518),
.Y(n_918)
);

AO21x1_ASAP7_75t_L g919 ( 
.A1(n_685),
.A2(n_264),
.B(n_274),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_684),
.B(n_272),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_708),
.A2(n_416),
.B(n_530),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_708),
.A2(n_416),
.B(n_530),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_732),
.B(n_518),
.Y(n_923)
);

BUFx2_ASAP7_75t_L g924 ( 
.A(n_697),
.Y(n_924)
);

AOI21x1_ASAP7_75t_L g925 ( 
.A1(n_756),
.A2(n_620),
.B(n_607),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_747),
.Y(n_926)
);

INVx1_ASAP7_75t_SL g927 ( 
.A(n_697),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_702),
.B(n_522),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_665),
.A2(n_607),
.B(n_522),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_654),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_684),
.B(n_304),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_750),
.B(n_540),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_667),
.A2(n_416),
.B(n_602),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_690),
.A2(n_326),
.B1(n_601),
.B2(n_573),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_690),
.B(n_308),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_670),
.A2(n_416),
.B(n_602),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_702),
.B(n_540),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_679),
.A2(n_602),
.B(n_530),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_700),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_681),
.A2(n_602),
.B(n_530),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_648),
.B(n_560),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_761),
.B(n_277),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_648),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_799),
.B(n_742),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_683),
.A2(n_580),
.B(n_601),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_673),
.Y(n_946)
);

AO21x1_ASAP7_75t_L g947 ( 
.A1(n_692),
.A2(n_321),
.B(n_262),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_686),
.A2(n_576),
.B(n_566),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_742),
.B(n_310),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_687),
.A2(n_602),
.B(n_597),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_694),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_752),
.A2(n_566),
.B1(n_591),
.B2(n_586),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_715),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_719),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_752),
.B(n_560),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_751),
.B(n_311),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_L g957 ( 
.A1(n_758),
.A2(n_573),
.B1(n_591),
.B2(n_586),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_751),
.B(n_575),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_692),
.B(n_575),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_705),
.A2(n_597),
.B(n_580),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_756),
.A2(n_597),
.B(n_576),
.Y(n_961)
);

BUFx4f_ASAP7_75t_L g962 ( 
.A(n_723),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_758),
.A2(n_324),
.B1(n_319),
.B2(n_323),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_643),
.A2(n_597),
.B(n_442),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_710),
.A2(n_713),
.B(n_709),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_647),
.A2(n_597),
.B(n_442),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_706),
.B(n_445),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_713),
.A2(n_597),
.B(n_436),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_698),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_725),
.A2(n_432),
.B(n_436),
.Y(n_970)
);

O2A1O1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_760),
.A2(n_454),
.B(n_453),
.C(n_452),
.Y(n_971)
);

NOR2x2_ASAP7_75t_L g972 ( 
.A(n_645),
.B(n_277),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_780),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_706),
.B(n_454),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_759),
.B(n_231),
.Y(n_975)
);

HB1xp67_ASAP7_75t_L g976 ( 
.A(n_727),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_707),
.B(n_453),
.Y(n_977)
);

AO21x1_ASAP7_75t_L g978 ( 
.A1(n_707),
.A2(n_262),
.B(n_321),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_730),
.A2(n_432),
.B(n_436),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_743),
.A2(n_765),
.B(n_754),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_SL g981 ( 
.A(n_721),
.B(n_270),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_737),
.A2(n_432),
.B(n_452),
.Y(n_982)
);

HB1xp67_ASAP7_75t_L g983 ( 
.A(n_727),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_759),
.B(n_782),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_767),
.A2(n_449),
.B(n_445),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_785),
.B(n_449),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_789),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_733),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_792),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_771),
.A2(n_466),
.B(n_317),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_724),
.A2(n_315),
.B1(n_312),
.B2(n_466),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_855),
.A2(n_741),
.B(n_796),
.C(n_793),
.Y(n_992)
);

AOI22xp33_ASAP7_75t_L g993 ( 
.A1(n_894),
.A2(n_935),
.B1(n_956),
.B2(n_949),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_867),
.B(n_779),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_867),
.B(n_726),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_915),
.B(n_794),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_826),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_846),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_820),
.B(n_729),
.Y(n_999)
);

XNOR2xp5_ASAP7_75t_L g1000 ( 
.A(n_807),
.B(n_729),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_969),
.Y(n_1001)
);

NOR2x1_ASAP7_75t_R g1002 ( 
.A(n_807),
.B(n_231),
.Y(n_1002)
);

CKINVDCx14_ASAP7_75t_R g1003 ( 
.A(n_832),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_821),
.B(n_698),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_935),
.B(n_795),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_949),
.A2(n_777),
.B(n_773),
.C(n_720),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_956),
.A2(n_669),
.B1(n_723),
.B2(n_781),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_969),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_926),
.B(n_723),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_973),
.B(n_723),
.Y(n_1010)
);

INVx4_ASAP7_75t_L g1011 ( 
.A(n_846),
.Y(n_1011)
);

A2O1A1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_920),
.A2(n_735),
.B(n_746),
.C(n_764),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_920),
.B(n_774),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_987),
.B(n_723),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_989),
.B(n_753),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_944),
.B(n_774),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_821),
.B(n_774),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_984),
.A2(n_774),
.B1(n_763),
.B2(n_698),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_931),
.A2(n_829),
.B(n_809),
.C(n_916),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_829),
.A2(n_763),
.B1(n_698),
.B2(n_776),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_931),
.A2(n_776),
.B(n_466),
.C(n_270),
.Y(n_1021)
);

O2A1O1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_916),
.A2(n_270),
.B(n_277),
.C(n_18),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_902),
.B(n_763),
.Y(n_1023)
);

CKINVDCx16_ASAP7_75t_R g1024 ( 
.A(n_832),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_826),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_R g1026 ( 
.A(n_896),
.B(n_763),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_909),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_828),
.B(n_17),
.Y(n_1028)
);

O2A1O1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_900),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_900),
.A2(n_20),
.B(n_22),
.C(n_26),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_813),
.A2(n_163),
.B1(n_140),
.B2(n_131),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_803),
.B(n_129),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_869),
.B(n_22),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_841),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_942),
.B(n_26),
.Y(n_1035)
);

AOI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_975),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_814),
.A2(n_125),
.B1(n_122),
.B2(n_119),
.Y(n_1037)
);

INVx4_ASAP7_75t_L g1038 ( 
.A(n_863),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_924),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_890),
.A2(n_30),
.B(n_32),
.C(n_37),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_927),
.B(n_111),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_801),
.B(n_109),
.Y(n_1042)
);

OAI21xp33_ASAP7_75t_L g1043 ( 
.A1(n_810),
.A2(n_40),
.B(n_41),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_808),
.A2(n_40),
.B(n_41),
.C(n_42),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_882),
.B(n_43),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_801),
.B(n_100),
.Y(n_1046)
);

BUFx12f_ASAP7_75t_L g1047 ( 
.A(n_896),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_823),
.B(n_43),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_890),
.A2(n_45),
.B(n_46),
.C(n_50),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_801),
.B(n_95),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_859),
.A2(n_94),
.B(n_92),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_880),
.B(n_50),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_885),
.B(n_52),
.Y(n_1053)
);

OAI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_908),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_849),
.B(n_85),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_849),
.B(n_80),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_895),
.A2(n_54),
.B(n_55),
.C(n_58),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_SL g1058 ( 
.A1(n_895),
.A2(n_67),
.B(n_70),
.C(n_68),
.Y(n_1058)
);

INVx4_ASAP7_75t_L g1059 ( 
.A(n_863),
.Y(n_1059)
);

AOI21xp33_ASAP7_75t_L g1060 ( 
.A1(n_906),
.A2(n_59),
.B(n_60),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_864),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_SL g1062 ( 
.A1(n_876),
.A2(n_79),
.B(n_63),
.C(n_64),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_858),
.B(n_60),
.Y(n_1063)
);

NOR2xp67_ASAP7_75t_L g1064 ( 
.A(n_909),
.B(n_976),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_975),
.A2(n_919),
.B1(n_947),
.B2(n_978),
.Y(n_1065)
);

OAI22x1_ASAP7_75t_L g1066 ( 
.A1(n_988),
.A2(n_939),
.B1(n_972),
.B2(n_983),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_SL g1067 ( 
.A(n_939),
.B(n_862),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_884),
.A2(n_834),
.B(n_974),
.C(n_977),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_859),
.A2(n_805),
.B(n_840),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_962),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_873),
.B(n_830),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_876),
.A2(n_877),
.B(n_871),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_967),
.B(n_804),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_899),
.B(n_825),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_817),
.A2(n_951),
.B1(n_836),
.B2(n_835),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_831),
.A2(n_827),
.B(n_843),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_848),
.B(n_850),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_853),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_865),
.Y(n_1079)
);

AO22x1_ASAP7_75t_L g1080 ( 
.A1(n_899),
.A2(n_963),
.B1(n_883),
.B2(n_875),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_881),
.B(n_904),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_804),
.B(n_847),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_986),
.B(n_958),
.Y(n_1083)
);

O2A1O1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_808),
.A2(n_854),
.B(n_857),
.C(n_991),
.Y(n_1084)
);

O2A1O1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_959),
.A2(n_898),
.B(n_879),
.C(n_990),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_923),
.B(n_847),
.Y(n_1086)
);

AOI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_899),
.A2(n_843),
.B1(n_856),
.B2(n_943),
.Y(n_1087)
);

O2A1O1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_879),
.A2(n_806),
.B(n_937),
.C(n_928),
.Y(n_1088)
);

NAND2x1p5_ASAP7_75t_L g1089 ( 
.A(n_962),
.B(n_943),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_981),
.B(n_816),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_816),
.B(n_818),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_818),
.B(n_934),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_918),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_886),
.A2(n_955),
.B(n_812),
.C(n_980),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_955),
.A2(n_838),
.B(n_932),
.C(n_815),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_819),
.A2(n_844),
.B(n_833),
.Y(n_1096)
);

OAI21xp33_ASAP7_75t_SL g1097 ( 
.A1(n_932),
.A2(n_964),
.B(n_966),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_910),
.B(n_911),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_930),
.B(n_946),
.Y(n_1099)
);

AND2x6_ASAP7_75t_L g1100 ( 
.A(n_887),
.B(n_930),
.Y(n_1100)
);

INVx2_ASAP7_75t_SL g1101 ( 
.A(n_946),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_953),
.B(n_954),
.Y(n_1102)
);

BUFx2_ASAP7_75t_L g1103 ( 
.A(n_972),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_954),
.B(n_872),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_941),
.B(n_868),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_917),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_860),
.B(n_866),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_893),
.B(n_844),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_889),
.A2(n_897),
.B(n_870),
.C(n_874),
.Y(n_1109)
);

OAI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_952),
.A2(n_957),
.B1(n_802),
.B2(n_914),
.Y(n_1110)
);

NAND2x1p5_ASAP7_75t_L g1111 ( 
.A(n_837),
.B(n_861),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_929),
.B(n_945),
.Y(n_1112)
);

BUFx10_ASAP7_75t_L g1113 ( 
.A(n_892),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_907),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_R g1115 ( 
.A(n_845),
.B(n_925),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_948),
.B(n_965),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_822),
.A2(n_824),
.B(n_811),
.Y(n_1117)
);

INVxp67_ASAP7_75t_L g1118 ( 
.A(n_982),
.Y(n_1118)
);

NOR3xp33_ASAP7_75t_SL g1119 ( 
.A(n_905),
.B(n_878),
.C(n_842),
.Y(n_1119)
);

NOR2xp67_ASAP7_75t_SL g1120 ( 
.A(n_839),
.B(n_903),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_901),
.A2(n_851),
.B(n_852),
.Y(n_1121)
);

OAI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_891),
.A2(n_960),
.B(n_985),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_971),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_970),
.B(n_979),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_912),
.A2(n_913),
.B(n_921),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_888),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_961),
.B(n_922),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_938),
.B(n_940),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_950),
.A2(n_933),
.B(n_936),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_968),
.B(n_926),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_869),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_859),
.A2(n_520),
.B(n_495),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_935),
.A2(n_956),
.B(n_949),
.C(n_931),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_926),
.B(n_973),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_926),
.B(n_973),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_944),
.A2(n_984),
.B1(n_926),
.B2(n_829),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_826),
.Y(n_1137)
);

OR2x2_ASAP7_75t_L g1138 ( 
.A(n_915),
.B(n_902),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_859),
.A2(n_520),
.B(n_495),
.Y(n_1139)
);

CKINVDCx20_ASAP7_75t_R g1140 ( 
.A(n_807),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_926),
.B(n_973),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_915),
.B(n_672),
.Y(n_1142)
);

O2A1O1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_855),
.A2(n_894),
.B(n_949),
.C(n_935),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_SL g1144 ( 
.A1(n_1143),
.A2(n_1044),
.B(n_1051),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1133),
.A2(n_1116),
.B(n_1132),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1005),
.B(n_1136),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_993),
.A2(n_1068),
.B(n_1019),
.Y(n_1147)
);

AO31x2_ASAP7_75t_L g1148 ( 
.A1(n_1094),
.A2(n_1095),
.A3(n_1128),
.B(n_1109),
.Y(n_1148)
);

INVx6_ASAP7_75t_L g1149 ( 
.A(n_1047),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_1070),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1117),
.A2(n_1125),
.B(n_1129),
.Y(n_1151)
);

BUFx10_ASAP7_75t_L g1152 ( 
.A(n_1033),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1005),
.B(n_1134),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_993),
.A2(n_1097),
.B(n_1072),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1121),
.A2(n_1069),
.B(n_1122),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_SL g1156 ( 
.A1(n_1013),
.A2(n_1085),
.B(n_1020),
.Y(n_1156)
);

O2A1O1Ixp33_ASAP7_75t_SL g1157 ( 
.A1(n_1040),
.A2(n_1057),
.B(n_1049),
.C(n_1060),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_997),
.Y(n_1158)
);

OAI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_994),
.A2(n_995),
.B1(n_1135),
.B2(n_1141),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1139),
.A2(n_1076),
.B(n_1083),
.Y(n_1160)
);

BUFx12f_ASAP7_75t_L g1161 ( 
.A(n_1034),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_L g1162 ( 
.A1(n_994),
.A2(n_1045),
.B1(n_1053),
.B2(n_1048),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1078),
.Y(n_1163)
);

AO31x2_ASAP7_75t_L g1164 ( 
.A1(n_1127),
.A2(n_1006),
.A3(n_1108),
.B(n_1106),
.Y(n_1164)
);

NOR2xp67_ASAP7_75t_L g1165 ( 
.A(n_1138),
.B(n_1090),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1110),
.A2(n_1112),
.B(n_1016),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1035),
.B(n_1039),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1110),
.A2(n_1130),
.B(n_1118),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_1131),
.Y(n_1169)
);

BUFx4_ASAP7_75t_SL g1170 ( 
.A(n_1140),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1074),
.B(n_999),
.Y(n_1171)
);

O2A1O1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1073),
.A2(n_1043),
.B(n_1084),
.C(n_1063),
.Y(n_1172)
);

O2A1O1Ixp5_ASAP7_75t_SL g1173 ( 
.A1(n_1126),
.A2(n_1092),
.B(n_1118),
.C(n_1123),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1075),
.A2(n_1108),
.B(n_1096),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_992),
.A2(n_1071),
.B(n_1088),
.C(n_1021),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_SL g1176 ( 
.A1(n_1036),
.A2(n_1029),
.B(n_1030),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1022),
.A2(n_1010),
.B(n_1014),
.C(n_1009),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1065),
.A2(n_1012),
.B(n_1127),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1105),
.A2(n_1018),
.B(n_1107),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_1142),
.B(n_1039),
.Y(n_1180)
);

AO31x2_ASAP7_75t_L g1181 ( 
.A1(n_1124),
.A2(n_1104),
.A3(n_1086),
.B(n_1037),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1032),
.A2(n_1042),
.B1(n_1046),
.B2(n_1050),
.Y(n_1182)
);

OA22x2_ASAP7_75t_L g1183 ( 
.A1(n_1066),
.A2(n_1103),
.B1(n_1000),
.B2(n_1079),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1081),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_1026),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1065),
.A2(n_1119),
.B(n_1087),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1098),
.A2(n_1093),
.B(n_1080),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1077),
.B(n_996),
.Y(n_1188)
);

OR2x2_ASAP7_75t_L g1189 ( 
.A(n_1052),
.B(n_1023),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1119),
.A2(n_1007),
.B(n_1100),
.Y(n_1190)
);

OAI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1007),
.A2(n_1100),
.B(n_1099),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1111),
.A2(n_1089),
.B(n_1102),
.Y(n_1192)
);

AO31x2_ASAP7_75t_L g1193 ( 
.A1(n_1031),
.A2(n_1077),
.A3(n_1091),
.B(n_1137),
.Y(n_1193)
);

OAI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1100),
.A2(n_1015),
.B(n_1061),
.Y(n_1194)
);

CKINVDCx20_ASAP7_75t_R g1195 ( 
.A(n_1024),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1101),
.B(n_1025),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_999),
.B(n_1028),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1004),
.A2(n_1017),
.B(n_1001),
.Y(n_1198)
);

AOI31xp67_ASAP7_75t_L g1199 ( 
.A1(n_1041),
.A2(n_1120),
.A3(n_1058),
.B(n_1056),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1114),
.A2(n_1055),
.B(n_1082),
.Y(n_1200)
);

O2A1O1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1054),
.A2(n_1062),
.B(n_1036),
.C(n_1067),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1008),
.A2(n_1115),
.B(n_1100),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1064),
.A2(n_1113),
.B(n_1070),
.Y(n_1203)
);

CKINVDCx20_ASAP7_75t_R g1204 ( 
.A(n_1003),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_998),
.B(n_1011),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1011),
.A2(n_1038),
.B(n_1059),
.Y(n_1206)
);

OA21x2_ASAP7_75t_L g1207 ( 
.A1(n_1054),
.A2(n_1070),
.B(n_1038),
.Y(n_1207)
);

AOI21xp33_ASAP7_75t_L g1208 ( 
.A1(n_1002),
.A2(n_1059),
.B(n_1027),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1005),
.B(n_1133),
.Y(n_1209)
);

BUFx12f_ASAP7_75t_L g1210 ( 
.A(n_1047),
.Y(n_1210)
);

BUFx2_ASAP7_75t_L g1211 ( 
.A(n_1131),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1005),
.B(n_1134),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1133),
.A2(n_663),
.B(n_859),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1133),
.A2(n_663),
.B(n_859),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1133),
.A2(n_1143),
.B(n_993),
.C(n_1005),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_993),
.A2(n_1133),
.B1(n_1005),
.B2(n_1019),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_997),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1133),
.A2(n_663),
.B(n_859),
.Y(n_1218)
);

AOI31xp67_ASAP7_75t_L g1219 ( 
.A1(n_1075),
.A2(n_1116),
.A3(n_769),
.B(n_1092),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1078),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1078),
.Y(n_1221)
);

NOR2xp67_ASAP7_75t_L g1222 ( 
.A(n_1138),
.B(n_828),
.Y(n_1222)
);

BUFx4_ASAP7_75t_SL g1223 ( 
.A(n_1140),
.Y(n_1223)
);

NAND2xp33_ASAP7_75t_L g1224 ( 
.A(n_1133),
.B(n_993),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1005),
.B(n_1133),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1133),
.A2(n_663),
.B(n_859),
.Y(n_1226)
);

NAND3xp33_ASAP7_75t_L g1227 ( 
.A(n_993),
.B(n_1133),
.C(n_949),
.Y(n_1227)
);

O2A1O1Ixp5_ASAP7_75t_SL g1228 ( 
.A1(n_1060),
.A2(n_894),
.B(n_855),
.C(n_769),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1133),
.A2(n_993),
.B(n_1143),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_1133),
.A2(n_806),
.A3(n_1094),
.B(n_1095),
.Y(n_1230)
);

AO32x2_ASAP7_75t_L g1231 ( 
.A1(n_1136),
.A2(n_1018),
.A3(n_1020),
.B1(n_898),
.B2(n_957),
.Y(n_1231)
);

INVx3_ASAP7_75t_SL g1232 ( 
.A(n_1024),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_997),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1005),
.B(n_1134),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1133),
.A2(n_663),
.B(n_859),
.Y(n_1235)
);

AOI211x1_ASAP7_75t_L g1236 ( 
.A1(n_1134),
.A2(n_738),
.B(n_1141),
.C(n_1135),
.Y(n_1236)
);

OAI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1133),
.A2(n_993),
.B(n_1143),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1133),
.A2(n_663),
.B(n_859),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_998),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1005),
.B(n_1133),
.Y(n_1240)
);

A2O1A1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1133),
.A2(n_1143),
.B(n_993),
.C(n_1005),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_998),
.Y(n_1242)
);

CKINVDCx11_ASAP7_75t_R g1243 ( 
.A(n_1140),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1133),
.A2(n_663),
.B(n_859),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1078),
.Y(n_1245)
);

AOI221xp5_ASAP7_75t_SL g1246 ( 
.A1(n_1133),
.A2(n_993),
.B1(n_1143),
.B2(n_1054),
.C(n_808),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1133),
.A2(n_993),
.B(n_1143),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1133),
.A2(n_993),
.B(n_1143),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1133),
.A2(n_993),
.B(n_1143),
.Y(n_1249)
);

AO31x2_ASAP7_75t_L g1250 ( 
.A1(n_1133),
.A2(n_806),
.A3(n_1094),
.B(n_1095),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1074),
.B(n_999),
.Y(n_1251)
);

AO31x2_ASAP7_75t_L g1252 ( 
.A1(n_1133),
.A2(n_806),
.A3(n_1094),
.B(n_1095),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_997),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1133),
.A2(n_663),
.B(n_859),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_997),
.Y(n_1255)
);

AOI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_993),
.A2(n_1133),
.B1(n_949),
.B2(n_956),
.Y(n_1256)
);

O2A1O1Ixp5_ASAP7_75t_L g1257 ( 
.A1(n_1133),
.A2(n_949),
.B(n_956),
.C(n_935),
.Y(n_1257)
);

AO21x2_ASAP7_75t_L g1258 ( 
.A1(n_1133),
.A2(n_1117),
.B(n_1110),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1074),
.B(n_999),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1048),
.B(n_902),
.Y(n_1260)
);

A2O1A1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1133),
.A2(n_1143),
.B(n_993),
.C(n_1005),
.Y(n_1261)
);

INVxp67_ASAP7_75t_SL g1262 ( 
.A(n_1138),
.Y(n_1262)
);

AOI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1120),
.A2(n_1080),
.B(n_1069),
.Y(n_1263)
);

NOR2xp67_ASAP7_75t_SL g1264 ( 
.A(n_1047),
.B(n_862),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_997),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1133),
.A2(n_663),
.B(n_859),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1117),
.A2(n_1125),
.B(n_1129),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_997),
.Y(n_1268)
);

NOR2xp67_ASAP7_75t_L g1269 ( 
.A(n_1138),
.B(n_828),
.Y(n_1269)
);

O2A1O1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1133),
.A2(n_1143),
.B(n_1019),
.C(n_956),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1078),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1133),
.B(n_666),
.Y(n_1272)
);

CKINVDCx11_ASAP7_75t_R g1273 ( 
.A(n_1140),
.Y(n_1273)
);

O2A1O1Ixp33_ASAP7_75t_SL g1274 ( 
.A1(n_1133),
.A2(n_1019),
.B(n_1143),
.C(n_894),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1117),
.A2(n_1125),
.B(n_1129),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_997),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_SL g1277 ( 
.A1(n_1143),
.A2(n_1044),
.B(n_1051),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1005),
.B(n_1133),
.Y(n_1278)
);

AOI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_993),
.A2(n_1133),
.B1(n_949),
.B2(n_956),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1117),
.A2(n_1125),
.B(n_1129),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_993),
.A2(n_1133),
.B1(n_949),
.B2(n_956),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1133),
.B(n_666),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1078),
.Y(n_1283)
);

A2O1A1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1133),
.A2(n_1143),
.B(n_993),
.C(n_1005),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1005),
.B(n_1133),
.Y(n_1285)
);

NOR2xp67_ASAP7_75t_L g1286 ( 
.A(n_1138),
.B(n_828),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1224),
.A2(n_1227),
.B1(n_1216),
.B2(n_1272),
.Y(n_1287)
);

OAI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1256),
.A2(n_1279),
.B1(n_1281),
.B2(n_1225),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_SL g1289 ( 
.A1(n_1282),
.A2(n_1216),
.B1(n_1248),
.B2(n_1249),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1260),
.B(n_1167),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1159),
.B(n_1153),
.Y(n_1291)
);

BUFx3_ASAP7_75t_L g1292 ( 
.A(n_1185),
.Y(n_1292)
);

BUFx2_ASAP7_75t_SL g1293 ( 
.A(n_1204),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1158),
.Y(n_1294)
);

INVx4_ASAP7_75t_L g1295 ( 
.A(n_1239),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1212),
.B(n_1234),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1162),
.A2(n_1225),
.B1(n_1285),
.B2(n_1240),
.Y(n_1297)
);

INVx6_ASAP7_75t_L g1298 ( 
.A(n_1239),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_1273),
.Y(n_1299)
);

CKINVDCx20_ASAP7_75t_R g1300 ( 
.A(n_1195),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1220),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_SL g1302 ( 
.A1(n_1229),
.A2(n_1247),
.B1(n_1237),
.B2(n_1248),
.Y(n_1302)
);

BUFx12f_ASAP7_75t_L g1303 ( 
.A(n_1210),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1221),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1245),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1229),
.A2(n_1249),
.B1(n_1237),
.B2(n_1247),
.Y(n_1306)
);

AOI21xp33_ASAP7_75t_L g1307 ( 
.A1(n_1270),
.A2(n_1257),
.B(n_1209),
.Y(n_1307)
);

INVx8_ASAP7_75t_L g1308 ( 
.A(n_1161),
.Y(n_1308)
);

BUFx8_ASAP7_75t_SL g1309 ( 
.A(n_1211),
.Y(n_1309)
);

NAND2x1p5_ASAP7_75t_L g1310 ( 
.A(n_1203),
.B(n_1207),
.Y(n_1310)
);

CKINVDCx6p67_ASAP7_75t_R g1311 ( 
.A(n_1232),
.Y(n_1311)
);

BUFx12f_ASAP7_75t_L g1312 ( 
.A(n_1149),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1271),
.Y(n_1313)
);

AND2x4_ASAP7_75t_SL g1314 ( 
.A(n_1171),
.B(n_1251),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1209),
.A2(n_1240),
.B1(n_1285),
.B2(n_1278),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_1170),
.Y(n_1316)
);

BUFx4f_ASAP7_75t_SL g1317 ( 
.A(n_1169),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1278),
.A2(n_1147),
.B1(n_1146),
.B2(n_1154),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1283),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1239),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1215),
.A2(n_1261),
.B1(n_1284),
.B2(n_1241),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1188),
.A2(n_1165),
.B1(n_1182),
.B2(n_1197),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1147),
.A2(n_1146),
.B1(n_1154),
.B2(n_1190),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1217),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1222),
.A2(n_1286),
.B1(n_1269),
.B2(n_1184),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1190),
.A2(n_1258),
.B1(n_1144),
.B2(n_1277),
.Y(n_1326)
);

CKINVDCx11_ASAP7_75t_R g1327 ( 
.A(n_1152),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1233),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1253),
.Y(n_1329)
);

CKINVDCx20_ASAP7_75t_R g1330 ( 
.A(n_1149),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1255),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1262),
.A2(n_1175),
.B1(n_1180),
.B2(n_1236),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_SL g1333 ( 
.A1(n_1152),
.A2(n_1183),
.B1(n_1258),
.B2(n_1186),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1186),
.A2(n_1168),
.B1(n_1166),
.B2(n_1178),
.Y(n_1334)
);

BUFx2_ASAP7_75t_SL g1335 ( 
.A(n_1242),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1178),
.A2(n_1191),
.B1(n_1174),
.B2(n_1183),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1242),
.Y(n_1337)
);

CKINVDCx11_ASAP7_75t_R g1338 ( 
.A(n_1223),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1191),
.A2(n_1174),
.B1(n_1189),
.B2(n_1226),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_SL g1340 ( 
.A1(n_1200),
.A2(n_1207),
.B1(n_1171),
.B2(n_1259),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1265),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1268),
.Y(n_1342)
);

INVx3_ASAP7_75t_SL g1343 ( 
.A(n_1251),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_1259),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1213),
.A2(n_1254),
.B1(n_1244),
.B2(n_1235),
.Y(n_1345)
);

BUFx3_ASAP7_75t_L g1346 ( 
.A(n_1150),
.Y(n_1346)
);

BUFx12f_ASAP7_75t_L g1347 ( 
.A(n_1264),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1276),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_SL g1349 ( 
.A(n_1208),
.Y(n_1349)
);

BUFx2_ASAP7_75t_SL g1350 ( 
.A(n_1205),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_1202),
.Y(n_1351)
);

INVx1_ASAP7_75t_SL g1352 ( 
.A(n_1196),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_SL g1353 ( 
.A1(n_1214),
.A2(n_1266),
.B1(n_1218),
.B2(n_1238),
.Y(n_1353)
);

NAND2x1p5_ASAP7_75t_L g1354 ( 
.A(n_1198),
.B(n_1192),
.Y(n_1354)
);

INVx3_ASAP7_75t_L g1355 ( 
.A(n_1164),
.Y(n_1355)
);

OAI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1176),
.A2(n_1196),
.B1(n_1194),
.B2(n_1187),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1145),
.A2(n_1246),
.B1(n_1194),
.B2(n_1274),
.Y(n_1357)
);

CKINVDCx11_ASAP7_75t_R g1358 ( 
.A(n_1208),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1164),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_SL g1360 ( 
.A1(n_1246),
.A2(n_1201),
.B1(n_1157),
.B2(n_1172),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1164),
.B(n_1179),
.Y(n_1361)
);

INVx6_ASAP7_75t_L g1362 ( 
.A(n_1206),
.Y(n_1362)
);

OAI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1160),
.A2(n_1228),
.B1(n_1156),
.B2(n_1263),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1148),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1219),
.Y(n_1365)
);

OAI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1231),
.A2(n_1173),
.B1(n_1230),
.B2(n_1252),
.Y(n_1366)
);

CKINVDCx11_ASAP7_75t_R g1367 ( 
.A(n_1199),
.Y(n_1367)
);

CKINVDCx20_ASAP7_75t_R g1368 ( 
.A(n_1177),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_1230),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_1230),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1231),
.A2(n_1193),
.B1(n_1181),
.B2(n_1250),
.Y(n_1371)
);

BUFx4f_ASAP7_75t_SL g1372 ( 
.A(n_1250),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1155),
.A2(n_1151),
.B1(n_1275),
.B2(n_1267),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1252),
.Y(n_1374)
);

BUFx4_ASAP7_75t_SL g1375 ( 
.A(n_1193),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1181),
.B(n_1280),
.Y(n_1376)
);

BUFx6f_ASAP7_75t_L g1377 ( 
.A(n_1231),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1162),
.A2(n_993),
.B1(n_1133),
.B2(n_1256),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1163),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1158),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1162),
.A2(n_993),
.B1(n_1133),
.B2(n_1256),
.Y(n_1381)
);

CKINVDCx8_ASAP7_75t_R g1382 ( 
.A(n_1185),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1163),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1163),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1224),
.A2(n_1227),
.B1(n_993),
.B2(n_1216),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1163),
.Y(n_1386)
);

CKINVDCx6p67_ASAP7_75t_R g1387 ( 
.A(n_1243),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1163),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1239),
.Y(n_1389)
);

BUFx6f_ASAP7_75t_L g1390 ( 
.A(n_1239),
.Y(n_1390)
);

INVx4_ASAP7_75t_L g1391 ( 
.A(n_1239),
.Y(n_1391)
);

OAI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1256),
.A2(n_1279),
.B1(n_1281),
.B2(n_1227),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1224),
.A2(n_1227),
.B1(n_993),
.B2(n_1216),
.Y(n_1393)
);

AOI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1256),
.A2(n_993),
.B1(n_1133),
.B2(n_935),
.Y(n_1394)
);

INVx1_ASAP7_75t_SL g1395 ( 
.A(n_1211),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1163),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1162),
.A2(n_993),
.B1(n_1133),
.B2(n_1256),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1163),
.Y(n_1398)
);

BUFx12f_ASAP7_75t_L g1399 ( 
.A(n_1243),
.Y(n_1399)
);

CKINVDCx11_ASAP7_75t_R g1400 ( 
.A(n_1243),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1163),
.Y(n_1401)
);

CKINVDCx11_ASAP7_75t_R g1402 ( 
.A(n_1243),
.Y(n_1402)
);

OAI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1256),
.A2(n_1279),
.B1(n_1281),
.B2(n_1227),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_SL g1404 ( 
.A1(n_1272),
.A2(n_1282),
.B1(n_1227),
.B2(n_935),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1224),
.A2(n_1227),
.B1(n_993),
.B2(n_1216),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1162),
.A2(n_993),
.B1(n_1133),
.B2(n_1256),
.Y(n_1406)
);

CKINVDCx11_ASAP7_75t_R g1407 ( 
.A(n_1243),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1163),
.Y(n_1408)
);

INVx6_ASAP7_75t_L g1409 ( 
.A(n_1239),
.Y(n_1409)
);

BUFx12f_ASAP7_75t_L g1410 ( 
.A(n_1243),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1224),
.A2(n_1227),
.B1(n_993),
.B2(n_1216),
.Y(n_1411)
);

INVx5_ASAP7_75t_L g1412 ( 
.A(n_1239),
.Y(n_1412)
);

INVx5_ASAP7_75t_L g1413 ( 
.A(n_1239),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1170),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1354),
.A2(n_1373),
.B(n_1376),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1369),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1364),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1351),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1374),
.Y(n_1419)
);

BUFx2_ASAP7_75t_L g1420 ( 
.A(n_1370),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1359),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1365),
.Y(n_1422)
);

OAI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1394),
.A2(n_1404),
.B(n_1289),
.Y(n_1423)
);

NAND2x1_ASAP7_75t_L g1424 ( 
.A(n_1362),
.B(n_1345),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1377),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1377),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1368),
.A2(n_1397),
.B1(n_1406),
.B2(n_1381),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1355),
.Y(n_1428)
);

NAND2x1_ASAP7_75t_L g1429 ( 
.A(n_1362),
.B(n_1345),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1361),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1318),
.B(n_1302),
.Y(n_1431)
);

AO21x2_ASAP7_75t_L g1432 ( 
.A1(n_1363),
.A2(n_1403),
.B(n_1392),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1354),
.Y(n_1433)
);

O2A1O1Ixp33_ASAP7_75t_SL g1434 ( 
.A1(n_1378),
.A2(n_1291),
.B(n_1403),
.C(n_1392),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1372),
.Y(n_1435)
);

OAI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1306),
.A2(n_1385),
.B(n_1411),
.Y(n_1436)
);

OAI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1306),
.A2(n_1385),
.B(n_1393),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1296),
.B(n_1352),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1371),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1310),
.Y(n_1440)
);

INVx2_ASAP7_75t_SL g1441 ( 
.A(n_1412),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1321),
.B(n_1334),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1357),
.A2(n_1326),
.B(n_1334),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1375),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1357),
.A2(n_1326),
.B(n_1287),
.Y(n_1445)
);

AOI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1393),
.A2(n_1411),
.B1(n_1405),
.B2(n_1287),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1292),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1405),
.A2(n_1288),
.B1(n_1336),
.B2(n_1323),
.Y(n_1448)
);

AO21x2_ASAP7_75t_L g1449 ( 
.A1(n_1363),
.A2(n_1366),
.B(n_1307),
.Y(n_1449)
);

INVx2_ASAP7_75t_SL g1450 ( 
.A(n_1412),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1301),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1315),
.A2(n_1339),
.B(n_1318),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1322),
.B(n_1297),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1304),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1305),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1313),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_1362),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1336),
.B(n_1323),
.Y(n_1458)
);

INVxp67_ASAP7_75t_L g1459 ( 
.A(n_1290),
.Y(n_1459)
);

OAI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1288),
.A2(n_1360),
.B(n_1353),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1319),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1379),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1333),
.A2(n_1349),
.B1(n_1358),
.B2(n_1332),
.Y(n_1463)
);

A2O1A1Ixp33_ASAP7_75t_L g1464 ( 
.A1(n_1339),
.A2(n_1325),
.B(n_1340),
.C(n_1314),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1383),
.Y(n_1465)
);

NAND2x1_ASAP7_75t_L g1466 ( 
.A(n_1384),
.B(n_1386),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1388),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1396),
.Y(n_1468)
);

INVx4_ASAP7_75t_SL g1469 ( 
.A(n_1349),
.Y(n_1469)
);

AO21x2_ASAP7_75t_L g1470 ( 
.A1(n_1366),
.A2(n_1356),
.B(n_1408),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1294),
.B(n_1380),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1398),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1356),
.A2(n_1341),
.B(n_1342),
.Y(n_1473)
);

AOI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1401),
.A2(n_1329),
.B(n_1324),
.Y(n_1474)
);

INVx3_ASAP7_75t_L g1475 ( 
.A(n_1367),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1328),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1331),
.B(n_1348),
.Y(n_1477)
);

OA21x2_ASAP7_75t_L g1478 ( 
.A1(n_1395),
.A2(n_1344),
.B(n_1350),
.Y(n_1478)
);

OA21x2_ASAP7_75t_L g1479 ( 
.A1(n_1412),
.A2(n_1413),
.B(n_1346),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1413),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1413),
.A2(n_1335),
.B(n_1389),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1343),
.B(n_1311),
.Y(n_1482)
);

INVx1_ASAP7_75t_SL g1483 ( 
.A(n_1298),
.Y(n_1483)
);

INVxp67_ASAP7_75t_SL g1484 ( 
.A(n_1390),
.Y(n_1484)
);

INVxp67_ASAP7_75t_L g1485 ( 
.A(n_1309),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1320),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_1312),
.Y(n_1487)
);

NOR2x1_ASAP7_75t_R g1488 ( 
.A(n_1338),
.B(n_1407),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1347),
.A2(n_1293),
.B1(n_1327),
.B2(n_1317),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1343),
.B(n_1314),
.Y(n_1490)
);

OAI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1446),
.A2(n_1387),
.B1(n_1410),
.B2(n_1382),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1472),
.Y(n_1492)
);

AO32x2_ASAP7_75t_L g1493 ( 
.A1(n_1470),
.A2(n_1295),
.A3(n_1391),
.B1(n_1317),
.B2(n_1409),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_1487),
.Y(n_1494)
);

AOI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1427),
.A2(n_1330),
.B1(n_1300),
.B2(n_1299),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1416),
.B(n_1420),
.Y(n_1496)
);

AND2x6_ASAP7_75t_L g1497 ( 
.A(n_1435),
.B(n_1337),
.Y(n_1497)
);

O2A1O1Ixp33_ASAP7_75t_SL g1498 ( 
.A1(n_1460),
.A2(n_1410),
.B(n_1402),
.C(n_1400),
.Y(n_1498)
);

INVx2_ASAP7_75t_SL g1499 ( 
.A(n_1482),
.Y(n_1499)
);

OA21x2_ASAP7_75t_L g1500 ( 
.A1(n_1443),
.A2(n_1415),
.B(n_1445),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1459),
.B(n_1316),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1447),
.B(n_1414),
.Y(n_1502)
);

AOI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1446),
.A2(n_1312),
.B1(n_1303),
.B2(n_1399),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1447),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1448),
.A2(n_1308),
.B1(n_1463),
.B2(n_1453),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1451),
.Y(n_1506)
);

OAI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1423),
.A2(n_1434),
.B(n_1460),
.Y(n_1507)
);

BUFx10_ASAP7_75t_L g1508 ( 
.A(n_1488),
.Y(n_1508)
);

AOI221xp5_ASAP7_75t_L g1509 ( 
.A1(n_1436),
.A2(n_1437),
.B1(n_1431),
.B2(n_1432),
.C(n_1458),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1472),
.Y(n_1510)
);

AO32x2_ASAP7_75t_L g1511 ( 
.A1(n_1470),
.A2(n_1450),
.A3(n_1441),
.B1(n_1449),
.B2(n_1432),
.Y(n_1511)
);

AND2x2_ASAP7_75t_SL g1512 ( 
.A(n_1442),
.B(n_1478),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_SL g1513 ( 
.A(n_1488),
.B(n_1485),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1424),
.A2(n_1429),
.B(n_1432),
.Y(n_1514)
);

O2A1O1Ixp33_ASAP7_75t_L g1515 ( 
.A1(n_1442),
.A2(n_1438),
.B(n_1464),
.C(n_1458),
.Y(n_1515)
);

NAND4xp25_ASAP7_75t_L g1516 ( 
.A(n_1473),
.B(n_1489),
.C(n_1477),
.D(n_1462),
.Y(n_1516)
);

OA21x2_ASAP7_75t_L g1517 ( 
.A1(n_1452),
.A2(n_1422),
.B(n_1473),
.Y(n_1517)
);

AO21x1_ASAP7_75t_L g1518 ( 
.A1(n_1466),
.A2(n_1444),
.B(n_1477),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1476),
.B(n_1471),
.Y(n_1519)
);

INVxp67_ASAP7_75t_L g1520 ( 
.A(n_1478),
.Y(n_1520)
);

A2O1A1Ixp33_ASAP7_75t_L g1521 ( 
.A1(n_1424),
.A2(n_1429),
.B(n_1475),
.C(n_1430),
.Y(n_1521)
);

A2O1A1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1475),
.A2(n_1430),
.B(n_1439),
.C(n_1466),
.Y(n_1522)
);

A2O1A1Ixp33_ASAP7_75t_L g1523 ( 
.A1(n_1475),
.A2(n_1439),
.B(n_1457),
.C(n_1481),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_1487),
.Y(n_1524)
);

OAI211xp5_ASAP7_75t_SL g1525 ( 
.A1(n_1482),
.A2(n_1457),
.B(n_1490),
.C(n_1465),
.Y(n_1525)
);

OAI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1457),
.A2(n_1478),
.B(n_1474),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1476),
.B(n_1471),
.Y(n_1527)
);

AO21x1_ASAP7_75t_L g1528 ( 
.A1(n_1444),
.A2(n_1454),
.B(n_1456),
.Y(n_1528)
);

AOI221xp5_ASAP7_75t_L g1529 ( 
.A1(n_1449),
.A2(n_1475),
.B1(n_1470),
.B2(n_1454),
.C(n_1467),
.Y(n_1529)
);

AOI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1469),
.A2(n_1490),
.B1(n_1449),
.B2(n_1483),
.Y(n_1530)
);

AOI221x1_ASAP7_75t_SL g1531 ( 
.A1(n_1456),
.A2(n_1467),
.B1(n_1462),
.B2(n_1465),
.C(n_1417),
.Y(n_1531)
);

OAI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1474),
.A2(n_1440),
.B(n_1484),
.Y(n_1532)
);

NAND3xp33_ASAP7_75t_SL g1533 ( 
.A(n_1507),
.B(n_1483),
.C(n_1486),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1506),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1509),
.B(n_1455),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1509),
.B(n_1461),
.Y(n_1536)
);

BUFx2_ASAP7_75t_L g1537 ( 
.A(n_1493),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1512),
.B(n_1426),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1512),
.B(n_1425),
.Y(n_1539)
);

OAI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1503),
.A2(n_1418),
.B1(n_1480),
.B2(n_1479),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1505),
.A2(n_1469),
.B1(n_1418),
.B2(n_1421),
.Y(n_1541)
);

INVxp67_ASAP7_75t_L g1542 ( 
.A(n_1519),
.Y(n_1542)
);

NAND2x1p5_ASAP7_75t_SL g1543 ( 
.A(n_1499),
.B(n_1433),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1492),
.Y(n_1544)
);

CKINVDCx14_ASAP7_75t_R g1545 ( 
.A(n_1508),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1531),
.B(n_1510),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1528),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1527),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1520),
.B(n_1468),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1491),
.A2(n_1468),
.B1(n_1461),
.B2(n_1479),
.Y(n_1550)
);

INVx5_ASAP7_75t_L g1551 ( 
.A(n_1497),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1517),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1530),
.B(n_1419),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1517),
.B(n_1422),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1493),
.B(n_1428),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1518),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1532),
.Y(n_1557)
);

NOR2x1_ASAP7_75t_SL g1558 ( 
.A(n_1551),
.B(n_1504),
.Y(n_1558)
);

INVxp67_ASAP7_75t_L g1559 ( 
.A(n_1556),
.Y(n_1559)
);

AO21x2_ASAP7_75t_L g1560 ( 
.A1(n_1547),
.A2(n_1526),
.B(n_1514),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1549),
.Y(n_1561)
);

BUFx2_ASAP7_75t_L g1562 ( 
.A(n_1537),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1535),
.A2(n_1491),
.B1(n_1516),
.B2(n_1529),
.Y(n_1563)
);

AO21x2_ASAP7_75t_L g1564 ( 
.A1(n_1547),
.A2(n_1514),
.B(n_1522),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1542),
.B(n_1557),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1542),
.B(n_1529),
.Y(n_1566)
);

OAI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1533),
.A2(n_1515),
.B(n_1521),
.Y(n_1567)
);

INVx3_ASAP7_75t_L g1568 ( 
.A(n_1552),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1534),
.Y(n_1569)
);

INVx5_ASAP7_75t_L g1570 ( 
.A(n_1551),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1534),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1554),
.Y(n_1572)
);

BUFx3_ASAP7_75t_L g1573 ( 
.A(n_1551),
.Y(n_1573)
);

INVxp67_ASAP7_75t_L g1574 ( 
.A(n_1556),
.Y(n_1574)
);

AOI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1550),
.A2(n_1533),
.B1(n_1541),
.B2(n_1498),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1535),
.A2(n_1515),
.B1(n_1521),
.B2(n_1522),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1557),
.B(n_1500),
.Y(n_1577)
);

INVxp67_ASAP7_75t_L g1578 ( 
.A(n_1546),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1555),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1551),
.B(n_1523),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1555),
.B(n_1511),
.Y(n_1581)
);

BUFx2_ASAP7_75t_L g1582 ( 
.A(n_1543),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1569),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1578),
.B(n_1546),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1568),
.Y(n_1585)
);

BUFx2_ASAP7_75t_L g1586 ( 
.A(n_1573),
.Y(n_1586)
);

BUFx6f_ASAP7_75t_L g1587 ( 
.A(n_1570),
.Y(n_1587)
);

INVxp33_ASAP7_75t_L g1588 ( 
.A(n_1567),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1569),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1562),
.B(n_1553),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1571),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1559),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1562),
.B(n_1538),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1562),
.B(n_1553),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1578),
.B(n_1548),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1565),
.B(n_1548),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1581),
.B(n_1538),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1563),
.A2(n_1536),
.B1(n_1550),
.B2(n_1495),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1581),
.B(n_1539),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1571),
.Y(n_1600)
);

INVx4_ASAP7_75t_L g1601 ( 
.A(n_1570),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1579),
.B(n_1539),
.Y(n_1602)
);

INVx1_ASAP7_75t_SL g1603 ( 
.A(n_1565),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1559),
.B(n_1544),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1563),
.A2(n_1536),
.B1(n_1496),
.B2(n_1525),
.Y(n_1605)
);

BUFx2_ASAP7_75t_L g1606 ( 
.A(n_1573),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1583),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_R g1608 ( 
.A(n_1584),
.B(n_1575),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1586),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1584),
.B(n_1574),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1583),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1603),
.B(n_1574),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1603),
.B(n_1566),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1588),
.B(n_1545),
.Y(n_1614)
);

INVx1_ASAP7_75t_SL g1615 ( 
.A(n_1586),
.Y(n_1615)
);

BUFx2_ASAP7_75t_L g1616 ( 
.A(n_1587),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1586),
.B(n_1582),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1585),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1595),
.B(n_1566),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1601),
.B(n_1558),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1595),
.B(n_1561),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1601),
.B(n_1558),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1606),
.B(n_1582),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1597),
.B(n_1558),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1585),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1597),
.B(n_1580),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1583),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1606),
.B(n_1582),
.Y(n_1628)
);

OAI31xp33_ASAP7_75t_L g1629 ( 
.A1(n_1588),
.A2(n_1576),
.A3(n_1498),
.B(n_1540),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1589),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1585),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1606),
.B(n_1572),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1585),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1590),
.B(n_1577),
.Y(n_1634)
);

INVx2_ASAP7_75t_SL g1635 ( 
.A(n_1587),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1591),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1597),
.B(n_1580),
.Y(n_1637)
);

AOI21xp33_ASAP7_75t_L g1638 ( 
.A1(n_1598),
.A2(n_1576),
.B(n_1567),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_L g1639 ( 
.A(n_1598),
.B(n_1508),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1600),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1600),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1601),
.B(n_1573),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1624),
.B(n_1597),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1632),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1638),
.B(n_1605),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1607),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1638),
.B(n_1605),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1619),
.B(n_1593),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1607),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1611),
.Y(n_1650)
);

INVx2_ASAP7_75t_SL g1651 ( 
.A(n_1635),
.Y(n_1651)
);

NAND2xp67_ASAP7_75t_L g1652 ( 
.A(n_1617),
.B(n_1501),
.Y(n_1652)
);

NOR2x1_ASAP7_75t_L g1653 ( 
.A(n_1616),
.B(n_1601),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1611),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1619),
.B(n_1593),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1627),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1610),
.B(n_1592),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1610),
.B(n_1613),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1613),
.B(n_1590),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1627),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1609),
.B(n_1592),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1635),
.B(n_1601),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1632),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1624),
.B(n_1593),
.Y(n_1664)
);

INVxp67_ASAP7_75t_L g1665 ( 
.A(n_1614),
.Y(n_1665)
);

INVx1_ASAP7_75t_SL g1666 ( 
.A(n_1609),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1632),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1630),
.Y(n_1668)
);

INVx2_ASAP7_75t_SL g1669 ( 
.A(n_1635),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1626),
.B(n_1599),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1626),
.B(n_1599),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1637),
.B(n_1599),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1637),
.B(n_1602),
.Y(n_1673)
);

O2A1O1Ixp5_ASAP7_75t_R g1674 ( 
.A1(n_1608),
.A2(n_1604),
.B(n_1596),
.C(n_1587),
.Y(n_1674)
);

NOR2x1_ASAP7_75t_L g1675 ( 
.A(n_1616),
.B(n_1601),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1615),
.B(n_1590),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1639),
.B(n_1596),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1642),
.B(n_1602),
.Y(n_1678)
);

NAND2xp33_ASAP7_75t_L g1679 ( 
.A(n_1645),
.B(n_1608),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1678),
.B(n_1642),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1651),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1651),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1647),
.A2(n_1575),
.B1(n_1580),
.B2(n_1642),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1669),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1678),
.B(n_1642),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1646),
.Y(n_1686)
);

AND2x4_ASAP7_75t_SL g1687 ( 
.A(n_1662),
.B(n_1587),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1646),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1649),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1649),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1650),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1664),
.B(n_1642),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1650),
.Y(n_1693)
);

AOI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1665),
.A2(n_1580),
.B1(n_1564),
.B2(n_1560),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1669),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1654),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1652),
.B(n_1615),
.Y(n_1697)
);

AOI211x1_ASAP7_75t_L g1698 ( 
.A1(n_1674),
.A2(n_1623),
.B(n_1628),
.C(n_1617),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1652),
.B(n_1658),
.Y(n_1699)
);

O2A1O1Ixp33_ASAP7_75t_L g1700 ( 
.A1(n_1674),
.A2(n_1629),
.B(n_1612),
.C(n_1623),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1654),
.Y(n_1701)
);

AOI22xp33_ASAP7_75t_SL g1702 ( 
.A1(n_1677),
.A2(n_1587),
.B1(n_1629),
.B2(n_1580),
.Y(n_1702)
);

OAI221xp5_ASAP7_75t_L g1703 ( 
.A1(n_1658),
.A2(n_1587),
.B1(n_1612),
.B2(n_1628),
.C(n_1617),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1666),
.A2(n_1594),
.B1(n_1587),
.B2(n_1580),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1686),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1686),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1680),
.B(n_1670),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1680),
.B(n_1685),
.Y(n_1708)
);

AOI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1679),
.A2(n_1702),
.B1(n_1683),
.B2(n_1685),
.Y(n_1709)
);

OAI322xp33_ASAP7_75t_L g1710 ( 
.A1(n_1700),
.A2(n_1699),
.A3(n_1666),
.B1(n_1703),
.B2(n_1697),
.C1(n_1657),
.C2(n_1694),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1687),
.B(n_1653),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1679),
.B(n_1670),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1681),
.B(n_1661),
.Y(n_1713)
);

AOI22x1_ASAP7_75t_SL g1714 ( 
.A1(n_1681),
.A2(n_1682),
.B1(n_1695),
.B2(n_1684),
.Y(n_1714)
);

INVx1_ASAP7_75t_SL g1715 ( 
.A(n_1687),
.Y(n_1715)
);

INVx2_ASAP7_75t_SL g1716 ( 
.A(n_1692),
.Y(n_1716)
);

INVxp67_ASAP7_75t_L g1717 ( 
.A(n_1682),
.Y(n_1717)
);

NOR2x1p5_ASAP7_75t_L g1718 ( 
.A(n_1684),
.B(n_1657),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1688),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1695),
.B(n_1648),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1698),
.B(n_1661),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_L g1722 ( 
.A(n_1692),
.B(n_1513),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1688),
.Y(n_1723)
);

AOI221xp5_ASAP7_75t_L g1724 ( 
.A1(n_1704),
.A2(n_1676),
.B1(n_1655),
.B2(n_1659),
.C(n_1628),
.Y(n_1724)
);

AOI221x1_ASAP7_75t_SL g1725 ( 
.A1(n_1721),
.A2(n_1701),
.B1(n_1696),
.B2(n_1693),
.C(n_1691),
.Y(n_1725)
);

INVx2_ASAP7_75t_SL g1726 ( 
.A(n_1711),
.Y(n_1726)
);

AOI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1716),
.A2(n_1708),
.B1(n_1722),
.B2(n_1714),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1711),
.Y(n_1728)
);

O2A1O1Ixp33_ASAP7_75t_L g1729 ( 
.A1(n_1710),
.A2(n_1690),
.B(n_1689),
.C(n_1676),
.Y(n_1729)
);

AOI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1721),
.A2(n_1675),
.B(n_1653),
.Y(n_1730)
);

INVxp67_ASAP7_75t_L g1731 ( 
.A(n_1712),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1718),
.B(n_1717),
.Y(n_1732)
);

NAND2xp33_ASAP7_75t_SL g1733 ( 
.A(n_1713),
.B(n_1659),
.Y(n_1733)
);

BUFx6f_ASAP7_75t_L g1734 ( 
.A(n_1713),
.Y(n_1734)
);

O2A1O1Ixp33_ASAP7_75t_L g1735 ( 
.A1(n_1715),
.A2(n_1690),
.B(n_1689),
.C(n_1675),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1734),
.Y(n_1736)
);

NOR3xp33_ASAP7_75t_SL g1737 ( 
.A(n_1732),
.B(n_1724),
.C(n_1706),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1726),
.B(n_1728),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1734),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1731),
.B(n_1725),
.Y(n_1740)
);

NAND3xp33_ASAP7_75t_SL g1741 ( 
.A(n_1729),
.B(n_1709),
.C(n_1715),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1733),
.B(n_1720),
.Y(n_1742)
);

NAND3xp33_ASAP7_75t_SL g1743 ( 
.A(n_1727),
.B(n_1707),
.C(n_1705),
.Y(n_1743)
);

NOR3xp33_ASAP7_75t_L g1744 ( 
.A(n_1735),
.B(n_1723),
.C(n_1719),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1730),
.B(n_1644),
.Y(n_1745)
);

NOR3xp33_ASAP7_75t_L g1746 ( 
.A(n_1743),
.B(n_1662),
.C(n_1644),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1738),
.B(n_1671),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1736),
.Y(n_1748)
);

OAI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1737),
.A2(n_1740),
.B1(n_1742),
.B2(n_1739),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1741),
.B(n_1662),
.Y(n_1750)
);

A2O1A1Ixp33_ASAP7_75t_SL g1751 ( 
.A1(n_1750),
.A2(n_1744),
.B(n_1644),
.C(n_1663),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1749),
.B(n_1745),
.Y(n_1752)
);

OAI221xp5_ASAP7_75t_L g1753 ( 
.A1(n_1746),
.A2(n_1747),
.B1(n_1748),
.B2(n_1587),
.C(n_1663),
.Y(n_1753)
);

OAI211xp5_ASAP7_75t_SL g1754 ( 
.A1(n_1749),
.A2(n_1667),
.B(n_1663),
.C(n_1656),
.Y(n_1754)
);

A2O1A1Ixp33_ASAP7_75t_SL g1755 ( 
.A1(n_1750),
.A2(n_1667),
.B(n_1656),
.C(n_1668),
.Y(n_1755)
);

AOI221xp5_ASAP7_75t_L g1756 ( 
.A1(n_1749),
.A2(n_1662),
.B1(n_1667),
.B2(n_1660),
.C(n_1668),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1752),
.Y(n_1757)
);

XNOR2x1_ASAP7_75t_L g1758 ( 
.A(n_1751),
.B(n_1753),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1756),
.B(n_1664),
.Y(n_1759)
);

AOI22xp5_ASAP7_75t_SL g1760 ( 
.A1(n_1755),
.A2(n_1620),
.B1(n_1622),
.B2(n_1623),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1754),
.Y(n_1761)
);

INVx1_ASAP7_75t_SL g1762 ( 
.A(n_1758),
.Y(n_1762)
);

AOI221xp5_ASAP7_75t_L g1763 ( 
.A1(n_1761),
.A2(n_1660),
.B1(n_1620),
.B2(n_1622),
.C(n_1587),
.Y(n_1763)
);

NAND3x1_ASAP7_75t_SL g1764 ( 
.A(n_1760),
.B(n_1643),
.C(n_1673),
.Y(n_1764)
);

AOI221xp5_ASAP7_75t_L g1765 ( 
.A1(n_1762),
.A2(n_1759),
.B1(n_1757),
.B2(n_1620),
.C(n_1622),
.Y(n_1765)
);

OAI22x1_ASAP7_75t_L g1766 ( 
.A1(n_1765),
.A2(n_1764),
.B1(n_1763),
.B2(n_1620),
.Y(n_1766)
);

OA22x2_ASAP7_75t_L g1767 ( 
.A1(n_1766),
.A2(n_1622),
.B1(n_1620),
.B2(n_1643),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1766),
.A2(n_1622),
.B1(n_1673),
.B2(n_1671),
.Y(n_1768)
);

OAI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1768),
.A2(n_1634),
.B1(n_1641),
.B2(n_1640),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1767),
.B(n_1672),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_SL g1771 ( 
.A1(n_1770),
.A2(n_1494),
.B1(n_1524),
.B2(n_1634),
.Y(n_1771)
);

OAI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1769),
.A2(n_1672),
.B(n_1621),
.Y(n_1772)
);

OA21x2_ASAP7_75t_L g1773 ( 
.A1(n_1772),
.A2(n_1625),
.B(n_1618),
.Y(n_1773)
);

OAI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1773),
.A2(n_1771),
.B(n_1621),
.Y(n_1774)
);

OAI22xp33_ASAP7_75t_SL g1775 ( 
.A1(n_1774),
.A2(n_1641),
.B1(n_1640),
.B2(n_1636),
.Y(n_1775)
);

OAI221xp5_ASAP7_75t_R g1776 ( 
.A1(n_1775),
.A2(n_1618),
.B1(n_1625),
.B2(n_1631),
.C(n_1633),
.Y(n_1776)
);

AOI211xp5_ASAP7_75t_L g1777 ( 
.A1(n_1776),
.A2(n_1494),
.B(n_1524),
.C(n_1502),
.Y(n_1777)
);


endmodule