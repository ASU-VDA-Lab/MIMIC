module fake_jpeg_14601_n_84 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_84);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_84;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx5_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx8_ASAP7_75t_SL g11 ( 
.A(n_5),
.Y(n_11)
);

OR2x2_ASAP7_75t_L g12 ( 
.A(n_3),
.B(n_5),
.Y(n_12)
);

BUFx4f_ASAP7_75t_SL g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_2),
.B(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_23),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_12),
.B(n_1),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_1),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_10),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_10),
.B1(n_15),
.B2(n_20),
.Y(n_32)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_28),
.Y(n_39)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_7),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_9),
.Y(n_31)
);

AOI21xp33_ASAP7_75t_L g48 ( 
.A1(n_32),
.A2(n_23),
.B(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_18),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_30),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_14),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_25),
.A2(n_15),
.B1(n_18),
.B2(n_20),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_21),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_44),
.B(n_23),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_48),
.B1(n_41),
.B2(n_14),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_54),
.B(n_55),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_49),
.B(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

AND2x4_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_33),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_30),
.Y(n_55)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_21),
.Y(n_64)
);

AO21x1_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_62),
.B(n_55),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_46),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_39),
.B(n_29),
.C(n_42),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_64),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_61),
.A2(n_54),
.B1(n_52),
.B2(n_55),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_66),
.Y(n_71)
);

XNOR2x1_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_46),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_67),
.A2(n_47),
.B1(n_50),
.B2(n_51),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_69),
.A2(n_62),
.B1(n_63),
.B2(n_56),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_58),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_68),
.C(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_74),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_75),
.A2(n_73),
.B(n_47),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_13),
.C(n_67),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_72),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_76),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_80),
.A2(n_13),
.B(n_51),
.Y(n_82)
);

BUFx24_ASAP7_75t_SL g83 ( 
.A(n_82),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_83),
.B(n_81),
.Y(n_84)
);


endmodule