module fake_jpeg_2907_n_596 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_596);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_596;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_17),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g167 ( 
.A(n_56),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_18),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_57),
.B(n_63),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_25),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_58),
.B(n_74),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_19),
.B(n_18),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_66),
.Y(n_144)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_67),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_68),
.B(n_92),
.Y(n_151)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_69),
.Y(n_149)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_70),
.Y(n_131)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_71),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_72),
.Y(n_168)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_75),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_76),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_25),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_77),
.B(n_90),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_78),
.Y(n_177)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_80),
.Y(n_159)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_81),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_82),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_43),
.Y(n_83)
);

NAND2xp33_ASAP7_75t_SL g190 ( 
.A(n_83),
.B(n_120),
.Y(n_190)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_84),
.Y(n_191)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_85),
.Y(n_189)
);

INVx2_ASAP7_75t_R g86 ( 
.A(n_39),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_86),
.B(n_33),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_88),
.Y(n_163)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_89),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_25),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_91),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_15),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_93),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_43),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_94),
.B(n_109),
.Y(n_162)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_95),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_96),
.Y(n_173)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_97),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_100),
.Y(n_192)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_101),
.Y(n_203)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_31),
.Y(n_102)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_102),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_37),
.B(n_0),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_103),
.B(n_107),
.Y(n_152)
);

BUFx24_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

BUFx2_ASAP7_75t_SL g138 ( 
.A(n_104),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_106),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_54),
.B(n_0),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_29),
.Y(n_108)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_108),
.Y(n_169)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_37),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_53),
.B(n_0),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_110),
.B(n_8),
.Y(n_198)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_111),
.Y(n_158)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_112),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_35),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_113),
.B(n_114),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_35),
.Y(n_114)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_26),
.Y(n_115)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_115),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_44),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_116),
.B(n_117),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_44),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_118),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_44),
.Y(n_119)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

BUFx24_ASAP7_75t_L g120 ( 
.A(n_26),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_29),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_121),
.B(n_123),
.Y(n_220)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_26),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_122),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_47),
.Y(n_123)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_52),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_124),
.Y(n_212)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_125),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_47),
.Y(n_126)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_126),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_47),
.B1(n_52),
.B2(n_36),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_129),
.A2(n_132),
.B1(n_136),
.B2(n_139),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_59),
.A2(n_34),
.B1(n_27),
.B2(n_41),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_L g135 ( 
.A1(n_67),
.A2(n_34),
.B1(n_27),
.B2(n_41),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_135),
.A2(n_175),
.B1(n_196),
.B2(n_202),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_62),
.A2(n_38),
.B1(n_36),
.B2(n_33),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_122),
.A2(n_55),
.B1(n_46),
.B2(n_38),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_143),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_125),
.A2(n_64),
.B1(n_79),
.B2(n_84),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_147),
.B(n_133),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_73),
.A2(n_55),
.B1(n_46),
.B2(n_32),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_150),
.A2(n_172),
.B1(n_182),
.B2(n_187),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_74),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_156),
.B(n_204),
.Y(n_223)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_86),
.A2(n_32),
.B(n_23),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_157),
.B(n_216),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_106),
.A2(n_55),
.B1(n_23),
.B2(n_2),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_99),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_118),
.B(n_1),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_179),
.B(n_186),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_75),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_65),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_184),
.A2(n_206),
.B1(n_182),
.B2(n_187),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_111),
.B(n_4),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_89),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_112),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_188),
.A2(n_218),
.B1(n_138),
.B2(n_201),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_66),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_93),
.Y(n_197)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_198),
.B(n_214),
.Y(n_278)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_100),
.Y(n_199)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_199),
.Y(n_242)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_60),
.Y(n_200)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_200),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_72),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_76),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_78),
.A2(n_9),
.B1(n_13),
.B2(n_15),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_104),
.B(n_70),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_208),
.B(n_217),
.Y(n_284)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_82),
.Y(n_209)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_209),
.Y(n_254)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_126),
.Y(n_211)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_211),
.Y(n_258)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_87),
.Y(n_213)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_213),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_105),
.B(n_13),
.Y(n_214)
);

OAI21xp33_ASAP7_75t_L g216 ( 
.A1(n_120),
.A2(n_13),
.B(n_104),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_88),
.B(n_98),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_108),
.A2(n_69),
.B1(n_80),
.B2(n_85),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_91),
.Y(n_219)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_219),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_115),
.B(n_96),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_119),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_212),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_222),
.Y(n_352)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_174),
.Y(n_224)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_224),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_162),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_225),
.B(n_240),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_226),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_142),
.B(n_124),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_227),
.B(n_237),
.Y(n_306)
);

INVx3_ASAP7_75t_SL g228 ( 
.A(n_181),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_228),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_128),
.Y(n_233)
);

INVx8_ASAP7_75t_L g312 ( 
.A(n_233),
.Y(n_312)
);

INVxp33_ASAP7_75t_L g234 ( 
.A(n_190),
.Y(n_234)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_234),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_157),
.A2(n_135),
.B1(n_136),
.B2(n_132),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_235),
.A2(n_260),
.B1(n_274),
.B2(n_231),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_210),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_236),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_176),
.B(n_56),
.Y(n_237)
);

AND2x2_ASAP7_75t_SL g238 ( 
.A(n_179),
.B(n_120),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_238),
.Y(n_324)
);

OAI32xp33_ASAP7_75t_L g239 ( 
.A1(n_152),
.A2(n_56),
.A3(n_151),
.B1(n_143),
.B2(n_153),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_239),
.A2(n_234),
.B(n_230),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_208),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_149),
.Y(n_241)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_241),
.Y(n_357)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_128),
.Y(n_243)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_243),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_244),
.A2(n_253),
.B1(n_271),
.B2(n_229),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_180),
.B(n_203),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_245),
.B(n_249),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_183),
.B(n_215),
.C(n_127),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_247),
.B(n_276),
.C(n_238),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_141),
.B(n_216),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_248),
.B(n_261),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_195),
.B(n_220),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_205),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_250),
.B(n_256),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_166),
.A2(n_169),
.B1(n_185),
.B2(n_171),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_251),
.B(n_295),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_184),
.A2(n_206),
.B1(n_139),
.B2(n_150),
.Y(n_253)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_134),
.Y(n_255)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_255),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_155),
.B(n_130),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_159),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_257),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_158),
.B(n_154),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_145),
.B(n_178),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_262),
.B(n_277),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_131),
.B(n_191),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_263),
.B(n_274),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_161),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_264),
.B(n_265),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_159),
.Y(n_265)
);

INVx8_ASAP7_75t_L g266 ( 
.A(n_134),
.Y(n_266)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_266),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_189),
.Y(n_267)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_267),
.Y(n_356)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_149),
.Y(n_268)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_268),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_131),
.B(n_192),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_269),
.B(n_281),
.Y(n_332)
);

OA22x2_ASAP7_75t_L g318 ( 
.A1(n_270),
.A2(n_246),
.B1(n_251),
.B2(n_241),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_194),
.A2(n_188),
.B1(n_218),
.B2(n_164),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_137),
.Y(n_272)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_272),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_137),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_273),
.A2(n_298),
.B1(n_300),
.B2(n_302),
.Y(n_320)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_191),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_275),
.B(n_286),
.Y(n_341)
);

AND2x2_ASAP7_75t_SL g276 ( 
.A(n_165),
.B(n_192),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_164),
.B(n_207),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_148),
.B(n_163),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_279),
.B(n_290),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_189),
.Y(n_280)
);

INVx13_ASAP7_75t_L g340 ( 
.A(n_280),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_167),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_165),
.B(n_160),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_282),
.B(n_283),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_167),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_140),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_285),
.B(n_291),
.Y(n_347)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_146),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_172),
.A2(n_163),
.B1(n_148),
.B2(n_193),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_287),
.A2(n_272),
.B1(n_298),
.B2(n_257),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_193),
.B(n_170),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_171),
.B(n_133),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_167),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_292),
.B(n_294),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_146),
.B(n_173),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_293),
.B(n_297),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_173),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_144),
.B(n_168),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_144),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_296),
.B(n_299),
.Y(n_338)
);

BUFx4f_ASAP7_75t_SL g297 ( 
.A(n_168),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_170),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_181),
.B(n_177),
.Y(n_299)
);

INVx8_ASAP7_75t_L g300 ( 
.A(n_177),
.Y(n_300)
);

INVx6_ASAP7_75t_L g301 ( 
.A(n_128),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_301),
.B(n_273),
.Y(n_339)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_145),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_304),
.B(n_316),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_259),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_308),
.B(n_313),
.C(n_328),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_310),
.A2(n_343),
.B1(n_349),
.B2(n_358),
.Y(n_363)
);

MAJx2_ASAP7_75t_L g313 ( 
.A(n_259),
.B(n_278),
.C(n_238),
.Y(n_313)
);

OAI32xp33_ASAP7_75t_L g316 ( 
.A1(n_248),
.A2(n_239),
.A3(n_278),
.B1(n_229),
.B2(n_261),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_317),
.B(n_313),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_318),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_321),
.A2(n_322),
.B1(n_326),
.B2(n_348),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_260),
.A2(n_296),
.B1(n_253),
.B2(n_279),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_244),
.A2(n_271),
.B1(n_287),
.B2(n_229),
.Y(n_326)
);

A2O1A1O1Ixp25_ASAP7_75t_L g327 ( 
.A1(n_277),
.A2(n_247),
.B(n_225),
.C(n_250),
.D(n_262),
.Y(n_327)
);

NOR3xp33_ASAP7_75t_L g396 ( 
.A(n_327),
.B(n_324),
.C(n_304),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_224),
.B(n_223),
.C(n_276),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_276),
.B(n_263),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_336),
.B(n_222),
.C(n_324),
.Y(n_378)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_339),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_290),
.A2(n_282),
.B1(n_285),
.B2(n_264),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_265),
.A2(n_293),
.B1(n_263),
.B2(n_280),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_346),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_254),
.A2(n_289),
.B1(n_288),
.B2(n_258),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_302),
.A2(n_289),
.B1(n_288),
.B2(n_258),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_254),
.B(n_252),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_350),
.B(n_275),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_293),
.A2(n_228),
.B1(n_297),
.B2(n_266),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_353),
.A2(n_354),
.B1(n_236),
.B2(n_267),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_228),
.A2(n_297),
.B1(n_300),
.B2(n_233),
.Y(n_354)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_357),
.Y(n_360)
);

INVx3_ASAP7_75t_SL g426 ( 
.A(n_360),
.Y(n_426)
);

INVx8_ASAP7_75t_L g364 ( 
.A(n_305),
.Y(n_364)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_364),
.Y(n_415)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_365),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_350),
.Y(n_367)
);

CKINVDCx14_ASAP7_75t_R g436 ( 
.A(n_367),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_368),
.B(n_376),
.Y(n_420)
);

OR2x2_ASAP7_75t_L g369 ( 
.A(n_307),
.B(n_286),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_369),
.A2(n_399),
.B(n_402),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_317),
.A2(n_232),
.B(n_242),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_371),
.A2(n_315),
.B(n_320),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_326),
.A2(n_252),
.B1(n_232),
.B2(n_242),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_373),
.A2(n_400),
.B1(n_353),
.B2(n_348),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_321),
.A2(n_243),
.B1(n_255),
.B2(n_301),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_374),
.A2(n_349),
.B1(n_337),
.B2(n_345),
.Y(n_417)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_303),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_375),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_319),
.B(n_268),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_325),
.B(n_294),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_377),
.B(n_380),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_378),
.B(n_401),
.C(n_315),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_308),
.B(n_306),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_303),
.Y(n_381)
);

INVx2_ASAP7_75t_SL g435 ( 
.A(n_381),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_319),
.B(n_325),
.Y(n_382)
);

OAI21xp33_ASAP7_75t_L g416 ( 
.A1(n_382),
.A2(n_385),
.B(n_388),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_330),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_383),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_329),
.B(n_314),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_384),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_342),
.B(n_316),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_341),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_386),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_329),
.B(n_311),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_387),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_351),
.B(n_334),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_342),
.B(n_327),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_389),
.B(n_390),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_338),
.B(n_343),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_391),
.B(n_403),
.Y(n_414)
);

BUFx16f_ASAP7_75t_L g392 ( 
.A(n_340),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_392),
.Y(n_430)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_341),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_393),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_341),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_394),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g395 ( 
.A(n_335),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_395),
.Y(n_409)
);

A2O1A1Ixp33_ASAP7_75t_L g432 ( 
.A1(n_396),
.A2(n_312),
.B(n_389),
.C(n_401),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_328),
.B(n_338),
.Y(n_397)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_397),
.B(n_398),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_336),
.B(n_347),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_332),
.B(n_309),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_333),
.A2(n_309),
.B1(n_358),
.B2(n_307),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_309),
.B(n_333),
.C(n_344),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_344),
.A2(n_318),
.B(n_355),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_339),
.B(n_344),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_404),
.B(n_438),
.Y(n_471)
);

AO21x1_ASAP7_75t_SL g405 ( 
.A1(n_391),
.A2(n_318),
.B(n_354),
.Y(n_405)
);

A2O1A1Ixp33_ASAP7_75t_SL g467 ( 
.A1(n_405),
.A2(n_418),
.B(n_364),
.C(n_437),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_410),
.A2(n_369),
.B(n_368),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_362),
.A2(n_318),
.B1(n_345),
.B2(n_337),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_413),
.A2(n_417),
.B1(n_421),
.B2(n_440),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_385),
.A2(n_359),
.B(n_356),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_379),
.A2(n_323),
.B1(n_357),
.B2(n_359),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_422),
.B(n_425),
.C(n_427),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_366),
.B(n_323),
.C(n_356),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_366),
.B(n_370),
.C(n_390),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_362),
.A2(n_312),
.B1(n_331),
.B2(n_352),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_428),
.B(n_437),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_366),
.B(n_352),
.C(n_340),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_431),
.B(n_378),
.C(n_372),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_432),
.B(n_371),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_363),
.A2(n_382),
.B1(n_367),
.B2(n_400),
.Y(n_437)
);

AO22x1_ASAP7_75t_SL g438 ( 
.A1(n_379),
.A2(n_374),
.B1(n_361),
.B2(n_363),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_438),
.B(n_365),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_361),
.A2(n_376),
.B1(n_377),
.B2(n_402),
.Y(n_440)
);

OAI21xp33_ASAP7_75t_L g477 ( 
.A1(n_441),
.A2(n_465),
.B(n_466),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_408),
.B(n_370),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_442),
.B(n_451),
.Y(n_475)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_435),
.Y(n_443)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_443),
.Y(n_476)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_435),
.Y(n_444)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_444),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_436),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_445),
.B(n_456),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_429),
.A2(n_440),
.B1(n_436),
.B2(n_438),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_446),
.A2(n_453),
.B1(n_413),
.B2(n_434),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_431),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_447),
.B(n_452),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_407),
.B(n_388),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_448),
.B(n_449),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_407),
.B(n_383),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_408),
.B(n_397),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_435),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_429),
.A2(n_373),
.B1(n_398),
.B2(n_372),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_455),
.B(n_458),
.C(n_462),
.Y(n_488)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_420),
.Y(n_456)
);

AOI322xp5_ASAP7_75t_L g457 ( 
.A1(n_416),
.A2(n_380),
.A3(n_403),
.B1(n_394),
.B2(n_399),
.C1(n_393),
.C2(n_386),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_457),
.A2(n_464),
.B(n_409),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_427),
.B(n_381),
.C(n_375),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_423),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_459),
.B(n_467),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_460),
.A2(n_470),
.B1(n_471),
.B2(n_434),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_461),
.A2(n_433),
.B(n_405),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_422),
.B(n_369),
.C(n_360),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_414),
.B(n_392),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_463),
.B(n_410),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_406),
.A2(n_395),
.B(n_392),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_411),
.B(n_395),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_439),
.B(n_364),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_419),
.B(n_424),
.Y(n_468)
);

OAI21xp33_ASAP7_75t_L g499 ( 
.A1(n_468),
.A2(n_453),
.B(n_474),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_426),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_469),
.Y(n_479)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_423),
.Y(n_470)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_415),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_472),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_425),
.B(n_419),
.C(n_432),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_474),
.B(n_406),
.C(n_418),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_442),
.B(n_419),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_478),
.B(n_483),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_482),
.B(n_467),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_451),
.B(n_424),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_454),
.B(n_414),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_485),
.B(n_493),
.Y(n_511)
);

INVx3_ASAP7_75t_SL g487 ( 
.A(n_471),
.Y(n_487)
);

INVx13_ASAP7_75t_L g524 ( 
.A(n_487),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_489),
.B(n_464),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_454),
.B(n_418),
.C(n_412),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_490),
.B(n_497),
.C(n_447),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_469),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_492),
.B(n_498),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_458),
.B(n_420),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_494),
.A2(n_467),
.B1(n_443),
.B2(n_444),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_495),
.B(n_504),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_496),
.A2(n_461),
.B(n_450),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_462),
.B(n_433),
.C(n_438),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_446),
.Y(n_498)
);

CKINVDCx14_ASAP7_75t_R g505 ( 
.A(n_499),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_471),
.A2(n_421),
.B1(n_417),
.B2(n_404),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_500),
.A2(n_501),
.B1(n_473),
.B2(n_450),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_460),
.A2(n_428),
.B1(n_415),
.B2(n_409),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_502),
.B(n_467),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_463),
.B(n_455),
.Y(n_504)
);

CKINVDCx16_ASAP7_75t_R g506 ( 
.A(n_491),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_506),
.B(n_516),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_507),
.B(n_509),
.C(n_514),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_484),
.B(n_430),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_508),
.B(n_525),
.Y(n_538)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_512),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_481),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_513),
.A2(n_519),
.B1(n_523),
.B2(n_528),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_475),
.B(n_470),
.C(n_459),
.Y(n_514)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_515),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_475),
.B(n_485),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_518),
.A2(n_520),
.B1(n_503),
.B2(n_487),
.Y(n_541)
);

INVx5_ASAP7_75t_L g519 ( 
.A(n_477),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_500),
.A2(n_467),
.B1(n_452),
.B2(n_426),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_521),
.B(n_526),
.Y(n_532)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_522),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_486),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_488),
.B(n_430),
.C(n_426),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_488),
.B(n_504),
.C(n_490),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_486),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_523),
.B(n_479),
.Y(n_530)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_530),
.Y(n_562)
);

INVx13_ASAP7_75t_L g533 ( 
.A(n_524),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_SL g557 ( 
.A(n_533),
.B(n_536),
.Y(n_557)
);

NOR3xp33_ASAP7_75t_SL g536 ( 
.A(n_519),
.B(n_503),
.C(n_502),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_517),
.B(n_476),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_539),
.B(n_540),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_525),
.B(n_476),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_541),
.A2(n_547),
.B1(n_494),
.B2(n_515),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_505),
.B(n_497),
.Y(n_542)
);

OA21x2_ASAP7_75t_SL g558 ( 
.A1(n_542),
.A2(n_545),
.B(n_480),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_513),
.A2(n_496),
.B1(n_480),
.B2(n_512),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_543),
.B(n_546),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_507),
.B(n_483),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_522),
.Y(n_546)
);

FAx1_ASAP7_75t_SL g547 ( 
.A(n_518),
.B(n_489),
.CI(n_478),
.CON(n_547),
.SN(n_547)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_537),
.B(n_526),
.C(n_511),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_548),
.B(n_549),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_537),
.B(n_511),
.C(n_516),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_L g550 ( 
.A1(n_529),
.A2(n_522),
.B(n_520),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_L g563 ( 
.A1(n_550),
.A2(n_541),
.B(n_544),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_545),
.B(n_514),
.C(n_510),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_553),
.B(n_555),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_542),
.B(n_527),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_554),
.B(n_561),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_540),
.B(n_510),
.C(n_509),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_556),
.B(n_559),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g567 ( 
.A(n_558),
.B(n_560),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_531),
.B(n_493),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_532),
.B(n_501),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_532),
.B(n_527),
.C(n_495),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_563),
.B(n_524),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_548),
.B(n_538),
.C(n_535),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_566),
.B(n_569),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_549),
.B(n_538),
.C(n_535),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_557),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_570),
.B(n_551),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_562),
.A2(n_534),
.B1(n_546),
.B2(n_544),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_571),
.A2(n_550),
.B1(n_562),
.B2(n_555),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_557),
.B(n_539),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_SL g582 ( 
.A(n_573),
.B(n_574),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_556),
.B(n_529),
.C(n_530),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g575 ( 
.A1(n_574),
.A2(n_553),
.B(n_552),
.Y(n_575)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_575),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_576),
.B(n_579),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_567),
.A2(n_551),
.B1(n_558),
.B2(n_554),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g587 ( 
.A(n_577),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_580),
.B(n_581),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_564),
.B(n_561),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_582),
.B(n_572),
.Y(n_583)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_583),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_584),
.B(n_578),
.C(n_569),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_588),
.B(n_589),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_SL g589 ( 
.A(n_586),
.B(n_566),
.Y(n_589)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_590),
.A2(n_587),
.B(n_565),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_L g593 ( 
.A1(n_591),
.A2(n_587),
.B(n_585),
.Y(n_593)
);

O2A1O1Ixp33_ASAP7_75t_SL g594 ( 
.A1(n_593),
.A2(n_592),
.B(n_577),
.C(n_533),
.Y(n_594)
);

AOI322xp5_ASAP7_75t_L g595 ( 
.A1(n_594),
.A2(n_533),
.A3(n_563),
.B1(n_536),
.B2(n_571),
.C1(n_568),
.C2(n_580),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g596 ( 
.A(n_595),
.B(n_576),
.Y(n_596)
);


endmodule