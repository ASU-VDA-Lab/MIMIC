module fake_jpeg_2916_n_71 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_71);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_71;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_21),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_30),
.B(n_25),
.C(n_26),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_26),
.Y(n_31)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_35),
.B(n_38),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_25),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_29),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_20),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_17),
.C(n_15),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_37),
.B1(n_2),
.B2(n_3),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_50),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_37),
.B(n_2),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_42),
.B(n_5),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_6),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_49),
.B1(n_46),
.B2(n_52),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_14),
.C(n_5),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_55),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_1),
.C(n_6),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_56),
.Y(n_63)
);

BUFx24_ASAP7_75t_SL g62 ( 
.A(n_58),
.Y(n_62)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_61),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_57),
.C(n_8),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_65),
.A2(n_60),
.B1(n_57),
.B2(n_63),
.Y(n_66)
);

AOI31xp67_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_64),
.A3(n_8),
.B(n_9),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_67),
.A2(n_7),
.B(n_10),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

OAI321xp33_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_7),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C(n_64),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_11),
.Y(n_71)
);


endmodule