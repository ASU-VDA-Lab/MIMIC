module real_aes_15807_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_635;
wire n_287;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_856;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_478;
wire n_356;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_875;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_880;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_891;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_899;
wire n_526;
wire n_637;
wire n_155;
wire n_653;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_0), .Y(n_218) );
AND2x4_ASAP7_75t_L g896 ( .A(n_1), .B(n_897), .Y(n_896) );
BUFx3_ASAP7_75t_L g149 ( .A(n_2), .Y(n_149) );
INVx1_ASAP7_75t_L g897 ( .A(n_3), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_4), .B(n_859), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_5), .B(n_158), .Y(n_157) );
OR2x2_ASAP7_75t_L g115 ( .A(n_6), .B(n_22), .Y(n_115) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_7), .Y(n_139) );
AOI22xp5_ASAP7_75t_L g853 ( .A1(n_8), .A2(n_53), .B1(n_854), .B2(n_855), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_8), .Y(n_854) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_9), .B(n_138), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_10), .B(n_138), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_11), .B(n_186), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_12), .A2(n_82), .B1(n_138), .B2(n_140), .Y(n_237) );
OAI21x1_ASAP7_75t_L g131 ( .A1(n_13), .A2(n_36), .B(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_14), .B(n_579), .Y(n_578) );
OAI21xp5_ASAP7_75t_L g871 ( .A1(n_15), .A2(n_872), .B(n_883), .Y(n_871) );
INVx1_ASAP7_75t_L g886 ( .A(n_15), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_16), .B(n_176), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_17), .Y(n_601) );
AO32x2_ASAP7_75t_L g234 ( .A1(n_18), .A2(n_129), .A3(n_130), .B1(n_235), .B2(n_238), .Y(n_234) );
AO32x1_ASAP7_75t_L g256 ( .A1(n_18), .A2(n_129), .A3(n_130), .B1(n_235), .B2(n_238), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_19), .B(n_564), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_20), .B(n_129), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_21), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_23), .A2(n_43), .B1(n_145), .B2(n_176), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g236 ( .A1(n_24), .A2(n_90), .B1(n_140), .B2(n_146), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_25), .B(n_160), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g604 ( .A(n_26), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_27), .B(n_193), .Y(n_247) );
OAI22xp5_ASAP7_75t_L g874 ( .A1(n_28), .A2(n_62), .B1(n_875), .B2(n_876), .Y(n_874) );
INVx1_ASAP7_75t_L g876 ( .A(n_28), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_29), .A2(n_64), .B1(n_146), .B2(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_30), .B(n_138), .Y(n_553) );
INVx2_ASAP7_75t_L g110 ( .A(n_31), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_32), .B(n_142), .Y(n_574) );
BUFx3_ASAP7_75t_L g113 ( .A(n_33), .Y(n_113) );
INVx1_ASAP7_75t_L g882 ( .A(n_33), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_34), .B(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_35), .B(n_531), .Y(n_580) );
AND2x2_ASAP7_75t_L g606 ( .A(n_37), .B(n_531), .Y(n_606) );
CKINVDCx5p33_ASAP7_75t_R g889 ( .A(n_38), .Y(n_889) );
CKINVDCx5p33_ASAP7_75t_R g213 ( .A(n_39), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_40), .B(n_192), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_41), .B(n_564), .Y(n_632) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_42), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_44), .B(n_543), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_45), .A2(n_77), .B1(n_192), .B2(n_193), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_46), .B(n_227), .Y(n_635) );
A2O1A1Ixp33_ASAP7_75t_L g599 ( .A1(n_47), .A2(n_177), .B(n_216), .C(n_600), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g137 ( .A1(n_48), .A2(n_79), .B1(n_138), .B2(n_140), .Y(n_137) );
INVx1_ASAP7_75t_L g132 ( .A(n_49), .Y(n_132) );
AND2x4_ASAP7_75t_L g134 ( .A(n_50), .B(n_135), .Y(n_134) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_51), .A2(n_52), .B1(n_145), .B2(n_146), .Y(n_566) );
INVxp67_ASAP7_75t_SL g855 ( .A(n_53), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_54), .B(n_129), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_55), .B(n_531), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g605 ( .A(n_56), .Y(n_605) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_57), .B(n_146), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_58), .B(n_140), .Y(n_156) );
INVx1_ASAP7_75t_L g135 ( .A(n_59), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_60), .B(n_129), .Y(n_165) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_61), .A2(n_216), .B(n_217), .C(n_219), .Y(n_215) );
INVx1_ASAP7_75t_SL g875 ( .A(n_62), .Y(n_875) );
NAND3xp33_ASAP7_75t_L g164 ( .A(n_63), .B(n_140), .C(n_162), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_65), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_66), .B(n_129), .Y(n_557) );
AND2x2_ASAP7_75t_L g221 ( .A(n_67), .B(n_222), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_68), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_69), .B(n_512), .Y(n_631) );
NAND3xp33_ASAP7_75t_L g575 ( .A(n_70), .B(n_142), .C(n_176), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_71), .A2(n_94), .B1(n_138), .B2(n_192), .Y(n_196) );
INVx2_ASAP7_75t_L g143 ( .A(n_72), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_73), .B(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_74), .B(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_75), .B(n_195), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_76), .B(n_138), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_78), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_80), .B(n_180), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_81), .A2(n_89), .B1(n_563), .B2(n_564), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_83), .B(n_138), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_84), .B(n_162), .Y(n_161) );
NAND2xp33_ASAP7_75t_SL g529 ( .A(n_85), .B(n_158), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_86), .B(n_174), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g144 ( .A1(n_87), .A2(n_101), .B1(n_145), .B2(n_146), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_88), .B(n_193), .Y(n_244) );
INVx1_ASAP7_75t_L g497 ( .A(n_91), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g880 ( .A(n_91), .B(n_881), .Y(n_880) );
OAI22x1_ASAP7_75t_L g851 ( .A1(n_92), .A2(n_852), .B1(n_853), .B2(n_856), .Y(n_851) );
INVx1_ASAP7_75t_L g856 ( .A(n_92), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_93), .B(n_186), .Y(n_250) );
NAND2xp33_ASAP7_75t_L g513 ( .A(n_95), .B(n_158), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_96), .B(n_531), .Y(n_636) );
NAND3xp33_ASAP7_75t_L g526 ( .A(n_97), .B(n_158), .C(n_195), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_98), .B(n_512), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_99), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g634 ( .A(n_100), .B(n_564), .Y(n_634) );
O2A1O1Ixp33_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_866), .B(n_891), .C(n_899), .Y(n_102) );
NAND2xp33_ASAP7_75t_L g103 ( .A(n_104), .B(n_858), .Y(n_103) );
INVxp33_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
NOR2xp67_ASAP7_75t_L g105 ( .A(n_106), .B(n_116), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
BUFx12f_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x6_ASAP7_75t_SL g108 ( .A(n_109), .B(n_111), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g862 ( .A(n_110), .B(n_863), .Y(n_862) );
INVx3_ASAP7_75t_L g870 ( .A(n_110), .Y(n_870) );
NOR2xp33_ASAP7_75t_L g912 ( .A(n_110), .B(n_890), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_114), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
NOR2x1_ASAP7_75t_L g865 ( .A(n_113), .B(n_115), .Y(n_865) );
AND2x6_ASAP7_75t_SL g879 ( .A(n_114), .B(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OAI21xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_851), .B(n_857), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NAND2xp33_ASAP7_75t_SL g857 ( .A(n_118), .B(n_851), .Y(n_857) );
OAI22x1_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_493), .B1(n_498), .B2(n_849), .Y(n_118) );
XOR2xp5_ASAP7_75t_L g873 ( .A(n_119), .B(n_874), .Y(n_873) );
AND2x4_ASAP7_75t_L g119 ( .A(n_120), .B(n_394), .Y(n_119) );
AND4x1_ASAP7_75t_L g120 ( .A(n_121), .B(n_316), .C(n_349), .D(n_380), .Y(n_120) );
NOR2xp33_ASAP7_75t_L g121 ( .A(n_122), .B(n_283), .Y(n_121) );
OAI221xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_202), .B1(n_251), .B2(n_261), .C(n_270), .Y(n_122) );
AOI21xp33_ASAP7_75t_L g388 ( .A1(n_123), .A2(n_373), .B(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_166), .Y(n_124) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_150), .Y(n_125) );
INVx2_ASAP7_75t_L g269 ( .A(n_126), .Y(n_269) );
AND2x2_ASAP7_75t_L g279 ( .A(n_126), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g315 ( .A(n_126), .B(n_188), .Y(n_315) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g304 ( .A(n_127), .Y(n_304) );
AOI31xp67_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_133), .A3(n_136), .B(n_147), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx4_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_130), .B(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g169 ( .A(n_130), .Y(n_169) );
BUFx3_ASAP7_75t_L g189 ( .A(n_130), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_130), .B(n_231), .Y(n_230) );
INVx2_ASAP7_75t_SL g241 ( .A(n_130), .Y(n_241) );
AND2x4_ASAP7_75t_SL g518 ( .A(n_130), .B(n_133), .Y(n_518) );
INVx1_ASAP7_75t_SL g522 ( .A(n_130), .Y(n_522) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g153 ( .A(n_131), .Y(n_153) );
OAI21x1_ASAP7_75t_L g154 ( .A1(n_133), .A2(n_155), .B(n_159), .Y(n_154) );
OAI21x1_ASAP7_75t_L g170 ( .A1(n_133), .A2(n_171), .B(n_178), .Y(n_170) );
OAI21x1_ASAP7_75t_L g523 ( .A1(n_133), .A2(n_524), .B(n_527), .Y(n_523) );
OAI21x1_ASAP7_75t_L g536 ( .A1(n_133), .A2(n_537), .B(n_540), .Y(n_536) );
OAI21x1_ASAP7_75t_L g550 ( .A1(n_133), .A2(n_551), .B(n_554), .Y(n_550) );
OAI21x1_ASAP7_75t_L g572 ( .A1(n_133), .A2(n_573), .B(n_576), .Y(n_572) );
OAI21x1_ASAP7_75t_L g629 ( .A1(n_133), .A2(n_630), .B(n_633), .Y(n_629) );
BUFx10_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g198 ( .A(n_134), .Y(n_198) );
INVx1_ASAP7_75t_L g220 ( .A(n_134), .Y(n_220) );
AO31x2_ASAP7_75t_L g224 ( .A1(n_134), .A2(n_189), .A3(n_225), .B(n_230), .Y(n_224) );
BUFx10_ASAP7_75t_L g568 ( .A(n_134), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_141), .B1(n_142), .B2(n_144), .Y(n_136) );
INVx3_ASAP7_75t_L g249 ( .A(n_138), .Y(n_249) );
OAI21xp5_ASAP7_75t_L g524 ( .A1(n_138), .A2(n_525), .B(n_526), .Y(n_524) );
INVx1_ASAP7_75t_L g579 ( .A(n_138), .Y(n_579) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g140 ( .A(n_139), .Y(n_140) );
INVx1_ASAP7_75t_L g145 ( .A(n_139), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_139), .Y(n_146) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_139), .Y(n_158) );
INVx1_ASAP7_75t_L g174 ( .A(n_139), .Y(n_174) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_139), .Y(n_176) );
INVx1_ASAP7_75t_L g192 ( .A(n_139), .Y(n_192) );
INVx1_ASAP7_75t_L g216 ( .A(n_139), .Y(n_216) );
INVx3_ASAP7_75t_L g512 ( .A(n_139), .Y(n_512) );
INVx1_ASAP7_75t_L g565 ( .A(n_139), .Y(n_565) );
INVx2_ASAP7_75t_SL g193 ( .A(n_140), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_140), .B(n_601), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g190 ( .A1(n_141), .A2(n_191), .B1(n_194), .B2(n_196), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_141), .A2(n_226), .B1(n_228), .B2(n_229), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_141), .A2(n_247), .B(n_248), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_141), .A2(n_562), .B1(n_566), .B2(n_567), .Y(n_561) );
INVx6_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_142), .A2(n_156), .B(n_157), .Y(n_155) );
OAI22xp5_ASAP7_75t_L g235 ( .A1(n_142), .A2(n_177), .B1(n_236), .B2(n_237), .Y(n_235) );
O2A1O1Ixp5_ASAP7_75t_L g537 ( .A1(n_142), .A2(n_173), .B(n_538), .C(n_539), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_142), .A2(n_555), .B(n_556), .Y(n_554) );
BUFx8_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g163 ( .A(n_143), .Y(n_163) );
INVx2_ASAP7_75t_L g182 ( .A(n_143), .Y(n_182) );
INVx1_ASAP7_75t_L g195 ( .A(n_143), .Y(n_195) );
INVx1_ASAP7_75t_L g183 ( .A(n_145), .Y(n_183) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_145), .A2(n_176), .B1(n_212), .B2(n_213), .Y(n_211) );
INVx2_ASAP7_75t_L g160 ( .A(n_146), .Y(n_160) );
INVx2_ASAP7_75t_L g563 ( .A(n_146), .Y(n_563) );
OAI21xp5_ASAP7_75t_L g573 ( .A1(n_146), .A2(n_574), .B(n_575), .Y(n_573) );
OAI22xp33_ASAP7_75t_L g603 ( .A1(n_146), .A2(n_512), .B1(n_604), .B2(n_605), .Y(n_603) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g290 ( .A(n_150), .B(n_280), .Y(n_290) );
OR2x2_ASAP7_75t_L g399 ( .A(n_150), .B(n_168), .Y(n_399) );
OAI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_154), .B(n_165), .Y(n_150) );
OAI21x1_ASAP7_75t_L g268 ( .A1(n_151), .A2(n_154), .B(n_165), .Y(n_268) );
OAI21x1_ASAP7_75t_L g535 ( .A1(n_151), .A2(n_536), .B(n_544), .Y(n_535) );
OAI21xp5_ASAP7_75t_L g617 ( .A1(n_151), .A2(n_536), .B(n_544), .Y(n_617) );
OAI21x1_ASAP7_75t_L g628 ( .A1(n_151), .A2(n_629), .B(n_636), .Y(n_628) );
OAI21xp33_ASAP7_75t_SL g654 ( .A1(n_151), .A2(n_629), .B(n_636), .Y(n_654) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g531 ( .A(n_152), .Y(n_531) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g187 ( .A(n_153), .Y(n_187) );
INVx2_ASAP7_75t_L g201 ( .A(n_153), .Y(n_201) );
INVx2_ASAP7_75t_L g543 ( .A(n_158), .Y(n_543) );
OAI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_164), .Y(n_159) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
BUFx4f_ASAP7_75t_L g177 ( .A(n_163), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_166), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
OR2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_188), .Y(n_167) );
INVx1_ASAP7_75t_L g264 ( .A(n_168), .Y(n_264) );
INVx2_ASAP7_75t_SL g341 ( .A(n_168), .Y(n_341) );
BUFx2_ASAP7_75t_L g371 ( .A(n_168), .Y(n_371) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_185), .Y(n_168) );
OA21x2_ASAP7_75t_L g280 ( .A1(n_169), .A2(n_170), .B(n_185), .Y(n_280) );
OAI21x1_ASAP7_75t_L g549 ( .A1(n_169), .A2(n_550), .B(n_557), .Y(n_549) );
OA21x2_ASAP7_75t_L g571 ( .A1(n_169), .A2(n_572), .B(n_580), .Y(n_571) );
OAI21x1_ASAP7_75t_L g587 ( .A1(n_169), .A2(n_550), .B(n_557), .Y(n_587) );
OAI21x1_ASAP7_75t_L g616 ( .A1(n_169), .A2(n_572), .B(n_580), .Y(n_616) );
O2A1O1Ixp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_175), .C(n_177), .Y(n_171) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g227 ( .A(n_176), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_177), .A2(n_511), .B(n_513), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_177), .A2(n_528), .B(n_529), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_177), .A2(n_552), .B(n_553), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_177), .A2(n_631), .B(n_632), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_181), .B1(n_183), .B2(n_184), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_180), .A2(n_541), .B(n_542), .Y(n_540) );
INVx2_ASAP7_75t_SL g180 ( .A(n_181), .Y(n_180) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_181), .A2(n_515), .B1(n_516), .B2(n_517), .Y(n_514) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
BUFx3_ASAP7_75t_L g219 ( .A(n_182), .Y(n_219) );
INVx2_ASAP7_75t_L g208 ( .A(n_186), .Y(n_208) );
NOR2xp67_ASAP7_75t_SL g596 ( .A(n_186), .B(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AO31x2_ASAP7_75t_L g560 ( .A1(n_187), .A2(n_561), .A3(n_568), .B(n_569), .Y(n_560) );
AND2x2_ASAP7_75t_L g263 ( .A(n_188), .B(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g282 ( .A(n_188), .Y(n_282) );
OR2x2_ASAP7_75t_L g302 ( .A(n_188), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g343 ( .A(n_188), .Y(n_343) );
INVx1_ASAP7_75t_L g354 ( .A(n_188), .Y(n_354) );
AND2x2_ASAP7_75t_L g361 ( .A(n_188), .B(n_303), .Y(n_361) );
AO31x2_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .A3(n_197), .B(n_199), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_192), .B(n_218), .Y(n_217) );
INVx1_ASAP7_75t_SL g194 ( .A(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g214 ( .A(n_195), .Y(n_214) );
INVx2_ASAP7_75t_SL g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_SL g238 ( .A(n_198), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
INVx2_ASAP7_75t_L g222 ( .A(n_201), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_201), .B(n_570), .Y(n_569) );
HB1xp67_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NAND2x1p5_ASAP7_75t_L g203 ( .A(n_204), .B(n_232), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_205), .B(n_223), .Y(n_204) );
INVx1_ASAP7_75t_L g275 ( .A(n_205), .Y(n_275) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_206), .Y(n_287) );
INVx1_ASAP7_75t_L g296 ( .A(n_206), .Y(n_296) );
INVx1_ASAP7_75t_L g335 ( .A(n_206), .Y(n_335) );
AND2x2_ASAP7_75t_L g365 ( .A(n_206), .B(n_224), .Y(n_365) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g259 ( .A(n_207), .Y(n_259) );
AOI21x1_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_221), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_215), .B(n_220), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_211), .B(n_214), .Y(n_210) );
AOI21x1_ASAP7_75t_L g576 ( .A1(n_214), .A2(n_577), .B(n_578), .Y(n_576) );
INVx1_ASAP7_75t_L g516 ( .A(n_216), .Y(n_516) );
INVx2_ASAP7_75t_L g229 ( .A(n_219), .Y(n_229) );
INVx2_ASAP7_75t_L g567 ( .A(n_219), .Y(n_567) );
INVx1_ASAP7_75t_L g271 ( .A(n_223), .Y(n_271) );
AND2x4_ASAP7_75t_L g320 ( .A(n_223), .B(n_234), .Y(n_320) );
AND2x2_ASAP7_75t_L g330 ( .A(n_223), .B(n_259), .Y(n_330) );
INVx1_ASAP7_75t_L g391 ( .A(n_223), .Y(n_391) );
INVx3_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
OR2x2_ASAP7_75t_L g277 ( .A(n_224), .B(n_256), .Y(n_277) );
AND2x2_ASAP7_75t_L g295 ( .A(n_224), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g311 ( .A(n_224), .B(n_256), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_224), .B(n_239), .Y(n_420) );
AOI21x1_ASAP7_75t_L g243 ( .A1(n_229), .A2(n_244), .B(n_245), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g633 ( .A1(n_229), .A2(n_634), .B(n_635), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_232), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_239), .Y(n_232) );
OR2x2_ASAP7_75t_L g437 ( .A(n_233), .B(n_239), .Y(n_437) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g384 ( .A(n_234), .Y(n_384) );
AND2x2_ASAP7_75t_L g409 ( .A(n_234), .B(n_239), .Y(n_409) );
OAI21x1_ASAP7_75t_L g242 ( .A1(n_238), .A2(n_243), .B(n_246), .Y(n_242) );
INVx3_ASAP7_75t_L g260 ( .A(n_239), .Y(n_260) );
AND2x2_ASAP7_75t_L g286 ( .A(n_239), .B(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g308 ( .A(n_239), .Y(n_308) );
INVx1_ASAP7_75t_L g322 ( .A(n_239), .Y(n_322) );
INVx1_ASAP7_75t_L g332 ( .A(n_239), .Y(n_332) );
BUFx2_ASAP7_75t_L g427 ( .A(n_239), .Y(n_427) );
OR2x2_ASAP7_75t_L g455 ( .A(n_239), .B(n_259), .Y(n_455) );
INVxp67_ASAP7_75t_L g472 ( .A(n_239), .Y(n_472) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
OAI21x1_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_250), .Y(n_240) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_257), .Y(n_252) );
AND2x4_ASAP7_75t_L g285 ( .A(n_253), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_253), .B(n_365), .Y(n_446) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g273 ( .A(n_255), .B(n_260), .Y(n_273) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_255), .Y(n_297) );
INVx1_ASAP7_75t_L g421 ( .A(n_255), .Y(n_421) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g334 ( .A(n_256), .Y(n_334) );
AND2x2_ASAP7_75t_L g348 ( .A(n_257), .B(n_311), .Y(n_348) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
INVx1_ASAP7_75t_L g310 ( .A(n_259), .Y(n_310) );
OR2x2_ASAP7_75t_L g368 ( .A(n_259), .B(n_334), .Y(n_368) );
INVx1_ASAP7_75t_L g431 ( .A(n_259), .Y(n_431) );
AND2x2_ASAP7_75t_L g374 ( .A(n_260), .B(n_320), .Y(n_374) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x4_ASAP7_75t_L g262 ( .A(n_263), .B(n_265), .Y(n_262) );
AND2x2_ASAP7_75t_L g377 ( .A(n_263), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_269), .Y(n_265) );
AND2x2_ASAP7_75t_L g281 ( .A(n_266), .B(n_282), .Y(n_281) );
NAND2x1p5_ASAP7_75t_L g326 ( .A(n_266), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g300 ( .A(n_267), .Y(n_300) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g379 ( .A(n_268), .B(n_304), .Y(n_379) );
AND2x2_ASAP7_75t_L g342 ( .A(n_269), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g413 ( .A(n_269), .Y(n_413) );
A2O1A1Ixp33_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_272), .B(n_274), .C(n_278), .Y(n_270) );
INVx1_ASAP7_75t_L g405 ( .A(n_272), .Y(n_405) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x4_ASAP7_75t_L g401 ( .A(n_273), .B(n_365), .Y(n_401) );
INVx1_ASAP7_75t_L g492 ( .A(n_273), .Y(n_492) );
INVx1_ASAP7_75t_L g457 ( .A(n_274), .Y(n_457) );
AND2x4_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
AND2x2_ASAP7_75t_L g490 ( .A(n_275), .B(n_409), .Y(n_490) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g307 ( .A(n_277), .B(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g462 ( .A(n_277), .B(n_427), .Y(n_462) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
INVxp67_ASAP7_75t_L g352 ( .A(n_279), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_279), .B(n_314), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_279), .B(n_281), .Y(n_444) );
INVx1_ASAP7_75t_L g327 ( .A(n_280), .Y(n_327) );
INVx2_ASAP7_75t_SL g292 ( .A(n_282), .Y(n_292) );
OR2x2_ASAP7_75t_L g321 ( .A(n_282), .B(n_322), .Y(n_321) );
OAI221xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_288), .B1(n_293), .B2(n_298), .C(n_305), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NOR2xp33_ASAP7_75t_SL g329 ( .A(n_285), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g357 ( .A(n_287), .Y(n_357) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx1_ASAP7_75t_L g414 ( .A(n_290), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_290), .B(n_292), .Y(n_452) );
OR2x2_ASAP7_75t_L g434 ( .A(n_291), .B(n_424), .Y(n_434) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g403 ( .A(n_292), .B(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g450 ( .A(n_292), .B(n_379), .Y(n_450) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
AND2x2_ASAP7_75t_L g385 ( .A(n_295), .B(n_308), .Y(n_385) );
BUFx2_ASAP7_75t_L g411 ( .A(n_295), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_299), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g314 ( .A(n_300), .Y(n_314) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g387 ( .A(n_302), .Y(n_387) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OAI21xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_309), .B(n_312), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g364 ( .A(n_308), .Y(n_364) );
INVxp67_ASAP7_75t_SL g367 ( .A(n_308), .Y(n_367) );
OR2x2_ASAP7_75t_L g477 ( .A(n_308), .B(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g438 ( .A(n_309), .Y(n_438) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_L g346 ( .A(n_310), .Y(n_346) );
AND2x2_ASAP7_75t_L g473 ( .A(n_311), .B(n_346), .Y(n_473) );
INVx2_ASAP7_75t_SL g478 ( .A(n_311), .Y(n_478) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx2_ASAP7_75t_L g360 ( .A(n_314), .Y(n_360) );
AND2x4_ASAP7_75t_L g336 ( .A(n_315), .B(n_325), .Y(n_336) );
INVx2_ASAP7_75t_L g400 ( .A(n_315), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_315), .B(n_341), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_315), .B(n_371), .Y(n_487) );
AOI221x1_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_323), .B1(n_328), .B2(n_336), .C(n_337), .Y(n_316) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
INVx2_ASAP7_75t_L g456 ( .A(n_319), .Y(n_456) );
AOI21xp33_ASAP7_75t_L g463 ( .A1(n_319), .A2(n_464), .B(n_466), .Y(n_463) );
INVx3_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g345 ( .A(n_320), .B(n_346), .Y(n_345) );
BUFx2_ASAP7_75t_L g376 ( .A(n_320), .Y(n_376) );
AND2x4_ASAP7_75t_L g430 ( .A(n_320), .B(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g390 ( .A(n_322), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI32xp33_ASAP7_75t_L g435 ( .A1(n_324), .A2(n_433), .A3(n_436), .B1(n_438), .B2(n_439), .Y(n_435) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_325), .B(n_342), .Y(n_458) );
AND2x2_ASAP7_75t_L g474 ( .A(n_325), .B(n_354), .Y(n_474) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_329), .B(n_331), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_330), .B(n_472), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g406 ( .A1(n_331), .A2(n_407), .B(n_410), .C(n_412), .Y(n_406) );
NAND2x1p5_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx1_ASAP7_75t_L g355 ( .A(n_333), .Y(n_355) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
OAI21xp33_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_344), .B(n_347), .Y(n_337) );
OAI21xp33_ASAP7_75t_L g372 ( .A1(n_338), .A2(n_373), .B(n_375), .Y(n_372) );
INVx2_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_342), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_341), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_345), .A2(n_418), .B1(n_422), .B2(n_423), .Y(n_417) );
AND2x2_ASAP7_75t_L g484 ( .A(n_345), .B(n_472), .Y(n_484) );
NOR2xp33_ASAP7_75t_SL g349 ( .A(n_350), .B(n_372), .Y(n_349) );
OAI221xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_355), .B1(n_356), .B2(n_358), .C(n_362), .Y(n_350) );
AOI21xp33_ASAP7_75t_L g460 ( .A1(n_351), .A2(n_461), .B(n_462), .Y(n_460) );
OR2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
AND2x2_ASAP7_75t_L g443 ( .A(n_357), .B(n_409), .Y(n_443) );
INVxp67_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
AOI31xp33_ASAP7_75t_L g380 ( .A1(n_360), .A2(n_381), .A3(n_386), .B(n_388), .Y(n_380) );
AND2x2_ASAP7_75t_L g480 ( .A(n_360), .B(n_387), .Y(n_480) );
AND2x2_ASAP7_75t_L g369 ( .A(n_361), .B(n_370), .Y(n_369) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_361), .Y(n_433) );
INVx1_ASAP7_75t_L g467 ( .A(n_361), .Y(n_467) );
OAI21xp33_ASAP7_75t_SL g362 ( .A1(n_363), .A2(n_366), .B(n_369), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVx2_ASAP7_75t_L g393 ( .A(n_365), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_365), .B(n_492), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_366), .A2(n_449), .B(n_451), .Y(n_448) );
NOR2x1p5_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
O2A1O1Ixp33_ASAP7_75t_L g389 ( .A1(n_368), .A2(n_383), .B(n_390), .C(n_392), .Y(n_389) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g402 ( .A(n_371), .B(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g422 ( .A(n_371), .B(n_378), .Y(n_422) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g404 ( .A(n_379), .Y(n_404) );
INVx1_ASAP7_75t_L g440 ( .A(n_379), .Y(n_440) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_385), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_385), .A2(n_402), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g461 ( .A(n_385), .Y(n_461) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NOR2x1_ASAP7_75t_L g394 ( .A(n_395), .B(n_447), .Y(n_394) );
NAND3xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_415), .C(n_425), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_401), .B1(n_402), .B2(n_405), .C(n_406), .Y(n_396) );
INVx3_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_403), .A2(n_470), .B1(n_473), .B2(n_474), .Y(n_469) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
BUFx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
OR2x2_ASAP7_75t_L g466 ( .A(n_414), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
INVx1_ASAP7_75t_L g465 ( .A(n_420), .Y(n_465) );
INVx2_ASAP7_75t_L g445 ( .A(n_422), .Y(n_445) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AOI211xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_428), .B(n_435), .C(n_441), .Y(n_425) );
BUFx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OAI21xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_432), .B(n_434), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g436 ( .A(n_431), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g479 ( .A(n_436), .Y(n_479) );
OAI22xp33_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_444), .B1(n_445), .B2(n_446), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND4xp75_ASAP7_75t_L g447 ( .A(n_448), .B(n_459), .C(n_468), .D(n_481), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OAI22xp33_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B1(n_457), .B2(n_458), .Y(n_451) );
NAND2x1_ASAP7_75t_SL g453 ( .A(n_454), .B(n_456), .Y(n_453) );
INVx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_463), .Y(n_459) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_475), .Y(n_468) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
OAI21xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_479), .B(n_480), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_484), .B1(n_485), .B2(n_488), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVxp67_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_491), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g494 ( .A(n_495), .Y(n_494) );
BUFx8_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g850 ( .A(n_496), .Y(n_850) );
AND2x2_ASAP7_75t_L g864 ( .A(n_496), .B(n_865), .Y(n_864) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_781), .Y(n_499) );
NAND4xp25_ASAP7_75t_L g500 ( .A(n_501), .B(n_656), .C(n_696), .D(n_745), .Y(n_500) );
NOR2xp67_ASAP7_75t_L g501 ( .A(n_502), .B(n_607), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_532), .B1(n_581), .B2(n_590), .Y(n_502) );
INVx1_ASAP7_75t_L g777 ( .A(n_503), .Y(n_777) );
INVx1_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_504), .B(n_626), .Y(n_693) );
AND2x2_ASAP7_75t_L g724 ( .A(n_504), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_519), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_505), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g648 ( .A(n_505), .Y(n_648) );
AND2x2_ASAP7_75t_L g823 ( .A(n_505), .B(n_691), .Y(n_823) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx2_ASAP7_75t_L g592 ( .A(n_506), .Y(n_592) );
AND2x2_ASAP7_75t_L g676 ( .A(n_506), .B(n_638), .Y(n_676) );
AND2x2_ASAP7_75t_L g720 ( .A(n_506), .B(n_627), .Y(n_720) );
OR2x2_ASAP7_75t_L g738 ( .A(n_506), .B(n_739), .Y(n_738) );
INVx4_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g642 ( .A(n_507), .B(n_627), .Y(n_642) );
BUFx2_ASAP7_75t_L g699 ( .A(n_507), .Y(n_699) );
OR2x2_ASAP7_75t_L g707 ( .A(n_507), .B(n_665), .Y(n_707) );
INVx1_ASAP7_75t_L g762 ( .A(n_507), .Y(n_762) );
AND2x4_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
OAI21x1_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_514), .B(n_518), .Y(n_509) );
AND2x2_ASAP7_75t_L g593 ( .A(n_519), .B(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g701 ( .A(n_519), .B(n_678), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_519), .B(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g739 ( .A(n_520), .Y(n_739) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_520), .Y(n_744) );
AND2x2_ASAP7_75t_L g761 ( .A(n_520), .B(n_762), .Y(n_761) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g651 ( .A(n_521), .B(n_595), .Y(n_651) );
INVx1_ASAP7_75t_L g665 ( .A(n_521), .Y(n_665) );
OAI21x1_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B(n_530), .Y(n_521) );
NAND2x1_ASAP7_75t_L g532 ( .A(n_533), .B(n_545), .Y(n_532) );
AND2x4_ASAP7_75t_L g826 ( .A(n_533), .B(n_754), .Y(n_826) );
INVxp67_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
INVxp67_ASAP7_75t_SL g589 ( .A(n_534), .Y(n_589) );
BUFx3_ASAP7_75t_L g622 ( .A(n_534), .Y(n_622) );
INVx1_ASAP7_75t_L g686 ( .A(n_534), .Y(n_686) );
AND2x2_ASAP7_75t_L g689 ( .A(n_534), .B(n_548), .Y(n_689) );
AND2x2_ASAP7_75t_L g714 ( .A(n_534), .B(n_571), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_534), .Y(n_717) );
AND2x2_ASAP7_75t_L g749 ( .A(n_534), .B(n_616), .Y(n_749) );
INVx3_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x4_ASAP7_75t_L g545 ( .A(n_546), .B(n_558), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g658 ( .A(n_547), .B(n_644), .Y(n_658) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g684 ( .A(n_549), .B(n_671), .Y(n_684) );
AND2x2_ASAP7_75t_L g713 ( .A(n_549), .B(n_560), .Y(n_713) );
OR2x2_ASAP7_75t_L g809 ( .A(n_549), .B(n_560), .Y(n_809) );
AND2x2_ASAP7_75t_L g688 ( .A(n_558), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g837 ( .A(n_558), .Y(n_837) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_559), .Y(n_583) );
OR2x2_ASAP7_75t_L g771 ( .A(n_559), .B(n_585), .Y(n_771) );
INVx1_ASAP7_75t_L g793 ( .A(n_559), .Y(n_793) );
OR2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_571), .Y(n_559) );
AND2x2_ASAP7_75t_L g611 ( .A(n_560), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g644 ( .A(n_560), .B(n_616), .Y(n_644) );
INVx1_ASAP7_75t_L g671 ( .A(n_560), .Y(n_671) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_560), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_560), .B(n_571), .Y(n_758) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_567), .B(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g597 ( .A(n_568), .Y(n_597) );
AND2x2_ASAP7_75t_L g695 ( .A(n_571), .B(n_617), .Y(n_695) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NOR3x1_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .C(n_588), .Y(n_582) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_585), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g643 ( .A(n_585), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g694 ( .A(n_585), .B(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g734 ( .A(n_585), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_585), .B(n_757), .Y(n_789) );
INVx3_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NOR2xp67_ASAP7_75t_L g730 ( .A(n_586), .B(n_670), .Y(n_730) );
AND2x2_ASAP7_75t_L g754 ( .A(n_586), .B(n_616), .Y(n_754) );
BUFx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g612 ( .A(n_587), .Y(n_612) );
BUFx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g765 ( .A(n_589), .B(n_644), .Y(n_765) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_592), .B(n_651), .Y(n_830) );
AND2x4_ASAP7_75t_L g822 ( .A(n_593), .B(n_823), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_593), .B(n_642), .Y(n_836) );
INVx2_ASAP7_75t_L g638 ( .A(n_594), .Y(n_638) );
INVx1_ASAP7_75t_L g641 ( .A(n_594), .Y(n_641) );
INVx2_ASAP7_75t_L g726 ( .A(n_594), .Y(n_726) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g710 ( .A(n_595), .Y(n_710) );
AOI21x1_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_598), .B(n_606), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_602), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_645), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_623), .B1(n_639), .B2(n_643), .Y(n_608) );
OAI21xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_613), .B(n_618), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g673 ( .A(n_611), .B(n_622), .Y(n_673) );
AND2x2_ASAP7_75t_L g833 ( .A(n_611), .B(n_714), .Y(n_833) );
BUFx2_ASAP7_75t_L g704 ( .A(n_612), .Y(n_704) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
BUFx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g703 ( .A(n_615), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
INVx1_ASAP7_75t_L g620 ( .A(n_616), .Y(n_620) );
INVx1_ASAP7_75t_L g670 ( .A(n_616), .Y(n_670) );
INVx1_ASAP7_75t_L g795 ( .A(n_617), .Y(n_795) );
AOI31xp33_ASAP7_75t_L g813 ( .A1(n_618), .A2(n_814), .A3(n_815), .B(n_816), .Y(n_813) );
OR2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_619), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_620), .B(n_713), .Y(n_812) );
INVx2_ASAP7_75t_L g840 ( .A(n_620), .Y(n_840) );
INVxp67_ASAP7_75t_SL g655 ( .A(n_621), .Y(n_655) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g668 ( .A(n_622), .B(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_622), .B(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g798 ( .A(n_622), .B(n_758), .Y(n_798) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_637), .Y(n_624) );
INVx1_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g709 ( .A(n_627), .B(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g678 ( .A(n_628), .Y(n_678) );
AND2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_641), .Y(n_662) );
INVx1_ASAP7_75t_L g702 ( .A(n_641), .Y(n_702) );
INVx1_ASAP7_75t_L g682 ( .A(n_642), .Y(n_682) );
AND2x2_ASAP7_75t_L g743 ( .A(n_642), .B(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g799 ( .A(n_642), .B(n_726), .Y(n_799) );
OAI21xp5_ASAP7_75t_L g715 ( .A1(n_643), .A2(n_716), .B(n_718), .Y(n_715) );
OR2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_655), .Y(n_645) );
NAND3x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_649), .C(n_652), .Y(n_646) );
BUFx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g817 ( .A(n_648), .B(n_737), .Y(n_817) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NOR2x1_ASAP7_75t_SL g770 ( .A(n_650), .B(n_682), .Y(n_770) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g690 ( .A(n_651), .B(n_691), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_652), .B(n_767), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_652), .B(n_761), .Y(n_788) );
NOR2xp33_ASAP7_75t_L g834 ( .A(n_652), .B(n_761), .Y(n_834) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
BUFx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g737 ( .A(n_654), .B(n_710), .Y(n_737) );
AND2x2_ASAP7_75t_L g657 ( .A(n_655), .B(n_658), .Y(n_657) );
AOI221x1_ASAP7_75t_SL g656 ( .A1(n_657), .A2(n_659), .B1(n_666), .B2(n_675), .C(n_679), .Y(n_656) );
AOI32xp33_ASAP7_75t_L g838 ( .A1(n_658), .A2(n_839), .A3(n_844), .B1(n_845), .B2(n_847), .Y(n_838) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_660), .B(n_663), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_663), .B(n_817), .Y(n_816) );
BUFx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVxp67_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g677 ( .A(n_665), .B(n_678), .Y(n_677) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_665), .Y(n_681) );
OR2x2_ASAP7_75t_L g794 ( .A(n_665), .B(n_795), .Y(n_794) );
NAND3xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_672), .C(n_674), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AND2x4_ASAP7_75t_L g716 ( .A(n_669), .B(n_717), .Y(n_716) );
AND2x4_ASAP7_75t_L g733 ( .A(n_669), .B(n_734), .Y(n_733) );
AND2x4_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_672), .A2(n_769), .B1(n_771), .B2(n_772), .Y(n_768) );
INVx3_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
INVx1_ASAP7_75t_L g846 ( .A(n_676), .Y(n_846) );
INVx2_ASAP7_75t_L g691 ( .A(n_678), .Y(n_691) );
OAI21xp33_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_683), .B(n_687), .Y(n_679) );
OR2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
INVx1_ASAP7_75t_L g815 ( .A(n_684), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_685), .B(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_690), .B1(n_692), .B2(n_694), .Y(n_687) );
AND2x4_ASAP7_75t_L g784 ( .A(n_690), .B(n_699), .Y(n_784) );
INVx1_ASAP7_75t_L g843 ( .A(n_691), .Y(n_843) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g722 ( .A(n_695), .B(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_695), .B(n_808), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_695), .B(n_723), .Y(n_814) );
AOI211x1_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_703), .B(n_705), .C(n_731), .Y(n_696) );
AND2x4_ASAP7_75t_L g697 ( .A(n_698), .B(n_700), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OR3x2_ASAP7_75t_L g806 ( .A(n_699), .B(n_701), .C(n_702), .Y(n_806) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_700), .A2(n_722), .B1(n_724), .B2(n_727), .Y(n_721) );
NOR2x1p5_ASAP7_75t_SL g700 ( .A(n_701), .B(n_702), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_701), .A2(n_840), .B1(n_841), .B2(n_842), .Y(n_839) );
INVx2_ASAP7_75t_L g723 ( .A(n_704), .Y(n_723) );
OAI211xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_711), .B(n_715), .C(n_721), .Y(n_705) );
OR2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_713), .B(n_717), .Y(n_728) );
INVx1_ASAP7_75t_L g755 ( .A(n_713), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_713), .B(n_820), .Y(n_828) );
OAI32xp33_ASAP7_75t_L g803 ( .A1(n_714), .A2(n_759), .A3(n_804), .B1(n_806), .B2(n_807), .Y(n_803) );
INVx1_ASAP7_75t_L g820 ( .A(n_714), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_714), .B(n_734), .Y(n_824) );
NAND2xp5_ASAP7_75t_SL g786 ( .A(n_717), .B(n_751), .Y(n_786) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g764 ( .A(n_723), .B(n_749), .Y(n_764) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g773 ( .A(n_726), .B(n_774), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
INVx1_ASAP7_75t_L g741 ( .A(n_729), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_735), .B1(n_740), .B2(n_742), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
OR2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_738), .Y(n_735) );
INVx1_ASAP7_75t_L g779 ( .A(n_736), .Y(n_779) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g760 ( .A(n_737), .B(n_761), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_737), .B(n_744), .Y(n_848) );
INVx1_ASAP7_75t_SL g774 ( .A(n_738), .Y(n_774) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx3_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NOR3xp33_ASAP7_75t_L g745 ( .A(n_746), .B(n_768), .C(n_775), .Y(n_745) );
OAI21xp33_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_759), .B(n_763), .Y(n_746) );
NOR2xp33_ASAP7_75t_SL g747 ( .A(n_748), .B(n_752), .Y(n_747) );
INVxp67_ASAP7_75t_L g780 ( .A(n_748), .Y(n_780) );
AND2x2_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
INVx1_ASAP7_75t_L g805 ( .A(n_750), .Y(n_805) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
NAND3xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_755), .C(n_756), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g767 ( .A(n_761), .Y(n_767) );
OAI21xp33_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_765), .B(n_766), .Y(n_763) );
INVx1_ASAP7_75t_L g776 ( .A(n_764), .Y(n_776) );
OAI221xp5_ASAP7_75t_L g819 ( .A1(n_769), .A2(n_820), .B1(n_821), .B2(n_824), .C(n_825), .Y(n_819) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
OAI32xp33_ASAP7_75t_L g775 ( .A1(n_772), .A2(n_776), .A3(n_777), .B1(n_778), .B2(n_780), .Y(n_775) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
OAI221xp5_ASAP7_75t_L g787 ( .A1(n_778), .A2(n_788), .B1(n_789), .B2(n_790), .C(n_796), .Y(n_787) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
NAND3xp33_ASAP7_75t_L g781 ( .A(n_782), .B(n_800), .C(n_818), .Y(n_781) );
AOI21xp5_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_785), .B(n_787), .Y(n_782) );
AOI211x1_ASAP7_75t_L g800 ( .A1(n_783), .A2(n_801), .B(n_803), .C(n_810), .Y(n_800) );
HB1xp67_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVxp67_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
NOR2x1_ASAP7_75t_SL g791 ( .A(n_792), .B(n_794), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g802 ( .A(n_793), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_797), .B(n_799), .Y(n_796) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
AO21x1_ASAP7_75t_L g810 ( .A1(n_799), .A2(n_811), .B(n_813), .Y(n_810) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVxp67_ASAP7_75t_SL g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g844 ( .A(n_815), .Y(n_844) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_819), .B(n_831), .Y(n_818) );
INVx3_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
OAI21xp33_ASAP7_75t_SL g825 ( .A1(n_826), .A2(n_827), .B(n_829), .Y(n_825) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_832), .B(n_838), .Y(n_831) );
AOI21xp5_ASAP7_75t_L g832 ( .A1(n_833), .A2(n_834), .B(n_835), .Y(n_832) );
NOR2xp67_ASAP7_75t_L g835 ( .A(n_836), .B(n_837), .Y(n_835) );
INVx1_ASAP7_75t_L g841 ( .A(n_840), .Y(n_841) );
INVxp67_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
BUFx12f_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx3_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx6_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
BUFx10_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVxp67_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_868), .B(n_871), .Y(n_867) );
CKINVDCx11_ASAP7_75t_R g868 ( .A(n_869), .Y(n_868) );
BUFx6f_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
NOR2xp33_ASAP7_75t_L g906 ( .A(n_870), .B(n_907), .Y(n_906) );
INVxp67_ASAP7_75t_SL g909 ( .A(n_871), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_873), .B(n_877), .Y(n_872) );
INVx1_ASAP7_75t_L g884 ( .A(n_873), .Y(n_884) );
INVx4_ASAP7_75t_L g887 ( .A(n_877), .Y(n_887) );
BUFx12f_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx4_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx3_ASAP7_75t_L g890 ( .A(n_879), .Y(n_890) );
INVx5_ASAP7_75t_L g898 ( .A(n_879), .Y(n_898) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
AOI21xp5_ASAP7_75t_L g883 ( .A1(n_884), .A2(n_885), .B(n_888), .Y(n_883) );
NOR2xp33_ASAP7_75t_L g885 ( .A(n_886), .B(n_887), .Y(n_885) );
OAI22xp5_ASAP7_75t_L g899 ( .A1(n_886), .A2(n_900), .B1(n_909), .B2(n_910), .Y(n_899) );
NOR2xp33_ASAP7_75t_L g888 ( .A(n_889), .B(n_890), .Y(n_888) );
OR2x6_ASAP7_75t_L g904 ( .A(n_890), .B(n_905), .Y(n_904) );
CKINVDCx20_ASAP7_75t_R g891 ( .A(n_892), .Y(n_891) );
CKINVDCx20_ASAP7_75t_R g892 ( .A(n_893), .Y(n_892) );
CKINVDCx5p33_ASAP7_75t_R g893 ( .A(n_894), .Y(n_893) );
CKINVDCx16_ASAP7_75t_R g894 ( .A(n_895), .Y(n_894) );
AND2x2_ASAP7_75t_L g895 ( .A(n_896), .B(n_898), .Y(n_895) );
INVx2_ASAP7_75t_SL g908 ( .A(n_896), .Y(n_908) );
CKINVDCx20_ASAP7_75t_R g900 ( .A(n_901), .Y(n_900) );
CKINVDCx20_ASAP7_75t_R g901 ( .A(n_902), .Y(n_901) );
INVx8_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
CKINVDCx20_ASAP7_75t_R g903 ( .A(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
OR2x4_ASAP7_75t_L g911 ( .A(n_907), .B(n_912), .Y(n_911) );
BUFx2_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx4_ASAP7_75t_SL g910 ( .A(n_911), .Y(n_910) );
endmodule