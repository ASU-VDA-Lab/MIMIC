module real_aes_1521_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_314;
wire n_252;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_0), .B(n_125), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_1), .A2(n_33), .B1(n_753), .B2(n_754), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_1), .Y(n_753) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_2), .A2(n_134), .B(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_3), .B(n_774), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_4), .B(n_125), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_5), .B(n_141), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_6), .B(n_141), .Y(n_545) );
INVx1_ASAP7_75t_L g132 ( .A(n_7), .Y(n_132) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_8), .A2(n_104), .B1(n_766), .B2(n_767), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_9), .B(n_141), .Y(n_512) );
CKINVDCx16_ASAP7_75t_R g774 ( .A(n_10), .Y(n_774) );
NAND2xp33_ASAP7_75t_L g522 ( .A(n_11), .B(n_143), .Y(n_522) );
AND2x2_ASAP7_75t_L g162 ( .A(n_12), .B(n_150), .Y(n_162) );
AND2x2_ASAP7_75t_L g171 ( .A(n_13), .B(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g147 ( .A(n_14), .Y(n_147) );
AOI221x1_ASAP7_75t_L g475 ( .A1(n_15), .A2(n_28), .B1(n_125), .B2(n_134), .C(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_16), .B(n_141), .Y(n_180) );
CKINVDCx16_ASAP7_75t_R g453 ( .A(n_17), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_18), .B(n_125), .Y(n_518) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_19), .A2(n_150), .B(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_20), .B(n_145), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_21), .B(n_141), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_22), .B(n_460), .Y(n_459) );
AO21x1_ASAP7_75t_L g540 ( .A1(n_23), .A2(n_125), .B(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_24), .B(n_125), .Y(n_205) );
INVx1_ASAP7_75t_L g457 ( .A(n_25), .Y(n_457) );
NOR2xp33_ASAP7_75t_SL g771 ( .A(n_25), .B(n_458), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_26), .A2(n_92), .B1(n_125), .B2(n_235), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g110 ( .A1(n_27), .A2(n_111), .B1(n_445), .B2(n_447), .Y(n_110) );
INVx1_ASAP7_75t_L g447 ( .A(n_27), .Y(n_447) );
NAND2x1_ASAP7_75t_L g485 ( .A(n_29), .B(n_141), .Y(n_485) );
NAND2x1_ASAP7_75t_L g511 ( .A(n_30), .B(n_143), .Y(n_511) );
OR2x2_ASAP7_75t_L g148 ( .A(n_31), .B(n_89), .Y(n_148) );
OA21x2_ASAP7_75t_L g151 ( .A1(n_31), .A2(n_89), .B(n_147), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_32), .B(n_143), .Y(n_506) );
CKINVDCx16_ASAP7_75t_R g754 ( .A(n_33), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_34), .B(n_141), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_35), .Y(n_761) );
AO21x2_ASAP7_75t_L g175 ( .A1(n_36), .A2(n_172), .B(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_37), .B(n_143), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_38), .A2(n_134), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_39), .B(n_141), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_40), .A2(n_134), .B(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g131 ( .A(n_41), .B(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g135 ( .A(n_41), .B(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g243 ( .A(n_41), .Y(n_243) );
OR2x6_ASAP7_75t_L g455 ( .A(n_42), .B(n_456), .Y(n_455) );
NOR3xp33_ASAP7_75t_L g772 ( .A(n_42), .B(n_453), .C(n_773), .Y(n_772) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_43), .B(n_125), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_44), .B(n_125), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_45), .B(n_141), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_46), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_47), .B(n_143), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_48), .B(n_125), .Y(n_124) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_49), .A2(n_134), .B(n_167), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_50), .A2(n_134), .B(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_51), .B(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_52), .B(n_143), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_53), .B(n_125), .Y(n_177) );
INVx1_ASAP7_75t_L g128 ( .A(n_54), .Y(n_128) );
INVx1_ASAP7_75t_L g138 ( .A(n_54), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_55), .B(n_141), .Y(n_169) );
OAI22xp5_ASAP7_75t_L g113 ( .A1(n_56), .A2(n_63), .B1(n_114), .B2(n_115), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_56), .Y(n_114) );
AND2x2_ASAP7_75t_L g196 ( .A(n_57), .B(n_145), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_58), .B(n_143), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_59), .B(n_141), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_60), .B(n_143), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_61), .A2(n_134), .B(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_62), .B(n_125), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_63), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_64), .B(n_125), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_65), .A2(n_134), .B(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g211 ( .A(n_66), .B(n_146), .Y(n_211) );
AO21x1_ASAP7_75t_L g542 ( .A1(n_67), .A2(n_134), .B(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_68), .B(n_125), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_69), .B(n_143), .Y(n_202) );
OAI22xp5_ASAP7_75t_SL g750 ( .A1(n_70), .A2(n_751), .B1(n_752), .B2(n_755), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_70), .Y(n_755) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_71), .B(n_125), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_72), .B(n_143), .Y(n_181) );
AOI22xp5_ASAP7_75t_L g240 ( .A1(n_73), .A2(n_97), .B1(n_134), .B2(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_74), .B(n_141), .Y(n_208) );
AND2x2_ASAP7_75t_L g496 ( .A(n_75), .B(n_146), .Y(n_496) );
INVx1_ASAP7_75t_L g130 ( .A(n_76), .Y(n_130) );
INVx1_ASAP7_75t_L g136 ( .A(n_76), .Y(n_136) );
AND2x2_ASAP7_75t_L g514 ( .A(n_77), .B(n_172), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_78), .B(n_143), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_79), .A2(n_134), .B(n_200), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g133 ( .A1(n_80), .A2(n_134), .B(n_139), .Y(n_133) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_81), .A2(n_134), .B(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g191 ( .A(n_82), .B(n_146), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_83), .B(n_145), .Y(n_232) );
INVx1_ASAP7_75t_L g458 ( .A(n_84), .Y(n_458) );
AND2x2_ASAP7_75t_L g500 ( .A(n_85), .B(n_172), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_86), .B(n_125), .Y(n_531) );
AND2x2_ASAP7_75t_L g149 ( .A(n_87), .B(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g541 ( .A(n_88), .B(n_182), .Y(n_541) );
AND2x2_ASAP7_75t_L g488 ( .A(n_90), .B(n_172), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_91), .B(n_143), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_93), .B(n_141), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_94), .B(n_143), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_95), .A2(n_134), .B(n_528), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_96), .A2(n_134), .B(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_98), .B(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_99), .B(n_141), .Y(n_505) );
BUFx2_ASAP7_75t_L g210 ( .A(n_100), .Y(n_210) );
BUFx2_ASAP7_75t_L g108 ( .A(n_101), .Y(n_108) );
INVx1_ASAP7_75t_SL g765 ( .A(n_101), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_102), .A2(n_134), .B(n_520), .Y(n_519) );
AO21x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_109), .B(n_462), .Y(n_104) );
BUFx3_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
HB1xp67_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OAI21xp5_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_448), .B(n_459), .Y(n_109) );
NAND2x1_ASAP7_75t_L g111 ( .A(n_112), .B(n_442), .Y(n_111) );
INVx1_ASAP7_75t_L g446 ( .A(n_112), .Y(n_446) );
NAND2x1p5_ASAP7_75t_L g112 ( .A(n_113), .B(n_116), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_113), .Y(n_444) );
INVx4_ASAP7_75t_L g443 ( .A(n_116), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_116), .A2(n_466), .B1(n_747), .B2(n_757), .Y(n_756) );
AND2x4_ASAP7_75t_L g116 ( .A(n_117), .B(n_350), .Y(n_116) );
NOR3xp33_ASAP7_75t_SL g117 ( .A(n_118), .B(n_273), .C(n_308), .Y(n_117) );
OAI211xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_173), .B(n_225), .C(n_263), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_152), .Y(n_120) );
AND2x2_ASAP7_75t_L g256 ( .A(n_121), .B(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_121), .B(n_262), .Y(n_296) );
AND2x2_ASAP7_75t_L g321 ( .A(n_121), .B(n_276), .Y(n_321) );
INVx4_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx2_ASAP7_75t_L g228 ( .A(n_122), .Y(n_228) );
OR2x2_ASAP7_75t_L g259 ( .A(n_122), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g267 ( .A(n_122), .B(n_163), .Y(n_267) );
AND2x2_ASAP7_75t_L g275 ( .A(n_122), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g302 ( .A(n_122), .B(n_303), .Y(n_302) );
NOR2x1_ASAP7_75t_L g313 ( .A(n_122), .B(n_305), .Y(n_313) );
AND2x4_ASAP7_75t_L g330 ( .A(n_122), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g368 ( .A(n_122), .Y(n_368) );
AND2x4_ASAP7_75t_SL g373 ( .A(n_122), .B(n_153), .Y(n_373) );
OR2x6_ASAP7_75t_L g122 ( .A(n_123), .B(n_149), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_133), .B(n_145), .Y(n_123) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_131), .Y(n_125) );
AND2x4_ASAP7_75t_L g126 ( .A(n_127), .B(n_129), .Y(n_126) );
AND2x6_ASAP7_75t_L g143 ( .A(n_127), .B(n_136), .Y(n_143) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g141 ( .A(n_129), .B(n_138), .Y(n_141) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx5_ASAP7_75t_L g144 ( .A(n_131), .Y(n_144) );
AND2x2_ASAP7_75t_L g137 ( .A(n_132), .B(n_138), .Y(n_137) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_132), .Y(n_238) );
AND2x6_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
BUFx3_ASAP7_75t_L g239 ( .A(n_135), .Y(n_239) );
INVx2_ASAP7_75t_L g245 ( .A(n_136), .Y(n_245) );
AND2x4_ASAP7_75t_L g241 ( .A(n_137), .B(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g237 ( .A(n_138), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_142), .B(n_144), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_143), .B(n_210), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_144), .A2(n_159), .B(n_160), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_144), .A2(n_168), .B(n_169), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_144), .A2(n_180), .B(n_181), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_144), .A2(n_188), .B(n_189), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_144), .A2(n_201), .B(n_202), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_144), .A2(n_208), .B(n_209), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_144), .A2(n_477), .B(n_478), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_144), .A2(n_485), .B(n_486), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_144), .A2(n_493), .B(n_494), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_144), .A2(n_505), .B(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_144), .A2(n_511), .B(n_512), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_144), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_144), .A2(n_529), .B(n_530), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_144), .A2(n_544), .B(n_545), .Y(n_543) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_145), .Y(n_155) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_145), .A2(n_234), .B(n_240), .Y(n_233) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_145), .A2(n_475), .B(n_479), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_145), .A2(n_502), .B(n_503), .Y(n_501) );
OA21x2_ASAP7_75t_L g581 ( .A1(n_145), .A2(n_475), .B(n_479), .Y(n_581) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_SL g146 ( .A(n_147), .B(n_148), .Y(n_146) );
AND2x4_ASAP7_75t_L g182 ( .A(n_147), .B(n_148), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_150), .A2(n_205), .B(n_206), .Y(n_204) );
BUFx4f_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx3_ASAP7_75t_L g164 ( .A(n_151), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_152), .B(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_152), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g152 ( .A(n_153), .B(n_163), .Y(n_152) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_153), .Y(n_268) );
INVx2_ASAP7_75t_L g304 ( .A(n_153), .Y(n_304) );
INVx1_ASAP7_75t_L g331 ( .A(n_153), .Y(n_331) );
AND2x2_ASAP7_75t_L g430 ( .A(n_153), .B(n_340), .Y(n_430) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_154), .Y(n_262) );
AND2x2_ASAP7_75t_L g276 ( .A(n_154), .B(n_163), .Y(n_276) );
AOI21x1_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_162), .Y(n_154) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_155), .A2(n_508), .B(n_514), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_157), .B(n_161), .Y(n_156) );
INVx2_ASAP7_75t_L g305 ( .A(n_163), .Y(n_305) );
INVx2_ASAP7_75t_L g340 ( .A(n_163), .Y(n_340) );
OR2x2_ASAP7_75t_L g425 ( .A(n_163), .B(n_257), .Y(n_425) );
AO21x2_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_165), .B(n_171), .Y(n_163) );
INVx4_ASAP7_75t_L g172 ( .A(n_164), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_166), .B(n_170), .Y(n_165) );
INVx3_ASAP7_75t_L g184 ( .A(n_172), .Y(n_184) );
AOI211xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_192), .B(n_212), .C(n_219), .Y(n_173) );
INVx2_ASAP7_75t_SL g314 ( .A(n_174), .Y(n_314) );
AND2x2_ASAP7_75t_L g320 ( .A(n_174), .B(n_193), .Y(n_320) );
AND2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_183), .Y(n_174) );
INVx1_ASAP7_75t_L g216 ( .A(n_175), .Y(n_216) );
INVx1_ASAP7_75t_L g222 ( .A(n_175), .Y(n_222) );
INVx2_ASAP7_75t_L g247 ( .A(n_175), .Y(n_247) );
AND2x2_ASAP7_75t_L g271 ( .A(n_175), .B(n_195), .Y(n_271) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_175), .Y(n_300) );
OR2x2_ASAP7_75t_L g380 ( .A(n_175), .B(n_203), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_182), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_182), .A2(n_198), .B(n_199), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_182), .A2(n_518), .B(n_519), .Y(n_517) );
INVx1_ASAP7_75t_SL g525 ( .A(n_182), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_182), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g246 ( .A(n_183), .B(n_247), .Y(n_246) );
NOR2x1_ASAP7_75t_SL g278 ( .A(n_183), .B(n_203), .Y(n_278) );
AO21x1_ASAP7_75t_SL g183 ( .A1(n_184), .A2(n_185), .B(n_191), .Y(n_183) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_184), .A2(n_185), .B(n_191), .Y(n_218) );
AO21x2_ASAP7_75t_L g481 ( .A1(n_184), .A2(n_482), .B(n_488), .Y(n_481) );
AO21x2_ASAP7_75t_L g489 ( .A1(n_184), .A2(n_490), .B(n_496), .Y(n_489) );
AO21x2_ASAP7_75t_L g548 ( .A1(n_184), .A2(n_490), .B(n_496), .Y(n_548) );
AO21x2_ASAP7_75t_L g573 ( .A1(n_184), .A2(n_482), .B(n_488), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_186), .B(n_190), .Y(n_185) );
INVxp67_ASAP7_75t_SL g192 ( .A(n_193), .Y(n_192) );
AND2x2_ASAP7_75t_L g292 ( .A(n_193), .B(n_215), .Y(n_292) );
AND2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_203), .Y(n_193) );
OR2x2_ASAP7_75t_L g224 ( .A(n_194), .B(n_203), .Y(n_224) );
BUFx2_ASAP7_75t_L g248 ( .A(n_194), .Y(n_248) );
NOR2xp67_ASAP7_75t_L g299 ( .A(n_194), .B(n_300), .Y(n_299) );
INVx4_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_195), .Y(n_251) );
AND2x2_ASAP7_75t_L g277 ( .A(n_195), .B(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g287 ( .A(n_195), .Y(n_287) );
NAND2x1_ASAP7_75t_L g325 ( .A(n_195), .B(n_203), .Y(n_325) );
OR2x2_ASAP7_75t_L g400 ( .A(n_195), .B(n_217), .Y(n_400) );
OR2x6_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
INVx2_ASAP7_75t_SL g213 ( .A(n_203), .Y(n_213) );
AND2x2_ASAP7_75t_L g272 ( .A(n_203), .B(n_217), .Y(n_272) );
AND2x2_ASAP7_75t_L g343 ( .A(n_203), .B(n_344), .Y(n_343) );
BUFx2_ASAP7_75t_L g364 ( .A(n_203), .Y(n_364) );
OR2x6_ASAP7_75t_L g203 ( .A(n_204), .B(n_211), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
INVx1_ASAP7_75t_SL g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g286 ( .A(n_215), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
BUFx2_ASAP7_75t_L g281 ( .A(n_216), .Y(n_281) );
AND2x2_ASAP7_75t_L g253 ( .A(n_217), .B(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g344 ( .A(n_217), .Y(n_344) );
INVx3_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_221), .B(n_223), .Y(n_220) );
OR2x2_ASAP7_75t_L g290 ( .A(n_221), .B(n_291), .Y(n_290) );
AND2x4_ASAP7_75t_SL g332 ( .A(n_221), .B(n_333), .Y(n_332) );
AOI322xp5_ASAP7_75t_L g369 ( .A1(n_221), .A2(n_248), .A3(n_370), .B1(n_372), .B2(n_375), .C1(n_377), .C2(n_379), .Y(n_369) );
AND2x2_ASAP7_75t_L g434 ( .A(n_221), .B(n_435), .Y(n_434) );
INVx3_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_222), .B(n_248), .Y(n_258) );
AOI322xp5_ASAP7_75t_L g309 ( .A1(n_223), .A2(n_310), .A3(n_314), .B1(n_315), .B2(n_318), .C1(n_320), .C2(n_321), .Y(n_309) );
INVx2_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
OR2x2_ASAP7_75t_L g361 ( .A(n_224), .B(n_314), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_224), .A2(n_421), .B1(n_423), .B2(n_426), .Y(n_420) );
OR2x2_ASAP7_75t_L g438 ( .A(n_224), .B(n_387), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_248), .B(n_249), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_229), .Y(n_226) );
AOI221xp5_ASAP7_75t_SL g288 ( .A1(n_227), .A2(n_264), .B1(n_289), .B2(n_292), .C(n_293), .Y(n_288) );
AND2x2_ASAP7_75t_L g315 ( .A(n_227), .B(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_228), .B(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g357 ( .A(n_228), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g386 ( .A(n_229), .Y(n_386) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_246), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_230), .B(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g328 ( .A(n_230), .Y(n_328) );
OR2x2_ASAP7_75t_L g335 ( .A(n_230), .B(n_336), .Y(n_335) );
INVx3_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g378 ( .A(n_231), .B(n_340), .Y(n_378) );
AND2x4_ASAP7_75t_L g231 ( .A(n_232), .B(n_233), .Y(n_231) );
AND2x4_ASAP7_75t_L g257 ( .A(n_232), .B(n_233), .Y(n_257) );
AND2x4_ASAP7_75t_L g235 ( .A(n_236), .B(n_239), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
NOR2x1p5_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
INVx3_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_246), .B(n_307), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_246), .B(n_287), .Y(n_383) );
INVx1_ASAP7_75t_L g387 ( .A(n_246), .Y(n_387) );
INVx1_ASAP7_75t_L g254 ( .A(n_247), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_255), .B1(n_258), .B2(n_259), .Y(n_249) );
OR2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
BUFx2_ASAP7_75t_SL g365 ( .A(n_253), .Y(n_365) );
AND2x2_ASAP7_75t_L g422 ( .A(n_254), .B(n_278), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_256), .B(n_285), .Y(n_284) );
NOR2xp33_ASAP7_75t_SL g294 ( .A(n_256), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_256), .B(n_415), .Y(n_414) );
BUFx3_ASAP7_75t_L g282 ( .A(n_257), .Y(n_282) );
INVx2_ASAP7_75t_L g312 ( .A(n_257), .Y(n_312) );
AND2x2_ASAP7_75t_L g355 ( .A(n_257), .B(n_339), .Y(n_355) );
INVx1_ASAP7_75t_L g269 ( .A(n_259), .Y(n_269) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
OAI21xp5_ASAP7_75t_SL g263 ( .A1(n_264), .A2(n_269), .B(n_270), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx1_ASAP7_75t_L g348 ( .A(n_267), .Y(n_348) );
INVx2_ASAP7_75t_L g336 ( .A(n_268), .Y(n_336) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
AND2x2_ASAP7_75t_L g333 ( .A(n_272), .B(n_287), .Y(n_333) );
OAI21xp5_ASAP7_75t_L g393 ( .A1(n_272), .A2(n_370), .B(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_274), .B(n_288), .Y(n_273) );
AOI32xp33_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_277), .A3(n_279), .B1(n_283), .B2(n_286), .Y(n_274) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_275), .Y(n_349) );
AOI221xp5_ASAP7_75t_L g381 ( .A1(n_275), .A2(n_364), .B1(n_382), .B2(n_384), .C(n_390), .Y(n_381) );
AND2x2_ASAP7_75t_L g401 ( .A(n_275), .B(n_282), .Y(n_401) );
BUFx2_ASAP7_75t_L g285 ( .A(n_276), .Y(n_285) );
INVx1_ASAP7_75t_L g410 ( .A(n_276), .Y(n_410) );
INVx1_ASAP7_75t_L g415 ( .A(n_276), .Y(n_415) );
INVx1_ASAP7_75t_SL g408 ( .A(n_277), .Y(n_408) );
INVx2_ASAP7_75t_L g291 ( .A(n_278), .Y(n_291) );
AND2x2_ASAP7_75t_L g403 ( .A(n_279), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
AND2x2_ASAP7_75t_L g375 ( .A(n_281), .B(n_376), .Y(n_375) );
OR2x2_ASAP7_75t_L g347 ( .A(n_282), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_282), .B(n_373), .Y(n_395) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g307 ( .A(n_287), .Y(n_307) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g297 ( .A(n_291), .B(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g306 ( .A(n_291), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g411 ( .A(n_292), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_297), .B1(n_301), .B2(n_306), .Y(n_293) );
INVx2_ASAP7_75t_SL g385 ( .A(n_295), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_295), .B(n_424), .Y(n_426) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_297), .A2(n_391), .B(n_392), .Y(n_390) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g342 ( .A(n_299), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g370 ( .A(n_302), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g317 ( .A(n_303), .Y(n_317) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_L g359 ( .A(n_305), .Y(n_359) );
INVx1_ASAP7_75t_L g404 ( .A(n_306), .Y(n_404) );
NAND3xp33_ASAP7_75t_L g308 ( .A(n_309), .B(n_322), .C(n_345), .Y(n_308) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
INVx2_ASAP7_75t_L g371 ( .A(n_311), .Y(n_371) );
AND2x2_ASAP7_75t_L g389 ( .A(n_311), .B(n_330), .Y(n_389) );
OR2x2_ASAP7_75t_L g428 ( .A(n_311), .B(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_312), .B(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g324 ( .A(n_314), .B(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g391 ( .A(n_317), .B(n_328), .Y(n_391) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_320), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g432 ( .A(n_320), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_326), .B1(n_330), .B2(n_332), .C(n_334), .Y(n_322) );
OAI21xp5_ASAP7_75t_L g345 ( .A1(n_323), .A2(n_346), .B(n_349), .Y(n_345) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx3_ASAP7_75t_L g376 ( .A(n_325), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_325), .B(n_419), .Y(n_418) );
INVxp33_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g337 ( .A(n_333), .Y(n_337) );
OAI22xp33_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_337), .B1(n_338), .B2(n_341), .Y(n_334) );
INVx2_ASAP7_75t_L g440 ( .A(n_336), .Y(n_440) );
BUFx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVxp67_ASAP7_75t_L g419 ( .A(n_344), .Y(n_419) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
NOR2x1_ASAP7_75t_L g350 ( .A(n_351), .B(n_396), .Y(n_350) );
NAND4xp25_ASAP7_75t_L g351 ( .A(n_352), .B(n_369), .C(n_381), .D(n_393), .Y(n_351) );
O2A1O1Ixp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_356), .B(n_360), .C(n_362), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g392 ( .A(n_355), .Y(n_392) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OAI21xp5_ASAP7_75t_L g362 ( .A1(n_357), .A2(n_363), .B(n_366), .Y(n_362) );
INVx2_ASAP7_75t_L g441 ( .A(n_358), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_359), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g374 ( .A(n_359), .Y(n_374) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
OR2x2_ASAP7_75t_L g436 ( .A(n_364), .B(n_400), .Y(n_436) );
INVxp67_ASAP7_75t_SL g407 ( .A(n_371), .Y(n_407) );
AND2x2_ASAP7_75t_SL g372 ( .A(n_373), .B(n_374), .Y(n_372) );
AND2x2_ASAP7_75t_L g377 ( .A(n_373), .B(n_378), .Y(n_377) );
AOI21xp5_ASAP7_75t_L g402 ( .A1(n_373), .A2(n_403), .B(n_405), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_373), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_SL g431 ( .A(n_373), .Y(n_431) );
INVxp67_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI22xp33_ASAP7_75t_SL g384 ( .A1(n_385), .A2(n_386), .B1(n_387), .B2(n_388), .Y(n_384) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND4xp25_ASAP7_75t_L g396 ( .A(n_397), .B(n_402), .C(n_412), .D(n_433), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_401), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_408), .B1(n_409), .B2(n_411), .Y(n_405) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AOI211xp5_ASAP7_75t_SL g412 ( .A1(n_413), .A2(n_416), .B(n_420), .C(n_427), .Y(n_412) );
INVxp67_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
AOI21xp33_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_431), .B(n_432), .Y(n_427) );
INVx1_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
OAI21xp5_ASAP7_75t_SL g433 ( .A1(n_434), .A2(n_437), .B(n_439), .Y(n_433) );
INVx1_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_443), .A2(n_444), .B(n_446), .Y(n_445) );
OAI22x1_ASAP7_75t_L g464 ( .A1(n_443), .A2(n_465), .B1(n_745), .B2(n_748), .Y(n_464) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVxp67_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx2_ASAP7_75t_R g451 ( .A(n_452), .Y(n_451) );
BUFx2_ASAP7_75t_L g461 ( .A(n_452), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
OR2x6_ASAP7_75t_SL g747 ( .A(n_453), .B(n_454), .Y(n_747) );
AND2x6_ASAP7_75t_SL g749 ( .A(n_453), .B(n_455), .Y(n_749) );
OR2x2_ASAP7_75t_L g764 ( .A(n_453), .B(n_455), .Y(n_764) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
AOI21xp5_ASAP7_75t_SL g462 ( .A1(n_459), .A2(n_463), .B(n_765), .Y(n_462) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AOI221xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_750), .B1(n_756), .B2(n_759), .C(n_760), .Y(n_463) );
INVx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x4_ASAP7_75t_L g466 ( .A(n_467), .B(n_657), .Y(n_466) );
AND4x1_ASAP7_75t_L g467 ( .A(n_468), .B(n_569), .C(n_596), .D(n_631), .Y(n_467) );
AOI221xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_497), .B1(n_534), .B2(n_549), .C(n_553), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_480), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_471), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OR2x2_ASAP7_75t_L g610 ( .A(n_472), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g665 ( .A(n_472), .B(n_620), .Y(n_665) );
BUFx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g568 ( .A(n_473), .B(n_489), .Y(n_568) );
AND2x4_ASAP7_75t_L g604 ( .A(n_473), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g618 ( .A(n_473), .B(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g535 ( .A(n_474), .Y(n_535) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_474), .Y(n_707) );
A2O1A1Ixp33_ASAP7_75t_SL g562 ( .A1(n_480), .A2(n_535), .B(n_563), .C(n_567), .Y(n_562) );
AND2x2_ASAP7_75t_L g583 ( .A(n_480), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_480), .B(n_535), .Y(n_723) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_489), .Y(n_480) );
INVx2_ASAP7_75t_L g603 ( .A(n_481), .Y(n_603) );
BUFx3_ASAP7_75t_L g619 ( .A(n_481), .Y(n_619) );
INVxp67_ASAP7_75t_L g623 ( .A(n_481), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_487), .Y(n_482) );
INVx2_ASAP7_75t_L g602 ( .A(n_489), .Y(n_602) );
AND2x2_ASAP7_75t_L g608 ( .A(n_489), .B(n_581), .Y(n_608) );
AND2x2_ASAP7_75t_L g634 ( .A(n_489), .B(n_603), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_491), .B(n_495), .Y(n_490) );
AOI211xp5_ASAP7_75t_L g631 ( .A1(n_497), .A2(n_632), .B(n_635), .C(n_645), .Y(n_631) );
AND2x2_ASAP7_75t_SL g497 ( .A(n_498), .B(n_515), .Y(n_497) );
OAI321xp33_ASAP7_75t_L g606 ( .A1(n_498), .A2(n_554), .A3(n_607), .B1(n_609), .B2(n_610), .C(n_612), .Y(n_606) );
AND2x2_ASAP7_75t_L g727 ( .A(n_498), .B(n_702), .Y(n_727) );
INVx1_ASAP7_75t_L g730 ( .A(n_498), .Y(n_730) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_507), .Y(n_498) );
INVx5_ASAP7_75t_L g552 ( .A(n_499), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_499), .B(n_566), .Y(n_565) );
NOR2x1_ASAP7_75t_SL g597 ( .A(n_499), .B(n_598), .Y(n_597) );
BUFx2_ASAP7_75t_L g642 ( .A(n_499), .Y(n_642) );
AND2x2_ASAP7_75t_L g744 ( .A(n_499), .B(n_516), .Y(n_744) );
OR2x6_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
AND2x2_ASAP7_75t_L g551 ( .A(n_507), .B(n_552), .Y(n_551) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_507), .Y(n_561) );
INVx4_ASAP7_75t_L g566 ( .A(n_507), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_513), .Y(n_508) );
INVx1_ASAP7_75t_L g609 ( .A(n_515), .Y(n_609) );
A2O1A1Ixp33_ASAP7_75t_R g712 ( .A1(n_515), .A2(n_551), .B(n_583), .C(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g732 ( .A(n_515), .B(n_557), .Y(n_732) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_523), .Y(n_515) );
INVx1_ASAP7_75t_L g550 ( .A(n_516), .Y(n_550) );
INVx2_ASAP7_75t_L g556 ( .A(n_516), .Y(n_556) );
OR2x2_ASAP7_75t_L g575 ( .A(n_516), .B(n_566), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_516), .B(n_598), .Y(n_644) );
BUFx3_ASAP7_75t_L g651 ( .A(n_516), .Y(n_651) );
INVx1_ASAP7_75t_L g614 ( .A(n_523), .Y(n_614) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_523), .Y(n_627) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g560 ( .A(n_524), .Y(n_560) );
INVx1_ASAP7_75t_L g669 ( .A(n_524), .Y(n_669) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_526), .B(n_532), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_525), .B(n_533), .Y(n_532) );
AO21x2_ASAP7_75t_L g598 ( .A1(n_525), .A2(n_526), .B(n_532), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_531), .Y(n_526) );
AND2x2_ASAP7_75t_L g570 ( .A(n_534), .B(n_571), .Y(n_570) );
OAI31xp33_ASAP7_75t_L g721 ( .A1(n_534), .A2(n_722), .A3(n_724), .B(n_727), .Y(n_721) );
INVx1_ASAP7_75t_SL g739 ( .A(n_534), .Y(n_739) );
AND2x4_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
AOI21xp33_ASAP7_75t_L g553 ( .A1(n_535), .A2(n_554), .B(n_562), .Y(n_553) );
NAND2x1_ASAP7_75t_L g633 ( .A(n_535), .B(n_634), .Y(n_633) );
INVx1_ASAP7_75t_SL g662 ( .A(n_535), .Y(n_662) );
INVx2_ASAP7_75t_L g611 ( .A(n_536), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_536), .B(n_594), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_536), .B(n_593), .Y(n_703) );
NOR2xp33_ASAP7_75t_SL g711 ( .A(n_536), .B(n_662), .Y(n_711) );
AND2x4_ASAP7_75t_L g536 ( .A(n_537), .B(n_548), .Y(n_536) );
AND2x2_ASAP7_75t_SL g580 ( .A(n_537), .B(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g591 ( .A(n_537), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g620 ( .A(n_537), .B(n_602), .Y(n_620) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx2_ASAP7_75t_L g584 ( .A(n_538), .Y(n_584) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g605 ( .A(n_539), .Y(n_605) );
OAI21x1_ASAP7_75t_SL g539 ( .A1(n_540), .A2(n_542), .B(n_546), .Y(n_539) );
INVx1_ASAP7_75t_L g547 ( .A(n_541), .Y(n_547) );
INVx2_ASAP7_75t_L g592 ( .A(n_548), .Y(n_592) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_548), .Y(n_652) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
INVx1_ASAP7_75t_L g588 ( .A(n_550), .Y(n_588) );
AND2x2_ASAP7_75t_L g667 ( .A(n_550), .B(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g578 ( .A(n_551), .B(n_572), .Y(n_578) );
INVx2_ASAP7_75t_SL g626 ( .A(n_551), .Y(n_626) );
INVx4_ASAP7_75t_L g557 ( .A(n_552), .Y(n_557) );
AND2x2_ASAP7_75t_L g655 ( .A(n_552), .B(n_598), .Y(n_655) );
AND2x2_ASAP7_75t_SL g673 ( .A(n_552), .B(n_668), .Y(n_673) );
NAND2x1p5_ASAP7_75t_L g690 ( .A(n_552), .B(n_566), .Y(n_690) );
INVx1_ASAP7_75t_L g696 ( .A(n_554), .Y(n_696) );
OR2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_558), .Y(n_554) );
INVx1_ASAP7_75t_L g615 ( .A(n_555), .Y(n_615) );
OR2x2_ASAP7_75t_L g628 ( .A(n_555), .B(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
OR2x2_ASAP7_75t_L g680 ( .A(n_556), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g710 ( .A(n_556), .B(n_598), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_557), .B(n_560), .Y(n_586) );
AND2x2_ASAP7_75t_L g678 ( .A(n_557), .B(n_668), .Y(n_678) );
AND2x4_ASAP7_75t_L g740 ( .A(n_557), .B(n_619), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
INVx2_ASAP7_75t_L g564 ( .A(n_559), .Y(n_564) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NOR2xp67_ASAP7_75t_SL g563 ( .A(n_564), .B(n_565), .Y(n_563) );
OAI322xp33_ASAP7_75t_SL g576 ( .A1(n_564), .A2(n_577), .A3(n_579), .B1(n_582), .B2(n_585), .C1(n_587), .C2(n_589), .Y(n_576) );
INVx1_ASAP7_75t_L g734 ( .A(n_564), .Y(n_734) );
OR2x2_ASAP7_75t_L g587 ( .A(n_565), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g613 ( .A(n_566), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_566), .B(n_614), .Y(n_629) );
INVx2_ASAP7_75t_L g656 ( .A(n_566), .Y(n_656) );
AND2x4_ASAP7_75t_L g668 ( .A(n_566), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_SL g671 ( .A(n_568), .B(n_584), .Y(n_671) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_574), .B(n_576), .Y(n_569) );
AND2x2_ASAP7_75t_L g637 ( .A(n_571), .B(n_604), .Y(n_637) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_572), .B(n_726), .Y(n_725) );
BUFx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g595 ( .A(n_573), .Y(n_595) );
AND2x4_ASAP7_75t_SL g677 ( .A(n_573), .B(n_592), .Y(n_677) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g585 ( .A(n_575), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_578), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g713 ( .A(n_580), .B(n_677), .Y(n_713) );
NOR4xp25_ASAP7_75t_L g717 ( .A(n_580), .B(n_594), .C(n_634), .D(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g594 ( .A(n_581), .B(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g630 ( .A(n_581), .B(n_605), .Y(n_630) );
AND2x4_ASAP7_75t_L g694 ( .A(n_581), .B(n_605), .Y(n_694) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_584), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
OR2x2_ASAP7_75t_L g683 ( .A(n_591), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g737 ( .A(n_591), .Y(n_737) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_592), .B(n_604), .Y(n_638) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
AOI211xp5_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_599), .B(n_606), .C(n_621), .Y(n_596) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_604), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_602), .B(n_605), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_603), .B(n_608), .Y(n_607) );
BUFx2_ASAP7_75t_L g685 ( .A(n_603), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_604), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g700 ( .A(n_604), .Y(n_700) );
OAI21xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_615), .B(n_616), .Y(n_612) );
AND2x4_ASAP7_75t_L g649 ( .A(n_613), .B(n_650), .Y(n_649) );
AND2x4_ASAP7_75t_L g743 ( .A(n_613), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
INVx1_ASAP7_75t_SL g647 ( .A(n_619), .Y(n_647) );
AND2x2_ASAP7_75t_L g706 ( .A(n_620), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g720 ( .A(n_620), .Y(n_720) );
O2A1O1Ixp33_ASAP7_75t_SL g621 ( .A1(n_622), .A2(n_624), .B(n_628), .C(n_630), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_622), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g698 ( .A(n_623), .B(n_699), .Y(n_698) );
OR2x2_ASAP7_75t_L g719 ( .A(n_623), .B(n_720), .Y(n_719) );
INVxp67_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
OR2x2_ASAP7_75t_L g708 ( .A(n_626), .B(n_650), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_629), .A2(n_636), .B1(n_638), .B2(n_639), .Y(n_635) );
INVx1_ASAP7_75t_SL g726 ( .A(n_630), .Y(n_726) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVxp67_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_641), .B(n_650), .Y(n_692) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVxp67_ASAP7_75t_SL g702 ( .A(n_644), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_648), .B1(n_652), .B2(n_653), .Y(n_645) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AOI21xp5_ASAP7_75t_SL g659 ( .A1(n_650), .A2(n_660), .B(n_663), .Y(n_659) );
AND2x2_ASAP7_75t_L g688 ( .A(n_650), .B(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND3x2_ASAP7_75t_L g654 ( .A(n_651), .B(n_655), .C(n_656), .Y(n_654) );
AND2x2_ASAP7_75t_L g716 ( .A(n_651), .B(n_673), .Y(n_716) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g701 ( .A(n_656), .B(n_702), .Y(n_701) );
NOR2xp67_ASAP7_75t_L g657 ( .A(n_658), .B(n_714), .Y(n_657) );
NAND4xp25_ASAP7_75t_L g658 ( .A(n_659), .B(n_674), .C(n_695), .D(n_712), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_666), .B1(n_670), .B2(n_672), .Y(n_663) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_666), .A2(n_680), .B1(n_700), .B2(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g681 ( .A(n_668), .Y(n_681) );
AOI21xp5_ASAP7_75t_L g741 ( .A1(n_670), .A2(n_693), .B(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx3_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_678), .B1(n_679), .B2(n_682), .C(n_686), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx2_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_691), .B1(n_692), .B2(n_693), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_689), .B(n_710), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_689), .B(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B1(n_701), .B2(n_703), .C(n_704), .Y(n_695) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_698), .B(n_700), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_708), .B1(n_709), .B2(n_711), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
OAI211xp5_ASAP7_75t_SL g729 ( .A1(n_710), .A2(n_730), .B(n_731), .C(n_733), .Y(n_729) );
OAI211xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_717), .B(n_721), .C(n_728), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
AOI221xp5_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_735), .B1(n_738), .B2(n_740), .C(n_741), .Y(n_728) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
CKINVDCx5p33_ASAP7_75t_R g745 ( .A(n_746), .Y(n_745) );
CKINVDCx11_ASAP7_75t_R g746 ( .A(n_747), .Y(n_746) );
INVx3_ASAP7_75t_SL g758 ( .A(n_748), .Y(n_758) );
CKINVDCx5p33_ASAP7_75t_R g748 ( .A(n_749), .Y(n_748) );
CKINVDCx12_ASAP7_75t_R g759 ( .A(n_750), .Y(n_759) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
CKINVDCx6p67_ASAP7_75t_R g757 ( .A(n_758), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
INVx2_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
INVx3_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx2_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
CKINVDCx16_ASAP7_75t_R g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_SL g770 ( .A(n_771), .B(n_772), .Y(n_770) );
endmodule