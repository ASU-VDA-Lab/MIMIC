module real_jpeg_3211_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_213;
wire n_167;
wire n_179;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_2),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_2),
.A2(n_39),
.B1(n_54),
.B2(n_55),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_2),
.A2(n_27),
.B1(n_30),
.B2(n_39),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_3),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_3),
.A2(n_29),
.B1(n_40),
.B2(n_42),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_4),
.A2(n_54),
.B(n_58),
.C(n_59),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_4),
.B(n_54),
.Y(n_58)
);

AO22x2_ASAP7_75t_L g59 ( 
.A1(n_4),
.A2(n_40),
.B1(n_42),
.B2(n_60),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

O2A1O1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_4),
.A2(n_12),
.B(n_54),
.C(n_180),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_8),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_8),
.A2(n_35),
.B1(n_40),
.B2(n_42),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_9),
.A2(n_40),
.B1(n_42),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_9),
.A2(n_49),
.B1(n_54),
.B2(n_55),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_9),
.A2(n_27),
.B1(n_30),
.B2(n_49),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_10),
.A2(n_69),
.B1(n_70),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_10),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_10),
.A2(n_54),
.B1(n_55),
.B2(n_128),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_10),
.A2(n_40),
.B1(n_42),
.B2(n_128),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_10),
.A2(n_27),
.B1(n_30),
.B2(n_128),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_11),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_11),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_11),
.A2(n_54),
.B1(n_55),
.B2(n_68),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_11),
.A2(n_40),
.B1(n_42),
.B2(n_68),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_11),
.A2(n_27),
.B1(n_30),
.B2(n_68),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_12),
.B(n_70),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_12),
.B(n_129),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_12),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_12),
.B(n_59),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_12),
.A2(n_54),
.B1(n_55),
.B2(n_181),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_12),
.B(n_27),
.C(n_45),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_12),
.A2(n_40),
.B1(n_42),
.B2(n_181),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_12),
.B(n_33),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_12),
.B(n_50),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_13),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_14),
.A2(n_54),
.B1(n_55),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_14),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_14),
.A2(n_62),
.B1(n_69),
.B2(n_70),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_14),
.A2(n_40),
.B1(n_42),
.B2(n_62),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_14),
.A2(n_27),
.B1(n_30),
.B2(n_62),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_15),
.A2(n_69),
.B1(n_70),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_15),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_15),
.A2(n_54),
.B1(n_55),
.B2(n_81),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_15),
.A2(n_40),
.B1(n_42),
.B2(n_81),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_15),
.A2(n_27),
.B1(n_30),
.B2(n_81),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_132),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_130),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_109),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_20),
.B(n_109),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_82),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_51),
.C(n_65),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_22),
.A2(n_23),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_24),
.A2(n_36),
.B1(n_37),
.B2(n_142),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_24),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_26),
.A2(n_33),
.B1(n_97),
.B2(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_32),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_27),
.A2(n_30),
.B1(n_45),
.B2(n_46),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_27),
.B(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_31),
.A2(n_32),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_31),
.A2(n_32),
.B1(n_156),
.B2(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_31),
.B(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_31),
.A2(n_212),
.B(n_213),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_31),
.A2(n_32),
.B1(n_212),
.B2(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_32),
.A2(n_171),
.B(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_32),
.B(n_185),
.Y(n_214)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_33),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_33),
.A2(n_184),
.B(n_241),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_43),
.B1(n_48),
.B2(n_50),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_38),
.A2(n_43),
.B1(n_50),
.B2(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_40),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_40),
.B(n_226),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g180 ( 
.A1(n_42),
.A2(n_60),
.B(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_43),
.A2(n_173),
.B(n_175),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_43),
.B(n_177),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_47),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_47),
.A2(n_86),
.B1(n_87),
.B2(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_47),
.A2(n_196),
.B(n_197),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_47),
.A2(n_197),
.B(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_47),
.A2(n_86),
.B1(n_174),
.B2(n_208),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_50),
.B(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_51),
.B(n_65),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_52),
.A2(n_63),
.B1(n_64),
.B2(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_52),
.A2(n_147),
.B(n_149),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_52),
.A2(n_149),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_53),
.B(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_53),
.A2(n_59),
.B1(n_148),
.B2(n_165),
.Y(n_193)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_55),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

AOI32xp33_ASAP7_75t_L g151 ( 
.A1(n_54),
.A2(n_69),
.A3(n_74),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_SL g153 ( 
.A(n_55),
.B(n_75),
.Y(n_153)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_59),
.B(n_125),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_61),
.A2(n_63),
.B(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_63),
.A2(n_124),
.B(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_71),
.B(n_78),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_67),
.A2(n_72),
.B1(n_127),
.B2(n_129),
.Y(n_126)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_69),
.A2(n_70),
.B1(n_74),
.B2(n_75),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_69),
.A2(n_71),
.B(n_181),
.C(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_103),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_77),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_101),
.B(n_102),
.Y(n_100)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_73),
.A2(n_102),
.B(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_79),
.B(n_189),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_92),
.B2(n_93),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_89),
.B(n_91),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_89),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_86),
.A2(n_176),
.B(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_105),
.B2(n_108),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_99),
.B1(n_100),
.B2(n_104),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_96),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_104),
.B1(n_106),
.B2(n_114),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_97),
.A2(n_181),
.B(n_214),
.Y(n_238)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_105),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_106),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.C(n_115),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_113),
.Y(n_135)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_122),
.C(n_126),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_117),
.B1(n_138),
.B2(n_140),
.Y(n_137)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_120),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_118),
.B(n_120),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_119),
.Y(n_196)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_122),
.A2(n_123),
.B1(n_126),
.B2(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI21x1_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_158),
.B(n_276),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_134),
.B(n_136),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_141),
.C(n_143),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_137),
.B(n_141),
.Y(n_261)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_138),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_143),
.B(n_261),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.C(n_150),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_144),
.B(n_146),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_150),
.B(n_264),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_151),
.A2(n_154),
.B1(n_155),
.B2(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_151),
.Y(n_200)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI31xp33_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_258),
.A3(n_268),
.B(n_273),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_202),
.B(n_257),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_186),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_161),
.B(n_186),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_172),
.C(n_178),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_162),
.B(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_167),
.C(n_170),
.Y(n_201)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_172),
.B(n_178),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_182),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_179),
.B(n_182),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_198),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_187),
.B(n_199),
.C(n_201),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_191),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_188),
.B(n_193),
.C(n_194),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_252),
.B(n_256),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_221),
.B(n_251),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_215),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_205),
.B(n_215),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.C(n_210),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_206),
.A2(n_207),
.B1(n_209),
.B2(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_210),
.A2(n_211),
.B1(n_230),
.B2(n_232),
.Y(n_229)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_220),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_217),
.B(n_219),
.C(n_220),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_233),
.B(n_250),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_229),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_229),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_224),
.A2(n_225),
.B1(n_227),
.B2(n_248),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_230),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_244),
.B(n_249),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_239),
.B(n_243),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_242),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_241),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_247),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_255),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_L g273 ( 
.A1(n_259),
.A2(n_274),
.B(n_275),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_262),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_265),
.C(n_266),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_270),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_265),
.Y(n_271)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_272),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_272),
.Y(n_274)
);


endmodule