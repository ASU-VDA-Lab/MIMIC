module fake_netlist_6_3358_n_1138 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1138);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1138;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_760;
wire n_741;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_1033;
wire n_607;
wire n_671;
wire n_726;
wire n_1052;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_955;
wire n_337;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1101;
wire n_1026;
wire n_443;
wire n_1099;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_1127;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_963;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_248;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_901;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_1078;
wire n_923;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_360;
wire n_977;
wire n_945;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_761;
wire n_428;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_842;
wire n_525;
wire n_1116;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_953;
wire n_1017;
wire n_1004;
wire n_886;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_986;
wire n_839;
wire n_734;
wire n_1088;
wire n_708;
wire n_196;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_1084;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_1121;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_984;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_981;
wire n_476;
wire n_880;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_982;
wire n_964;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_409;
wire n_345;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_1125;
wire n_275;
wire n_553;
wire n_652;
wire n_970;
wire n_849;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_882;
wire n_811;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_722;
wire n_688;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_956;
wire n_960;
wire n_841;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_1134;
wire n_332;
wire n_891;
wire n_336;
wire n_410;
wire n_398;
wire n_1129;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_43),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_80),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_106),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_179),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_101),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_23),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_77),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_128),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_17),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_191),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_115),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_175),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_176),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_61),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_97),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_81),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_4),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_155),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_79),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_32),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_50),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_130),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_54),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_168),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_183),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_78),
.Y(n_223)
);

BUFx10_ASAP7_75t_L g224 ( 
.A(n_99),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_178),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_20),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_129),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_60),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_24),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_188),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_24),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_169),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_1),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_0),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_6),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_38),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_75),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_164),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_31),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_102),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_181),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_143),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_89),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_1),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_171),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_105),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_87),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_67),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_3),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_17),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_121),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_39),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_12),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_34),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_14),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_124),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_63),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_165),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_15),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_190),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_103),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_30),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_166),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_46),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_194),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_119),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_96),
.Y(n_267)
);

INVxp67_ASAP7_75t_SL g268 ( 
.A(n_225),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_229),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_233),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_253),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_207),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_207),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_198),
.Y(n_274)
);

BUFx6f_ASAP7_75t_SL g275 ( 
.A(n_224),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_205),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_214),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_201),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_219),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_208),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_223),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_228),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_207),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_207),
.Y(n_284)
);

INVxp33_ASAP7_75t_L g285 ( 
.A(n_250),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_203),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_237),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_204),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_207),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_219),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_239),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g292 ( 
.A(n_213),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_264),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_267),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_260),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_260),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_234),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_261),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_207),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_261),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_262),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_262),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_226),
.Y(n_303)
);

INVxp33_ASAP7_75t_SL g304 ( 
.A(n_231),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_235),
.Y(n_305)
);

INVxp33_ASAP7_75t_SL g306 ( 
.A(n_244),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_255),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_241),
.Y(n_308)
);

NOR2xp67_ASAP7_75t_L g309 ( 
.A(n_213),
.B(n_0),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_212),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_259),
.Y(n_311)
);

INVxp33_ASAP7_75t_L g312 ( 
.A(n_212),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_212),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_217),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_212),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_249),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_310),
.Y(n_317)
);

NOR2x1_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_266),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_265),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_316),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_279),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_313),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_279),
.Y(n_323)
);

AND2x4_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_196),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_286),
.B(n_224),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_279),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_274),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_290),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_290),
.Y(n_329)
);

INVx5_ASAP7_75t_L g330 ( 
.A(n_272),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_312),
.B(n_197),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_276),
.Y(n_332)
);

AND2x4_ASAP7_75t_L g333 ( 
.A(n_280),
.B(n_263),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_269),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_268),
.B(n_232),
.Y(n_335)
);

OA21x2_ASAP7_75t_L g336 ( 
.A1(n_295),
.A2(n_200),
.B(n_199),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_270),
.Y(n_337)
);

INVx5_ASAP7_75t_L g338 ( 
.A(n_272),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_296),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_298),
.Y(n_340)
);

AND2x2_ASAP7_75t_SL g341 ( 
.A(n_314),
.B(n_232),
.Y(n_341)
);

AND2x4_ASAP7_75t_L g342 ( 
.A(n_281),
.B(n_258),
.Y(n_342)
);

AND2x6_ASAP7_75t_L g343 ( 
.A(n_273),
.B(n_29),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_300),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_301),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_302),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_273),
.Y(n_347)
);

BUFx12f_ASAP7_75t_L g348 ( 
.A(n_271),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_282),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_308),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_283),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_287),
.B(n_257),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_291),
.B(n_202),
.Y(n_353)
);

AND2x6_ASAP7_75t_L g354 ( 
.A(n_283),
.B(n_33),
.Y(n_354)
);

BUFx8_ASAP7_75t_L g355 ( 
.A(n_275),
.Y(n_355)
);

AND2x4_ASAP7_75t_L g356 ( 
.A(n_293),
.B(n_206),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_316),
.A2(n_236),
.B1(n_254),
.B2(n_252),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_284),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_284),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_294),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_289),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_278),
.B(n_209),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_277),
.B(n_210),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_289),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_299),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_299),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_278),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_307),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_307),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_297),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_275),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_R g372 ( 
.A(n_371),
.B(n_271),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_371),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_R g374 ( 
.A(n_348),
.B(n_288),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_360),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_360),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_317),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_334),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_317),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_370),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_334),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_355),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_355),
.Y(n_383)
);

NAND2xp33_ASAP7_75t_R g384 ( 
.A(n_320),
.B(n_304),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_355),
.Y(n_385)
);

NAND2xp33_ASAP7_75t_R g386 ( 
.A(n_320),
.B(n_304),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_358),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_355),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_R g389 ( 
.A(n_348),
.B(n_288),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_370),
.Y(n_390)
);

BUFx10_ASAP7_75t_L g391 ( 
.A(n_341),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_362),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_341),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_341),
.B(n_303),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_358),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_331),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_367),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_367),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_363),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_337),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_352),
.B(n_306),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_368),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_R g403 ( 
.A(n_368),
.B(n_303),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_317),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_369),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_369),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_357),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_337),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_363),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_R g410 ( 
.A(n_319),
.B(n_305),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_327),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_357),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_R g413 ( 
.A(n_319),
.B(n_305),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_317),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_325),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_327),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_332),
.Y(n_417)
);

BUFx10_ASAP7_75t_L g418 ( 
.A(n_333),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_335),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_332),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_349),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_349),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_335),
.Y(n_423)
);

OAI21x1_ASAP7_75t_L g424 ( 
.A1(n_347),
.A2(n_215),
.B(n_211),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_333),
.Y(n_425)
);

BUFx10_ASAP7_75t_L g426 ( 
.A(n_333),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_333),
.Y(n_427)
);

INVxp33_ASAP7_75t_L g428 ( 
.A(n_350),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_318),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_342),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_342),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_350),
.Y(n_432)
);

NOR2xp67_ASAP7_75t_L g433 ( 
.A(n_330),
.B(n_216),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_318),
.Y(n_434)
);

BUFx10_ASAP7_75t_L g435 ( 
.A(n_342),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_324),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_342),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_353),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_364),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_353),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_317),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_324),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_353),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_364),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_353),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_380),
.B(n_306),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_375),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_376),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_436),
.B(n_347),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_390),
.B(n_285),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_387),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_378),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_381),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_428),
.B(n_356),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_400),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_436),
.B(n_324),
.Y(n_456)
);

INVx5_ASAP7_75t_L g457 ( 
.A(n_379),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_387),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_374),
.Y(n_459)
);

NAND3xp33_ASAP7_75t_L g460 ( 
.A(n_399),
.B(n_356),
.C(n_336),
.Y(n_460)
);

INVx4_ASAP7_75t_L g461 ( 
.A(n_379),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_395),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_411),
.B(n_356),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_395),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_409),
.B(n_356),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_374),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_442),
.Y(n_467)
);

INVx8_ASAP7_75t_L g468 ( 
.A(n_425),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_442),
.B(n_324),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_392),
.B(n_218),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_408),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_439),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_444),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_423),
.B(n_311),
.Y(n_474)
);

AND2x6_ASAP7_75t_L g475 ( 
.A(n_416),
.B(n_351),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_432),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_421),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_422),
.B(n_339),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_379),
.Y(n_479)
);

BUFx12f_ASAP7_75t_L g480 ( 
.A(n_382),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_440),
.B(n_339),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_417),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_418),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_427),
.B(n_401),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_379),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_401),
.B(n_351),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_434),
.Y(n_487)
);

INVx4_ASAP7_75t_L g488 ( 
.A(n_420),
.Y(n_488)
);

INVx6_ASAP7_75t_L g489 ( 
.A(n_418),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_430),
.B(n_220),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_429),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_410),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_377),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_404),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_396),
.B(n_366),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_410),
.B(n_311),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_373),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_414),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_407),
.A2(n_344),
.B1(n_328),
.B2(n_336),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_441),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_431),
.B(n_366),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_424),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_397),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_413),
.B(n_344),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_398),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_413),
.B(n_336),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_426),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_402),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_437),
.Y(n_509)
);

AND2x2_ASAP7_75t_SL g510 ( 
.A(n_394),
.B(n_336),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_438),
.B(n_361),
.Y(n_511)
);

INVx5_ASAP7_75t_L g512 ( 
.A(n_426),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_419),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_383),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_389),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_405),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_403),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_403),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_435),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_406),
.Y(n_520)
);

NAND2xp33_ASAP7_75t_R g521 ( 
.A(n_412),
.B(n_2),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_435),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_433),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_443),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_445),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_415),
.B(n_221),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_391),
.Y(n_527)
);

BUFx4f_ASAP7_75t_L g528 ( 
.A(n_384),
.Y(n_528)
);

OAI22xp33_ASAP7_75t_L g529 ( 
.A1(n_393),
.A2(n_328),
.B1(n_345),
.B2(n_346),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_391),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_447),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_448),
.Y(n_532)
);

A2O1A1Ixp33_ASAP7_75t_L g533 ( 
.A1(n_465),
.A2(n_345),
.B(n_346),
.C(n_329),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_528),
.B(n_389),
.Y(n_534)
);

BUFx8_ASAP7_75t_L g535 ( 
.A(n_513),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_486),
.B(n_458),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_518),
.B(n_385),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_459),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_452),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_522),
.B(n_388),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_487),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_472),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_453),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_522),
.B(n_329),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_473),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g546 ( 
.A(n_450),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_446),
.B(n_372),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_491),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_510),
.A2(n_343),
.B1(n_354),
.B2(n_340),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_455),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_471),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_510),
.A2(n_343),
.B1(n_354),
.B2(n_340),
.Y(n_552)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_446),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_486),
.B(n_361),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_476),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_522),
.B(n_343),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_504),
.B(n_372),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_478),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_495),
.B(n_358),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_481),
.B(n_343),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_458),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_478),
.Y(n_562)
);

NOR2xp67_ASAP7_75t_L g563 ( 
.A(n_460),
.B(n_512),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_503),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_481),
.Y(n_565)
);

A2O1A1Ixp33_ASAP7_75t_L g566 ( 
.A1(n_465),
.A2(n_222),
.B(n_227),
.C(n_246),
.Y(n_566)
);

BUFx8_ASAP7_75t_L g567 ( 
.A(n_480),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g568 ( 
.A1(n_505),
.A2(n_386),
.B1(n_384),
.B2(n_247),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_528),
.B(n_230),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_449),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_449),
.Y(n_571)
);

AND2x6_ASAP7_75t_L g572 ( 
.A(n_506),
.B(n_361),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_518),
.B(n_275),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_516),
.B(n_238),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_495),
.B(n_359),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_507),
.B(n_343),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_494),
.Y(n_577)
);

AO22x2_ASAP7_75t_L g578 ( 
.A1(n_499),
.A2(n_386),
.B1(n_3),
.B2(n_4),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_494),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_482),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_477),
.Y(n_581)
);

AO22x2_ASAP7_75t_L g582 ( 
.A1(n_499),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_582)
);

NAND3xp33_ASAP7_75t_L g583 ( 
.A(n_456),
.B(n_242),
.C(n_240),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_454),
.B(n_501),
.Y(n_584)
);

NAND2x1p5_ASAP7_75t_L g585 ( 
.A(n_483),
.B(n_321),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_451),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_462),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_464),
.Y(n_588)
);

AND2x6_ASAP7_75t_L g589 ( 
.A(n_483),
.B(n_361),
.Y(n_589)
);

A2O1A1Ixp33_ASAP7_75t_L g590 ( 
.A1(n_501),
.A2(n_243),
.B(n_245),
.C(n_248),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_511),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_467),
.B(n_456),
.Y(n_592)
);

BUFx4f_ASAP7_75t_L g593 ( 
.A(n_527),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_520),
.A2(n_529),
.B1(n_484),
.B2(n_508),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_517),
.B(n_321),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_493),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_500),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_492),
.B(n_321),
.Y(n_598)
);

AOI21x1_ASAP7_75t_L g599 ( 
.A1(n_563),
.A2(n_469),
.B(n_502),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_584),
.B(n_511),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_591),
.B(n_529),
.Y(n_601)
);

CKINVDCx16_ASAP7_75t_R g602 ( 
.A(n_580),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_SL g603 ( 
.A(n_593),
.B(n_488),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_536),
.A2(n_469),
.B(n_457),
.Y(n_604)
);

INVxp67_ASAP7_75t_SL g605 ( 
.A(n_536),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_553),
.A2(n_467),
.B1(n_484),
.B2(n_489),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_593),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g608 ( 
.A(n_541),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_546),
.B(n_474),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_554),
.A2(n_457),
.B(n_523),
.Y(n_610)
);

AND2x4_ASAP7_75t_SL g611 ( 
.A(n_540),
.B(n_483),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_L g612 ( 
.A1(n_582),
.A2(n_467),
.B1(n_489),
.B2(n_527),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_542),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_546),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_570),
.B(n_470),
.Y(n_615)
);

O2A1O1Ixp33_ASAP7_75t_L g616 ( 
.A1(n_594),
.A2(n_470),
.B(n_526),
.C(n_490),
.Y(n_616)
);

OA22x2_ASAP7_75t_L g617 ( 
.A1(n_594),
.A2(n_548),
.B1(n_564),
.B2(n_565),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_571),
.B(n_463),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_561),
.B(n_463),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_557),
.B(n_483),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_535),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_554),
.A2(n_457),
.B(n_523),
.Y(n_622)
);

AO22x1_ASAP7_75t_L g623 ( 
.A1(n_547),
.A2(n_496),
.B1(n_466),
.B2(n_515),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_531),
.Y(n_624)
);

NAND3xp33_ASAP7_75t_L g625 ( 
.A(n_574),
.B(n_526),
.C(n_490),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_592),
.A2(n_457),
.B(n_461),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_L g627 ( 
.A1(n_549),
.A2(n_498),
.B(n_485),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_592),
.A2(n_461),
.B(n_559),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_532),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_598),
.B(n_488),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_539),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_575),
.A2(n_512),
.B(n_479),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_543),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_550),
.B(n_519),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_563),
.A2(n_512),
.B(n_338),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_558),
.B(n_527),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_545),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_552),
.A2(n_512),
.B(n_338),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_551),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_555),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_562),
.A2(n_530),
.B1(n_509),
.B2(n_525),
.Y(n_641)
);

AOI22x1_ASAP7_75t_L g642 ( 
.A1(n_586),
.A2(n_509),
.B1(n_527),
.B2(n_524),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_568),
.B(n_524),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_L g644 ( 
.A1(n_533),
.A2(n_475),
.B(n_354),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_560),
.A2(n_338),
.B(n_330),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_560),
.A2(n_489),
.B1(n_524),
.B2(n_525),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_556),
.A2(n_338),
.B(n_330),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_535),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_595),
.B(n_525),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_537),
.B(n_497),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_577),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_568),
.B(n_468),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_556),
.A2(n_576),
.B(n_583),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_589),
.Y(n_654)
);

CKINVDCx8_ASAP7_75t_R g655 ( 
.A(n_538),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_544),
.B(n_468),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_576),
.A2(n_338),
.B(n_330),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_579),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_583),
.A2(n_597),
.B1(n_596),
.B2(n_588),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_581),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_544),
.A2(n_338),
.B(n_330),
.Y(n_661)
);

OA22x2_ASAP7_75t_L g662 ( 
.A1(n_540),
.A2(n_521),
.B1(n_468),
.B2(n_514),
.Y(n_662)
);

NAND2x1p5_ASAP7_75t_L g663 ( 
.A(n_587),
.B(n_323),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_578),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_569),
.A2(n_330),
.B(n_359),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_605),
.B(n_573),
.Y(n_666)
);

OAI21xp33_ASAP7_75t_SL g667 ( 
.A1(n_617),
.A2(n_534),
.B(n_578),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_624),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_655),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_650),
.B(n_590),
.Y(n_670)
);

CKINVDCx8_ASAP7_75t_R g671 ( 
.A(n_602),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_609),
.B(n_566),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_600),
.B(n_572),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_630),
.B(n_582),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_614),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_629),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_631),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_649),
.B(n_585),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_608),
.B(n_567),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_607),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_625),
.B(n_567),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_625),
.A2(n_572),
.B1(n_475),
.B2(n_589),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_604),
.A2(n_572),
.B(n_359),
.Y(n_683)
);

NOR3xp33_ASAP7_75t_L g684 ( 
.A(n_623),
.B(n_521),
.C(n_256),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_662),
.B(n_323),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_603),
.B(n_251),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_601),
.B(n_572),
.Y(n_687)
);

O2A1O1Ixp33_ASAP7_75t_L g688 ( 
.A1(n_616),
.A2(n_322),
.B(n_323),
.C(n_326),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_615),
.B(n_589),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_648),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_618),
.B(n_589),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_603),
.B(n_340),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_610),
.A2(n_365),
.B(n_326),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_607),
.B(n_340),
.Y(n_694)
);

O2A1O1Ixp33_ASAP7_75t_L g695 ( 
.A1(n_643),
.A2(n_322),
.B(n_365),
.C(n_8),
.Y(n_695)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_622),
.A2(n_365),
.B(n_340),
.Y(n_696)
);

OR2x6_ASAP7_75t_L g697 ( 
.A(n_607),
.B(n_365),
.Y(n_697)
);

INVx4_ASAP7_75t_L g698 ( 
.A(n_611),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_656),
.Y(n_699)
);

O2A1O1Ixp33_ASAP7_75t_L g700 ( 
.A1(n_606),
.A2(n_5),
.B(n_7),
.C(n_8),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_633),
.B(n_475),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_654),
.Y(n_702)
);

NOR3xp33_ASAP7_75t_L g703 ( 
.A(n_646),
.B(n_475),
.C(n_354),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_639),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_653),
.A2(n_354),
.B(n_343),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_628),
.A2(n_354),
.B(n_343),
.Y(n_706)
);

AOI21xp33_ASAP7_75t_L g707 ( 
.A1(n_659),
.A2(n_7),
.B(n_9),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_654),
.Y(n_708)
);

NOR3xp33_ASAP7_75t_SL g709 ( 
.A(n_652),
.B(n_9),
.C(n_10),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_640),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_634),
.B(n_475),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_619),
.A2(n_354),
.B1(n_11),
.B2(n_12),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_613),
.Y(n_713)
);

INVx3_ASAP7_75t_SL g714 ( 
.A(n_620),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_637),
.Y(n_715)
);

OAI21x1_ASAP7_75t_SL g716 ( 
.A1(n_612),
.A2(n_36),
.B(n_35),
.Y(n_716)
);

O2A1O1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_612),
.A2(n_10),
.B(n_11),
.C(n_13),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_660),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_651),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_658),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_638),
.A2(n_40),
.B(n_37),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_641),
.B(n_13),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_664),
.B(n_14),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_663),
.Y(n_724)
);

A2O1A1Ixp33_ASAP7_75t_L g725 ( 
.A1(n_632),
.A2(n_15),
.B(n_16),
.C(n_18),
.Y(n_725)
);

INVx1_ASAP7_75t_SL g726 ( 
.A(n_675),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_671),
.Y(n_727)
);

BUFx2_ASAP7_75t_R g728 ( 
.A(n_669),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_704),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_722),
.A2(n_642),
.B1(n_636),
.B2(n_621),
.Y(n_730)
);

NAND2x1p5_ASAP7_75t_L g731 ( 
.A(n_698),
.B(n_626),
.Y(n_731)
);

INVx5_ASAP7_75t_L g732 ( 
.A(n_680),
.Y(n_732)
);

INVx5_ASAP7_75t_L g733 ( 
.A(n_680),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_698),
.B(n_680),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_690),
.Y(n_735)
);

INVx1_ASAP7_75t_SL g736 ( 
.A(n_699),
.Y(n_736)
);

INVx3_ASAP7_75t_SL g737 ( 
.A(n_681),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_670),
.B(n_663),
.Y(n_738)
);

INVx4_ASAP7_75t_L g739 ( 
.A(n_697),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_713),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_702),
.Y(n_741)
);

INVx3_ASAP7_75t_SL g742 ( 
.A(n_699),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_699),
.Y(n_743)
);

NOR2x1_ASAP7_75t_L g744 ( 
.A(n_666),
.B(n_627),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_679),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_720),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_668),
.Y(n_747)
);

INVx8_ASAP7_75t_L g748 ( 
.A(n_697),
.Y(n_748)
);

INVx5_ASAP7_75t_L g749 ( 
.A(n_702),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_714),
.Y(n_750)
);

BUFx12f_ASAP7_75t_L g751 ( 
.A(n_685),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_702),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_708),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_L g754 ( 
.A1(n_674),
.A2(n_687),
.B1(n_689),
.B2(n_678),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_718),
.Y(n_755)
);

INVx1_ASAP7_75t_SL g756 ( 
.A(n_676),
.Y(n_756)
);

INVx5_ASAP7_75t_L g757 ( 
.A(n_708),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_677),
.Y(n_758)
);

BUFx4_ASAP7_75t_SL g759 ( 
.A(n_710),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_719),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_709),
.B(n_627),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_708),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_715),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_723),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_724),
.Y(n_765)
);

INVx4_ASAP7_75t_L g766 ( 
.A(n_716),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_684),
.B(n_599),
.Y(n_767)
);

BUFx4_ASAP7_75t_SL g768 ( 
.A(n_667),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_688),
.Y(n_769)
);

CKINVDCx20_ASAP7_75t_R g770 ( 
.A(n_686),
.Y(n_770)
);

BUFx2_ASAP7_75t_L g771 ( 
.A(n_691),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_672),
.B(n_694),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_673),
.B(n_665),
.Y(n_773)
);

BUFx2_ASAP7_75t_SL g774 ( 
.A(n_692),
.Y(n_774)
);

CKINVDCx8_ASAP7_75t_R g775 ( 
.A(n_711),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_701),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_717),
.Y(n_777)
);

INVxp67_ASAP7_75t_SL g778 ( 
.A(n_695),
.Y(n_778)
);

INVx1_ASAP7_75t_SL g779 ( 
.A(n_707),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_700),
.B(n_635),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_725),
.B(n_16),
.Y(n_781)
);

INVx1_ASAP7_75t_SL g782 ( 
.A(n_712),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_682),
.B(n_705),
.Y(n_783)
);

NAND2x1p5_ASAP7_75t_L g784 ( 
.A(n_721),
.B(n_683),
.Y(n_784)
);

BUFx12f_ASAP7_75t_L g785 ( 
.A(n_703),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_693),
.Y(n_786)
);

BUFx2_ASAP7_75t_SL g787 ( 
.A(n_706),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_696),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_722),
.A2(n_644),
.B1(n_661),
.B2(n_657),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_680),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_680),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_704),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_680),
.Y(n_793)
);

NAND2x1p5_ASAP7_75t_L g794 ( 
.A(n_698),
.B(n_647),
.Y(n_794)
);

INVxp67_ASAP7_75t_L g795 ( 
.A(n_675),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_680),
.Y(n_796)
);

OAI21x1_ASAP7_75t_L g797 ( 
.A1(n_784),
.A2(n_644),
.B(n_645),
.Y(n_797)
);

AO21x2_ASAP7_75t_L g798 ( 
.A1(n_786),
.A2(n_18),
.B(n_19),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_786),
.A2(n_42),
.B(n_41),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_758),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_771),
.Y(n_801)
);

OAI21x1_ASAP7_75t_SL g802 ( 
.A1(n_781),
.A2(n_19),
.B(n_20),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_764),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_L g804 ( 
.A1(n_779),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_749),
.Y(n_805)
);

CKINVDCx6p67_ASAP7_75t_R g806 ( 
.A(n_735),
.Y(n_806)
);

OAI21x1_ASAP7_75t_L g807 ( 
.A1(n_773),
.A2(n_45),
.B(n_44),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_750),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_793),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_743),
.B(n_47),
.Y(n_810)
);

NOR2x1_ASAP7_75t_SL g811 ( 
.A(n_774),
.B(n_48),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_754),
.B(n_25),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_740),
.Y(n_813)
);

BUFx4f_ASAP7_75t_L g814 ( 
.A(n_742),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_747),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_744),
.B(n_26),
.Y(n_816)
);

OAI21x1_ASAP7_75t_L g817 ( 
.A1(n_783),
.A2(n_138),
.B(n_193),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_736),
.B(n_49),
.Y(n_818)
);

OAI21x1_ASAP7_75t_L g819 ( 
.A1(n_731),
.A2(n_139),
.B(n_192),
.Y(n_819)
);

OAI21x1_ASAP7_75t_L g820 ( 
.A1(n_780),
.A2(n_137),
.B(n_189),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_756),
.B(n_755),
.Y(n_821)
);

BUFx12f_ASAP7_75t_L g822 ( 
.A(n_793),
.Y(n_822)
);

OAI21x1_ASAP7_75t_L g823 ( 
.A1(n_769),
.A2(n_136),
.B(n_187),
.Y(n_823)
);

OA21x2_ASAP7_75t_L g824 ( 
.A1(n_769),
.A2(n_789),
.B(n_767),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_760),
.Y(n_825)
);

OAI21x1_ASAP7_75t_L g826 ( 
.A1(n_794),
.A2(n_135),
.B(n_186),
.Y(n_826)
);

OAI21x1_ASAP7_75t_L g827 ( 
.A1(n_760),
.A2(n_134),
.B(n_185),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_751),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_738),
.A2(n_788),
.B(n_767),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_729),
.Y(n_830)
);

OAI22xp33_ASAP7_75t_L g831 ( 
.A1(n_777),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_831)
);

AOI21x1_ASAP7_75t_L g832 ( 
.A1(n_761),
.A2(n_133),
.B(n_184),
.Y(n_832)
);

OAI21xp5_ASAP7_75t_L g833 ( 
.A1(n_778),
.A2(n_27),
.B(n_28),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_772),
.B(n_51),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_777),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_772),
.B(n_56),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_727),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_776),
.B(n_57),
.Y(n_838)
);

AOI21x1_ASAP7_75t_L g839 ( 
.A1(n_792),
.A2(n_765),
.B(n_734),
.Y(n_839)
);

BUFx2_ASAP7_75t_L g840 ( 
.A(n_793),
.Y(n_840)
);

BUFx12f_ASAP7_75t_L g841 ( 
.A(n_734),
.Y(n_841)
);

BUFx2_ASAP7_75t_SL g842 ( 
.A(n_732),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_763),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_741),
.Y(n_844)
);

BUFx3_ASAP7_75t_L g845 ( 
.A(n_732),
.Y(n_845)
);

OAI21xp33_ASAP7_75t_SL g846 ( 
.A1(n_766),
.A2(n_58),
.B(n_59),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_777),
.A2(n_195),
.B1(n_64),
.B2(n_65),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_787),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_770),
.A2(n_62),
.B1(n_66),
.B2(n_68),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_741),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_752),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_732),
.B(n_69),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_782),
.B(n_70),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_737),
.A2(n_182),
.B1(n_72),
.B2(n_73),
.Y(n_854)
);

NAND2x1_ASAP7_75t_L g855 ( 
.A(n_766),
.B(n_71),
.Y(n_855)
);

OAI221xp5_ASAP7_75t_L g856 ( 
.A1(n_730),
.A2(n_74),
.B1(n_76),
.B2(n_82),
.C(n_83),
.Y(n_856)
);

OAI21x1_ASAP7_75t_L g857 ( 
.A1(n_787),
.A2(n_84),
.B(n_85),
.Y(n_857)
);

OA21x2_ASAP7_75t_L g858 ( 
.A1(n_795),
.A2(n_86),
.B(n_88),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_774),
.B(n_90),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_825),
.Y(n_860)
);

BUFx2_ASAP7_75t_L g861 ( 
.A(n_848),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_801),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_839),
.Y(n_863)
);

OAI21x1_ASAP7_75t_L g864 ( 
.A1(n_797),
.A2(n_752),
.B(n_753),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_801),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_815),
.Y(n_866)
);

NAND2x1p5_ASAP7_75t_L g867 ( 
.A(n_824),
.B(n_749),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_806),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_830),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_845),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_848),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_824),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_845),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_812),
.A2(n_785),
.B1(n_745),
.B2(n_739),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_800),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_829),
.B(n_775),
.Y(n_876)
);

CKINVDCx20_ASAP7_75t_R g877 ( 
.A(n_808),
.Y(n_877)
);

AO21x2_ASAP7_75t_L g878 ( 
.A1(n_829),
.A2(n_768),
.B(n_739),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_813),
.Y(n_879)
);

AO21x1_ASAP7_75t_SL g880 ( 
.A1(n_833),
.A2(n_759),
.B(n_733),
.Y(n_880)
);

BUFx12f_ASAP7_75t_L g881 ( 
.A(n_822),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_798),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_833),
.B(n_726),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_821),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_798),
.Y(n_885)
);

AO21x2_ASAP7_75t_L g886 ( 
.A1(n_799),
.A2(n_733),
.B(n_749),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_812),
.B(n_746),
.Y(n_887)
);

CKINVDCx20_ASAP7_75t_R g888 ( 
.A(n_837),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_816),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_816),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_843),
.Y(n_891)
);

OAI22xp33_ASAP7_75t_L g892 ( 
.A1(n_803),
.A2(n_748),
.B1(n_733),
.B2(n_757),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_814),
.B(n_853),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_858),
.Y(n_894)
);

OAI21x1_ASAP7_75t_L g895 ( 
.A1(n_820),
.A2(n_762),
.B(n_753),
.Y(n_895)
);

BUFx12f_ASAP7_75t_L g896 ( 
.A(n_828),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_844),
.B(n_762),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_858),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_840),
.Y(n_899)
);

AO21x2_ASAP7_75t_L g900 ( 
.A1(n_799),
.A2(n_757),
.B(n_748),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_807),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_850),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_851),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_827),
.Y(n_904)
);

AOI21x1_ASAP7_75t_L g905 ( 
.A1(n_832),
.A2(n_859),
.B(n_855),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_823),
.Y(n_906)
);

OAI22xp33_ASAP7_75t_L g907 ( 
.A1(n_856),
.A2(n_757),
.B1(n_791),
.B2(n_790),
.Y(n_907)
);

OA21x2_ASAP7_75t_L g908 ( 
.A1(n_817),
.A2(n_796),
.B(n_92),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_857),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_834),
.B(n_91),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_856),
.A2(n_728),
.B(n_94),
.Y(n_911)
);

NAND2xp33_ASAP7_75t_R g912 ( 
.A(n_868),
.B(n_838),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_896),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_889),
.B(n_831),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_875),
.Y(n_915)
);

AND2x2_ASAP7_75t_SL g916 ( 
.A(n_884),
.B(n_814),
.Y(n_916)
);

AO31x2_ASAP7_75t_L g917 ( 
.A1(n_882),
.A2(n_811),
.A3(n_835),
.B(n_804),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_861),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_870),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_870),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_861),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_866),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_889),
.B(n_831),
.Y(n_923)
);

NAND2xp33_ASAP7_75t_R g924 ( 
.A(n_884),
.B(n_852),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_871),
.Y(n_925)
);

OR2x2_ASAP7_75t_L g926 ( 
.A(n_871),
.B(n_834),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_875),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_890),
.B(n_804),
.Y(n_928)
);

NAND2xp33_ASAP7_75t_R g929 ( 
.A(n_887),
.B(n_852),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_890),
.B(n_862),
.Y(n_930)
);

OA222x2_ASAP7_75t_L g931 ( 
.A1(n_872),
.A2(n_859),
.B1(n_836),
.B2(n_805),
.C1(n_853),
.C2(n_854),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_899),
.B(n_809),
.Y(n_932)
);

INVx3_ASAP7_75t_SL g933 ( 
.A(n_888),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_865),
.B(n_805),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_866),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_875),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_879),
.Y(n_937)
);

OR2x6_ASAP7_75t_L g938 ( 
.A(n_867),
.B(n_842),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_869),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_869),
.B(n_836),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_860),
.B(n_802),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_899),
.B(n_809),
.Y(n_942)
);

AND2x6_ASAP7_75t_L g943 ( 
.A(n_872),
.B(n_810),
.Y(n_943)
);

INVx8_ASAP7_75t_L g944 ( 
.A(n_881),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_915),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_933),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_918),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_938),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_925),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_927),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_925),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_918),
.B(n_872),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_921),
.B(n_872),
.Y(n_953)
);

NOR2x1_ASAP7_75t_SL g954 ( 
.A(n_938),
.B(n_878),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_936),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_921),
.B(n_867),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_934),
.B(n_867),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_942),
.B(n_894),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_944),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_930),
.B(n_891),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_919),
.B(n_894),
.Y(n_961)
);

OR2x2_ASAP7_75t_L g962 ( 
.A(n_930),
.B(n_882),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_926),
.B(n_902),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_937),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_940),
.B(n_879),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_919),
.B(n_920),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_920),
.B(n_898),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_957),
.B(n_916),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_949),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_949),
.Y(n_970)
);

NAND3xp33_ASAP7_75t_L g971 ( 
.A(n_960),
.B(n_883),
.C(n_911),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_956),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_959),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_954),
.A2(n_876),
.B(n_907),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_951),
.B(n_922),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_963),
.B(n_940),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_946),
.B(n_913),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_956),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_947),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_957),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_948),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_954),
.A2(n_893),
.B(n_878),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_948),
.A2(n_878),
.B(n_914),
.Y(n_983)
);

NOR3xp33_ASAP7_75t_L g984 ( 
.A(n_959),
.B(n_928),
.C(n_923),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_968),
.B(n_958),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_975),
.Y(n_986)
);

AOI211xp5_ASAP7_75t_L g987 ( 
.A1(n_971),
.A2(n_892),
.B(n_931),
.C(n_923),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_981),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_975),
.Y(n_989)
);

OR2x2_ASAP7_75t_L g990 ( 
.A(n_976),
.B(n_962),
.Y(n_990)
);

INVx3_ASAP7_75t_L g991 ( 
.A(n_973),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_969),
.Y(n_992)
);

AO21x2_ASAP7_75t_L g993 ( 
.A1(n_983),
.A2(n_951),
.B(n_952),
.Y(n_993)
);

NAND4xp25_ASAP7_75t_L g994 ( 
.A(n_971),
.B(n_874),
.C(n_928),
.D(n_914),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_970),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_979),
.B(n_962),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_985),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_991),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_992),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_991),
.B(n_977),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_987),
.B(n_974),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_988),
.B(n_984),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_995),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_990),
.B(n_972),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_997),
.B(n_1002),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_999),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_1003),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_1000),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_998),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_1000),
.Y(n_1010)
);

INVx1_ASAP7_75t_SL g1011 ( 
.A(n_1010),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_1006),
.Y(n_1012)
);

AOI33xp33_ASAP7_75t_L g1013 ( 
.A1(n_1009),
.A2(n_987),
.A3(n_1001),
.B1(n_997),
.B2(n_986),
.B3(n_989),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_1007),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_1010),
.Y(n_1015)
);

OR2x6_ASAP7_75t_L g1016 ( 
.A(n_1008),
.B(n_944),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1005),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1006),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_1006),
.Y(n_1019)
);

OR2x2_ASAP7_75t_L g1020 ( 
.A(n_1005),
.B(n_1001),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_1011),
.B(n_1004),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_1013),
.B(n_993),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_1016),
.B(n_973),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1017),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_1016),
.B(n_973),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1015),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1012),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1014),
.Y(n_1028)
);

NOR3xp33_ASAP7_75t_L g1029 ( 
.A(n_1024),
.B(n_1020),
.C(n_1019),
.Y(n_1029)
);

OR2x2_ASAP7_75t_L g1030 ( 
.A(n_1026),
.B(n_1018),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_1021),
.B(n_994),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_1023),
.B(n_913),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1022),
.B(n_994),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1022),
.B(n_993),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1027),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_1025),
.B(n_944),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_SL g1037 ( 
.A(n_1036),
.B(n_1028),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1029),
.B(n_996),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1030),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_1031),
.B(n_1033),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_1032),
.A2(n_912),
.B1(n_896),
.B2(n_913),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1035),
.B(n_978),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1039),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1038),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1042),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1040),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_1041),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_1037),
.B(n_1034),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_1039),
.B(n_980),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_1039),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1039),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_1051),
.B(n_877),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_1049),
.B(n_896),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_1048),
.A2(n_835),
.B(n_982),
.C(n_854),
.Y(n_1054)
);

NOR3xp33_ASAP7_75t_L g1055 ( 
.A(n_1044),
.B(n_910),
.C(n_818),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_1043),
.A2(n_941),
.B(n_910),
.Y(n_1056)
);

NAND3xp33_ASAP7_75t_L g1057 ( 
.A(n_1043),
.B(n_1050),
.C(n_1047),
.Y(n_1057)
);

NOR3xp33_ASAP7_75t_L g1058 ( 
.A(n_1046),
.B(n_849),
.C(n_941),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_1045),
.B(n_881),
.Y(n_1059)
);

AOI31xp33_ASAP7_75t_L g1060 ( 
.A1(n_1044),
.A2(n_847),
.A3(n_929),
.B(n_924),
.Y(n_1060)
);

OAI221xp5_ASAP7_75t_L g1061 ( 
.A1(n_1057),
.A2(n_847),
.B1(n_938),
.B2(n_846),
.C(n_870),
.Y(n_1061)
);

AOI222xp33_ASAP7_75t_L g1062 ( 
.A1(n_1059),
.A2(n_881),
.B1(n_885),
.B2(n_898),
.C1(n_953),
.C2(n_952),
.Y(n_1062)
);

OAI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_1052),
.A2(n_810),
.B(n_819),
.Y(n_1063)
);

AOI221xp5_ASAP7_75t_L g1064 ( 
.A1(n_1053),
.A2(n_885),
.B1(n_953),
.B2(n_961),
.C(n_967),
.Y(n_1064)
);

OAI211xp5_ASAP7_75t_SL g1065 ( 
.A1(n_1054),
.A2(n_880),
.B(n_901),
.C(n_965),
.Y(n_1065)
);

AOI221xp5_ASAP7_75t_L g1066 ( 
.A1(n_1056),
.A2(n_1058),
.B1(n_1060),
.B2(n_1055),
.C(n_967),
.Y(n_1066)
);

OAI211xp5_ASAP7_75t_L g1067 ( 
.A1(n_1057),
.A2(n_826),
.B(n_961),
.C(n_873),
.Y(n_1067)
);

AOI221xp5_ASAP7_75t_L g1068 ( 
.A1(n_1066),
.A2(n_966),
.B1(n_958),
.B2(n_873),
.C(n_955),
.Y(n_1068)
);

NOR3xp33_ASAP7_75t_L g1069 ( 
.A(n_1065),
.B(n_905),
.C(n_901),
.Y(n_1069)
);

AOI221x1_ASAP7_75t_L g1070 ( 
.A1(n_1063),
.A2(n_966),
.B1(n_809),
.B2(n_932),
.C(n_903),
.Y(n_1070)
);

OAI221xp5_ASAP7_75t_SL g1071 ( 
.A1(n_1067),
.A2(n_873),
.B1(n_880),
.B2(n_899),
.C(n_945),
.Y(n_1071)
);

NAND4xp75_ASAP7_75t_L g1072 ( 
.A(n_1064),
.B(n_908),
.C(n_897),
.D(n_903),
.Y(n_1072)
);

AOI211x1_ASAP7_75t_SL g1073 ( 
.A1(n_1062),
.A2(n_964),
.B(n_955),
.C(n_950),
.Y(n_1073)
);

AOI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_1061),
.A2(n_841),
.B1(n_932),
.B2(n_900),
.Y(n_1074)
);

AOI21xp33_ASAP7_75t_L g1075 ( 
.A1(n_1067),
.A2(n_901),
.B(n_900),
.Y(n_1075)
);

OAI221xp5_ASAP7_75t_L g1076 ( 
.A1(n_1066),
.A2(n_905),
.B1(n_908),
.B2(n_906),
.C(n_863),
.Y(n_1076)
);

XNOR2xp5_ASAP7_75t_L g1077 ( 
.A(n_1066),
.B(n_93),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1077),
.B(n_917),
.Y(n_1078)
);

AOI211xp5_ASAP7_75t_SL g1079 ( 
.A1(n_1071),
.A2(n_863),
.B(n_906),
.C(n_897),
.Y(n_1079)
);

OAI321xp33_ASAP7_75t_L g1080 ( 
.A1(n_1074),
.A2(n_809),
.A3(n_935),
.B1(n_939),
.B2(n_909),
.C(n_904),
.Y(n_1080)
);

NOR4xp75_ASAP7_75t_L g1081 ( 
.A(n_1076),
.B(n_863),
.C(n_906),
.D(n_100),
.Y(n_1081)
);

NAND4xp75_ASAP7_75t_L g1082 ( 
.A(n_1070),
.B(n_908),
.C(n_98),
.D(n_104),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_1069),
.B(n_917),
.Y(n_1083)
);

NOR3xp33_ASAP7_75t_L g1084 ( 
.A(n_1068),
.B(n_906),
.C(n_895),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1075),
.B(n_945),
.Y(n_1085)
);

NAND2xp33_ASAP7_75t_SL g1086 ( 
.A(n_1073),
.B(n_900),
.Y(n_1086)
);

AOI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_1072),
.A2(n_943),
.B1(n_886),
.B2(n_964),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1077),
.B(n_917),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1078),
.Y(n_1089)
);

NAND3x1_ASAP7_75t_SL g1090 ( 
.A(n_1085),
.B(n_95),
.C(n_107),
.Y(n_1090)
);

XNOR2xp5_ASAP7_75t_L g1091 ( 
.A(n_1081),
.B(n_108),
.Y(n_1091)
);

NAND2x1p5_ASAP7_75t_L g1092 ( 
.A(n_1083),
.B(n_908),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_1088),
.B(n_1084),
.Y(n_1093)
);

NOR4xp75_ASAP7_75t_L g1094 ( 
.A(n_1082),
.B(n_863),
.C(n_110),
.D(n_111),
.Y(n_1094)
);

OAI211xp5_ASAP7_75t_SL g1095 ( 
.A1(n_1079),
.A2(n_109),
.B(n_112),
.C(n_113),
.Y(n_1095)
);

NOR3xp33_ASAP7_75t_SL g1096 ( 
.A(n_1086),
.B(n_114),
.C(n_116),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_1087),
.B(n_950),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1080),
.B(n_886),
.Y(n_1098)
);

NOR3x1_ASAP7_75t_L g1099 ( 
.A(n_1078),
.B(n_895),
.C(n_118),
.Y(n_1099)
);

NOR4xp25_ASAP7_75t_L g1100 ( 
.A(n_1078),
.B(n_909),
.C(n_904),
.D(n_122),
.Y(n_1100)
);

NOR2x1p5_ASAP7_75t_L g1101 ( 
.A(n_1082),
.B(n_909),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1091),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_SL g1103 ( 
.A1(n_1089),
.A2(n_904),
.B1(n_879),
.B2(n_860),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_1096),
.Y(n_1104)
);

INVx1_ASAP7_75t_SL g1105 ( 
.A(n_1094),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_1101),
.B(n_886),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_1093),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1090),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1099),
.B(n_943),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_1097),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_1108),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1110),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1105),
.A2(n_1095),
.B1(n_1098),
.B2(n_1100),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1104),
.A2(n_1092),
.B1(n_860),
.B2(n_943),
.Y(n_1114)
);

XNOR2xp5_ASAP7_75t_L g1115 ( 
.A(n_1102),
.B(n_117),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1106),
.A2(n_1109),
.B(n_1107),
.Y(n_1116)
);

XNOR2x1_ASAP7_75t_L g1117 ( 
.A(n_1107),
.B(n_120),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1112),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1115),
.B(n_1103),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1117),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1118),
.Y(n_1121)
);

NOR2x1_ASAP7_75t_L g1122 ( 
.A(n_1121),
.B(n_1111),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_SL g1123 ( 
.A1(n_1122),
.A2(n_1116),
.B1(n_1120),
.B2(n_1113),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1123),
.A2(n_1119),
.B1(n_1114),
.B2(n_943),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1123),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_1123),
.A2(n_943),
.B1(n_864),
.B2(n_126),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1125),
.A2(n_123),
.B(n_125),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1124),
.A2(n_127),
.B1(n_131),
.B2(n_132),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1126),
.A2(n_140),
.B(n_141),
.Y(n_1129)
);

AOI222xp33_ASAP7_75t_SL g1130 ( 
.A1(n_1125),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.C1(n_146),
.C2(n_147),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_R g1131 ( 
.A1(n_1128),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1130),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1129),
.A2(n_154),
.B1(n_156),
.B2(n_157),
.Y(n_1133)
);

AOI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1127),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_1134)
);

AO21x2_ASAP7_75t_L g1135 ( 
.A1(n_1132),
.A2(n_161),
.B(n_162),
.Y(n_1135)
);

OA21x2_ASAP7_75t_L g1136 ( 
.A1(n_1134),
.A2(n_163),
.B(n_167),
.Y(n_1136)
);

AOI221xp5_ASAP7_75t_L g1137 ( 
.A1(n_1135),
.A2(n_1133),
.B1(n_1131),
.B2(n_172),
.C(n_173),
.Y(n_1137)
);

AOI211xp5_ASAP7_75t_L g1138 ( 
.A1(n_1137),
.A2(n_1136),
.B(n_170),
.C(n_174),
.Y(n_1138)
);


endmodule