module fake_jpeg_11964_n_105 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_105);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVxp67_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_52),
.Y(n_58)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_48)
);

NOR2x1_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_38),
.Y(n_60)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NAND2xp33_ASAP7_75t_SL g56 ( 
.A(n_50),
.B(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_46),
.B(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_5),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_60),
.B(n_8),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_61),
.Y(n_64)
);

OR2x2_ASAP7_75t_SL g62 ( 
.A(n_49),
.B(n_32),
.Y(n_62)
);

OR2x4_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_0),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_32),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_11),
.Y(n_76)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_38),
.B1(n_42),
.B2(n_4),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_76),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_42),
.B1(n_1),
.B2(n_4),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_71),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_55),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_72),
.C(n_19),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_70),
.B(n_73),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_59),
.B1(n_62),
.B2(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_9),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_75),
.Y(n_83)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_12),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_84),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_15),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_16),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_86),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_20),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_31),
.Y(n_95)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_90),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_93),
.A2(n_89),
.B(n_79),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_24),
.B(n_27),
.C(n_29),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_94),
.B(n_95),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_91),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_100),
.C(n_78),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_92),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_97),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_102),
.B(n_83),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_103),
.A2(n_80),
.B(n_90),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_88),
.Y(n_105)
);


endmodule