module fake_jpeg_5648_n_327 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_327);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_30),
.B(n_35),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_31),
.A2(n_26),
.B1(n_18),
.B2(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_6),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_26),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_12),
.Y(n_51)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_30),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_31),
.A2(n_13),
.B1(n_20),
.B2(n_27),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_45),
.A2(n_52),
.B1(n_22),
.B2(n_21),
.Y(n_78)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_51),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_31),
.A2(n_13),
.B1(n_20),
.B2(n_27),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_14),
.B1(n_18),
.B2(n_19),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_15),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_35),
.B1(n_30),
.B2(n_13),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_58),
.A2(n_22),
.B1(n_21),
.B2(n_17),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_48),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_64),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_33),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_69),
.Y(n_91)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_36),
.B1(n_35),
.B2(n_15),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_70),
.B1(n_43),
.B2(n_41),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_66),
.B(n_41),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_24),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_32),
.B(n_28),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_56),
.B(n_49),
.Y(n_80)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_11),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_42),
.A2(n_36),
.B1(n_32),
.B2(n_28),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_78),
.A2(n_50),
.B1(n_43),
.B2(n_42),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_83),
.B1(n_97),
.B2(n_98),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_46),
.B(n_44),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_82),
.B(n_66),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_63),
.B(n_66),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_75),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_85),
.B(n_73),
.Y(n_106)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_40),
.B1(n_22),
.B2(n_21),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_87),
.A2(n_67),
.B1(n_68),
.B2(n_57),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_94),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_47),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_72),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_47),
.B1(n_22),
.B2(n_21),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_70),
.A2(n_17),
.B1(n_24),
.B2(n_16),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_100),
.B1(n_60),
.B2(n_64),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_74),
.A2(n_17),
.B1(n_16),
.B2(n_8),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_67),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_62),
.Y(n_103)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_113),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_89),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_119),
.Y(n_129)
);

NOR2x1_ASAP7_75t_R g130 ( 
.A(n_106),
.B(n_104),
.Y(n_130)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_107),
.B(n_108),
.Y(n_144)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_110),
.A2(n_90),
.B(n_100),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_74),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_112),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_84),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_124),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_62),
.Y(n_116)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_117),
.A2(n_121),
.B1(n_85),
.B2(n_92),
.Y(n_137)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_101),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_89),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_88),
.A2(n_83),
.B1(n_91),
.B2(n_98),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_81),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_90),
.B1(n_68),
.B2(n_59),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_57),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_126),
.B(n_131),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_96),
.C(n_80),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_138),
.C(n_120),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_114),
.A2(n_96),
.B1(n_97),
.B2(n_82),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_120),
.B(n_109),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_L g134 ( 
.A1(n_111),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_134),
.A2(n_136),
.B1(n_137),
.B2(n_106),
.Y(n_159)
);

OA22x2_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_99),
.B1(n_77),
.B2(n_85),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_85),
.C(n_77),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_118),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_92),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_113),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_114),
.A2(n_122),
.B1(n_110),
.B2(n_109),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_101),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_142),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_112),
.Y(n_143)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_145),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_146),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_101),
.Y(n_147)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_59),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_121),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_149),
.A2(n_108),
.B(n_107),
.Y(n_171)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_102),
.Y(n_153)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_154),
.A2(n_157),
.B1(n_102),
.B2(n_95),
.Y(n_183)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_139),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_160),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_163),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_121),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_144),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_161),
.Y(n_185)
);

FAx1_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_136),
.CI(n_138),
.CON(n_193),
.SN(n_193)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_102),
.Y(n_166)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_150),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_167),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_137),
.A2(n_136),
.B1(n_131),
.B2(n_141),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_168),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_171),
.A2(n_95),
.B(n_16),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_108),
.C(n_107),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_148),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_129),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_174),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_175),
.B(n_135),
.Y(n_194)
);

NAND3xp33_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_123),
.C(n_71),
.Y(n_176)
);

AOI21xp33_ASAP7_75t_L g202 ( 
.A1(n_176),
.A2(n_17),
.B(n_16),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_133),
.B(n_140),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_132),
.Y(n_182)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_183),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_136),
.B1(n_129),
.B2(n_150),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_184),
.A2(n_204),
.B1(n_205),
.B2(n_177),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_132),
.Y(n_186)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_171),
.A2(n_149),
.B(n_136),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_158),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_143),
.Y(n_190)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_193),
.B(n_197),
.Y(n_213)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_201),
.C(n_163),
.Y(n_217)
);

XOR2x1_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_128),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_152),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_170),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_165),
.B(n_142),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_200),
.B(n_153),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_76),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_24),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_203),
.A2(n_174),
.B1(n_169),
.B2(n_156),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_164),
.A2(n_95),
.B1(n_61),
.B2(n_24),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_155),
.A2(n_9),
.B(n_10),
.Y(n_205)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_208),
.A2(n_209),
.B1(n_180),
.B2(n_204),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_181),
.A2(n_168),
.B1(n_159),
.B2(n_155),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_198),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_215),
.Y(n_234)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_228),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_198),
.Y(n_215)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_195),
.C(n_191),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_190),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_186),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_185),
.B(n_173),
.Y(n_220)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_220),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_197),
.A2(n_177),
.B1(n_170),
.B2(n_156),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_221),
.A2(n_226),
.B1(n_203),
.B2(n_187),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_185),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_222),
.B(n_223),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_199),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_189),
.A2(n_166),
.B1(n_161),
.B2(n_165),
.Y(n_226)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_179),
.B(n_167),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_179),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_238),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_230),
.B(n_216),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_192),
.Y(n_231)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_226),
.Y(n_232)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_232),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_221),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_246),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_201),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_209),
.A2(n_180),
.B1(n_196),
.B2(n_188),
.Y(n_239)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_245),
.C(n_218),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_224),
.A2(n_188),
.B1(n_196),
.B2(n_193),
.Y(n_241)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_192),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_242),
.B(n_205),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_243),
.A2(n_227),
.B1(n_225),
.B2(n_182),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_206),
.C(n_207),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_213),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_252),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_191),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_258),
.C(n_261),
.Y(n_273)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_234),
.Y(n_257)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_257),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_210),
.C(n_207),
.Y(n_258)
);

NOR2xp67_ASAP7_75t_SL g260 ( 
.A(n_235),
.B(n_224),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_260),
.A2(n_262),
.B(n_265),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_210),
.C(n_218),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_187),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_244),
.A2(n_225),
.B(n_193),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_266),
.A2(n_241),
.B1(n_239),
.B2(n_230),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_267),
.A2(n_24),
.B(n_71),
.Y(n_283)
);

BUFx24_ASAP7_75t_SL g268 ( 
.A(n_247),
.Y(n_268)
);

BUFx24_ASAP7_75t_SL g284 ( 
.A(n_268),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_275),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_249),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_271),
.A2(n_283),
.B(n_5),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_233),
.B1(n_248),
.B2(n_246),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_274),
.A2(n_277),
.B1(n_280),
.B2(n_7),
.Y(n_291)
);

OA21x2_ASAP7_75t_L g277 ( 
.A1(n_259),
.A2(n_243),
.B(n_227),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_252),
.B(n_235),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_282),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_157),
.C(n_154),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_281),
.C(n_71),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_255),
.A2(n_263),
.B1(n_254),
.B2(n_261),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_253),
.B(n_95),
.C(n_76),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_251),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_61),
.Y(n_285)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_285),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_256),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_288),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_287),
.A2(n_5),
.B1(n_12),
.B2(n_10),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_250),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_292),
.C(n_296),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_7),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_290),
.B(n_294),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_291),
.B(n_8),
.Y(n_302)
);

AOI21xp33_ASAP7_75t_L g292 ( 
.A1(n_269),
.A2(n_24),
.B(n_7),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_272),
.A2(n_7),
.B1(n_11),
.B2(n_10),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_279),
.A2(n_5),
.B(n_11),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_273),
.B(n_281),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_273),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_298),
.B(n_303),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_299),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_282),
.Y(n_303)
);

NOR2xp67_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_278),
.Y(n_305)
);

AND2x2_ASAP7_75t_SL g310 ( 
.A(n_305),
.B(n_288),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_308),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_289),
.A2(n_284),
.B1(n_4),
.B2(n_3),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_310),
.A2(n_312),
.B(n_315),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_295),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_301),
.B(n_4),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_313),
.A2(n_304),
.B1(n_302),
.B2(n_300),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_4),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_4),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_317),
.C(n_319),
.Y(n_321)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_309),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_318),
.A2(n_310),
.B(n_311),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_8),
.C(n_9),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_9),
.Y(n_323)
);

OAI321xp33_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_321),
.A3(n_9),
.B1(n_2),
.B2(n_1),
.C(n_0),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_324),
.A2(n_0),
.B(n_1),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_325),
.B(n_0),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_1),
.B1(n_2),
.B2(n_275),
.Y(n_327)
);


endmodule