module real_jpeg_3904_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_0),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_0),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_0),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_0),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_0),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_0),
.B(n_267),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_0),
.B(n_288),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_0),
.B(n_227),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_1),
.Y(n_101)
);

INVx8_ASAP7_75t_L g229 ( 
.A(n_1),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_1),
.Y(n_257)
);

BUFx5_ASAP7_75t_L g310 ( 
.A(n_1),
.Y(n_310)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_1),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_1),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_1),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_2),
.B(n_34),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_2),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_2),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_2),
.B(n_136),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_2),
.B(n_319),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_2),
.B(n_335),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_2),
.B(n_58),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_3),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_3),
.Y(n_112)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_3),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_3),
.Y(n_170)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_3),
.Y(n_194)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_3),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_4),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_4),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_4),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_4),
.B(n_303),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_4),
.B(n_267),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_4),
.B(n_344),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_4),
.B(n_369),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_4),
.B(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_5),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_5),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_5),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_5),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_5),
.B(n_172),
.Y(n_171)
);

AND2x2_ASAP7_75t_SL g226 ( 
.A(n_5),
.B(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_6),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_6),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_6),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g384 ( 
.A(n_6),
.Y(n_384)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_7),
.Y(n_479)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_8),
.Y(n_231)
);

BUFx5_ASAP7_75t_L g288 ( 
.A(n_8),
.Y(n_288)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_10),
.Y(n_482)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_11),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_11),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_11),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_12),
.B(n_193),
.Y(n_222)
);

NAND2x1p5_ASAP7_75t_L g263 ( 
.A(n_12),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_12),
.B(n_74),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_12),
.B(n_288),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_12),
.B(n_286),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_12),
.B(n_89),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_12),
.B(n_382),
.Y(n_381)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_14),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_14),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_14),
.B(n_50),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_14),
.B(n_211),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g283 ( 
.A(n_14),
.B(n_53),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_14),
.B(n_358),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_14),
.B(n_400),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_15),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_15),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_15),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_15),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_15),
.B(n_286),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_15),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_15),
.B(n_361),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_15),
.B(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_16),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_16),
.B(n_74),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_16),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_16),
.B(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g149 ( 
.A(n_16),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_17),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_17),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_17),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_17),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_17),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_17),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_18),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_18),
.B(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_18),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_18),
.B(n_327),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_18),
.B(n_50),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_18),
.B(n_65),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_18),
.B(n_384),
.Y(n_383)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_478),
.B(n_480),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_196),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_195),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_156),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_25),
.B(n_156),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_113),
.B2(n_155),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_79),
.C(n_96),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_28),
.B(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_48),
.C(n_61),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_29),
.A2(n_30),
.B1(n_48),
.B2(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_36),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_31),
.B(n_37),
.C(n_44),
.Y(n_126)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_44),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_42),
.Y(n_392)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_43),
.Y(n_150)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_43),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_47),
.Y(n_120)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_47),
.Y(n_189)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_48),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.C(n_56),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_49),
.B(n_56),
.Y(n_176)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_52),
.B(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g307 ( 
.A(n_55),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_59),
.Y(n_369)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_60),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_60),
.Y(n_286)
);

INVx5_ASAP7_75t_L g328 ( 
.A(n_60),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_61),
.B(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_68),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_62),
.B(n_70),
.C(n_73),
.Y(n_125)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_66),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_66),
.Y(n_382)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_67),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_73),
.B2(n_78),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_69),
.A2(n_70),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_69),
.B(n_117),
.C(n_121),
.Y(n_141)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_71),
.Y(n_355)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx5_ASAP7_75t_L g344 ( 
.A(n_72),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_73),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_99),
.C(n_102),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_73),
.A2(n_78),
.B1(n_99),
.B2(n_100),
.Y(n_164)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_75),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_76),
.Y(n_361)
);

INVx5_ASAP7_75t_L g401 ( 
.A(n_76),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_79),
.B(n_96),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_84),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_80),
.B(n_85),
.C(n_95),
.Y(n_139)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_91),
.B2(n_95),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_90),
.Y(n_273)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_105),
.C(n_109),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_97),
.A2(n_98),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_99),
.B(n_166),
.C(n_171),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_99),
.A2(n_100),
.B1(n_171),
.B2(n_217),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_101),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_102),
.B(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_104),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_105),
.A2(n_109),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_105),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_105),
.B(n_183),
.C(n_191),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_105),
.A2(n_180),
.B1(n_191),
.B2(n_192),
.Y(n_219)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_109),
.Y(n_181)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_127),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_125),
.C(n_126),
.Y(n_114)
);

FAx1_ASAP7_75t_SL g159 ( 
.A(n_115),
.B(n_125),
.CI(n_126),
.CON(n_159),
.SN(n_159)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_121),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_118),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_124),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_140),
.B2(n_154),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_139),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_152),
.B2(n_153),
.Y(n_140)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_146),
.B1(n_147),
.B2(n_151),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_143),
.Y(n_151)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.C(n_160),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_157),
.B(n_159),
.Y(n_474)
);

BUFx24_ASAP7_75t_SL g484 ( 
.A(n_159),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_160),
.B(n_474),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_177),
.C(n_182),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_161),
.A2(n_162),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.C(n_175),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_163),
.B(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_165),
.B(n_175),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_167),
.B(n_216),
.Y(n_215)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_171),
.Y(n_217)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_177),
.B(n_182),
.Y(n_240)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_219),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.C(n_190),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_190),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_186),
.B(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

AO21x1_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_471),
.B(n_476),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_290),
.B(n_470),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_241),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_200),
.B(n_241),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_234),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_201),
.B(n_235),
.C(n_238),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_218),
.C(n_220),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_202),
.B(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.C(n_215),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_203),
.B(n_456),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_205),
.A2(n_206),
.B1(n_215),
.B2(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.C(n_213),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_207),
.B(n_213),
.Y(n_446)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_210),
.B(n_446),
.Y(n_445)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_215),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_220),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_230),
.C(n_232),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_221),
.B(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.C(n_226),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_222),
.B(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_226),
.Y(n_253)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_230),
.B(n_232),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_238),
.Y(n_234)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.C(n_248),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_243),
.B(n_246),
.Y(n_466)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_248),
.B(n_466),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_274),
.C(n_277),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_250),
.B(n_459),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.C(n_261),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_251),
.A2(n_252),
.B1(n_437),
.B2(n_438),
.Y(n_436)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_254),
.A2(n_255),
.B(n_258),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_254),
.B(n_261),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx6_ASAP7_75t_SL g259 ( 
.A(n_260),
.Y(n_259)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.C(n_269),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_262),
.A2(n_263),
.B1(n_265),
.B2(n_266),
.Y(n_414)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

BUFx8_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx5_ASAP7_75t_L g335 ( 
.A(n_268),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_269),
.B(n_414),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_270),
.B(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g459 ( 
.A1(n_274),
.A2(n_275),
.B1(n_277),
.B2(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_277),
.Y(n_460)
);

MAJx2_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_287),
.C(n_289),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_279),
.B(n_448),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_283),
.C(n_284),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_280),
.B(n_426),
.Y(n_425)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_283),
.Y(n_427)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_287),
.B(n_289),
.Y(n_448)
);

AOI21x1_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_464),
.B(n_469),
.Y(n_290)
);

OAI21x1_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_451),
.B(n_463),
.Y(n_291)
);

AOI21x1_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_433),
.B(n_450),
.Y(n_292)
);

OAI21x1_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_407),
.B(n_432),
.Y(n_293)
);

AOI21x1_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_376),
.B(n_406),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_347),
.B(n_375),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_330),
.B(n_346),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_312),
.B(n_329),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_308),
.B(n_311),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_305),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_305),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_309),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_302),
.Y(n_313)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx8_ASAP7_75t_L g394 ( 
.A(n_307),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_314),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_321),
.B2(n_322),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_324),
.C(n_325),
.Y(n_345)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_317),
.B(n_318),
.Y(n_338)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_323),
.A2(n_324),
.B1(n_325),
.B2(n_326),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_345),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_331),
.B(n_345),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_339),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_338),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_333),
.B(n_338),
.C(n_349),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_336),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_334),
.B(n_336),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_339),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_340),
.B(n_365),
.C(n_366),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_342),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_343),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_350),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_348),
.B(n_350),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_363),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_351),
.B(n_364),
.C(n_367),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_352),
.B(n_354),
.C(n_356),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_356),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_357),
.A2(n_359),
.B1(n_360),
.B2(n_362),
.Y(n_356)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_357),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_359),
.B(n_362),
.Y(n_385)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_367),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_370),
.Y(n_367)
);

MAJx2_ASAP7_75t_L g404 ( 
.A(n_368),
.B(n_372),
.C(n_373),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_371),
.A2(n_372),
.B1(n_373),
.B2(n_374),
.Y(n_370)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_371),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_372),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_377),
.B(n_405),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_377),
.B(n_405),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_378),
.B(n_387),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_386),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_379),
.B(n_386),
.C(n_431),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_385),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_383),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_381),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_383),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_385),
.B(n_421),
.C(n_422),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_387),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_396),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_388),
.B(n_398),
.C(n_403),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_395),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_393),
.Y(n_389)
);

MAJx2_ASAP7_75t_L g418 ( 
.A(n_390),
.B(n_393),
.C(n_395),
.Y(n_418)
);

INVx6_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_398),
.B1(n_403),
.B2(n_404),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_402),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_399),
.B(n_402),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_404),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_430),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_408),
.B(n_430),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_419),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_410),
.B(n_411),
.C(n_419),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_412),
.A2(n_413),
.B1(n_415),
.B2(n_416),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_412),
.B(n_442),
.C(n_443),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_417),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_418),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_420),
.B(n_423),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_420),
.B(n_424),
.C(n_429),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_424),
.A2(n_425),
.B1(n_428),
.B2(n_429),
.Y(n_423)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_424),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_425),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_434),
.B(n_449),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_434),
.B(n_449),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_435),
.B(n_440),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_439),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_436),
.B(n_439),
.C(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_437),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_440),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_441),
.B(n_444),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_441),
.B(n_445),
.C(n_447),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_447),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_452),
.B(n_461),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_452),
.B(n_461),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_454),
.Y(n_452)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_453),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_458),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_455),
.B(n_458),
.C(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_465),
.B(n_467),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_465),
.B(n_467),
.Y(n_469)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_473),
.B(n_475),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_473),
.B(n_475),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx5_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx8_ASAP7_75t_L g481 ( 
.A(n_479),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_482),
.Y(n_480)
);


endmodule