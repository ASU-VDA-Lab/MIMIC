module real_jpeg_32772_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_313;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_0),
.Y(n_235)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_0),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_0),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_1),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_1),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_1),
.B(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_1),
.A2(n_7),
.B1(n_256),
.B2(n_258),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_1),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_1),
.B(n_439),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_1),
.B(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_1),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_2),
.A2(n_19),
.B(n_536),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_2),
.B(n_537),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_3),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_4),
.Y(n_88)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_5),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_5),
.Y(n_195)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_5),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_6),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_6),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_6),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_6),
.B(n_268),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_6),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_6),
.B(n_418),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_6),
.B(n_422),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_6),
.Y(n_446)
);

NAND2x1_ASAP7_75t_SL g36 ( 
.A(n_7),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_7),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_7),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_7),
.B(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_7),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_7),
.B(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_8),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_9),
.Y(n_150)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_9),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_9),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_10),
.B(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_10),
.B(n_285),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_10),
.B(n_299),
.Y(n_298)
);

NAND2x1_ASAP7_75t_L g308 ( 
.A(n_10),
.B(n_309),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_10),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_10),
.B(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_10),
.B(n_458),
.Y(n_457)
);

AND2x2_ASAP7_75t_SL g496 ( 
.A(n_10),
.B(n_497),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_11),
.B(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_R g94 ( 
.A(n_11),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_11),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_11),
.B(n_214),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_11),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_11),
.B(n_313),
.Y(n_312)
);

AND2x4_ASAP7_75t_L g345 ( 
.A(n_11),
.B(n_346),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_12),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_12),
.B(n_43),
.Y(n_42)
);

AND2x4_ASAP7_75t_SL g66 ( 
.A(n_12),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_12),
.B(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_12),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_12),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_12),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_12),
.B(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_13),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_14),
.Y(n_78)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_15),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_15),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_15),
.B(n_435),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_15),
.B(n_500),
.Y(n_499)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_16),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_16),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_16),
.Y(n_291)
);

AND2x2_ASAP7_75t_SL g26 ( 
.A(n_17),
.B(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_17),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_17),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_17),
.B(n_119),
.Y(n_118)
);

NAND2x1_ASAP7_75t_L g124 ( 
.A(n_17),
.B(n_125),
.Y(n_124)
);

NAND2x1p5_ASAP7_75t_L g153 ( 
.A(n_17),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_17),
.B(n_67),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_222),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_220),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_169),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_22),
.B(n_169),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_97),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_68),
.C(n_82),
.Y(n_23)
);

XNOR2x1_ASAP7_75t_L g171 ( 
.A(n_24),
.B(n_172),
.Y(n_171)
);

MAJx2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_40),
.C(n_54),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_25),
.B(n_40),
.Y(n_390)
);

XNOR2x1_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_R g116 ( 
.A(n_26),
.B(n_32),
.C(n_35),
.Y(n_116)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_31),
.A2(n_32),
.B1(n_206),
.B2(n_232),
.Y(n_425)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_32),
.A2(n_107),
.B(n_111),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_32),
.B(n_107),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_32),
.B(n_107),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_32),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_32),
.B(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_39),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_39),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_39),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_39),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_45),
.C(n_49),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

XNOR2x1_ASAP7_75t_L g197 ( 
.A(n_42),
.B(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22x1_ASAP7_75t_SL g198 ( 
.A1(n_45),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_198)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_48),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_48),
.Y(n_265)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_52),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_52),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_53),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_53),
.Y(n_441)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_54),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_61),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_55),
.A2(n_56),
.B1(n_267),
.B2(n_270),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_62),
.C(n_66),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_56),
.B(n_262),
.C(n_267),
.Y(n_323)
);

OR2x2_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_66),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_85),
.C(n_89),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_66),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_66),
.B(n_416),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_66),
.B(n_417),
.Y(n_489)
);

INVx4_ASAP7_75t_SL g247 ( 
.A(n_67),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_70),
.B(n_83),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_80),
.B2(n_81),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_76),
.B1(n_77),
.B2(n_79),
.Y(n_72)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_75),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_76),
.A2(n_77),
.B1(n_92),
.B2(n_93),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_84),
.C(n_92),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_77),
.B(n_142),
.C(n_143),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_78),
.Y(n_211)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_78),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_78),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

INVxp33_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_84),
.B(n_219),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_85),
.A2(n_134),
.B1(n_139),
.B2(n_140),
.Y(n_133)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_85),
.A2(n_140),
.B1(n_182),
.B2(n_184),
.Y(n_181)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_88),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_88),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_88),
.Y(n_502)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_89),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_89),
.A2(n_183),
.B1(n_275),
.B2(n_278),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_89),
.B(n_275),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx6_ASAP7_75t_L g420 ( 
.A(n_91),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_91),
.Y(n_473)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_144),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_129),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_115),
.C(n_117),
.Y(n_99)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_100),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_106),
.B(n_112),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_113),
.B(n_114),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_101),
.A2(n_102),
.B1(n_153),
.B2(n_160),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_101),
.B(n_165),
.C(n_166),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_101),
.A2(n_102),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_102),
.B(n_293),
.C(n_298),
.Y(n_304)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_104),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_107),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_111),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_117),
.Y(n_177)
);

XOR2x2_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_126),
.C(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_121),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_126),
.B2(n_128),
.Y(n_122)
);

MAJx2_ASAP7_75t_L g186 ( 
.A(n_123),
.B(n_187),
.C(n_190),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_123),
.A2(n_124),
.B1(n_188),
.B2(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_126),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_141),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_161),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_151),
.B2(n_152),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_146),
.A2(n_147),
.B1(n_308),
.B2(n_311),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_146),
.B(n_308),
.C(n_312),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_164),
.B1(n_167),
.B2(n_168),
.Y(n_161)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_162),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.C(n_178),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_171),
.B(n_174),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

INVxp33_ASAP7_75t_SL g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_179),
.B(n_400),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_199),
.C(n_217),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g386 ( 
.A(n_180),
.B(n_387),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_185),
.C(n_196),
.Y(n_180)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_181),
.Y(n_372)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_182),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_186),
.B(n_197),
.Y(n_373)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_188),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_190),
.B(n_325),
.Y(n_324)
);

NOR2xp67_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_195),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_199),
.A2(n_200),
.B1(n_217),
.B2(n_218),
.Y(n_387)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_209),
.C(n_212),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2x1_ASAP7_75t_L g364 ( 
.A(n_202),
.B(n_365),
.Y(n_364)
);

MAJx2_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_206),
.C(n_207),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_203),
.A2(n_206),
.B1(n_232),
.B2(n_339),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_203),
.Y(n_339)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_206),
.Y(n_232)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_207),
.Y(n_341)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_208),
.Y(n_300)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_210),
.B(n_213),
.Y(n_365)
);

INVxp33_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OA21x2_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_376),
.B(n_527),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_354),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_315),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g529 ( 
.A(n_227),
.B(n_315),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_271),
.C(n_301),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_228),
.B(n_404),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_243),
.Y(n_228)
);

MAJx2_ASAP7_75t_L g317 ( 
.A(n_229),
.B(n_244),
.C(n_261),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_233),
.C(n_236),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_230),
.A2(n_231),
.B1(n_411),
.B2(n_412),
.Y(n_410)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_233),
.A2(n_236),
.B1(n_237),
.B2(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_233),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_240),
.Y(n_310)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_261),
.Y(n_243)
);

OA21x2_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_248),
.B(n_254),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_253),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_254),
.A2(n_255),
.B1(n_343),
.B2(n_344),
.Y(n_342)
);

INVxp33_ASAP7_75t_SL g254 ( 
.A(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_255),
.B(n_368),
.C(n_369),
.Y(n_367)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_266),
.Y(n_261)
);

NOR2x1_ASAP7_75t_R g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_276),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_263),
.B(n_472),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_263),
.B(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_272),
.B(n_302),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_279),
.C(n_292),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_273),
.A2(n_274),
.B1(n_279),
.B2(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_275),
.Y(n_278)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_279),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_284),
.C(n_287),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_280),
.A2(n_281),
.B1(n_287),
.B2(n_288),
.Y(n_512)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_284),
.B(n_512),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx8_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_292),
.B(n_408),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_296),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_306),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_304),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_305),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_306),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_312),
.Y(n_306)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_308),
.Y(n_311)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_327),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_317),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_318),
.B(n_328),
.C(n_375),
.Y(n_374)
);

XNOR2x1_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_322),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

MAJx2_ASAP7_75t_L g362 ( 
.A(n_321),
.B(n_323),
.C(n_324),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_335),
.Y(n_328)
);

OA21x2_ASAP7_75t_L g356 ( 
.A1(n_329),
.A2(n_357),
.B(n_358),
.Y(n_356)
);

OAI21x1_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_333),
.B(n_334),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_332),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_342),
.B1(n_352),
.B2(n_353),
.Y(n_335)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_336),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_337),
.A2(n_338),
.B1(n_340),
.B2(n_341),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_342),
.Y(n_352)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_349),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_345),
.Y(n_368)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_349),
.Y(n_369)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_352),
.B(n_353),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_352),
.B(n_353),
.Y(n_358)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_354),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_374),
.Y(n_354)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_355),
.B(n_374),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_359),
.Y(n_355)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_356),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_371),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_360),
.Y(n_382)
);

OAI22x1_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_362),
.B1(n_363),
.B2(n_370),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_362),
.B(n_393),
.C(n_394),
.Y(n_392)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_363),
.Y(n_370)
);

XNOR2x1_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_366),
.Y(n_363)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_364),
.Y(n_394)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_367),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_371),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_401),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_377),
.A2(n_528),
.B(n_532),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_383),
.B1(n_395),
.B2(n_398),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_379),
.B(n_384),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_381),
.C(n_382),
.Y(n_379)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_388),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_386),
.B(n_392),
.C(n_397),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_392),
.Y(n_388)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_389),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_391),
.Y(n_389)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

NOR2x1_ASAP7_75t_L g533 ( 
.A(n_396),
.B(n_399),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_396),
.B(n_399),
.Y(n_535)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_399),
.Y(n_398)
);

AO21x1_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_426),
.B(n_526),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_403),
.B(n_405),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_403),
.B(n_405),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_410),
.C(n_414),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_406),
.A2(n_407),
.B1(n_523),
.B2(n_524),
.Y(n_522)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_410),
.B(n_414),
.Y(n_524)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_421),
.C(n_424),
.Y(n_414)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_415),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g418 ( 
.A(n_419),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_421),
.A2(n_424),
.B1(n_425),
.B2(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_421),
.Y(n_516)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_520),
.B(n_525),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_428),
.A2(n_504),
.B(n_519),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_482),
.B(n_503),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_430),
.A2(n_464),
.B(n_481),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_431),
.B(n_455),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_431),
.B(n_455),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_433),
.B1(n_442),
.B2(n_443),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g433 ( 
.A(n_434),
.B(n_438),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_434),
.B(n_438),
.C(n_442),
.Y(n_483)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_444),
.A2(n_445),
.B1(n_450),
.B2(n_451),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_445),
.B(n_450),
.Y(n_487)
);

NOR2x1_ASAP7_75t_SL g445 ( 
.A(n_446),
.B(n_447),
.Y(n_445)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_449),
.Y(n_470)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_454),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_460),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_456),
.A2(n_457),
.B1(n_460),
.B2(n_461),
.Y(n_479)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

BUFx4f_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_465),
.A2(n_474),
.B(n_480),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_466),
.B(n_471),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_468),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_467),
.B(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_479),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_475),
.B(n_479),
.Y(n_480)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_484),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_483),
.B(n_484),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_490),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_486),
.A2(n_487),
.B1(n_488),
.B2(n_489),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_486),
.B(n_489),
.C(n_490),
.Y(n_505)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_494),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_491),
.B(n_496),
.C(n_498),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_493),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_495),
.A2(n_496),
.B1(n_498),
.B2(n_499),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx5_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx5_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_506),
.Y(n_504)
);

NOR2xp67_ASAP7_75t_L g519 ( 
.A(n_505),
.B(n_506),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_507),
.A2(n_513),
.B1(n_517),
.B2(n_518),
.Y(n_506)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_507),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_508),
.A2(n_509),
.B1(n_510),
.B2(n_511),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_509),
.B(n_510),
.C(n_518),
.Y(n_521)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_513),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_515),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_522),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_521),
.B(n_522),
.Y(n_525)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g528 ( 
.A1(n_529),
.A2(n_530),
.B(n_531),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_533),
.A2(n_534),
.B(n_535),
.Y(n_532)
);


endmodule