module fake_jpeg_30068_n_234 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_234);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_234;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_40),
.B(n_44),
.Y(n_80)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_20),
.B(n_0),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_50),
.Y(n_91)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_28),
.B(n_1),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_56),
.Y(n_85)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_21),
.B(n_26),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_65),
.Y(n_70)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_23),
.B(n_3),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

NAND2xp33_ASAP7_75t_SL g72 ( 
.A(n_62),
.B(n_36),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_29),
.B(n_4),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_30),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_17),
.B(n_10),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_35),
.Y(n_75)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_61),
.A2(n_19),
.B1(n_37),
.B2(n_31),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_67),
.A2(n_45),
.B(n_39),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_90),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_33),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_75),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_41),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_83),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_17),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_41),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_88),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_50),
.A2(n_36),
.B1(n_37),
.B2(n_31),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_87),
.A2(n_59),
.B1(n_57),
.B2(n_55),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_43),
.B(n_33),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_36),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_34),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_47),
.B(n_13),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_9),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_80),
.B(n_58),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_98),
.B(n_112),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_85),
.B(n_14),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_99),
.B(n_105),
.Y(n_131)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_101),
.Y(n_144)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_70),
.B(n_15),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_72),
.A2(n_34),
.B(n_15),
.C(n_7),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_115),
.Y(n_129)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_121),
.B(n_69),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_67),
.B(n_46),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_42),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_116),
.Y(n_148)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_78),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_48),
.Y(n_116)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_94),
.B(n_60),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_100),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_123),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_34),
.Y(n_123)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_124),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_68),
.B(n_39),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_126),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_112),
.A2(n_71),
.B1(n_76),
.B2(n_89),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_128),
.A2(n_130),
.B1(n_135),
.B2(n_141),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_98),
.A2(n_87),
.B1(n_71),
.B2(n_86),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_110),
.A2(n_86),
.B1(n_82),
.B2(n_97),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_116),
.B1(n_117),
.B2(n_121),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_142),
.A2(n_145),
.B1(n_144),
.B2(n_148),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_120),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_149),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_101),
.A2(n_97),
.B1(n_81),
.B2(n_66),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_117),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_151),
.B(n_152),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_117),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_126),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_155),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_131),
.B(n_102),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_159),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_102),
.C(n_111),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_157),
.A2(n_145),
.B1(n_150),
.B2(n_133),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_111),
.B(n_69),
.Y(n_158)
);

OAI21x1_ASAP7_75t_L g173 ( 
.A1(n_158),
.A2(n_167),
.B(n_169),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_105),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_104),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_165),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_107),
.Y(n_162)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_162),
.Y(n_172)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_99),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_166),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_133),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_114),
.C(n_119),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_106),
.B(n_109),
.Y(n_167)
);

AND2x6_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_103),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_138),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_134),
.A2(n_124),
.B(n_103),
.Y(n_169)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

BUFx2_ASAP7_75t_SL g179 ( 
.A(n_170),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_139),
.B(n_108),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_136),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_161),
.A2(n_139),
.B1(n_150),
.B2(n_118),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_180),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_153),
.B(n_164),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_177),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_162),
.A2(n_138),
.B1(n_136),
.B2(n_146),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_173),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_186),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_169),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_157),
.Y(n_199)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

AO22x1_ASAP7_75t_L g189 ( 
.A1(n_173),
.A2(n_162),
.B1(n_158),
.B2(n_168),
.Y(n_189)
);

AO21x1_ASAP7_75t_L g209 ( 
.A1(n_189),
.A2(n_172),
.B(n_175),
.Y(n_209)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_181),
.B(n_155),
.Y(n_191)
);

NAND3xp33_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_184),
.C(n_177),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_192),
.B(n_194),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_152),
.C(n_151),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_184),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_198),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_156),
.C(n_166),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_199),
.B(n_200),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_161),
.C(n_167),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_208),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_195),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_209),
.Y(n_210)
);

BUFx24_ASAP7_75t_SL g208 ( 
.A(n_193),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_204),
.Y(n_212)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_212),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_181),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_214),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_202),
.B(n_198),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_209),
.A2(n_197),
.B(n_189),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_215),
.B(n_192),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_187),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_203),
.C(n_182),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_217),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_210),
.A2(n_172),
.B(n_195),
.C(n_186),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_SL g224 ( 
.A1(n_219),
.A2(n_127),
.B(n_124),
.C(n_108),
.Y(n_224)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_194),
.C(n_200),
.Y(n_220)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_222),
.C(n_127),
.Y(n_226)
);

AOI322xp5_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_211),
.A3(n_176),
.B1(n_180),
.B2(n_179),
.C1(n_170),
.C2(n_146),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_223),
.A2(n_219),
.B(n_217),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_226),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_225),
.B(n_221),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_227),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_229),
.A2(n_220),
.B(n_6),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_228),
.C(n_6),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_232),
.A2(n_230),
.B1(n_5),
.B2(n_39),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_5),
.C(n_218),
.Y(n_234)
);


endmodule