module fake_ariane_2740_n_552 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_552);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_552;

wire n_295;
wire n_356;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_516;
wire n_332;
wire n_294;
wire n_197;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_205;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_424;
wire n_528;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_462;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_264;
wire n_198;
wire n_232;
wire n_441;
wire n_385;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_399;
wire n_520;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_500;
wire n_336;
wire n_315;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_487;
wire n_167;
wire n_422;
wire n_269;
wire n_158;
wire n_259;
wire n_446;
wire n_405;
wire n_169;
wire n_173;
wire n_242;
wire n_309;
wire n_331;
wire n_320;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_247;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_518;
wire n_439;
wire n_222;
wire n_478;
wire n_510;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_330;
wire n_400;
wire n_282;
wire n_328;
wire n_368;
wire n_277;
wire n_301;
wire n_248;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_427;
wire n_497;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_511;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_334;
wire n_192;
wire n_488;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_440;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_459;
wire n_321;
wire n_221;
wire n_361;
wire n_458;
wire n_383;
wire n_237;
wire n_175;
wire n_453;
wire n_491;
wire n_181;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_236;
wire n_281;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_464;
wire n_546;
wire n_297;
wire n_503;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_217;
wire n_452;
wire n_178;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_343;
wire n_414;
wire n_287;
wire n_302;
wire n_380;
wire n_284;
wire n_448;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_278;
wire n_255;
wire n_450;
wire n_257;
wire n_451;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_182;
wire n_482;
wire n_316;
wire n_196;
wire n_407;
wire n_254;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_234;
wire n_492;
wire n_280;
wire n_252;
wire n_215;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_540;
wire n_216;
wire n_544;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_195;
wire n_213;
wire n_304;
wire n_509;
wire n_306;
wire n_313;
wire n_430;
wire n_493;
wire n_203;
wire n_378;
wire n_436;
wire n_375;
wire n_324;
wire n_337;
wire n_437;
wire n_274;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_292;
wire n_174;
wire n_275;
wire n_204;
wire n_521;
wire n_496;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_494;
wire n_263;
wire n_434;
wire n_360;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_425;
wire n_431;
wire n_508;
wire n_411;
wire n_484;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_408;
wire n_322;
wire n_251;
wire n_506;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_359;
wire n_531;

INVxp67_ASAP7_75t_SL g158 ( 
.A(n_4),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_140),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_36),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_90),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_62),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_79),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_69),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_102),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_118),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_17),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_146),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_27),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_72),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_80),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_73),
.Y(n_174)
);

INVxp33_ASAP7_75t_SL g175 ( 
.A(n_74),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_139),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_2),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_3),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_106),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_58),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_96),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_123),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_31),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_6),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_117),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

BUFx2_ASAP7_75t_SL g189 ( 
.A(n_52),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_61),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_103),
.Y(n_191)
);

INVxp67_ASAP7_75t_SL g192 ( 
.A(n_55),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_50),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_1),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_42),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_9),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_70),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_104),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_86),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_49),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_84),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_14),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_0),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_115),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_64),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_46),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_135),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_18),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_154),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_125),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_110),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_32),
.Y(n_213)
);

INVxp67_ASAP7_75t_SL g214 ( 
.A(n_141),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_33),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_78),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_127),
.Y(n_217)
);

INVxp33_ASAP7_75t_SL g218 ( 
.A(n_16),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_155),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_6),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_20),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_85),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_51),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_89),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_29),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_97),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_5),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_54),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_105),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_5),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_10),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_56),
.Y(n_232)
);

INVxp33_ASAP7_75t_L g233 ( 
.A(n_67),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_81),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_120),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_119),
.Y(n_236)
);

INVxp67_ASAP7_75t_SL g237 ( 
.A(n_157),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_28),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_88),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_83),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_99),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_194),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_0),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

AND2x4_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_1),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_177),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_201),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_236),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_158),
.Y(n_251)
);

AND2x4_ASAP7_75t_L g252 ( 
.A(n_205),
.B(n_2),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_178),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_205),
.B(n_3),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_162),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_186),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_203),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_201),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_164),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_165),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_166),
.B(n_4),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_168),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_159),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_171),
.B(n_232),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_169),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_196),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_172),
.Y(n_268)
);

AND2x4_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_7),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_174),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_180),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_181),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_160),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_161),
.B(n_7),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_188),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_190),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_191),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_193),
.B(n_8),
.Y(n_278)
);

AND2x4_ASAP7_75t_L g279 ( 
.A(n_182),
.B(n_195),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_167),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_175),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_256),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_264),
.Y(n_283)
);

CKINVDCx8_ASAP7_75t_R g284 ( 
.A(n_280),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_242),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_265),
.B(n_161),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_243),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_244),
.B(n_187),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_256),
.B(n_250),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_246),
.A2(n_237),
.B1(n_218),
.B2(n_189),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_255),
.B(n_237),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_198),
.Y(n_292)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_243),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_247),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_243),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_245),
.Y(n_296)
);

INVxp67_ASAP7_75t_SL g297 ( 
.A(n_251),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_253),
.B(n_187),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_274),
.A2(n_211),
.B1(n_170),
.B2(n_222),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_R g300 ( 
.A(n_273),
.B(n_185),
.Y(n_300)
);

AND3x1_ASAP7_75t_L g301 ( 
.A(n_262),
.B(n_240),
.C(n_238),
.Y(n_301)
);

AND2x4_ASAP7_75t_L g302 ( 
.A(n_250),
.B(n_252),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_200),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_243),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_260),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_253),
.B(n_183),
.Y(n_306)
);

AND2x6_ASAP7_75t_SL g307 ( 
.A(n_246),
.B(n_204),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_269),
.B(n_183),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_252),
.B(n_197),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_261),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_263),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_273),
.B(n_199),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_258),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_279),
.B(n_197),
.Y(n_314)
);

INVx4_ASAP7_75t_SL g315 ( 
.A(n_269),
.Y(n_315)
);

BUFx10_ASAP7_75t_L g316 ( 
.A(n_279),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_270),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_249),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_249),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_249),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_275),
.B(n_202),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_302),
.B(n_315),
.Y(n_322)
);

OR2x6_ASAP7_75t_L g323 ( 
.A(n_299),
.B(n_267),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_305),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_310),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_298),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_313),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_290),
.B(n_274),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_290),
.B(n_262),
.Y(n_329)
);

NOR2xp67_ASAP7_75t_L g330 ( 
.A(n_313),
.B(n_268),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_283),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_254),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_311),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_315),
.B(n_276),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_315),
.B(n_277),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_284),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_317),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_299),
.A2(n_278),
.B1(n_213),
.B2(n_206),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_285),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_293),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_282),
.B(n_272),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_308),
.A2(n_278),
.B1(n_192),
.B2(n_214),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_296),
.Y(n_343)
);

INVx2_ASAP7_75t_SL g344 ( 
.A(n_316),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g345 ( 
.A(n_316),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_281),
.B(n_308),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_286),
.B(n_207),
.Y(n_347)
);

OAI221xp5_ASAP7_75t_L g348 ( 
.A1(n_297),
.A2(n_219),
.B1(n_208),
.B2(n_216),
.C(n_235),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_289),
.B(n_249),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_287),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_306),
.B(n_163),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_283),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_297),
.B(n_259),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_301),
.B(n_291),
.Y(n_354)
);

NAND2x1p5_ASAP7_75t_L g355 ( 
.A(n_309),
.B(n_212),
.Y(n_355)
);

NOR3xp33_ASAP7_75t_L g356 ( 
.A(n_321),
.B(n_267),
.C(n_223),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_312),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_300),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_314),
.Y(n_359)
);

OR2x6_ASAP7_75t_L g360 ( 
.A(n_291),
.B(n_248),
.Y(n_360)
);

BUFx4f_ASAP7_75t_L g361 ( 
.A(n_294),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_292),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_307),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_292),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_303),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_288),
.B(n_259),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_303),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_327),
.Y(n_368)
);

CKINVDCx8_ASAP7_75t_R g369 ( 
.A(n_358),
.Y(n_369)
);

INVx2_ASAP7_75t_SL g370 ( 
.A(n_331),
.Y(n_370)
);

NAND2x1p5_ASAP7_75t_L g371 ( 
.A(n_352),
.B(n_293),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_352),
.B(n_248),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_346),
.A2(n_234),
.B1(n_215),
.B2(n_228),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_343),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_336),
.B(n_221),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_323),
.A2(n_338),
.B1(n_326),
.B2(n_360),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_324),
.Y(n_377)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_340),
.Y(n_378)
);

AO22x1_ASAP7_75t_L g379 ( 
.A1(n_356),
.A2(n_224),
.B1(n_226),
.B2(n_229),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_364),
.A2(n_231),
.B1(n_217),
.B2(n_209),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_365),
.A2(n_320),
.B(n_319),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_359),
.B(n_344),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_353),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_362),
.B(n_173),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_367),
.B(n_176),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_345),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_340),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_325),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_339),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_333),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_322),
.Y(n_391)
);

NOR2xp67_ASAP7_75t_L g392 ( 
.A(n_334),
.B(n_295),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_350),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_328),
.B(n_179),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_337),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_361),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_335),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_361),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_366),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_332),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_355),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_341),
.A2(n_318),
.B(n_304),
.Y(n_402)
);

INVx5_ASAP7_75t_L g403 ( 
.A(n_360),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_329),
.A2(n_342),
.B1(n_351),
.B2(n_354),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_355),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_347),
.B(n_184),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_360),
.B(n_225),
.Y(n_407)
);

A2O1A1Ixp33_ASAP7_75t_L g408 ( 
.A1(n_338),
.A2(n_210),
.B(n_259),
.C(n_8),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_323),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_393),
.Y(n_410)
);

OR2x2_ASAP7_75t_L g411 ( 
.A(n_372),
.B(n_357),
.Y(n_411)
);

AOI21x1_ASAP7_75t_L g412 ( 
.A1(n_402),
.A2(n_349),
.B(n_330),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_389),
.Y(n_413)
);

A2O1A1Ixp33_ASAP7_75t_L g414 ( 
.A1(n_394),
.A2(n_348),
.B(n_210),
.C(n_363),
.Y(n_414)
);

OAI21x1_ASAP7_75t_L g415 ( 
.A1(n_381),
.A2(n_210),
.B(n_11),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_396),
.B(n_323),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_384),
.A2(n_259),
.B1(n_9),
.B2(n_13),
.Y(n_417)
);

OAI21x1_ASAP7_75t_L g418 ( 
.A1(n_397),
.A2(n_12),
.B(n_15),
.Y(n_418)
);

OA21x2_ASAP7_75t_L g419 ( 
.A1(n_397),
.A2(n_19),
.B(n_21),
.Y(n_419)
);

OA21x2_ASAP7_75t_L g420 ( 
.A1(n_383),
.A2(n_22),
.B(n_23),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_389),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_377),
.Y(n_422)
);

AO21x1_ASAP7_75t_L g423 ( 
.A1(n_404),
.A2(n_156),
.B(n_25),
.Y(n_423)
);

NAND2xp33_ASAP7_75t_L g424 ( 
.A(n_398),
.B(n_387),
.Y(n_424)
);

OA21x2_ASAP7_75t_L g425 ( 
.A1(n_383),
.A2(n_24),
.B(n_26),
.Y(n_425)
);

OAI21x1_ASAP7_75t_L g426 ( 
.A1(n_393),
.A2(n_30),
.B(n_34),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_378),
.Y(n_427)
);

OAI21x1_ASAP7_75t_SL g428 ( 
.A1(n_373),
.A2(n_153),
.B(n_37),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_370),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_374),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_382),
.Y(n_431)
);

AO21x1_ASAP7_75t_L g432 ( 
.A1(n_380),
.A2(n_152),
.B(n_38),
.Y(n_432)
);

OAI21x1_ASAP7_75t_L g433 ( 
.A1(n_387),
.A2(n_35),
.B(n_39),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_382),
.B(n_40),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_385),
.A2(n_41),
.B(n_43),
.Y(n_435)
);

OAI21x1_ASAP7_75t_L g436 ( 
.A1(n_399),
.A2(n_44),
.B(n_45),
.Y(n_436)
);

O2A1O1Ixp33_ASAP7_75t_L g437 ( 
.A1(n_400),
.A2(n_47),
.B(n_48),
.C(n_53),
.Y(n_437)
);

CKINVDCx11_ASAP7_75t_R g438 ( 
.A(n_369),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_398),
.B(n_57),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_388),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_375),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_L g442 ( 
.A1(n_441),
.A2(n_376),
.B1(n_409),
.B2(n_407),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_L g443 ( 
.A1(n_416),
.A2(n_403),
.B1(n_375),
.B2(n_390),
.Y(n_443)
);

OAI21xp33_ASAP7_75t_L g444 ( 
.A1(n_413),
.A2(n_406),
.B(n_408),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_421),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_427),
.A2(n_378),
.B1(n_386),
.B2(n_395),
.Y(n_446)
);

AO31x2_ASAP7_75t_L g447 ( 
.A1(n_423),
.A2(n_399),
.A3(n_405),
.B(n_368),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_L g448 ( 
.A1(n_416),
.A2(n_403),
.B1(n_401),
.B2(n_391),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_410),
.Y(n_449)
);

AOI221xp5_ASAP7_75t_L g450 ( 
.A1(n_414),
.A2(n_379),
.B1(n_403),
.B2(n_371),
.C(n_391),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_431),
.B(n_391),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_424),
.A2(n_392),
.B(n_60),
.Y(n_452)
);

AOI221xp5_ASAP7_75t_L g453 ( 
.A1(n_414),
.A2(n_59),
.B1(n_63),
.B2(n_65),
.C(n_66),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_410),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_422),
.Y(n_455)
);

OAI221xp5_ASAP7_75t_L g456 ( 
.A1(n_431),
.A2(n_68),
.B1(n_71),
.B2(n_75),
.C(n_76),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_438),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_SL g458 ( 
.A1(n_434),
.A2(n_77),
.B1(n_82),
.B2(n_87),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_440),
.B(n_91),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_429),
.B(n_150),
.Y(n_460)
);

BUFx8_ASAP7_75t_L g461 ( 
.A(n_411),
.Y(n_461)
);

INVx5_ASAP7_75t_L g462 ( 
.A(n_427),
.Y(n_462)
);

OAI21x1_ASAP7_75t_L g463 ( 
.A1(n_415),
.A2(n_92),
.B(n_93),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_449),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_462),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_442),
.B(n_438),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_460),
.B(n_430),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_462),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_455),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_454),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_443),
.B(n_430),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_445),
.B(n_417),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_450),
.B(n_424),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_457),
.B(n_439),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_451),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_461),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_459),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_444),
.B(n_439),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_462),
.B(n_435),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_447),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_447),
.Y(n_481)
);

AOI211xp5_ASAP7_75t_L g482 ( 
.A1(n_474),
.A2(n_437),
.B(n_453),
.C(n_432),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_466),
.B(n_448),
.Y(n_483)
);

OAI31xp33_ASAP7_75t_L g484 ( 
.A1(n_478),
.A2(n_456),
.A3(n_446),
.B(n_437),
.Y(n_484)
);

NAND2xp33_ASAP7_75t_SL g485 ( 
.A(n_478),
.B(n_458),
.Y(n_485)
);

INVxp67_ASAP7_75t_SL g486 ( 
.A(n_464),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_467),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g488 ( 
.A(n_476),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_464),
.B(n_470),
.Y(n_489)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_470),
.B(n_447),
.Y(n_490)
);

NAND3xp33_ASAP7_75t_L g491 ( 
.A(n_472),
.B(n_435),
.C(n_425),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_469),
.B(n_425),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_471),
.B(n_420),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_480),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_468),
.B(n_433),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_475),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_481),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_475),
.B(n_420),
.Y(n_498)
);

AOI221x1_ASAP7_75t_L g499 ( 
.A1(n_479),
.A2(n_428),
.B1(n_452),
.B2(n_419),
.C(n_436),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_473),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_487),
.B(n_468),
.Y(n_501)
);

NAND4xp25_ASAP7_75t_SL g502 ( 
.A(n_482),
.B(n_484),
.C(n_491),
.D(n_483),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_489),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_496),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_497),
.Y(n_505)
);

NOR2xp67_ASAP7_75t_L g506 ( 
.A(n_500),
.B(n_479),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_486),
.B(n_465),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_488),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_497),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_486),
.B(n_465),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_495),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_490),
.B(n_473),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_493),
.B(n_477),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_492),
.B(n_465),
.Y(n_514)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_494),
.B(n_419),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_494),
.Y(n_516)
);

OR2x2_ASAP7_75t_L g517 ( 
.A(n_498),
.B(n_418),
.Y(n_517)
);

NAND3xp33_ASAP7_75t_L g518 ( 
.A(n_506),
.B(n_485),
.C(n_499),
.Y(n_518)
);

OAI31xp33_ASAP7_75t_L g519 ( 
.A1(n_502),
.A2(n_485),
.A3(n_498),
.B(n_495),
.Y(n_519)
);

OAI22xp33_ASAP7_75t_L g520 ( 
.A1(n_512),
.A2(n_495),
.B1(n_412),
.B2(n_463),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_504),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_506),
.B(n_426),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_507),
.B(n_94),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_505),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_503),
.B(n_95),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_519),
.B(n_510),
.Y(n_526)
);

AOI32xp33_ASAP7_75t_L g527 ( 
.A1(n_520),
.A2(n_502),
.A3(n_501),
.B1(n_525),
.B2(n_518),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_523),
.B(n_508),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_521),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_526),
.A2(n_514),
.B1(n_508),
.B2(n_511),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_527),
.B(n_513),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_529),
.Y(n_532)
);

NAND4xp75_ASAP7_75t_L g533 ( 
.A(n_531),
.B(n_528),
.C(n_522),
.D(n_516),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_530),
.B(n_517),
.Y(n_534)
);

OAI211xp5_ASAP7_75t_L g535 ( 
.A1(n_532),
.A2(n_522),
.B(n_515),
.C(n_524),
.Y(n_535)
);

NOR3xp33_ASAP7_75t_L g536 ( 
.A(n_533),
.B(n_509),
.C(n_100),
.Y(n_536)
);

O2A1O1Ixp33_ASAP7_75t_L g537 ( 
.A1(n_535),
.A2(n_509),
.B(n_101),
.C(n_107),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_534),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_98),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_537),
.A2(n_108),
.B(n_109),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_536),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_541),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_542)
);

NOR3xp33_ASAP7_75t_L g543 ( 
.A(n_539),
.B(n_114),
.C(n_121),
.Y(n_543)
);

NAND3xp33_ASAP7_75t_L g544 ( 
.A(n_543),
.B(n_540),
.C(n_124),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_542),
.Y(n_545)
);

AO22x1_ASAP7_75t_L g546 ( 
.A1(n_545),
.A2(n_122),
.B1(n_126),
.B2(n_128),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_546),
.B(n_544),
.Y(n_547)
);

AOI21xp33_ASAP7_75t_SL g548 ( 
.A1(n_546),
.A2(n_129),
.B(n_130),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_547),
.A2(n_131),
.B1(n_132),
.B2(n_136),
.Y(n_549)
);

AO21x1_ASAP7_75t_L g550 ( 
.A1(n_548),
.A2(n_138),
.B(n_142),
.Y(n_550)
);

AOI221xp5_ASAP7_75t_L g551 ( 
.A1(n_550),
.A2(n_143),
.B1(n_145),
.B2(n_147),
.C(n_148),
.Y(n_551)
);

NOR3xp33_ASAP7_75t_L g552 ( 
.A(n_551),
.B(n_549),
.C(n_149),
.Y(n_552)
);


endmodule