module fake_netlist_1_9172_n_38 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_38);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
BUFx3_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_4), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_6), .Y(n_13) );
NOR2xp33_ASAP7_75t_R g14 ( .A(n_0), .B(n_2), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_7), .Y(n_15) );
NAND2xp33_ASAP7_75t_SL g16 ( .A(n_4), .B(n_8), .Y(n_16) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_8), .Y(n_17) );
O2A1O1Ixp5_ASAP7_75t_L g18 ( .A1(n_16), .A2(n_0), .B(n_1), .C(n_2), .Y(n_18) );
AOI21xp5_ASAP7_75t_L g19 ( .A1(n_11), .A2(n_0), .B(n_1), .Y(n_19) );
INVx5_ASAP7_75t_L g20 ( .A(n_11), .Y(n_20) );
O2A1O1Ixp33_ASAP7_75t_L g21 ( .A1(n_17), .A2(n_1), .B(n_2), .C(n_3), .Y(n_21) );
AOI22xp33_ASAP7_75t_L g22 ( .A1(n_11), .A2(n_3), .B1(n_5), .B2(n_7), .Y(n_22) );
INVxp67_ASAP7_75t_L g23 ( .A(n_19), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_20), .Y(n_24) );
OR2x2_ASAP7_75t_L g25 ( .A(n_22), .B(n_17), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_23), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
NOR2xp33_ASAP7_75t_L g28 ( .A(n_25), .B(n_13), .Y(n_28) );
OAI211xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_21), .B(n_14), .C(n_16), .Y(n_29) );
NAND2xp5_ASAP7_75t_SL g30 ( .A(n_26), .B(n_18), .Y(n_30) );
OAI211xp5_ASAP7_75t_SL g31 ( .A1(n_29), .A2(n_27), .B(n_26), .C(n_12), .Y(n_31) );
OA21x2_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_24), .B(n_13), .Y(n_32) );
AOI222xp33_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_12), .B1(n_15), .B2(n_11), .C1(n_14), .C2(n_20), .Y(n_33) );
NAND3xp33_ASAP7_75t_L g34 ( .A(n_32), .B(n_15), .C(n_11), .Y(n_34) );
NAND4xp25_ASAP7_75t_L g35 ( .A(n_32), .B(n_5), .C(n_9), .D(n_10), .Y(n_35) );
OAI22xp5_ASAP7_75t_SL g36 ( .A1(n_34), .A2(n_32), .B1(n_10), .B2(n_9), .Y(n_36) );
OAI22xp5_ASAP7_75t_L g37 ( .A1(n_33), .A2(n_20), .B1(n_12), .B2(n_34), .Y(n_37) );
AOI22xp5_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_20), .B1(n_35), .B2(n_36), .Y(n_38) );
endmodule