module fake_jpeg_9812_n_48 (n_3, n_2, n_1, n_0, n_4, n_5, n_48);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_48;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

OR2x2_ASAP7_75t_L g8 ( 
.A(n_2),
.B(n_3),
.Y(n_8)
);

INVx13_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_2),
.B(n_5),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx2_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_8),
.B(n_0),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_15),
.B(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_0),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_18),
.A2(n_22),
.B(n_1),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_12),
.A2(n_13),
.B1(n_9),
.B2(n_14),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_19),
.A2(n_14),
.B1(n_6),
.B2(n_9),
.Y(n_24)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_21),
.B1(n_23),
.B2(n_6),
.Y(n_25)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_27),
.C(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_20),
.A2(n_21),
.B1(n_19),
.B2(n_23),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_18),
.A2(n_13),
.B1(n_7),
.B2(n_11),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_29),
.B(n_22),
.Y(n_31)
);

NAND3xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_34),
.C(n_24),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_22),
.Y(n_34)
);

AOI21x1_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_11),
.B(n_4),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_30),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_27),
.C(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_37),
.B(n_4),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_32),
.A2(n_17),
.B1(n_28),
.B2(n_22),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_38),
.A2(n_11),
.B1(n_28),
.B2(n_4),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_41),
.C(n_36),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_42),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_39),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_47),
.A2(n_37),
.B1(n_45),
.B2(n_5),
.Y(n_48)
);


endmodule