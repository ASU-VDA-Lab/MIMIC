module fake_netlist_1_8912_n_25 (n_1, n_2, n_4, n_3, n_5, n_0, n_25);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_25;
wire n_20;
wire n_23;
wire n_8;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_6;
wire n_7;
BUFx6f_ASAP7_75t_L g6 ( .A(n_5), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_4), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_2), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_2), .Y(n_9) );
BUFx2_ASAP7_75t_L g10 ( .A(n_1), .Y(n_10) );
AND2x2_ASAP7_75t_L g11 ( .A(n_0), .B(n_3), .Y(n_11) );
INVx2_ASAP7_75t_SL g12 ( .A(n_0), .Y(n_12) );
AND2x2_ASAP7_75t_L g13 ( .A(n_10), .B(n_1), .Y(n_13) );
OAI21x1_ASAP7_75t_L g14 ( .A1(n_7), .A2(n_11), .B(n_9), .Y(n_14) );
AO31x2_ASAP7_75t_L g15 ( .A1(n_9), .A2(n_8), .A3(n_12), .B(n_6), .Y(n_15) );
INVx4_ASAP7_75t_L g16 ( .A(n_6), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_14), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_15), .Y(n_18) );
AND2x2_ASAP7_75t_L g19 ( .A(n_13), .B(n_6), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_17), .Y(n_21) );
NOR2xp33_ASAP7_75t_L g22 ( .A(n_20), .B(n_18), .Y(n_22) );
NAND2x1p5_ASAP7_75t_L g23 ( .A(n_22), .B(n_21), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
AOI21xp5_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_16), .B(n_15), .Y(n_25) );
endmodule