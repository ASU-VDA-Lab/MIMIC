module fake_jpeg_31855_n_332 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g83 ( 
.A(n_42),
.Y(n_83)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_25),
.Y(n_44)
);

CKINVDCx12_ASAP7_75t_R g87 ( 
.A(n_44),
.Y(n_87)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_32),
.B(n_10),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_68),
.Y(n_84)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

CKINVDCx6p67_ASAP7_75t_R g114 ( 
.A(n_48),
.Y(n_114)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_50),
.Y(n_120)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_51),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_59),
.Y(n_79)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx5_ASAP7_75t_SL g92 ( 
.A(n_54),
.Y(n_92)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_22),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_69),
.Y(n_85)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_64),
.Y(n_98)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_10),
.Y(n_68)
);

INVx6_ASAP7_75t_SL g69 ( 
.A(n_37),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_15),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_72),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_23),
.B(n_9),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_29),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_37),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_74),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_16),
.B(n_9),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_76),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_35),
.B1(n_18),
.B2(n_33),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_86),
.A2(n_97),
.B1(n_105),
.B2(n_126),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_88),
.B(n_125),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_21),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_91),
.B(n_95),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_55),
.B(n_16),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_93),
.B(n_100),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_21),
.Y(n_95)
);

AO22x2_ASAP7_75t_L g97 ( 
.A1(n_60),
.A2(n_39),
.B1(n_35),
.B2(n_18),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_66),
.A2(n_39),
.B1(n_24),
.B2(n_33),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_99),
.A2(n_102),
.B1(n_117),
.B2(n_119),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_48),
.B(n_29),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_38),
.B1(n_28),
.B2(n_23),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_54),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_107),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_43),
.A2(n_38),
.B1(n_28),
.B2(n_24),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_54),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_59),
.B(n_27),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_108),
.B(n_113),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_53),
.B(n_27),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_110),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_59),
.B(n_7),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_58),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_116),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_45),
.B(n_7),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_11),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_115),
.B(n_118),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_53),
.B(n_2),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_64),
.A2(n_0),
.B1(n_4),
.B2(n_6),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_6),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_62),
.A2(n_0),
.B1(n_6),
.B2(n_12),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g125 ( 
.A1(n_42),
.A2(n_12),
.B(n_13),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_75),
.A2(n_65),
.B1(n_63),
.B2(n_56),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_48),
.A2(n_0),
.B1(n_12),
.B2(n_13),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_117),
.B1(n_119),
.B2(n_83),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_87),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_153),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_14),
.C(n_78),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_134),
.B(n_156),
.Y(n_203)
);

INVx4_ASAP7_75t_SL g136 ( 
.A(n_114),
.Y(n_136)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_136),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_86),
.B(n_14),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_139),
.B(n_140),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_86),
.B(n_97),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_96),
.B(n_88),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_141),
.B(n_150),
.Y(n_185)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_142),
.Y(n_198)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

BUFx4f_ASAP7_75t_SL g197 ( 
.A(n_143),
.Y(n_197)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_144),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_84),
.B(n_86),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_145),
.Y(n_212)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_146),
.Y(n_204)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_147),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_97),
.B(n_105),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_149),
.B(n_152),
.Y(n_190)
);

FAx1_ASAP7_75t_SL g150 ( 
.A(n_99),
.B(n_97),
.CI(n_78),
.CON(n_150),
.SN(n_150)
);

AND2x4_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_127),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

INVx3_ASAP7_75t_SL g154 ( 
.A(n_104),
.Y(n_154)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_94),
.B1(n_112),
.B2(n_135),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_90),
.B(n_129),
.C(n_123),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_90),
.B(n_123),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_163),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_79),
.Y(n_159)
);

INVxp33_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_77),
.Y(n_160)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_104),
.A2(n_82),
.B1(n_92),
.B2(n_126),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_161),
.A2(n_170),
.B1(n_140),
.B2(n_152),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_77),
.Y(n_162)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_85),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_164),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_106),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_166),
.Y(n_194)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_81),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_81),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_168),
.Y(n_200)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_98),
.A2(n_122),
.B1(n_83),
.B2(n_126),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_170),
.A2(n_149),
.B(n_174),
.Y(n_186)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_173),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_121),
.B(n_122),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_121),
.B(n_94),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_175),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_92),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_181),
.A2(n_183),
.B1(n_186),
.B2(n_193),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_145),
.A2(n_112),
.B1(n_137),
.B2(n_150),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_130),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_151),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_188),
.A2(n_142),
.B1(n_146),
.B2(n_154),
.Y(n_219)
);

AO22x1_ASAP7_75t_L g189 ( 
.A1(n_137),
.A2(n_150),
.B1(n_139),
.B2(n_152),
.Y(n_189)
);

AO22x1_ASAP7_75t_L g215 ( 
.A1(n_189),
.A2(n_183),
.B1(n_186),
.B2(n_184),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_137),
.A2(n_152),
.B1(n_161),
.B2(n_176),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_134),
.B(n_157),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_201),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_163),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_156),
.B(n_159),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_207),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_133),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_158),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_178),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_213),
.Y(n_246)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_214),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_215),
.B(n_226),
.Y(n_262)
);

NOR4xp25_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_131),
.C(n_173),
.D(n_136),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_216),
.Y(n_253)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_217),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_219),
.A2(n_196),
.B1(n_202),
.B2(n_204),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_153),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_221),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_147),
.B1(n_162),
.B2(n_160),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_177),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_225),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_200),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_223),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_153),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_227),
.Y(n_249)
);

AND2x6_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_143),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_184),
.B(n_189),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_195),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_211),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_231),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_181),
.A2(n_190),
.B1(n_212),
.B2(n_195),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_191),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_207),
.Y(n_231)
);

AND2x6_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_203),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_233),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_205),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_206),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_236),
.Y(n_255)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_180),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_235),
.B(n_240),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_197),
.B(n_182),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_188),
.A2(n_180),
.B1(n_202),
.B2(n_198),
.Y(n_237)
);

BUFx4f_ASAP7_75t_SL g247 ( 
.A(n_237),
.Y(n_247)
);

NOR2xp67_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_197),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_230),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_210),
.B(n_178),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_241),
.B(n_209),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_215),
.A2(n_210),
.B(n_196),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_243),
.A2(n_263),
.B(n_215),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_191),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_226),
.C(n_220),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_254),
.A2(n_221),
.B1(n_217),
.B2(n_214),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_258),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_218),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_219),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_241),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_209),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_264),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_197),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_240),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_213),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_266),
.B(n_271),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_267),
.A2(n_279),
.B(n_280),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_218),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_268),
.B(n_273),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_252),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_272),
.A2(n_245),
.B1(n_256),
.B2(n_264),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_232),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_257),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_274),
.B(n_276),
.Y(n_293)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_275),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_252),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_277),
.B(n_278),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_239),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_243),
.A2(n_225),
.B(n_224),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_246),
.B(n_223),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_281),
.B(n_249),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_235),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_265),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_229),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_283),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_246),
.A2(n_244),
.B1(n_245),
.B2(n_242),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_284),
.A2(n_253),
.B1(n_279),
.B2(n_254),
.Y(n_289)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_285),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_255),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_286),
.B(n_292),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_280),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_291),
.A2(n_274),
.B1(n_262),
.B2(n_260),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_279),
.A2(n_253),
.B1(n_247),
.B2(n_262),
.Y(n_292)
);

NAND3xp33_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_216),
.C(n_269),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_249),
.Y(n_297)
);

AO21x1_ASAP7_75t_L g308 ( 
.A1(n_297),
.A2(n_270),
.B(n_267),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_273),
.C(n_268),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_301),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_278),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_307),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g303 ( 
.A(n_288),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_303),
.B(n_297),
.Y(n_318)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_304),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_309),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_290),
.A2(n_295),
.B(n_287),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_308),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_276),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_291),
.A2(n_247),
.B1(n_260),
.B2(n_272),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_298),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_313),
.B(n_317),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_298),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_318),
.A2(n_285),
.B(n_270),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_320),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_299),
.C(n_307),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_314),
.A2(n_289),
.B1(n_315),
.B2(n_312),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_321),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_SL g322 ( 
.A(n_315),
.B(n_290),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_322),
.A2(n_311),
.B(n_300),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_292),
.B1(n_308),
.B2(n_247),
.Y(n_324)
);

A2O1A1Ixp33_ASAP7_75t_SL g328 ( 
.A1(n_324),
.A2(n_247),
.B(n_326),
.C(n_327),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_325),
.A2(n_316),
.B(n_320),
.Y(n_329)
);

OAI21x1_ASAP7_75t_L g330 ( 
.A1(n_328),
.A2(n_329),
.B(n_326),
.Y(n_330)
);

AOI21x1_ASAP7_75t_SL g331 ( 
.A1(n_330),
.A2(n_248),
.B(n_198),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_248),
.Y(n_332)
);


endmodule