module real_aes_1067_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_769;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_756;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g238 ( .A(n_0), .B(n_159), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_1), .B(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_2), .B(n_143), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_3), .B(n_161), .Y(n_489) );
INVx1_ASAP7_75t_L g150 ( .A(n_4), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_5), .B(n_143), .Y(n_142) );
NAND2xp33_ASAP7_75t_SL g229 ( .A(n_6), .B(n_149), .Y(n_229) );
INVx1_ASAP7_75t_L g210 ( .A(n_7), .Y(n_210) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_8), .Y(n_113) );
AND2x2_ASAP7_75t_L g137 ( .A(n_9), .B(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g491 ( .A(n_10), .B(n_200), .Y(n_491) );
AND2x2_ASAP7_75t_L g499 ( .A(n_11), .B(n_226), .Y(n_499) );
INVx2_ASAP7_75t_L g139 ( .A(n_12), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_13), .B(n_161), .Y(n_508) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_14), .Y(n_106) );
AOI221x1_ASAP7_75t_L g223 ( .A1(n_15), .A2(n_152), .B1(n_224), .B2(n_226), .C(n_228), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_16), .B(n_143), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_17), .B(n_143), .Y(n_522) );
INVx1_ASAP7_75t_L g109 ( .A(n_18), .Y(n_109) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_19), .A2(n_87), .B1(n_143), .B2(n_211), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_20), .A2(n_769), .B1(n_771), .B2(n_774), .Y(n_770) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_21), .A2(n_152), .B(n_157), .Y(n_151) );
AOI221xp5_ASAP7_75t_SL g187 ( .A1(n_22), .A2(n_37), .B1(n_143), .B2(n_152), .C(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_23), .B(n_159), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g788 ( .A(n_24), .Y(n_788) );
OR2x2_ASAP7_75t_L g140 ( .A(n_25), .B(n_86), .Y(n_140) );
OA21x2_ASAP7_75t_L g201 ( .A1(n_25), .A2(n_86), .B(n_139), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_26), .B(n_161), .Y(n_199) );
INVxp67_ASAP7_75t_L g222 ( .A(n_27), .Y(n_222) );
AND2x2_ASAP7_75t_L g183 ( .A(n_28), .B(n_173), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_29), .A2(n_152), .B(n_237), .Y(n_236) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_30), .A2(n_226), .B(n_504), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_31), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_32), .B(n_161), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_33), .A2(n_152), .B(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_34), .B(n_161), .Y(n_517) );
AND2x2_ASAP7_75t_L g149 ( .A(n_35), .B(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g153 ( .A(n_35), .B(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g218 ( .A(n_35), .Y(n_218) );
OR2x6_ASAP7_75t_L g107 ( .A(n_36), .B(n_108), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_38), .B(n_143), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_39), .A2(n_79), .B1(n_152), .B2(n_216), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_40), .B(n_161), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_41), .B(n_143), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_42), .B(n_159), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_43), .A2(n_152), .B(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g241 ( .A(n_44), .B(n_173), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_45), .B(n_159), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_46), .B(n_173), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_47), .B(n_143), .Y(n_505) );
INVx1_ASAP7_75t_L g146 ( .A(n_48), .Y(n_146) );
INVx1_ASAP7_75t_L g156 ( .A(n_48), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_49), .B(n_161), .Y(n_497) );
AND2x2_ASAP7_75t_L g533 ( .A(n_50), .B(n_173), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_51), .B(n_143), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_52), .B(n_159), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_53), .B(n_159), .Y(n_516) );
AND2x2_ASAP7_75t_L g174 ( .A(n_54), .B(n_173), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_55), .B(n_143), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_56), .B(n_161), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_57), .B(n_143), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_58), .A2(n_152), .B(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_59), .B(n_159), .Y(n_170) );
AND2x2_ASAP7_75t_SL g202 ( .A(n_60), .B(n_138), .Y(n_202) );
AND2x2_ASAP7_75t_L g528 ( .A(n_61), .B(n_138), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_62), .A2(n_152), .B(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_63), .B(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_SL g254 ( .A(n_64), .B(n_200), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_65), .B(n_159), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_66), .B(n_159), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_67), .A2(n_90), .B1(n_152), .B2(n_216), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_68), .B(n_161), .Y(n_525) );
INVx1_ASAP7_75t_L g148 ( .A(n_69), .Y(n_148) );
INVx1_ASAP7_75t_L g154 ( .A(n_69), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_70), .B(n_159), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g781 ( .A1(n_71), .A2(n_130), .B1(n_782), .B2(n_783), .Y(n_781) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_71), .Y(n_782) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_72), .A2(n_152), .B(n_537), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_73), .A2(n_152), .B(n_479), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_74), .A2(n_152), .B(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g519 ( .A(n_75), .B(n_138), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_76), .B(n_173), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_77), .B(n_143), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_78), .A2(n_81), .B1(n_143), .B2(n_211), .Y(n_252) );
INVx1_ASAP7_75t_L g110 ( .A(n_80), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_82), .B(n_159), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_83), .B(n_159), .Y(n_190) );
AND2x2_ASAP7_75t_L g482 ( .A(n_84), .B(n_200), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_85), .A2(n_152), .B(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_88), .B(n_161), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_89), .A2(n_152), .B(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_91), .B(n_161), .Y(n_480) );
INVxp67_ASAP7_75t_L g225 ( .A(n_92), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_93), .B(n_143), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_94), .B(n_161), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_95), .A2(n_152), .B(n_197), .Y(n_196) );
BUFx2_ASAP7_75t_L g527 ( .A(n_96), .Y(n_527) );
BUFx2_ASAP7_75t_L g119 ( .A(n_97), .Y(n_119) );
BUFx2_ASAP7_75t_SL g779 ( .A(n_97), .Y(n_779) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_98), .Y(n_769) );
AOI21xp33_ASAP7_75t_SL g99 ( .A1(n_100), .A2(n_114), .B(n_787), .Y(n_99) );
INVx2_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
INVx4_ASAP7_75t_R g101 ( .A(n_102), .Y(n_101) );
INVx2_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g789 ( .A(n_103), .Y(n_789) );
NAND2xp5_ASAP7_75t_SL g103 ( .A(n_104), .B(n_111), .Y(n_103) );
INVx3_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
BUFx2_ASAP7_75t_L g775 ( .A(n_105), .Y(n_775) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_106), .B(n_125), .Y(n_124) );
AND2x6_ASAP7_75t_SL g467 ( .A(n_106), .B(n_107), .Y(n_467) );
OR2x6_ASAP7_75t_SL g768 ( .A(n_106), .B(n_125), .Y(n_768) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_107), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OA21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_127), .B(n_776), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_120), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVxp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g780 ( .A1(n_121), .A2(n_781), .B(n_784), .Y(n_780) );
NOR2xp33_ASAP7_75t_SL g121 ( .A(n_122), .B(n_126), .Y(n_121) );
HB1xp67_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
BUFx3_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
BUFx2_ASAP7_75t_R g786 ( .A(n_124), .Y(n_786) );
OAI21xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_769), .B(n_770), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OAI22x1_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_464), .B1(n_468), .B2(n_768), .Y(n_129) );
INVx4_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_131), .A2(n_464), .B1(n_469), .B2(n_772), .Y(n_771) );
HB1xp67_ASAP7_75t_L g783 ( .A(n_131), .Y(n_783) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_375), .Y(n_131) );
NOR3xp33_ASAP7_75t_L g132 ( .A(n_133), .B(n_297), .C(n_347), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_264), .Y(n_133) );
AOI221xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_184), .B1(n_203), .B2(n_246), .C(n_256), .Y(n_134) );
INVx1_ASAP7_75t_SL g346 ( .A(n_135), .Y(n_346) );
AND2x4_ASAP7_75t_SL g135 ( .A(n_136), .B(n_164), .Y(n_135) );
INVx2_ASAP7_75t_L g268 ( .A(n_136), .Y(n_268) );
OR2x2_ASAP7_75t_L g290 ( .A(n_136), .B(n_281), .Y(n_290) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_136), .Y(n_305) );
INVx5_ASAP7_75t_L g312 ( .A(n_136), .Y(n_312) );
AND2x4_ASAP7_75t_L g318 ( .A(n_136), .B(n_176), .Y(n_318) );
AND2x2_ASAP7_75t_SL g321 ( .A(n_136), .B(n_248), .Y(n_321) );
OR2x2_ASAP7_75t_L g330 ( .A(n_136), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g337 ( .A(n_136), .B(n_165), .Y(n_337) );
AND2x2_ASAP7_75t_L g438 ( .A(n_136), .B(n_175), .Y(n_438) );
OR2x6_ASAP7_75t_L g136 ( .A(n_137), .B(n_141), .Y(n_136) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_138), .Y(n_173) );
AND2x2_ASAP7_75t_SL g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x4_ASAP7_75t_L g163 ( .A(n_139), .B(n_140), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_151), .B(n_163), .Y(n_141) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_149), .Y(n_143) );
INVx1_ASAP7_75t_L g230 ( .A(n_144), .Y(n_230) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
AND2x6_ASAP7_75t_L g159 ( .A(n_145), .B(n_154), .Y(n_159) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x4_ASAP7_75t_L g161 ( .A(n_147), .B(n_156), .Y(n_161) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx5_ASAP7_75t_L g162 ( .A(n_149), .Y(n_162) );
AND2x2_ASAP7_75t_L g155 ( .A(n_150), .B(n_156), .Y(n_155) );
HB1xp67_ASAP7_75t_L g214 ( .A(n_150), .Y(n_214) );
AND2x6_ASAP7_75t_L g152 ( .A(n_153), .B(n_155), .Y(n_152) );
BUFx3_ASAP7_75t_L g215 ( .A(n_153), .Y(n_215) );
INVx2_ASAP7_75t_L g220 ( .A(n_154), .Y(n_220) );
AND2x4_ASAP7_75t_L g216 ( .A(n_155), .B(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g213 ( .A(n_156), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_160), .B(n_162), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_159), .B(n_527), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_162), .A2(n_169), .B(n_170), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_162), .A2(n_180), .B(n_181), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_162), .A2(n_189), .B(n_190), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_162), .A2(n_198), .B(n_199), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_162), .A2(n_238), .B(n_239), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_162), .A2(n_480), .B(n_481), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_162), .A2(n_488), .B(n_489), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_162), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_162), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_162), .A2(n_516), .B(n_517), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_162), .A2(n_525), .B(n_526), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_162), .A2(n_538), .B(n_539), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_163), .B(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_163), .B(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_163), .B(n_225), .Y(n_224) );
NOR3xp33_ASAP7_75t_L g228 ( .A(n_163), .B(n_229), .C(n_230), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_163), .A2(n_505), .B(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_163), .A2(n_535), .B(n_536), .Y(n_534) );
INVx3_ASAP7_75t_SL g289 ( .A(n_164), .Y(n_289) );
AND2x2_ASAP7_75t_L g333 ( .A(n_164), .B(n_248), .Y(n_333) );
OAI21xp5_ASAP7_75t_L g336 ( .A1(n_164), .A2(n_337), .B(n_338), .Y(n_336) );
AND2x2_ASAP7_75t_L g374 ( .A(n_164), .B(n_312), .Y(n_374) );
AND2x4_ASAP7_75t_L g164 ( .A(n_165), .B(n_175), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_165), .B(n_176), .Y(n_255) );
OR2x2_ASAP7_75t_L g259 ( .A(n_165), .B(n_176), .Y(n_259) );
INVx1_ASAP7_75t_L g267 ( .A(n_165), .Y(n_267) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_165), .Y(n_279) );
INVx2_ASAP7_75t_L g287 ( .A(n_165), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_165), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g396 ( .A(n_165), .B(n_281), .Y(n_396) );
AND2x2_ASAP7_75t_L g411 ( .A(n_165), .B(n_248), .Y(n_411) );
AO21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_172), .B(n_174), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_167), .B(n_171), .Y(n_166) );
AO21x2_ASAP7_75t_L g176 ( .A1(n_172), .A2(n_177), .B(n_183), .Y(n_176) );
AO21x2_ASAP7_75t_L g331 ( .A1(n_172), .A2(n_177), .B(n_183), .Y(n_331) );
AOI21x1_ASAP7_75t_L g484 ( .A1(n_172), .A2(n_485), .B(n_491), .Y(n_484) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_173), .Y(n_172) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_173), .A2(n_187), .B(n_191), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_173), .A2(n_477), .B(n_478), .Y(n_476) );
AO21x2_ASAP7_75t_L g559 ( .A1(n_173), .A2(n_560), .B(n_561), .Y(n_559) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g280 ( .A(n_176), .B(n_281), .Y(n_280) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_176), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_178), .B(n_182), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_184), .B(n_404), .Y(n_403) );
NOR2x1p5_ASAP7_75t_L g184 ( .A(n_185), .B(n_192), .Y(n_184) );
BUFx3_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g232 ( .A(n_186), .B(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_186), .B(n_193), .Y(n_262) );
INVx1_ASAP7_75t_L g272 ( .A(n_186), .Y(n_272) );
INVx2_ASAP7_75t_L g295 ( .A(n_186), .Y(n_295) );
INVx2_ASAP7_75t_L g301 ( .A(n_186), .Y(n_301) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_186), .Y(n_371) );
OR2x2_ASAP7_75t_L g402 ( .A(n_186), .B(n_193), .Y(n_402) );
OR2x2_ASAP7_75t_L g418 ( .A(n_192), .B(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
AND2x4_ASAP7_75t_SL g206 ( .A(n_193), .B(n_207), .Y(n_206) );
AND2x4_ASAP7_75t_L g244 ( .A(n_193), .B(n_245), .Y(n_244) );
OR2x2_ASAP7_75t_L g282 ( .A(n_193), .B(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g294 ( .A(n_193), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g307 ( .A(n_193), .B(n_273), .Y(n_307) );
OR2x2_ASAP7_75t_L g315 ( .A(n_193), .B(n_207), .Y(n_315) );
INVx2_ASAP7_75t_L g342 ( .A(n_193), .Y(n_342) );
INVx1_ASAP7_75t_L g360 ( .A(n_193), .Y(n_360) );
NOR2xp33_ASAP7_75t_R g393 ( .A(n_193), .B(n_233), .Y(n_393) );
OR2x6_ASAP7_75t_L g193 ( .A(n_194), .B(n_202), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_200), .Y(n_194) );
INVx2_ASAP7_75t_SL g250 ( .A(n_200), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_200), .A2(n_522), .B(n_523), .Y(n_521) );
BUFx4f_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx3_ASAP7_75t_L g227 ( .A(n_201), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_204), .B(n_242), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g284 ( .A1(n_204), .A2(n_285), .B1(n_288), .B2(n_291), .Y(n_284) );
OR2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_231), .Y(n_204) );
INVx1_ASAP7_75t_SL g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g299 ( .A(n_206), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g334 ( .A(n_206), .B(n_335), .Y(n_334) );
AND2x4_ASAP7_75t_L g413 ( .A(n_206), .B(n_391), .Y(n_413) );
INVx3_ASAP7_75t_L g245 ( .A(n_207), .Y(n_245) );
AND2x4_ASAP7_75t_L g273 ( .A(n_207), .B(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_207), .B(n_233), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_207), .B(n_295), .Y(n_340) );
AND2x2_ASAP7_75t_L g345 ( .A(n_207), .B(n_342), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_207), .B(n_232), .Y(n_382) );
INVx1_ASAP7_75t_L g452 ( .A(n_207), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_207), .B(n_370), .Y(n_463) );
AND2x4_ASAP7_75t_L g207 ( .A(n_208), .B(n_223), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_211), .B1(n_216), .B2(n_221), .Y(n_208) );
AND2x4_ASAP7_75t_L g211 ( .A(n_212), .B(n_215), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
NOR2x1p5_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
INVx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx3_ASAP7_75t_L g512 ( .A(n_226), .Y(n_512) );
INVx4_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AOI21x1_ASAP7_75t_L g234 ( .A1(n_227), .A2(n_235), .B(n_241), .Y(n_234) );
AO21x2_ASAP7_75t_L g492 ( .A1(n_227), .A2(n_493), .B(n_499), .Y(n_492) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g243 ( .A(n_233), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_233), .B(n_245), .Y(n_263) );
INVx2_ASAP7_75t_L g274 ( .A(n_233), .Y(n_274) );
AND2x2_ASAP7_75t_L g300 ( .A(n_233), .B(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g316 ( .A(n_233), .B(n_295), .Y(n_316) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_233), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_233), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g405 ( .A(n_233), .Y(n_405) );
INVx3_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_240), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_243), .B(n_272), .Y(n_283) );
AOI221x1_ASAP7_75t_SL g377 ( .A1(n_244), .A2(n_378), .B1(n_381), .B2(n_383), .C(n_387), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_244), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g435 ( .A(n_244), .B(n_300), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_244), .B(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g366 ( .A(n_245), .B(n_294), .Y(n_366) );
AND2x2_ASAP7_75t_L g404 ( .A(n_245), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_255), .Y(n_247) );
AND2x2_ASAP7_75t_L g257 ( .A(n_248), .B(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g352 ( .A(n_248), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_248), .B(n_268), .Y(n_357) );
AND2x4_ASAP7_75t_L g386 ( .A(n_248), .B(n_287), .Y(n_386) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_248), .B(n_318), .Y(n_422) );
OR2x2_ASAP7_75t_L g440 ( .A(n_248), .B(n_371), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_248), .B(n_331), .Y(n_450) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g281 ( .A(n_249), .Y(n_281) );
AOI21x1_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_251), .B(n_254), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
INVx1_ASAP7_75t_L g306 ( .A(n_255), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_255), .A2(n_314), .B1(n_317), .B2(n_319), .Y(n_313) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_260), .Y(n_256) );
INVx2_ASAP7_75t_L g269 ( .A(n_257), .Y(n_269) );
AND2x2_ASAP7_75t_L g408 ( .A(n_258), .B(n_268), .Y(n_408) );
AND2x2_ASAP7_75t_L g454 ( .A(n_258), .B(n_321), .Y(n_454) );
AND2x2_ASAP7_75t_L g459 ( .A(n_258), .B(n_310), .Y(n_459) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AOI32xp33_ASAP7_75t_L g428 ( .A1(n_260), .A2(n_330), .A3(n_410), .B1(n_429), .B2(n_431), .Y(n_428) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
INVx1_ASAP7_75t_L g296 ( .A(n_263), .Y(n_296) );
AOI211xp5_ASAP7_75t_SL g264 ( .A1(n_265), .A2(n_270), .B(n_275), .C(n_284), .Y(n_264) );
OAI21xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_268), .B(n_269), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_267), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_268), .B(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g448 ( .A(n_268), .Y(n_448) );
AND2x2_ASAP7_75t_L g358 ( .A(n_270), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_SL g270 ( .A(n_271), .B(n_273), .Y(n_270) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_271), .Y(n_458) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVxp67_ASAP7_75t_SL g327 ( .A(n_272), .Y(n_327) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_272), .Y(n_427) );
INVx1_ASAP7_75t_L g324 ( .A(n_273), .Y(n_324) );
AND2x2_ASAP7_75t_L g390 ( .A(n_273), .B(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_273), .B(n_401), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_276), .B(n_282), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OAI21xp33_ASAP7_75t_L g356 ( .A1(n_277), .A2(n_357), .B(n_358), .Y(n_356) );
AND2x2_ASAP7_75t_SL g277 ( .A(n_278), .B(n_280), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g286 ( .A(n_281), .B(n_287), .Y(n_286) );
BUFx2_ASAP7_75t_L g310 ( .A(n_281), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_286), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g417 ( .A(n_286), .Y(n_417) );
AND2x2_ASAP7_75t_L g447 ( .A(n_286), .B(n_448), .Y(n_447) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_287), .Y(n_424) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_289), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_SL g364 ( .A(n_290), .Y(n_364) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x4_ASAP7_75t_L g292 ( .A(n_293), .B(n_296), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g323 ( .A(n_294), .B(n_324), .Y(n_323) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_295), .Y(n_391) );
AND2x2_ASAP7_75t_L g400 ( .A(n_296), .B(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_320), .Y(n_297) );
AOI221xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_302), .B1(n_307), .B2(n_308), .C(n_313), .Y(n_298) );
INVx1_ASAP7_75t_L g419 ( .A(n_300), .Y(n_419) );
INVxp33_ASAP7_75t_SL g451 ( .A(n_300), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g397 ( .A1(n_302), .A2(n_398), .B(n_406), .Y(n_397) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_304), .B(n_306), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_306), .B(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g319 ( .A(n_307), .Y(n_319) );
AND2x2_ASAP7_75t_L g354 ( .A(n_307), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g373 ( .A(n_307), .B(n_374), .Y(n_373) );
AOI22xp33_ASAP7_75t_SL g434 ( .A1(n_307), .A2(n_435), .B1(n_436), .B2(n_439), .Y(n_434) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
OR2x2_ASAP7_75t_L g329 ( .A(n_310), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_310), .B(n_318), .Y(n_368) );
AND2x4_ASAP7_75t_L g385 ( .A(n_312), .B(n_331), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_312), .B(n_386), .Y(n_432) );
AND2x2_ASAP7_75t_L g444 ( .A(n_312), .B(n_396), .Y(n_444) );
NAND2xp33_ASAP7_75t_L g429 ( .A(n_314), .B(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx1_ASAP7_75t_SL g372 ( .A(n_315), .Y(n_372) );
INVx1_ASAP7_75t_L g443 ( .A(n_316), .Y(n_443) );
INVx2_ASAP7_75t_SL g395 ( .A(n_318), .Y(n_395) );
AOI211xp5_ASAP7_75t_SL g320 ( .A1(n_321), .A2(n_322), .B(n_325), .C(n_343), .Y(n_320) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OAI211xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_329), .B(n_332), .C(n_336), .Y(n_325) );
OR2x6_ASAP7_75t_SL g326 ( .A(n_327), .B(n_328), .Y(n_326) );
INVx1_ASAP7_75t_L g355 ( .A(n_327), .Y(n_355) );
INVx1_ASAP7_75t_SL g380 ( .A(n_330), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_330), .B(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_335), .B(n_345), .Y(n_344) );
INVx2_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
OAI22xp33_ASAP7_75t_L g421 ( .A1(n_339), .A2(n_422), .B1(n_423), .B2(n_425), .Y(n_421) );
OR2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
OAI211xp5_ASAP7_75t_SL g347 ( .A1(n_348), .A2(n_353), .B(n_356), .C(n_361), .Y(n_347) );
INVxp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AOI221xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_365), .B1(n_367), .B2(n_369), .C(n_373), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AOI222xp33_ASAP7_75t_L g453 ( .A1(n_372), .A2(n_454), .B1(n_455), .B2(n_459), .C1(n_460), .C2(n_462), .Y(n_453) );
INVx2_ASAP7_75t_L g388 ( .A(n_374), .Y(n_388) );
NOR3xp33_ASAP7_75t_L g375 ( .A(n_376), .B(n_414), .C(n_433), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_397), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVxp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_385), .B(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_386), .B(n_448), .Y(n_461) );
OAI22xp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B1(n_392), .B2(n_394), .Y(n_387) );
INVx1_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
INVxp33_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_395), .B(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_403), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_403), .A2(n_407), .B1(n_409), .B2(n_412), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
CKINVDCx16_ASAP7_75t_R g412 ( .A(n_413), .Y(n_412) );
OAI211xp5_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_418), .B(n_420), .C(n_428), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVxp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NAND3xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_441), .C(n_453), .Y(n_433) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OAI21xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_445), .B(n_452), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_449), .B(n_451), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
CKINVDCx11_ASAP7_75t_R g464 ( .A(n_465), .Y(n_464) );
INVx3_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g466 ( .A(n_467), .Y(n_466) );
INVx5_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x4_ASAP7_75t_L g469 ( .A(n_470), .B(n_672), .Y(n_469) );
NOR3xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_597), .C(n_633), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_571), .Y(n_471) );
AOI211xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_500), .B(n_529), .C(n_554), .Y(n_472) );
AND2x2_ASAP7_75t_L g662 ( .A(n_473), .B(n_531), .Y(n_662) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_483), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_474), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g695 ( .A(n_474), .B(n_577), .Y(n_695) );
AND2x2_ASAP7_75t_L g711 ( .A(n_474), .B(n_546), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_474), .B(n_721), .Y(n_720) );
NAND2x1p5_ASAP7_75t_L g744 ( .A(n_474), .B(n_745), .Y(n_744) );
INVx4_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x4_ASAP7_75t_SL g541 ( .A(n_475), .B(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g566 ( .A(n_475), .Y(n_566) );
AND2x2_ASAP7_75t_L g613 ( .A(n_475), .B(n_556), .Y(n_613) );
AND2x2_ASAP7_75t_L g632 ( .A(n_475), .B(n_483), .Y(n_632) );
BUFx2_ASAP7_75t_L g637 ( .A(n_475), .Y(n_637) );
AND2x2_ASAP7_75t_L g681 ( .A(n_475), .B(n_492), .Y(n_681) );
AND2x4_ASAP7_75t_L g753 ( .A(n_475), .B(n_754), .Y(n_753) );
NOR2x1_ASAP7_75t_L g765 ( .A(n_475), .B(n_545), .Y(n_765) );
OR2x6_ASAP7_75t_L g475 ( .A(n_476), .B(n_482), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_483), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g684 ( .A(n_483), .Y(n_684) );
BUFx2_ASAP7_75t_L g733 ( .A(n_483), .Y(n_733) );
INVx1_ASAP7_75t_L g755 ( .A(n_483), .Y(n_755) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_492), .Y(n_483) );
INVx3_ASAP7_75t_L g542 ( .A(n_484), .Y(n_542) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_484), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_486), .B(n_490), .Y(n_485) );
INVx2_ASAP7_75t_L g545 ( .A(n_492), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_492), .B(n_542), .Y(n_546) );
INVx2_ASAP7_75t_L g621 ( .A(n_492), .Y(n_621) );
OR2x2_ASAP7_75t_L g628 ( .A(n_492), .B(n_577), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_498), .Y(n_493) );
AND2x2_ASAP7_75t_L g583 ( .A(n_500), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g617 ( .A(n_500), .B(n_580), .Y(n_617) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_510), .Y(n_500) );
AND2x2_ASAP7_75t_L g653 ( .A(n_501), .B(n_552), .Y(n_653) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g610 ( .A(n_502), .B(n_511), .Y(n_610) );
AND2x2_ASAP7_75t_L g729 ( .A(n_502), .B(n_520), .Y(n_729) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g551 ( .A(n_503), .Y(n_551) );
INVx1_ASAP7_75t_L g569 ( .A(n_503), .Y(n_569) );
AND2x2_ASAP7_75t_L g625 ( .A(n_503), .B(n_511), .Y(n_625) );
AND2x2_ASAP7_75t_L g630 ( .A(n_503), .B(n_532), .Y(n_630) );
OR2x2_ASAP7_75t_L g693 ( .A(n_503), .B(n_520), .Y(n_693) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_503), .Y(n_702) );
AND2x2_ASAP7_75t_L g531 ( .A(n_510), .B(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g570 ( .A(n_510), .Y(n_570) );
NOR2x1_ASAP7_75t_SL g510 ( .A(n_511), .B(n_520), .Y(n_510) );
AO21x1_ASAP7_75t_SL g511 ( .A1(n_512), .A2(n_513), .B(n_519), .Y(n_511) );
AO21x2_ASAP7_75t_L g553 ( .A1(n_512), .A2(n_513), .B(n_519), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_518), .Y(n_513) );
AND2x2_ASAP7_75t_L g548 ( .A(n_520), .B(n_549), .Y(n_548) );
INVx2_ASAP7_75t_SL g596 ( .A(n_520), .Y(n_596) );
NAND2x1_ASAP7_75t_L g606 ( .A(n_520), .B(n_532), .Y(n_606) );
OR2x2_ASAP7_75t_L g611 ( .A(n_520), .B(n_549), .Y(n_611) );
BUFx2_ASAP7_75t_L g667 ( .A(n_520), .Y(n_667) );
AND2x2_ASAP7_75t_L g703 ( .A(n_520), .B(n_582), .Y(n_703) );
AND2x2_ASAP7_75t_L g714 ( .A(n_520), .B(n_552), .Y(n_714) );
OR2x6_ASAP7_75t_L g520 ( .A(n_521), .B(n_528), .Y(n_520) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_540), .B1(n_546), .B2(n_547), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_531), .A2(n_711), .B1(n_761), .B2(n_766), .Y(n_760) );
INVx4_ASAP7_75t_L g549 ( .A(n_532), .Y(n_549) );
INVx2_ASAP7_75t_L g580 ( .A(n_532), .Y(n_580) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_532), .Y(n_651) );
OR2x2_ASAP7_75t_L g666 ( .A(n_532), .B(n_552), .Y(n_666) );
OR2x2_ASAP7_75t_SL g692 ( .A(n_532), .B(n_693), .Y(n_692) );
OR2x6_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
AND2x2_ASAP7_75t_SL g540 ( .A(n_541), .B(n_543), .Y(n_540) );
INVx2_ASAP7_75t_SL g573 ( .A(n_541), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_541), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g641 ( .A(n_541), .B(n_589), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_541), .B(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g563 ( .A(n_542), .Y(n_563) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_542), .Y(n_588) );
AND2x2_ASAP7_75t_L g644 ( .A(n_542), .B(n_621), .Y(n_644) );
INVx1_ASAP7_75t_L g754 ( .A(n_542), .Y(n_754) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_544), .B(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_544), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g562 ( .A(n_545), .B(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_546), .B(n_695), .Y(n_694) );
AOI321xp33_ASAP7_75t_L g716 ( .A1(n_547), .A2(n_618), .A3(n_686), .B1(n_717), .B2(n_718), .C(n_722), .Y(n_716) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
INVxp67_ASAP7_75t_SL g615 ( .A(n_548), .Y(n_615) );
AND2x2_ASAP7_75t_L g640 ( .A(n_548), .B(n_569), .Y(n_640) );
AND2x2_ASAP7_75t_L g715 ( .A(n_548), .B(n_625), .Y(n_715) );
INVx1_ASAP7_75t_L g584 ( .A(n_549), .Y(n_584) );
BUFx2_ASAP7_75t_L g594 ( .A(n_549), .Y(n_594) );
NOR2xp67_ASAP7_75t_L g701 ( .A(n_549), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g639 ( .A(n_550), .Y(n_639) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
BUFx2_ASAP7_75t_L g646 ( .A(n_551), .Y(n_646) );
INVx2_ASAP7_75t_L g582 ( .A(n_552), .Y(n_582) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_552), .Y(n_605) );
INVx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AOI21xp33_ASAP7_75t_SL g554 ( .A1(n_555), .A2(n_564), .B(n_567), .Y(n_554) );
NOR2xp67_ASAP7_75t_L g698 ( .A(n_555), .B(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_562), .Y(n_556) );
INVx3_ASAP7_75t_L g589 ( .A(n_557), .Y(n_589) );
AND2x2_ASAP7_75t_L g620 ( .A(n_557), .B(n_621), .Y(n_620) );
AND2x4_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
AND2x4_ASAP7_75t_L g577 ( .A(n_558), .B(n_559), .Y(n_577) );
INVx1_ASAP7_75t_L g660 ( .A(n_562), .Y(n_660) );
INVx1_ASAP7_75t_SL g745 ( .A(n_563), .Y(n_745) );
INVxp33_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_566), .B(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g671 ( .A(n_566), .B(n_628), .Y(n_671) );
OR2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
AND2x2_ASAP7_75t_L g675 ( .A(n_568), .B(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_568), .B(n_690), .Y(n_689) );
INVx3_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_569), .B(n_606), .Y(n_661) );
NOR4xp25_ASAP7_75t_L g756 ( .A(n_569), .B(n_600), .C(n_757), .D(n_758), .Y(n_756) );
OR2x2_ASAP7_75t_L g724 ( .A(n_570), .B(n_725), .Y(n_724) );
AOI221xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_578), .B1(n_583), .B2(n_585), .C(n_590), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
AND2x2_ASAP7_75t_L g599 ( .A(n_574), .B(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g636 ( .A(n_575), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g656 ( .A(n_576), .Y(n_656) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
BUFx3_ASAP7_75t_L g679 ( .A(n_577), .Y(n_679) );
AND2x2_ASAP7_75t_L g686 ( .A(n_577), .B(n_687), .Y(n_686) );
INVxp67_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
OR2x2_ASAP7_75t_L g623 ( .A(n_580), .B(n_624), .Y(n_623) );
INVxp67_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_582), .B(n_596), .Y(n_595) );
INVxp67_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
INVx2_ASAP7_75t_L g600 ( .A(n_587), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_587), .B(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g592 ( .A(n_589), .Y(n_592) );
OAI321xp33_ASAP7_75t_L g704 ( .A1(n_589), .A2(n_697), .A3(n_705), .B1(n_710), .B2(n_712), .C(n_716), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
OR2x2_ASAP7_75t_L g659 ( .A(n_592), .B(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
INVx1_ASAP7_75t_L g759 ( .A(n_595), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_596), .B(n_639), .Y(n_638) );
NAND2xp33_ASAP7_75t_SL g739 ( .A(n_596), .B(n_610), .Y(n_739) );
OAI211xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_601), .B(n_612), .C(n_616), .Y(n_597) );
INVxp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NOR2x1_ASAP7_75t_L g601 ( .A(n_602), .B(n_607), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g708 ( .A(n_605), .Y(n_708) );
INVx3_ASAP7_75t_L g647 ( .A(n_606), .Y(n_647) );
OR2x2_ASAP7_75t_L g750 ( .A(n_606), .B(n_624), .Y(n_750) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_608), .A2(n_692), .B1(n_694), .B2(n_696), .Y(n_691) );
OR2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_SL g690 ( .A(n_611), .Y(n_690) );
OR2x2_ASAP7_75t_L g767 ( .A(n_611), .B(n_624), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AOI21xp5_ASAP7_75t_SL g616 ( .A1(n_617), .A2(n_618), .B(n_622), .Y(n_616) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_620), .B(n_637), .Y(n_736) );
AND2x2_ASAP7_75t_L g742 ( .A(n_620), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g687 ( .A(n_621), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_626), .B1(n_629), .B2(n_631), .Y(n_622) );
A2O1A1Ixp33_ASAP7_75t_L g668 ( .A1(n_624), .A2(n_667), .B(n_669), .C(n_671), .Y(n_668) );
INVx2_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_627), .B(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_627), .B(n_719), .Y(n_741) );
INVx2_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g713 ( .A(n_630), .B(n_714), .Y(n_713) );
INVx2_ASAP7_75t_SL g631 ( .A(n_632), .Y(n_631) );
A2O1A1Ixp33_ASAP7_75t_L g663 ( .A1(n_632), .A2(n_664), .B(n_667), .C(n_668), .Y(n_663) );
NAND3xp33_ASAP7_75t_SL g633 ( .A(n_634), .B(n_648), .C(n_663), .Y(n_633) );
AOI222xp33_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_638), .B1(n_640), .B2(n_641), .C1(n_642), .C2(n_645), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g697 ( .A(n_637), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_637), .B(n_670), .Y(n_723) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_SL g657 ( .A(n_644), .Y(n_657) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
OR2x2_ASAP7_75t_L g762 ( .A(n_646), .B(n_679), .Y(n_762) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_647), .A2(n_738), .B1(n_740), .B2(n_742), .Y(n_737) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_654), .B1(n_658), .B2(n_661), .C(n_662), .Y(n_648) );
INVx2_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AOI21xp5_ASAP7_75t_SL g722 ( .A1(n_655), .A2(n_723), .B(n_724), .Y(n_722) );
OR2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
INVx2_ASAP7_75t_L g670 ( .A(n_656), .Y(n_670) );
AND2x2_ASAP7_75t_L g764 ( .A(n_656), .B(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g748 ( .A(n_660), .Y(n_748) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OR2x2_ASAP7_75t_L g677 ( .A(n_666), .B(n_667), .Y(n_677) );
INVx1_ASAP7_75t_L g730 ( .A(n_666), .Y(n_730) );
NOR3xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_704), .C(n_726), .Y(n_672) );
OAI211xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_678), .B(n_680), .C(n_685), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
OAI21xp33_ASAP7_75t_L g680 ( .A1(n_675), .A2(n_681), .B(n_682), .Y(n_680) );
INVx1_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AOI211xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_688), .B(n_691), .C(n_698), .Y(n_685) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g709 ( .A(n_692), .Y(n_709) );
INVxp67_ASAP7_75t_SL g734 ( .A(n_693), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_695), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g757 ( .A(n_695), .Y(n_757) );
AND2x2_ASAP7_75t_L g747 ( .A(n_697), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g717 ( .A(n_699), .Y(n_717) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_703), .Y(n_700) );
INVx1_ASAP7_75t_L g725 ( .A(n_701), .Y(n_725) );
INVx2_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
AND2x4_ASAP7_75t_L g706 ( .A(n_707), .B(n_709), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_715), .Y(n_712) );
AOI221xp5_ASAP7_75t_L g746 ( .A1(n_713), .A2(n_747), .B1(n_749), .B2(n_751), .C(n_756), .Y(n_746) );
OAI21xp33_ASAP7_75t_SL g761 ( .A1(n_718), .A2(n_762), .B(n_763), .Y(n_761) );
INVx2_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NAND4xp25_ASAP7_75t_L g726 ( .A(n_727), .B(n_737), .C(n_746), .D(n_760), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_731), .B1(n_734), .B2(n_735), .Y(n_727) );
AND2x4_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVxp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_755), .Y(n_751) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
CKINVDCx11_ASAP7_75t_R g773 ( .A(n_768), .Y(n_773) );
INVx1_ASAP7_75t_SL g772 ( .A(n_773), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_777), .B(n_780), .Y(n_776) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
CKINVDCx5p33_ASAP7_75t_R g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_SL g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_SL g785 ( .A(n_786), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_788), .B(n_789), .Y(n_787) );
endmodule