module fake_jpeg_21_n_585 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_585);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_585;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_387;
wire n_270;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_54),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_19),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_56),
.B(n_60),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_20),
.B(n_19),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_57),
.B(n_66),
.Y(n_111)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_33),
.B(n_0),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_32),
.Y(n_64)
);

INVx6_ASAP7_75t_SL g110 ( 
.A(n_64),
.Y(n_110)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_65),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_48),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_1),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_68),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_20),
.B(n_1),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_69),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_72),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_33),
.B(n_1),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_73),
.B(n_81),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_32),
.Y(n_74)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_74),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_2),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_75),
.B(n_79),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_76),
.Y(n_149)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_78),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_48),
.Y(n_79)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_80),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_3),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_82),
.Y(n_157)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_84),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_25),
.B(n_3),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_85),
.B(n_87),
.Y(n_136)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_34),
.B(n_4),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_88),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_89),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_23),
.Y(n_91)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

BUFx10_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_93),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_94),
.Y(n_141)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_95),
.Y(n_161)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx6_ASAP7_75t_SL g135 ( 
.A(n_96),
.Y(n_135)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

BUFx8_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

CKINVDCx9p33_ASAP7_75t_R g117 ( 
.A(n_98),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_34),
.B(n_4),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_99),
.B(n_106),
.Y(n_143)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

OR2x2_ASAP7_75t_SL g103 ( 
.A(n_32),
.B(n_4),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_104),
.Y(n_131)
);

INVx4_ASAP7_75t_SL g104 ( 
.A(n_21),
.Y(n_104)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_35),
.B(n_5),
.Y(n_106)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_32),
.Y(n_107)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_108),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_62),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_115),
.B(n_142),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_64),
.A2(n_74),
.B1(n_98),
.B2(n_104),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_123),
.A2(n_126),
.B1(n_137),
.B2(n_163),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_75),
.B(n_51),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_124),
.B(n_140),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_98),
.A2(n_48),
.B1(n_39),
.B2(n_46),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_107),
.A2(n_39),
.B1(n_38),
.B2(n_50),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_67),
.B(n_52),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_91),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_51),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_144),
.B(n_145),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_54),
.B(n_35),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_63),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_150),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_58),
.B(n_47),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_78),
.B(n_47),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_160),
.Y(n_181)
);

NAND2xp33_ASAP7_75t_SL g159 ( 
.A(n_84),
.B(n_28),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_93),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_65),
.B(n_28),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_70),
.A2(n_50),
.B1(n_46),
.B2(n_38),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_162),
.A2(n_72),
.B1(n_76),
.B2(n_88),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_77),
.A2(n_39),
.B1(n_46),
.B2(n_50),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_95),
.B(n_52),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_173),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_69),
.B(n_40),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_174),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_175),
.A2(n_233),
.B1(n_236),
.B2(n_164),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_117),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_176),
.Y(n_254)
);

AO22x1_ASAP7_75t_L g177 ( 
.A1(n_110),
.A2(n_96),
.B1(n_102),
.B2(n_80),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_178),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_113),
.B(n_71),
.C(n_90),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_179),
.B(n_209),
.C(n_153),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_117),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_182),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_183),
.Y(n_263)
);

INVx11_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_184),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_131),
.A2(n_94),
.B1(n_89),
.B2(n_82),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_185),
.A2(n_199),
.B1(n_213),
.B2(n_225),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_123),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_186),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_131),
.A2(n_129),
.B1(n_163),
.B2(n_126),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_187),
.A2(n_219),
.B1(n_221),
.B2(n_118),
.Y(n_247)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_188),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_140),
.B(n_31),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_189),
.B(n_190),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_140),
.B(n_31),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_132),
.Y(n_191)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_191),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_155),
.A2(n_31),
.B1(n_28),
.B2(n_40),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_194),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_155),
.A2(n_40),
.B1(n_42),
.B2(n_24),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_195),
.A2(n_210),
.B1(n_216),
.B2(n_218),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_133),
.B(n_105),
.Y(n_196)
);

AND2x2_ASAP7_75t_SL g250 ( 
.A(n_196),
.B(n_167),
.Y(n_250)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_197),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_172),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_198),
.B(n_200),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_136),
.A2(n_100),
.B1(n_46),
.B2(n_36),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_135),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_201),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_122),
.B(n_42),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_202),
.B(n_206),
.Y(n_261)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_203),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_135),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_204),
.B(n_217),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_130),
.B(n_42),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_138),
.Y(n_207)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_207),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_111),
.B(n_133),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_208),
.B(n_228),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_120),
.B(n_36),
.C(n_38),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_152),
.A2(n_24),
.B1(n_52),
.B2(n_49),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_132),
.Y(n_211)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_211),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_143),
.A2(n_50),
.B1(n_38),
.B2(n_92),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_165),
.Y(n_214)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_214),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_151),
.Y(n_215)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_215),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_152),
.A2(n_41),
.B1(n_24),
.B2(n_22),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_127),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_116),
.A2(n_44),
.B1(n_41),
.B2(n_22),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_137),
.A2(n_44),
.B1(n_41),
.B2(n_22),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_139),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_220),
.Y(n_258)
);

O2A1O1Ixp33_ASAP7_75t_SL g221 ( 
.A1(n_125),
.A2(n_30),
.B(n_49),
.C(n_44),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_161),
.Y(n_222)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_222),
.Y(n_269)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_168),
.Y(n_223)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_223),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_170),
.B(n_61),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_232),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_114),
.A2(n_92),
.B1(n_55),
.B2(n_49),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_165),
.Y(n_227)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_227),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_134),
.B(n_55),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_121),
.Y(n_229)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_229),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_138),
.A2(n_30),
.B1(n_27),
.B2(n_8),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_234),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_114),
.A2(n_30),
.B1(n_27),
.B2(n_8),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_231),
.A2(n_235),
.B1(n_141),
.B2(n_118),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_139),
.B(n_6),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_121),
.A2(n_30),
.B1(n_7),
.B2(n_9),
.Y(n_233)
);

O2A1O1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_112),
.A2(n_30),
.B(n_9),
.C(n_11),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_148),
.A2(n_30),
.B1(n_9),
.B2(n_11),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_148),
.A2(n_6),
.B1(n_11),
.B2(n_12),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_188),
.A2(n_170),
.B1(n_164),
.B2(n_149),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_239),
.A2(n_274),
.B1(n_289),
.B2(n_184),
.Y(n_342)
);

MAJx2_ASAP7_75t_L g240 ( 
.A(n_192),
.B(n_134),
.C(n_157),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_240),
.B(n_286),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_109),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_243),
.B(n_276),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_247),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_250),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_252),
.A2(n_253),
.B1(n_267),
.B2(n_278),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_175),
.A2(n_128),
.B1(n_146),
.B2(n_149),
.Y(n_253)
);

FAx1_ASAP7_75t_SL g257 ( 
.A(n_181),
.B(n_119),
.CI(n_112),
.CON(n_257),
.SN(n_257)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_257),
.B(n_271),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_205),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_262),
.B(n_265),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_182),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_196),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_266),
.B(n_200),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_212),
.A2(n_146),
.B1(n_128),
.B2(n_141),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_192),
.B(n_167),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_199),
.A2(n_213),
.B1(n_185),
.B2(n_183),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_180),
.B(n_109),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_212),
.A2(n_157),
.B1(n_151),
.B2(n_168),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_280),
.A2(n_284),
.B1(n_287),
.B2(n_177),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_193),
.A2(n_156),
.B1(n_167),
.B2(n_119),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_181),
.B(n_119),
.Y(n_286)
);

OAI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_180),
.A2(n_153),
.B1(n_156),
.B2(n_13),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_226),
.B(n_11),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_288),
.B(n_176),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_183),
.A2(n_153),
.B1(n_13),
.B2(n_14),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_292),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_189),
.B(n_12),
.Y(n_292)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_264),
.Y(n_296)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_296),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_297),
.B(n_318),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_256),
.A2(n_186),
.B(n_221),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_299),
.A2(n_302),
.B(n_313),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_242),
.A2(n_233),
.B1(n_235),
.B2(n_236),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_300),
.A2(n_310),
.B1(n_314),
.B2(n_323),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_256),
.A2(n_221),
.B(n_190),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_268),
.Y(n_303)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_303),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_261),
.B(n_206),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_304),
.B(n_309),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_246),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_305),
.B(n_311),
.Y(n_370)
);

BUFx12f_ASAP7_75t_L g307 ( 
.A(n_275),
.Y(n_307)
);

INVx8_ASAP7_75t_L g351 ( 
.A(n_307),
.Y(n_351)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_237),
.B(n_226),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_308),
.A2(n_248),
.B(n_255),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_261),
.B(n_202),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_242),
.A2(n_179),
.B1(n_225),
.B2(n_177),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_246),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_263),
.A2(n_249),
.B(n_281),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_274),
.A2(n_209),
.B1(n_228),
.B2(n_231),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_264),
.Y(n_315)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_315),
.Y(n_364)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_269),
.Y(n_316)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_316),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_241),
.B(n_217),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_317),
.B(n_319),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_241),
.B(n_198),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_269),
.Y(n_320)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_320),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_283),
.B(n_197),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_321),
.B(n_327),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_246),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_322),
.B(n_338),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_252),
.A2(n_223),
.B1(n_215),
.B2(n_196),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_250),
.Y(n_324)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_324),
.Y(n_374)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_285),
.Y(n_325)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_325),
.Y(n_384)
);

OAI32xp33_ASAP7_75t_L g327 ( 
.A1(n_283),
.A2(n_203),
.A3(n_222),
.B1(n_174),
.B2(n_234),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_237),
.A2(n_215),
.B1(n_191),
.B2(n_211),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_328),
.A2(n_293),
.B1(n_297),
.B2(n_323),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_240),
.B(n_229),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_329),
.B(n_332),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_247),
.A2(n_230),
.B1(n_229),
.B2(n_227),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_330),
.A2(n_342),
.B1(n_278),
.B2(n_267),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_331),
.B(n_339),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_292),
.B(n_227),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_259),
.Y(n_333)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_333),
.Y(n_389)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_259),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_334),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_286),
.B(n_214),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_335),
.B(n_336),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_290),
.B(n_214),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_238),
.B(n_207),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_337),
.B(n_251),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_260),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_262),
.B(n_245),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_250),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_340),
.B(n_344),
.Y(n_349)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_268),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_341),
.B(n_343),
.Y(n_359)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_255),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_285),
.B(n_12),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_348),
.A2(n_310),
.B1(n_314),
.B2(n_308),
.Y(n_397)
);

OR2x2_ASAP7_75t_L g353 ( 
.A(n_302),
.B(n_257),
.Y(n_353)
);

A2O1A1Ixp33_ASAP7_75t_SL g413 ( 
.A1(n_353),
.A2(n_356),
.B(n_383),
.C(n_341),
.Y(n_413)
);

INVx2_ASAP7_75t_R g354 ( 
.A(n_313),
.Y(n_354)
);

INVxp33_ASAP7_75t_L g423 ( 
.A(n_354),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_299),
.A2(n_249),
.B(n_281),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_355),
.A2(n_367),
.B(n_382),
.Y(n_409)
);

O2A1O1Ixp33_ASAP7_75t_SL g356 ( 
.A1(n_306),
.A2(n_244),
.B(n_277),
.C(n_257),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_306),
.A2(n_244),
.B1(n_263),
.B2(n_253),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_358),
.A2(n_368),
.B1(n_378),
.B2(n_328),
.Y(n_411)
);

A2O1A1Ixp33_ASAP7_75t_L g360 ( 
.A1(n_329),
.A2(n_266),
.B(n_244),
.C(n_265),
.Y(n_360)
);

OAI21xp33_ASAP7_75t_L g392 ( 
.A1(n_360),
.A2(n_387),
.B(n_312),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_294),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_362),
.B(n_371),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_330),
.A2(n_284),
.B1(n_342),
.B2(n_325),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_300),
.A2(n_280),
.B1(n_289),
.B2(n_258),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_369),
.A2(n_321),
.B1(n_319),
.B2(n_295),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_317),
.B(n_258),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_326),
.Y(n_376)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_376),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_339),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_377),
.B(n_379),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_293),
.A2(n_282),
.B1(n_270),
.B2(n_275),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_337),
.Y(n_379)
);

O2A1O1Ixp33_ASAP7_75t_L g383 ( 
.A1(n_327),
.A2(n_248),
.B(n_273),
.C(n_254),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_385),
.B(n_386),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_308),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_305),
.A2(n_273),
.B1(n_272),
.B2(n_291),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_301),
.B(n_251),
.C(n_272),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_388),
.B(n_298),
.C(n_336),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_390),
.B(n_395),
.C(n_403),
.Y(n_433)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_347),
.Y(n_391)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_391),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_392),
.A2(n_396),
.B1(n_397),
.B2(n_404),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_362),
.B(n_338),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_393),
.B(n_394),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_377),
.B(n_380),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_381),
.B(n_298),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_359),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_398),
.B(n_399),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_380),
.B(n_376),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_359),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_400),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_350),
.B(n_301),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_401),
.B(n_412),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_381),
.B(n_335),
.C(n_324),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_346),
.A2(n_295),
.B1(n_304),
.B2(n_309),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_346),
.A2(n_312),
.B1(n_334),
.B2(n_333),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_405),
.A2(n_416),
.B1(n_424),
.B2(n_352),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_388),
.B(n_343),
.C(n_320),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_407),
.B(n_408),
.C(n_415),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_350),
.B(n_374),
.C(n_357),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_357),
.A2(n_296),
.B(n_316),
.Y(n_410)
);

AO21x1_ASAP7_75t_L g448 ( 
.A1(n_410),
.A2(n_413),
.B(n_354),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_411),
.A2(n_366),
.B1(n_360),
.B2(n_358),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_361),
.B(n_332),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_375),
.B(n_315),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_369),
.A2(n_366),
.B1(n_348),
.B2(n_361),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_375),
.B(n_303),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_417),
.B(n_426),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_372),
.B(n_307),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_418),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_371),
.B(n_322),
.Y(n_419)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_419),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_379),
.B(n_311),
.Y(n_420)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_420),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_384),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_421),
.Y(n_450)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_389),
.Y(n_422)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_422),
.Y(n_459)
);

OAI21xp33_ASAP7_75t_L g424 ( 
.A1(n_349),
.A2(n_291),
.B(n_282),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_345),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_425),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_374),
.B(n_270),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_370),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_427),
.Y(n_434)
);

XOR2x2_ASAP7_75t_L g429 ( 
.A(n_395),
.B(n_382),
.Y(n_429)
);

XNOR2x1_ASAP7_75t_L g475 ( 
.A(n_429),
.B(n_413),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_416),
.A2(n_366),
.B1(n_386),
.B2(n_368),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_441),
.A2(n_445),
.B1(n_446),
.B2(n_453),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_420),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_442),
.B(n_423),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_443),
.A2(n_455),
.B1(n_413),
.B2(n_383),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_402),
.B(n_385),
.Y(n_444)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_444),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_397),
.A2(n_353),
.B1(n_355),
.B2(n_378),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_396),
.A2(n_353),
.B1(n_356),
.B2(n_383),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_448),
.A2(n_462),
.B(n_443),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_402),
.B(n_370),
.Y(n_449)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_449),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_390),
.B(n_372),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_451),
.B(n_460),
.C(n_407),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_406),
.B(n_389),
.Y(n_452)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_452),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_411),
.A2(n_410),
.B1(n_405),
.B2(n_406),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_419),
.B(n_352),
.Y(n_456)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_456),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_414),
.B(n_373),
.Y(n_458)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_458),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_401),
.B(n_354),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_415),
.B(n_364),
.Y(n_461)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_461),
.Y(n_488)
);

OA21x2_ASAP7_75t_L g462 ( 
.A1(n_413),
.A2(n_356),
.B(n_408),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_463),
.B(n_475),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_444),
.B(n_417),
.Y(n_464)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_464),
.Y(n_494)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_465),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_449),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_467),
.B(n_473),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_433),
.B(n_403),
.C(n_426),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_468),
.B(n_470),
.C(n_471),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_455),
.A2(n_442),
.B1(n_440),
.B2(n_437),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_469),
.A2(n_484),
.B1(n_487),
.B2(n_441),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_433),
.B(n_423),
.C(n_404),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_447),
.B(n_412),
.C(n_409),
.Y(n_471)
);

CKINVDCx14_ASAP7_75t_R g473 ( 
.A(n_457),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_439),
.B(n_428),
.Y(n_476)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_476),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_447),
.B(n_409),
.C(n_365),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_478),
.B(n_486),
.C(n_489),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_456),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_479),
.B(n_482),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_480),
.A2(n_491),
.B(n_448),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_452),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_430),
.B(n_365),
.Y(n_483)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_483),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_451),
.B(n_429),
.C(n_435),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_440),
.A2(n_373),
.B1(n_364),
.B2(n_363),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_435),
.B(n_363),
.C(n_384),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_430),
.B(n_307),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_490),
.B(n_279),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_448),
.A2(n_351),
.B(n_307),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_481),
.A2(n_437),
.B1(n_458),
.B2(n_436),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_492),
.B(n_500),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_476),
.B(n_432),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_495),
.B(n_501),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_468),
.B(n_454),
.C(n_460),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_498),
.B(n_502),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_499),
.A2(n_491),
.B(n_465),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_489),
.B(n_432),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_463),
.B(n_454),
.C(n_438),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_470),
.B(n_461),
.C(n_462),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_503),
.B(n_510),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_467),
.B(n_431),
.Y(n_507)
);

OAI221xp5_ASAP7_75t_L g535 ( 
.A1(n_507),
.A2(n_466),
.B1(n_490),
.B2(n_474),
.C(n_487),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_469),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_508),
.B(n_472),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_484),
.A2(n_445),
.B1(n_462),
.B2(n_446),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_509),
.B(n_512),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_478),
.B(n_434),
.C(n_450),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_481),
.A2(n_434),
.B1(n_431),
.B2(n_459),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_486),
.B(n_459),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_514),
.B(n_515),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_471),
.B(n_450),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_516),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_515),
.B(n_480),
.C(n_488),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_518),
.B(n_524),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_521),
.A2(n_500),
.B(n_505),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_496),
.B(n_497),
.C(n_514),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_SL g525 ( 
.A1(n_499),
.A2(n_479),
.B(n_482),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_SL g539 ( 
.A1(n_525),
.A2(n_529),
.B(n_533),
.Y(n_539)
);

OAI21xp33_ASAP7_75t_L g526 ( 
.A1(n_493),
.A2(n_488),
.B(n_472),
.Y(n_526)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_526),
.Y(n_537)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_527),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_509),
.A2(n_477),
.B(n_485),
.Y(n_529)
);

NOR3xp33_ASAP7_75t_L g530 ( 
.A(n_506),
.B(n_483),
.C(n_466),
.Y(n_530)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_530),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_496),
.B(n_475),
.C(n_464),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_532),
.B(n_497),
.C(n_502),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_511),
.A2(n_477),
.B(n_485),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_516),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_534),
.B(n_492),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_535),
.A2(n_351),
.B1(n_279),
.B2(n_254),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_536),
.B(n_543),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_524),
.B(n_510),
.C(n_503),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_538),
.B(n_540),
.C(n_536),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_528),
.B(n_523),
.C(n_518),
.Y(n_540)
);

AOI21x1_ASAP7_75t_L g541 ( 
.A1(n_525),
.A2(n_504),
.B(n_513),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g564 ( 
.A1(n_541),
.A2(n_546),
.B(n_549),
.Y(n_564)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_542),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_519),
.A2(n_512),
.B1(n_494),
.B2(n_474),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_532),
.B(n_505),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_545),
.B(n_547),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_519),
.A2(n_522),
.B1(n_517),
.B2(n_531),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_523),
.B(n_498),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_548),
.B(n_16),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_522),
.A2(n_351),
.B1(n_14),
.B2(n_15),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_552),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_537),
.A2(n_533),
.B(n_521),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_553),
.A2(n_539),
.B(n_546),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_554),
.B(n_555),
.Y(n_567)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_544),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_538),
.B(n_520),
.C(n_529),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_556),
.B(n_557),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_541),
.Y(n_557)
);

AOI322xp5_ASAP7_75t_L g558 ( 
.A1(n_550),
.A2(n_13),
.A3(n_14),
.B1(n_15),
.B2(n_16),
.C1(n_17),
.C2(n_539),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_558),
.A2(n_559),
.B1(n_551),
.B2(n_552),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_561),
.B(n_549),
.Y(n_573)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_543),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_563),
.B(n_540),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_L g574 ( 
.A1(n_566),
.A2(n_553),
.B(n_562),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_554),
.B(n_548),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_568),
.B(n_565),
.Y(n_578)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_562),
.Y(n_570)
);

AO21x1_ASAP7_75t_L g575 ( 
.A1(n_570),
.A2(n_572),
.B(n_564),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_571),
.B(n_573),
.Y(n_577)
);

NAND3xp33_ASAP7_75t_L g579 ( 
.A(n_574),
.B(n_575),
.C(n_576),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_570),
.B(n_556),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_578),
.B(n_560),
.C(n_567),
.Y(n_580)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_580),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_577),
.B(n_569),
.C(n_560),
.Y(n_581)
);

AOI321xp33_ASAP7_75t_L g582 ( 
.A1(n_581),
.A2(n_564),
.A3(n_565),
.B1(n_545),
.B2(n_559),
.C(n_17),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_SL g584 ( 
.A1(n_582),
.A2(n_579),
.B(n_17),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_584),
.B(n_583),
.Y(n_585)
);


endmodule