module fake_jpeg_1438_n_691 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_691);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_691;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_331;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_539;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_11),
.B(n_1),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_19),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_60),
.Y(n_150)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_62),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_63),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_64),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_46),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_65),
.B(n_69),
.Y(n_135)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_66),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_67),
.Y(n_178)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_68),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_9),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_25),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_70),
.B(n_51),
.Y(n_137)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_71),
.Y(n_146)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_72),
.Y(n_158)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_73),
.Y(n_148)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_74),
.Y(n_162)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_76),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_77),
.Y(n_195)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_79),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_32),
.Y(n_80)
);

HAxp5_ASAP7_75t_SL g217 ( 
.A(n_80),
.B(n_103),
.CON(n_217),
.SN(n_217)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_81),
.Y(n_165)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_82),
.Y(n_191)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_83),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_84),
.Y(n_179)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_85),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_86),
.Y(n_200)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_87),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_88),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_36),
.B(n_9),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_89),
.B(n_90),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_37),
.B(n_9),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_91),
.Y(n_171)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_92),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_93),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_37),
.B(n_12),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_94),
.B(n_96),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_95),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_23),
.B(n_19),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_98),
.Y(n_167)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_20),
.Y(n_99)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_99),
.Y(n_183)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_100),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_39),
.Y(n_101)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_101),
.Y(n_209)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_102),
.Y(n_185)
);

HAxp5_ASAP7_75t_SL g103 ( 
.A(n_23),
.B(n_0),
.CON(n_103),
.SN(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_21),
.Y(n_104)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_104),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_30),
.B(n_19),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_19),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_28),
.Y(n_106)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_106),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_28),
.Y(n_107)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_107),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_21),
.Y(n_108)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_108),
.Y(n_222)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_20),
.Y(n_109)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_109),
.Y(n_214)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_34),
.Y(n_110)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_110),
.Y(n_228)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

INVx4_ASAP7_75t_SL g112 ( 
.A(n_20),
.Y(n_112)
);

CKINVDCx6p67_ASAP7_75t_R g140 ( 
.A(n_112),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_29),
.Y(n_113)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_113),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_114),
.Y(n_227)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_115),
.Y(n_229)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_29),
.Y(n_116)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_116),
.Y(n_203)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_117),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_39),
.Y(n_118)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_118),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_29),
.Y(n_119)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_120),
.Y(n_206)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_121),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_39),
.Y(n_122)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_122),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_34),
.Y(n_123)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_123),
.Y(n_226)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_43),
.Y(n_124)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_124),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_39),
.Y(n_125)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

BUFx12_ASAP7_75t_L g126 ( 
.A(n_22),
.Y(n_126)
);

INVx6_ASAP7_75t_SL g221 ( 
.A(n_126),
.Y(n_221)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_44),
.Y(n_127)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

BUFx4f_ASAP7_75t_L g128 ( 
.A(n_33),
.Y(n_128)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_48),
.Y(n_129)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_44),
.Y(n_130)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_130),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_39),
.Y(n_131)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_131),
.Y(n_202)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_48),
.Y(n_132)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_132),
.Y(n_215)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_51),
.Y(n_133)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_133),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_137),
.B(n_186),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_58),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_142),
.B(n_163),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_67),
.A2(n_53),
.B1(n_30),
.B2(n_49),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_143),
.A2(n_168),
.B1(n_169),
.B2(n_176),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_147),
.B(n_160),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_60),
.A2(n_64),
.B1(n_62),
.B2(n_98),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_152),
.A2(n_181),
.B1(n_126),
.B2(n_2),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_87),
.B(n_57),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_101),
.B(n_58),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_80),
.B(n_57),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_164),
.B(n_170),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_63),
.A2(n_53),
.B1(n_49),
.B2(n_38),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_77),
.A2(n_40),
.B1(n_38),
.B2(n_52),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_113),
.B(n_26),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_119),
.B(n_26),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_172),
.B(n_213),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_101),
.B(n_40),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_173),
.B(n_177),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_86),
.A2(n_52),
.B1(n_22),
.B2(n_55),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_118),
.B(n_15),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_L g181 ( 
.A1(n_93),
.A2(n_54),
.B1(n_33),
.B2(n_44),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_95),
.A2(n_47),
.B1(n_54),
.B2(n_14),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_184),
.A2(n_189),
.B1(n_196),
.B2(n_122),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_118),
.B(n_13),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_63),
.B(n_13),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_187),
.B(n_190),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_128),
.A2(n_55),
.B1(n_22),
.B2(n_47),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_81),
.B(n_13),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_92),
.A2(n_55),
.B1(n_22),
.B2(n_47),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_84),
.B(n_13),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_197),
.B(n_212),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_103),
.B(n_47),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_199),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_61),
.B(n_14),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_120),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_83),
.B(n_18),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_100),
.B(n_18),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_218),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_78),
.B(n_17),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_223),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_106),
.B(n_17),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_110),
.B(n_17),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_225),
.Y(n_266)
);

BUFx4f_ASAP7_75t_SL g233 ( 
.A(n_221),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_233),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_154),
.Y(n_236)
);

INVx8_ASAP7_75t_L g370 ( 
.A(n_236),
.Y(n_370)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_237),
.Y(n_344)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_136),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_238),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_140),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_239),
.B(n_257),
.Y(n_323)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_157),
.Y(n_240)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_240),
.Y(n_363)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_206),
.Y(n_241)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_241),
.Y(n_325)
);

INVx8_ASAP7_75t_L g242 ( 
.A(n_188),
.Y(n_242)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_242),
.Y(n_321)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_159),
.Y(n_244)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_244),
.Y(n_334)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_139),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_245),
.B(n_246),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_140),
.Y(n_246)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_154),
.Y(n_247)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_247),
.Y(n_330)
);

OAI21xp33_ASAP7_75t_L g248 ( 
.A1(n_199),
.A2(n_16),
.B(n_15),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g380 ( 
.A(n_248),
.Y(n_380)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_150),
.Y(n_250)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_250),
.Y(n_332)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_165),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_252),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_143),
.A2(n_108),
.B1(n_114),
.B2(n_107),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_254),
.A2(n_300),
.B1(n_228),
.B2(n_161),
.Y(n_345)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_215),
.Y(n_256)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_256),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_140),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_165),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_258),
.Y(n_354)
);

INVx11_ASAP7_75t_L g259 ( 
.A(n_182),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_259),
.Y(n_357)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_134),
.Y(n_260)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_260),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_149),
.B(n_111),
.Y(n_261)
);

AND2x2_ASAP7_75t_SL g356 ( 
.A(n_261),
.B(n_281),
.Y(n_356)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_134),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_262),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_185),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_263),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_193),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_264),
.B(n_269),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_182),
.Y(n_268)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_268),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_193),
.Y(n_269)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_153),
.Y(n_270)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_270),
.Y(n_360)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_150),
.Y(n_271)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_271),
.Y(n_373)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_156),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_272),
.B(n_273),
.Y(n_364)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_155),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_167),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_274),
.B(n_275),
.Y(n_374)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_167),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_145),
.B(n_117),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_276),
.B(n_299),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_181),
.A2(n_82),
.B1(n_71),
.B2(n_76),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_277),
.A2(n_282),
.B1(n_284),
.B2(n_285),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_226),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_278),
.B(n_280),
.Y(n_379)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_153),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_230),
.B(n_127),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_219),
.A2(n_130),
.B1(n_131),
.B2(n_125),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_217),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_283),
.B(n_222),
.Y(n_327)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_211),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_179),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_286),
.A2(n_287),
.B1(n_289),
.B2(n_290),
.Y(n_362)
);

INVx8_ASAP7_75t_L g287 ( 
.A(n_188),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_166),
.B(n_174),
.Y(n_288)
);

AND2x4_ASAP7_75t_L g342 ( 
.A(n_288),
.B(n_296),
.Y(n_342)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_224),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_158),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_175),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_292),
.A2(n_293),
.B1(n_294),
.B2(n_298),
.Y(n_378)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_144),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_202),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_198),
.Y(n_295)
);

BUFx24_ASAP7_75t_SL g350 ( 
.A(n_295),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_180),
.B(n_0),
.Y(n_296)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_178),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_183),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_176),
.A2(n_203),
.B1(n_207),
.B2(n_229),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_148),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_307),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_162),
.B(n_214),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_222),
.C(n_146),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_219),
.A2(n_55),
.B1(n_22),
.B2(n_47),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_L g353 ( 
.A1(n_303),
.A2(n_306),
.B1(n_314),
.B2(n_231),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_209),
.Y(n_305)
);

NOR2x1_ASAP7_75t_L g329 ( 
.A(n_305),
.B(n_313),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_217),
.A2(n_55),
.B1(n_16),
.B2(n_15),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_138),
.B(n_0),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_178),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_308),
.B(n_309),
.Y(n_337)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_171),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_151),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_310),
.B(n_311),
.Y(n_343)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_195),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_135),
.A2(n_126),
.B1(n_16),
.B2(n_3),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_312),
.A2(n_248),
.B1(n_196),
.B2(n_307),
.Y(n_322)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_155),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_194),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_315),
.B(n_316),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_227),
.B(n_1),
.Y(n_316)
);

INVx8_ASAP7_75t_L g317 ( 
.A(n_192),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_317),
.A2(n_179),
.B1(n_208),
.B2(n_191),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_279),
.A2(n_168),
.B1(n_189),
.B2(n_200),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_318),
.A2(n_328),
.B1(n_331),
.B2(n_333),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_322),
.B(n_366),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_324),
.Y(n_385)
);

CKINVDCx14_ASAP7_75t_R g405 ( 
.A(n_327),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_276),
.A2(n_200),
.B1(n_195),
.B2(n_205),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_235),
.A2(n_198),
.B1(n_192),
.B2(n_205),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_314),
.A2(n_201),
.B1(n_161),
.B2(n_210),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_249),
.B(n_141),
.C(n_228),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_341),
.B(n_369),
.C(n_268),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_345),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_347),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_243),
.A2(n_201),
.B1(n_141),
.B2(n_208),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_351),
.A2(n_355),
.B1(n_361),
.B2(n_371),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_353),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_243),
.A2(n_231),
.B1(n_232),
.B2(n_191),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_253),
.A2(n_232),
.B1(n_146),
.B2(n_3),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_359),
.A2(n_375),
.B(n_252),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_253),
.A2(n_266),
.B1(n_316),
.B2(n_234),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_266),
.B(n_1),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_5),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_251),
.B(n_1),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_234),
.A2(n_297),
.B(n_302),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_367),
.A2(n_7),
.B(n_323),
.Y(n_426)
);

MAJx2_ASAP7_75t_L g369 ( 
.A(n_265),
.B(n_2),
.C(n_3),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_304),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_255),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_372),
.A2(n_376),
.B1(n_272),
.B2(n_240),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_267),
.A2(n_288),
.B(n_296),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_296),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_376)
);

OA22x2_ASAP7_75t_L g377 ( 
.A1(n_293),
.A2(n_294),
.B1(n_270),
.B2(n_280),
.Y(n_377)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_377),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_382),
.B(n_390),
.Y(n_436)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_343),
.Y(n_383)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_383),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_344),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_384),
.B(n_394),
.Y(n_464)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_343),
.Y(n_387)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_387),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_349),
.Y(n_388)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_388),
.Y(n_444)
);

OR2x2_ASAP7_75t_L g389 ( 
.A(n_327),
.B(n_291),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_389),
.A2(n_401),
.B(n_339),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_319),
.B(n_348),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_319),
.A2(n_261),
.B1(n_281),
.B2(n_302),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_392),
.A2(n_397),
.B1(n_422),
.B2(n_427),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_393),
.B(n_402),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_344),
.Y(n_394)
);

MAJx2_ASAP7_75t_L g395 ( 
.A(n_375),
.B(n_288),
.C(n_261),
.Y(n_395)
);

MAJx2_ASAP7_75t_L g467 ( 
.A(n_395),
.B(n_326),
.C(n_338),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_331),
.A2(n_274),
.B1(n_275),
.B2(n_271),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_396),
.A2(n_400),
.B1(n_410),
.B2(n_358),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_362),
.A2(n_281),
.B1(n_250),
.B2(n_308),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_337),
.Y(n_398)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_398),
.Y(n_457)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_337),
.Y(n_399)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_399),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_318),
.A2(n_311),
.B1(n_298),
.B2(n_237),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g401 ( 
.A(n_329),
.B(n_233),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_348),
.B(n_284),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_344),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_403),
.B(n_407),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_320),
.B(n_278),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_404),
.B(n_408),
.C(n_417),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_406),
.B(n_417),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_361),
.B(n_233),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_320),
.B(n_241),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_333),
.A2(n_317),
.B1(n_242),
.B2(n_287),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_367),
.B(n_313),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g433 ( 
.A(n_413),
.B(n_425),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_380),
.A2(n_365),
.B(n_342),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_415),
.A2(n_416),
.B(n_426),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_341),
.B(n_285),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_342),
.B(n_262),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_418),
.B(n_419),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_342),
.B(n_273),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_342),
.B(n_369),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_420),
.B(n_421),
.C(n_423),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_342),
.B(n_260),
.C(n_258),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_356),
.A2(n_247),
.B1(n_236),
.B2(n_244),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_356),
.B(n_305),
.C(n_259),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_366),
.B(n_7),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_424),
.B(n_376),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_350),
.B(n_368),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_356),
.A2(n_336),
.B1(n_322),
.B2(n_351),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_330),
.Y(n_428)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_428),
.Y(n_431)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_374),
.Y(n_429)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_429),
.Y(n_463)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_374),
.Y(n_430)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_430),
.Y(n_468)
);

AOI22x1_ASAP7_75t_L g432 ( 
.A1(n_414),
.A2(n_355),
.B1(n_328),
.B2(n_371),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_432),
.A2(n_452),
.B1(n_465),
.B2(n_469),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_401),
.A2(n_329),
.B(n_352),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_435),
.A2(n_449),
.B(n_451),
.Y(n_486)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_428),
.Y(n_438)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_438),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_428),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_442),
.B(n_454),
.Y(n_490)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_445),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_390),
.B(n_369),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_446),
.B(n_455),
.C(n_385),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_447),
.B(n_450),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_416),
.A2(n_329),
.B(n_359),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_383),
.B(n_356),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_415),
.A2(n_368),
.B(n_379),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_427),
.A2(n_372),
.B1(n_330),
.B2(n_321),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_387),
.B(n_398),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_453),
.B(n_456),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_426),
.Y(n_454)
);

AO22x1_ASAP7_75t_L g456 ( 
.A1(n_414),
.A2(n_377),
.B1(n_326),
.B2(n_364),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_459),
.A2(n_389),
.B(n_424),
.Y(n_500)
);

AO21x2_ASAP7_75t_L g461 ( 
.A1(n_381),
.A2(n_377),
.B(n_360),
.Y(n_461)
);

AO21x1_ASAP7_75t_L g511 ( 
.A1(n_461),
.A2(n_377),
.B(n_364),
.Y(n_511)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_399),
.Y(n_462)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_462),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_381),
.A2(n_391),
.B1(n_411),
.B2(n_409),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_404),
.B(n_324),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_466),
.B(n_467),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_391),
.A2(n_321),
.B1(n_360),
.B2(n_358),
.Y(n_469)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_429),
.Y(n_471)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_471),
.Y(n_484)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_430),
.Y(n_472)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_472),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_465),
.A2(n_448),
.B1(n_452),
.B2(n_461),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_473),
.A2(n_478),
.B1(n_482),
.B2(n_485),
.Y(n_533)
);

CKINVDCx14_ASAP7_75t_R g478 ( 
.A(n_451),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_481),
.B(n_493),
.C(n_507),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_456),
.A2(n_411),
.B1(n_405),
.B2(n_385),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_448),
.A2(n_412),
.B1(n_397),
.B2(n_386),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_464),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_487),
.B(n_495),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_436),
.B(n_408),
.Y(n_488)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_488),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_461),
.A2(n_412),
.B1(n_386),
.B2(n_406),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_489),
.A2(n_501),
.B1(n_508),
.B2(n_485),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_455),
.B(n_434),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_491),
.B(n_496),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_436),
.B(n_402),
.Y(n_492)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_492),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_440),
.B(n_420),
.C(n_395),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_461),
.A2(n_412),
.B1(n_400),
.B2(n_401),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_494),
.A2(n_498),
.B1(n_456),
.B2(n_457),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_453),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_434),
.B(n_466),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_441),
.A2(n_419),
.B(n_418),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_497),
.A2(n_500),
.B(n_509),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_461),
.A2(n_410),
.B1(n_423),
.B2(n_421),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_433),
.B(n_389),
.Y(n_499)
);

CKINVDCx14_ASAP7_75t_R g550 ( 
.A(n_499),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_439),
.A2(n_422),
.B1(n_392),
.B2(n_396),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_470),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_503),
.B(n_444),
.Y(n_520)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_462),
.Y(n_504)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_504),
.Y(n_526)
);

CKINVDCx14_ASAP7_75t_R g505 ( 
.A(n_433),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_505),
.B(n_468),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_440),
.B(n_382),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_506),
.B(n_446),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_467),
.B(n_338),
.C(n_346),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_439),
.A2(n_393),
.B1(n_403),
.B2(n_384),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_441),
.A2(n_347),
.B(n_339),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_459),
.A2(n_394),
.B(n_378),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_510),
.A2(n_377),
.B(n_335),
.Y(n_549)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_511),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_444),
.Y(n_512)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_512),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_491),
.B(n_450),
.C(n_458),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_515),
.B(n_523),
.C(n_524),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g574 ( 
.A1(n_518),
.A2(n_536),
.B1(n_501),
.B2(n_508),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_490),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_519),
.B(n_527),
.Y(n_567)
);

INVxp67_ASAP7_75t_SL g571 ( 
.A(n_520),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_496),
.B(n_458),
.C(n_457),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_525),
.A2(n_538),
.B1(n_547),
.B2(n_548),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_477),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_479),
.B(n_460),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_530),
.B(n_531),
.C(n_545),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_493),
.B(n_472),
.C(n_471),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_489),
.Y(n_532)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_532),
.Y(n_577)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_484),
.Y(n_534)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_534),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_495),
.B(n_468),
.Y(n_535)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_535),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_475),
.A2(n_437),
.B1(n_469),
.B2(n_445),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_SL g556 ( 
.A(n_537),
.B(n_541),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_473),
.A2(n_437),
.B1(n_435),
.B2(n_463),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_487),
.B(n_463),
.Y(n_539)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_539),
.Y(n_569)
);

OA21x2_ASAP7_75t_L g540 ( 
.A1(n_477),
.A2(n_494),
.B(n_475),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_540),
.B(n_511),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_503),
.B(n_334),
.Y(n_541)
);

CKINVDCx16_ASAP7_75t_R g542 ( 
.A(n_482),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_542),
.B(n_500),
.Y(n_572)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_484),
.Y(n_543)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_543),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_492),
.B(n_443),
.Y(n_544)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_544),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_481),
.B(n_443),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_479),
.B(n_449),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_546),
.B(n_506),
.C(n_486),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_476),
.A2(n_432),
.B1(n_447),
.B2(n_431),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_476),
.A2(n_432),
.B1(n_431),
.B2(n_438),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_L g562 ( 
.A1(n_549),
.A2(n_509),
.B(n_511),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g586 ( 
.A(n_551),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_SL g553 ( 
.A(n_546),
.B(n_507),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_SL g609 ( 
.A(n_553),
.B(n_581),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_516),
.B(n_504),
.Y(n_555)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_555),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_522),
.A2(n_486),
.B(n_510),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_SL g598 ( 
.A1(n_557),
.A2(n_562),
.B(n_549),
.Y(n_598)
);

NOR3xp33_ASAP7_75t_SL g558 ( 
.A(n_516),
.B(n_550),
.C(n_539),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_558),
.B(n_566),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_529),
.B(n_502),
.Y(n_561)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_561),
.Y(n_589)
);

XOR2xp5_ASAP7_75t_L g596 ( 
.A(n_563),
.B(n_514),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_529),
.B(n_502),
.Y(n_564)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_564),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_525),
.A2(n_483),
.B1(n_498),
.B2(n_497),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g600 ( 
.A1(n_565),
.A2(n_528),
.B1(n_513),
.B2(n_540),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_520),
.B(n_480),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_535),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_570),
.B(n_573),
.Y(n_594)
);

CKINVDCx14_ASAP7_75t_R g603 ( 
.A(n_572),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g573 ( 
.A(n_526),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_574),
.A2(n_575),
.B1(n_576),
.B2(n_579),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_532),
.A2(n_480),
.B1(n_488),
.B2(n_474),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_SL g576 ( 
.A1(n_518),
.A2(n_474),
.B1(n_370),
.B2(n_357),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g579 ( 
.A1(n_536),
.A2(n_370),
.B1(n_357),
.B2(n_340),
.Y(n_579)
);

NAND3xp33_ASAP7_75t_SL g580 ( 
.A(n_522),
.B(n_521),
.C(n_544),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_580),
.B(n_582),
.Y(n_608)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_534),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_521),
.B(n_374),
.Y(n_583)
);

CKINVDCx14_ASAP7_75t_R g606 ( 
.A(n_583),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_552),
.B(n_517),
.C(n_531),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_584),
.B(n_592),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_552),
.B(n_524),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_587),
.B(n_590),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_SL g588 ( 
.A1(n_574),
.A2(n_533),
.B1(n_538),
.B2(n_528),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_SL g624 ( 
.A1(n_588),
.A2(n_597),
.B1(n_605),
.B2(n_566),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_560),
.B(n_545),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_560),
.B(n_517),
.C(n_514),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_596),
.B(n_598),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_570),
.A2(n_540),
.B1(n_547),
.B2(n_548),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_SL g599 ( 
.A(n_567),
.B(n_515),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_599),
.B(n_556),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_600),
.A2(n_562),
.B1(n_551),
.B2(n_569),
.Y(n_617)
);

XOR2xp5_ASAP7_75t_L g601 ( 
.A(n_563),
.B(n_530),
.Y(n_601)
);

XOR2xp5_ASAP7_75t_L g626 ( 
.A(n_601),
.B(n_609),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_553),
.B(n_523),
.C(n_513),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_602),
.B(n_604),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_557),
.B(n_526),
.C(n_543),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_SL g605 ( 
.A1(n_569),
.A2(n_340),
.B1(n_349),
.B2(n_334),
.Y(n_605)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_555),
.B(n_364),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g623 ( 
.A(n_607),
.B(n_583),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_SL g611 ( 
.A1(n_597),
.A2(n_559),
.B1(n_565),
.B2(n_568),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_611),
.A2(n_615),
.B1(n_625),
.B2(n_629),
.Y(n_639)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_589),
.Y(n_614)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_614),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_SL g615 ( 
.A1(n_591),
.A2(n_559),
.B1(n_588),
.B2(n_568),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_587),
.B(n_575),
.C(n_577),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_L g632 ( 
.A(n_616),
.B(n_618),
.Y(n_632)
);

INVxp33_ASAP7_75t_L g636 ( 
.A(n_617),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_584),
.B(n_577),
.C(n_571),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_590),
.B(n_576),
.C(n_573),
.Y(n_620)
);

XNOR2xp5_ASAP7_75t_L g644 ( 
.A(n_620),
.B(n_628),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_SL g642 ( 
.A(n_621),
.B(n_622),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_595),
.B(n_558),
.Y(n_622)
);

XOR2xp5_ASAP7_75t_L g635 ( 
.A(n_623),
.B(n_607),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_SL g641 ( 
.A1(n_624),
.A2(n_600),
.B1(n_586),
.B2(n_591),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g625 ( 
.A(n_604),
.Y(n_625)
);

INVx6_ASAP7_75t_L g627 ( 
.A(n_603),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_SL g634 ( 
.A1(n_627),
.A2(n_585),
.B1(n_606),
.B2(n_605),
.Y(n_634)
);

XOR2xp5_ASAP7_75t_SL g628 ( 
.A(n_598),
.B(n_581),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_594),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_592),
.B(n_579),
.C(n_564),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g646 ( 
.A(n_630),
.B(n_586),
.C(n_578),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_SL g631 ( 
.A1(n_593),
.A2(n_561),
.B1(n_582),
.B2(n_578),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_631),
.A2(n_554),
.B1(n_332),
.B2(n_373),
.Y(n_648)
);

NAND2xp33_ASAP7_75t_R g633 ( 
.A(n_619),
.B(n_608),
.Y(n_633)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_633),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_634),
.B(n_638),
.Y(n_658)
);

XOR2xp5_ASAP7_75t_L g662 ( 
.A(n_635),
.B(n_325),
.Y(n_662)
);

XNOR2xp5_ASAP7_75t_L g638 ( 
.A(n_630),
.B(n_620),
.Y(n_638)
);

AOI31xp33_ASAP7_75t_L g640 ( 
.A1(n_618),
.A2(n_602),
.A3(n_556),
.B(n_609),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_640),
.B(n_647),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_641),
.B(n_643),
.Y(n_650)
);

XNOR2xp5_ASAP7_75t_L g643 ( 
.A(n_616),
.B(n_596),
.Y(n_643)
);

XNOR2xp5_ASAP7_75t_L g645 ( 
.A(n_612),
.B(n_601),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_645),
.B(n_646),
.Y(n_651)
);

BUFx24_ASAP7_75t_SL g647 ( 
.A(n_610),
.Y(n_647)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_648),
.Y(n_663)
);

MAJIxp5_ASAP7_75t_L g649 ( 
.A(n_613),
.B(n_554),
.C(n_332),
.Y(n_649)
);

MAJIxp5_ASAP7_75t_L g653 ( 
.A(n_649),
.B(n_628),
.C(n_619),
.Y(n_653)
);

XNOR2xp5_ASAP7_75t_L g667 ( 
.A(n_653),
.B(n_662),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_636),
.A2(n_615),
.B1(n_611),
.B2(n_617),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_SL g672 ( 
.A1(n_654),
.A2(n_643),
.B1(n_354),
.B2(n_363),
.Y(n_672)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_632),
.B(n_613),
.C(n_626),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_655),
.B(n_656),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_642),
.B(n_627),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_646),
.B(n_626),
.Y(n_657)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_657),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_638),
.B(n_623),
.Y(n_659)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_659),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_636),
.A2(n_373),
.B(n_325),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_660),
.A2(n_649),
.B(n_635),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_644),
.B(n_370),
.Y(n_664)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_664),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_652),
.B(n_639),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_665),
.B(n_671),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_SL g666 ( 
.A1(n_661),
.A2(n_641),
.B(n_637),
.Y(n_666)
);

MAJx2_ASAP7_75t_L g675 ( 
.A(n_666),
.B(n_658),
.C(n_663),
.Y(n_675)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_668),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_651),
.B(n_645),
.Y(n_671)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_672),
.Y(n_680)
);

XNOR2xp5_ASAP7_75t_L g685 ( 
.A(n_675),
.B(n_654),
.Y(n_685)
);

AOI21x1_ASAP7_75t_L g676 ( 
.A1(n_666),
.A2(n_658),
.B(n_650),
.Y(n_676)
);

NOR3xp33_ASAP7_75t_L g682 ( 
.A(n_676),
.B(n_677),
.C(n_681),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_673),
.A2(n_655),
.B(n_653),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_668),
.Y(n_681)
);

MAJIxp5_ASAP7_75t_L g683 ( 
.A(n_679),
.B(n_669),
.C(n_670),
.Y(n_683)
);

OAI21xp5_ASAP7_75t_L g687 ( 
.A1(n_683),
.A2(n_684),
.B(n_685),
.Y(n_687)
);

MAJIxp5_ASAP7_75t_L g684 ( 
.A(n_678),
.B(n_674),
.C(n_667),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_SL g686 ( 
.A1(n_682),
.A2(n_680),
.B(n_675),
.Y(n_686)
);

AOI21xp33_ASAP7_75t_L g688 ( 
.A1(n_686),
.A2(n_660),
.B(n_663),
.Y(n_688)
);

MAJIxp5_ASAP7_75t_L g689 ( 
.A(n_688),
.B(n_687),
.C(n_672),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_689),
.A2(n_667),
.B(n_662),
.Y(n_690)
);

MAJIxp5_ASAP7_75t_L g691 ( 
.A(n_690),
.B(n_354),
.C(n_363),
.Y(n_691)
);


endmodule