module real_jpeg_29648_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_176;
wire n_221;
wire n_166;
wire n_286;
wire n_288;
wire n_292;
wire n_300;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_173;
wire n_105;
wire n_299;
wire n_197;
wire n_115;
wire n_243;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_184;
wire n_164;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_305;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_304;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_262;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_295;
wire n_213;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_0),
.A2(n_34),
.B1(n_35),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_0),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_57),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_0),
.A2(n_57),
.B1(n_76),
.B2(n_77),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_0),
.A2(n_47),
.B1(n_50),
.B2(n_57),
.Y(n_116)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_1),
.Y(n_91)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_1),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_1),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_2),
.A2(n_38),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_2),
.A2(n_38),
.B1(n_47),
.B2(n_50),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_3),
.A2(n_76),
.B1(n_77),
.B2(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_3),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_155),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_3),
.A2(n_34),
.B1(n_35),
.B2(n_155),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_3),
.A2(n_47),
.B1(n_50),
.B2(n_155),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_40),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_4),
.A2(n_40),
.B1(n_47),
.B2(n_50),
.Y(n_143)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_6),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_6),
.B(n_72),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_6),
.B(n_29),
.Y(n_214)
);

AOI21xp33_ASAP7_75t_L g218 ( 
.A1(n_6),
.A2(n_29),
.B(n_214),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_174),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_6),
.A2(n_47),
.B(n_51),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_6),
.B(n_121),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_6),
.A2(n_88),
.B1(n_91),
.B2(n_262),
.Y(n_264)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_8),
.A2(n_76),
.B1(n_77),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_8),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_127),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_127),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_8),
.A2(n_47),
.B1(n_50),
.B2(n_127),
.Y(n_249)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_9),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_10),
.A2(n_44),
.B1(n_47),
.B2(n_50),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_10),
.A2(n_44),
.B1(n_76),
.B2(n_77),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_44),
.Y(n_151)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_12),
.A2(n_76),
.B1(n_77),
.B2(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_12),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_176),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_176),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_12),
.A2(n_47),
.B1(n_50),
.B2(n_176),
.Y(n_262)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx11_ASAP7_75t_SL g48 ( 
.A(n_15),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_131),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_129),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_104),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_19),
.B(n_104),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_85),
.B2(n_86),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_58),
.B2(n_59),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_23),
.A2(n_24),
.B(n_41),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_41),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_33),
.B1(n_36),
.B2(n_39),
.Y(n_24)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_25),
.B(n_69),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_25),
.A2(n_33),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_25),
.A2(n_33),
.B1(n_170),
.B2(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_25),
.A2(n_33),
.B1(n_200),
.B2(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_33),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_27),
.Y(n_213)
);

NAND2xp33_ASAP7_75t_SL g215 ( 
.A(n_27),
.B(n_35),
.Y(n_215)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_29),
.A2(n_30),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_29),
.B(n_73),
.Y(n_188)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_30),
.A2(n_80),
.B1(n_173),
.B2(n_188),
.Y(n_187)
);

AOI32xp33_ASAP7_75t_L g212 ( 
.A1(n_30),
.A2(n_34),
.A3(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_212)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_33),
.B(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_33),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_33),
.B(n_151),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_35),
.B1(n_49),
.B2(n_51),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_35),
.A2(n_49),
.B(n_174),
.C(n_241),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_37),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_39),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_52),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_42),
.A2(n_54),
.B(n_222),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_45),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_45),
.B(n_56),
.Y(n_100)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_54),
.B(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_46),
.A2(n_54),
.B1(n_99),
.B2(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_46),
.A2(n_52),
.B(n_119),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_46),
.A2(n_54),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_46),
.A2(n_54),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_46),
.A2(n_54),
.B1(n_221),
.B2(n_239),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_46),
.B(n_174),
.Y(n_260)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_47),
.Y(n_50)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_50),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_54),
.A2(n_99),
.B(n_100),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_54),
.A2(n_63),
.B(n_100),
.Y(n_167)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_70),
.B1(n_83),
.B2(n_84),
.Y(n_59)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B(n_68),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_66),
.A2(n_68),
.B(n_150),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_66),
.A2(n_184),
.B(n_185),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_70),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_75),
.B(n_78),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_82),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_71),
.A2(n_125),
.B1(n_126),
.B2(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_71),
.A2(n_125),
.B1(n_154),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_73),
.B(n_77),
.C(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_72),
.B(n_102),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_72),
.A2(n_79),
.B1(n_173),
.B2(n_175),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_77),
.Y(n_80)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

HAxp5_ASAP7_75t_SL g173 ( 
.A(n_77),
.B(n_174),
.CON(n_173),
.SN(n_173)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_102),
.B(n_103),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_97),
.B(n_101),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_101),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_87),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_87),
.A2(n_98),
.B1(n_108),
.B2(n_139),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_92),
.B(n_95),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_88),
.A2(n_143),
.B(n_144),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_88),
.A2(n_143),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_88),
.A2(n_117),
.B(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_88),
.A2(n_91),
.B1(n_254),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_89),
.A2(n_96),
.B(n_145),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_89),
.A2(n_93),
.B1(n_253),
.B2(n_255),
.Y(n_252)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_91),
.B(n_174),
.Y(n_266)
);

INVx5_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_96),
.Y(n_117)
);

INVx11_ASAP7_75t_L g191 ( 
.A(n_93),
.Y(n_191)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_98),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_101),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.C(n_110),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_105),
.B(n_109),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_110),
.A2(n_111),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_120),
.C(n_123),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_118),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_113),
.B(n_118),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_114),
.A2(n_190),
.B(n_191),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_120),
.A2(n_123),
.B1(n_124),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_120),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B(n_128),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_159),
.B(n_305),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_156),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_133),
.B(n_156),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_138),
.C(n_140),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_134),
.A2(n_135),
.B1(n_138),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_138),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_140),
.B(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_149),
.C(n_152),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_141),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_148),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_148),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_149),
.A2(n_152),
.B1(n_153),
.B2(n_295),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_149),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_299),
.B(n_304),
.Y(n_159)
);

O2A1O1Ixp33_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_204),
.B(n_285),
.C(n_298),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_192),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_162),
.B(n_192),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_177),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_164),
.B(n_165),
.C(n_177),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.C(n_172),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_172),
.B(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_175),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_186),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_182),
.B2(n_183),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_179),
.B(n_183),
.C(n_186),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_189),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.C(n_198),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_193),
.A2(n_194),
.B1(n_280),
.B2(n_282),
.Y(n_279)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_281),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_198),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.C(n_203),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_203),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_284),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_277),
.B(n_283),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_232),
.B(n_276),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_223),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_208),
.B(n_223),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_216),
.C(n_219),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_209),
.A2(n_210),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_212),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_228),
.B2(n_229),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_224),
.B(n_230),
.C(n_231),
.Y(n_278)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_270),
.B(n_275),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_250),
.B(n_269),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_242),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_235),
.B(n_242),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_240),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_236),
.A2(n_237),
.B1(n_240),
.B2(n_257),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_240),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_248),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_244),
.B(n_247),
.C(n_248),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_249),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_258),
.B(n_268),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_256),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_252),
.B(n_256),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_263),
.B(n_267),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_260),
.B(n_261),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_271),
.B(n_272),
.Y(n_275)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_278),
.B(n_279),
.Y(n_283)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_280),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_286),
.B(n_287),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_296),
.B2(n_297),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_293),
.C(n_297),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_296),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_300),
.B(n_301),
.Y(n_304)
);


endmodule