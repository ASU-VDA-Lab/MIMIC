module fake_jpeg_19748_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_10),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_21),
.B(n_9),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_39),
.B(n_44),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_32),
.Y(n_57)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_9),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_47),
.Y(n_75)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_19),
.B(n_9),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_50),
.B(n_30),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_56),
.B(n_61),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_57),
.B(n_90),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_44),
.B(n_19),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_59),
.B(n_74),
.Y(n_104)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_62),
.B(n_65),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_36),
.B1(n_25),
.B2(n_33),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_64),
.A2(n_80),
.B1(n_86),
.B2(n_89),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_29),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_29),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_67),
.B(n_69),
.Y(n_122)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_79),
.Y(n_124)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_30),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_40),
.A2(n_25),
.B1(n_36),
.B2(n_33),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_76),
.A2(n_77),
.B1(n_78),
.B2(n_83),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_40),
.A2(n_25),
.B1(n_36),
.B2(n_33),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_37),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_45),
.A2(n_36),
.B1(n_16),
.B2(n_37),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_81),
.B(n_82),
.Y(n_133)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_42),
.A2(n_16),
.B1(n_31),
.B2(n_18),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_41),
.A2(n_18),
.B1(n_20),
.B2(n_31),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_87),
.A2(n_24),
.B1(n_22),
.B2(n_28),
.Y(n_115)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_42),
.A2(n_20),
.B1(n_22),
.B2(n_27),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_27),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_34),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_91),
.Y(n_128)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_39),
.B(n_34),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_39),
.B(n_34),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_39),
.B(n_28),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_97),
.B(n_100),
.Y(n_127)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_41),
.B(n_27),
.C(n_35),
.Y(n_99)
);

FAx1_ASAP7_75t_SL g106 ( 
.A(n_99),
.B(n_22),
.CI(n_27),
.CON(n_106),
.SN(n_106)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_39),
.B(n_28),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_106),
.B(n_134),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

BUFx12_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_110),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_78),
.B1(n_58),
.B2(n_55),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_58),
.B1(n_55),
.B2(n_72),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_75),
.A2(n_22),
.B1(n_38),
.B2(n_17),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_126),
.Y(n_150)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_26),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_91),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_136),
.B(n_144),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_137),
.A2(n_141),
.B1(n_142),
.B2(n_159),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_108),
.B(n_66),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_143),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_114),
.A2(n_86),
.B1(n_80),
.B2(n_89),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_108),
.B(n_73),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_60),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_145),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_134),
.A2(n_106),
.B(n_128),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_147),
.A2(n_163),
.B(n_164),
.Y(n_173)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_149),
.B(n_157),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_63),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_151),
.B(n_152),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_104),
.B(n_77),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_96),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_166),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_127),
.B(n_11),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_109),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_115),
.A2(n_64),
.B1(n_75),
.B2(n_70),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_102),
.Y(n_160)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_161),
.Y(n_201)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_162),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_121),
.Y(n_163)
);

O2A1O1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_106),
.A2(n_92),
.B(n_61),
.C(n_54),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_112),
.B(n_53),
.Y(n_166)
);

AO21x1_ASAP7_75t_L g167 ( 
.A1(n_127),
.A2(n_22),
.B(n_68),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_94),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_116),
.A2(n_94),
.B1(n_24),
.B2(n_12),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_168),
.A2(n_141),
.B1(n_164),
.B2(n_135),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_26),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_107),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_124),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_SL g172 ( 
.A(n_152),
.B(n_151),
.C(n_140),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_172),
.B(n_175),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_161),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_111),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_176),
.A2(n_188),
.B(n_193),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_107),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_156),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_154),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_179),
.B(n_184),
.Y(n_220)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_182),
.Y(n_216)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_183),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_160),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_186),
.A2(n_105),
.B1(n_153),
.B2(n_121),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_189),
.Y(n_223)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_138),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_190),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_164),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_200),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_168),
.A2(n_111),
.B1(n_113),
.B2(n_117),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_199),
.A2(n_117),
.B1(n_158),
.B2(n_163),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_166),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_167),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_202),
.Y(n_233)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_138),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_204),
.Y(n_213)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_145),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_L g208 ( 
.A1(n_205),
.A2(n_156),
.B(n_167),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_229),
.Y(n_235)
);

AO21x1_ASAP7_75t_L g236 ( 
.A1(n_208),
.A2(n_205),
.B(n_196),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_186),
.A2(n_137),
.B1(n_169),
.B2(n_157),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_209),
.A2(n_219),
.B1(n_176),
.B2(n_188),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_211),
.A2(n_218),
.B1(n_226),
.B2(n_183),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_150),
.C(n_130),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_230),
.C(n_201),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_150),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_217),
.B(n_224),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_129),
.B1(n_130),
.B2(n_113),
.Y(n_218)
);

NOR2x1_ASAP7_75t_L g221 ( 
.A(n_172),
.B(n_162),
.Y(n_221)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_165),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_193),
.A2(n_105),
.B1(n_131),
.B2(n_139),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_181),
.B(n_139),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_231),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_165),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_228),
.B(n_232),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_173),
.B(n_131),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_173),
.B(n_120),
.C(n_110),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_181),
.B(n_26),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_120),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_110),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_191),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_239),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_237),
.A2(n_240),
.B1(n_245),
.B2(n_218),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_219),
.A2(n_185),
.B1(n_176),
.B2(n_171),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_212),
.B(n_174),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_241),
.B(n_221),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_214),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_252),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_243),
.B(n_244),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_187),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_209),
.A2(n_185),
.B1(n_171),
.B2(n_182),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_213),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_248),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_230),
.A2(n_194),
.B1(n_189),
.B2(n_177),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_249),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_233),
.A2(n_203),
.B1(n_190),
.B2(n_180),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_253),
.Y(n_267)
);

AOI221xp5_ASAP7_75t_L g252 ( 
.A1(n_221),
.A2(n_204),
.B1(n_180),
.B2(n_38),
.C(n_17),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_220),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_192),
.C(n_195),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_222),
.C(n_225),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_222),
.A2(n_195),
.B(n_110),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_233),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_231),
.Y(n_256)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_256),
.Y(n_260)
);

INVxp67_ASAP7_75t_SL g258 ( 
.A(n_253),
.Y(n_258)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_251),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_272),
.Y(n_278)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_247),
.Y(n_261)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_257),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_268),
.A2(n_257),
.B(n_246),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_269),
.A2(n_271),
.B1(n_266),
.B2(n_260),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_187),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_270),
.B(n_274),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_245),
.A2(n_226),
.B1(n_211),
.B2(n_213),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_247),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_254),
.C(n_239),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_238),
.B(n_223),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_276),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_242),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_263),
.Y(n_295)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_281),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_285),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_292),
.C(n_279),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_260),
.A2(n_276),
.B(n_272),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_288),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_269),
.A2(n_237),
.B1(n_240),
.B2(n_236),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_255),
.B(n_225),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_291),
.Y(n_293)
);

OAI21xp33_ASAP7_75t_L g290 ( 
.A1(n_259),
.A2(n_275),
.B(n_264),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_290),
.A2(n_265),
.B(n_223),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_210),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_235),
.C(n_249),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_301),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_266),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_298),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_261),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_304),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_302),
.C(n_285),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_265),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_235),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_283),
.C(n_288),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_278),
.B(n_271),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_277),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_308),
.C(n_312),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_282),
.C(n_284),
.Y(n_308)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_309),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_293),
.A2(n_210),
.B(n_216),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_310),
.A2(n_313),
.B(n_314),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_289),
.C(n_216),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_304),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_296),
.A2(n_287),
.B(n_13),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_303),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_11),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_301),
.C(n_315),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_321),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_294),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_295),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_323),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_192),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_324),
.B(n_328),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_322),
.A2(n_125),
.B(n_10),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_317),
.C(n_316),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_125),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_329),
.A2(n_331),
.B(n_327),
.Y(n_332)
);

AOI321xp33_ASAP7_75t_L g331 ( 
.A1(n_326),
.A2(n_318),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C(n_4),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_330),
.B(n_324),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_333),
.B(n_8),
.Y(n_334)
);


endmodule