module real_jpeg_812_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_120;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_1),
.A2(n_43),
.B1(n_44),
.B2(n_64),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_1),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_1),
.A2(n_22),
.B1(n_23),
.B2(n_64),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_1),
.A2(n_28),
.B1(n_30),
.B2(n_64),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_3),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_3),
.A2(n_22),
.B1(n_23),
.B2(n_66),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_3),
.A2(n_28),
.B1(n_30),
.B2(n_66),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_4),
.A2(n_22),
.B1(n_23),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_4),
.A2(n_28),
.B1(n_30),
.B2(n_36),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_5),
.A2(n_28),
.B1(n_30),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_6),
.A2(n_28),
.B1(n_30),
.B2(n_77),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_6),
.Y(n_77)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_10),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_10),
.B(n_70),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_10),
.A2(n_42),
.B(n_43),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_10),
.B(n_25),
.C(n_30),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_10),
.A2(n_22),
.B1(n_23),
.B2(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_10),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_10),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_10),
.B(n_52),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_10),
.B(n_88),
.Y(n_121)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_12),
.A2(n_22),
.B1(n_23),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_12),
.A2(n_28),
.B1(n_30),
.B2(n_33),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_91),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_89),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_79),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_17),
.B(n_79),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_58),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_37),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_31),
.B(n_34),
.Y(n_19)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_20),
.A2(n_88),
.B1(n_100),
.B2(n_102),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_20),
.A2(n_86),
.B1(n_88),
.B2(n_102),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_27),
.Y(n_20)
);

OAI22xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_21)
);

NAND3xp33_ASAP7_75t_L g46 ( 
.A(n_22),
.B(n_44),
.C(n_47),
.Y(n_46)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_22),
.A2(n_23),
.B1(n_39),
.B2(n_47),
.Y(n_62)
);

CKINVDCx6p67_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

A2O1A1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_23),
.A2(n_39),
.B(n_41),
.C(n_46),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_23),
.B(n_97),
.Y(n_96)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_25),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_30),
.B(n_115),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_32),
.A2(n_84),
.B1(n_85),
.B2(n_87),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_48),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_38),
.B(n_48),
.Y(n_80)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_43),
.B1(n_44),
.B2(n_47),
.Y(n_61)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_44),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_54),
.B(n_55),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_49),
.A2(n_51),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_50),
.B(n_56),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_50),
.A2(n_105),
.B(n_106),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_50),
.A2(n_52),
.B1(n_101),
.B2(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_50),
.A2(n_52),
.B1(n_117),
.B2(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_51),
.A2(n_76),
.B(n_78),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_51),
.B(n_54),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_52),
.B(n_56),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_67),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_62),
.B1(n_63),
.B2(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.C(n_83),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_80),
.B(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_81),
.B(n_83),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_130),
.B(n_134),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_111),
.B(n_129),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_103),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_103),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_95),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_108),
.C(n_109),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_105),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_123),
.B(n_128),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_118),
.B(n_122),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_121),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_127),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_131),
.B(n_132),
.Y(n_134)
);


endmodule