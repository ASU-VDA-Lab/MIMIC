module fake_jpeg_8266_n_53 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_53);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_53;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_0),
.B(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

INVxp33_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

FAx1_ASAP7_75t_SL g27 ( 
.A(n_21),
.B(n_0),
.CI(n_1),
.CON(n_27),
.SN(n_27)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_27),
.B(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_29),
.B(n_32),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_20),
.C(n_25),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_34),
.C(n_35),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_2),
.B1(n_5),
.B2(n_7),
.Y(n_34)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_41),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_30),
.A2(n_10),
.B(n_14),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_26),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_49),
.C(n_46),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_43),
.B(n_42),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_45),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_38),
.B(n_36),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_38),
.B(n_36),
.Y(n_53)
);


endmodule