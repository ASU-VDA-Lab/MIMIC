module fake_ibex_1300_n_2405 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_108, n_350, n_165, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_421, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_244, n_73, n_343, n_310, n_426, n_323, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_434, n_296, n_120, n_168, n_155, n_315, n_441, n_13, n_122, n_116, n_370, n_431, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_22, n_136, n_261, n_30, n_367, n_221, n_437, n_355, n_407, n_102, n_52, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_420, n_141, n_222, n_186, n_349, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_429, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_445, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_416, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_26, n_188, n_200, n_444, n_199, n_410, n_308, n_411, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_381, n_382, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_408, n_119, n_361, n_419, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_443, n_344, n_393, n_436, n_428, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_399, n_254, n_213, n_424, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_425, n_2405);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_108;
input n_350;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_434;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_116;
input n_370;
input n_431;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_367;
input n_221;
input n_437;
input n_355;
input n_407;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_141;
input n_222;
input n_186;
input n_349;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_429;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_416;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_26;
input n_188;
input n_200;
input n_444;
input n_199;
input n_410;
input n_308;
input n_411;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_381;
input n_382;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_419;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_443;
input n_344;
input n_393;
input n_436;
input n_428;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_399;
input n_254;
input n_213;
input n_424;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;
input n_425;

output n_2405;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_2201;
wire n_766;
wire n_2175;
wire n_2071;
wire n_1110;
wire n_1382;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_452;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_773;
wire n_2038;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_957;
wire n_1652;
wire n_969;
wire n_678;
wire n_1954;
wire n_2183;
wire n_1859;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_2276;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2139;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_884;
wire n_667;
wire n_2396;
wire n_850;
wire n_1971;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_557;
wire n_641;
wire n_1937;
wire n_2311;
wire n_527;
wire n_893;
wire n_1654;
wire n_496;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_2015;
wire n_1130;
wire n_1228;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_538;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2003;
wire n_1970;
wire n_1778;
wire n_448;
wire n_646;
wire n_466;
wire n_2347;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2362;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_2090;
wire n_666;
wire n_2260;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_793;
wire n_937;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_2393;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_2283;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_553;
wire n_554;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_2373;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_2275;
wire n_2189;
wire n_745;
wire n_2112;
wire n_447;
wire n_1753;
wire n_564;
wire n_562;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2171;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_1350;
wire n_451;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_579;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_2401;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2350;
wire n_1742;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_2203;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_455;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2256;
wire n_606;
wire n_737;
wire n_1571;
wire n_1980;
wire n_462;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2355;
wire n_1543;
wire n_823;
wire n_2233;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2377;
wire n_1591;
wire n_583;
wire n_2289;
wire n_2288;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2101;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_1831;
wire n_864;
wire n_608;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_846;
wire n_471;
wire n_1793;
wire n_1237;
wire n_2390;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_2375;
wire n_458;
wire n_1498;
wire n_2312;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_469;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_1589;
wire n_2204;
wire n_1210;
wire n_2319;
wire n_591;
wire n_1933;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2006;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_2358;
wire n_594;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_585;
wire n_1982;
wire n_2252;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_483;
wire n_1695;
wire n_1418;
wire n_2402;
wire n_1137;
wire n_660;
wire n_524;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_576;
wire n_1602;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_827;
wire n_607;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_2287;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_488;
wire n_705;
wire n_2142;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_472;
wire n_1704;
wire n_2160;
wire n_2234;
wire n_847;
wire n_1436;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_456;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_801;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_1836;
wire n_2398;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_650;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_517;
wire n_817;
wire n_2193;
wire n_2095;
wire n_555;
wire n_2395;
wire n_951;
wire n_2053;
wire n_468;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_502;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_863;
wire n_597;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_2376;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_2170;
wire n_1785;
wire n_486;
wire n_1870;
wire n_1405;
wire n_997;
wire n_2308;
wire n_1428;
wire n_2243;
wire n_2400;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_485;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_1925;
wire n_2106;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_890;
wire n_628;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_2298;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1845;
wire n_1104;
wire n_2205;
wire n_1011;
wire n_1667;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2064;
wire n_1679;
wire n_2342;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1997;
wire n_1894;
wire n_2110;
wire n_634;
wire n_961;
wire n_991;
wire n_1331;
wire n_1223;
wire n_1349;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_1629;
wire n_2011;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_2344;
wire n_2317;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_1099;
wire n_598;
wire n_2141;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2210;
wire n_1517;
wire n_690;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_2087;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_2380;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2120;
wire n_1037;
wire n_2031;
wire n_1899;
wire n_464;
wire n_1348;
wire n_838;
wire n_1289;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_2309;
wire n_842;
wire n_2274;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_636;
wire n_1259;
wire n_490;
wire n_2108;
wire n_595;
wire n_1001;
wire n_570;
wire n_2143;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_1538;
wire n_487;
wire n_454;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2351;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_1725;
wire n_2149;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_648;
wire n_571;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_473;
wire n_1241;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_1270;
wire n_834;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2012;
wire n_722;
wire n_2251;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_480;
wire n_2182;
wire n_1057;
wire n_1473;
wire n_516;
wire n_2125;
wire n_1403;
wire n_2181;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_950;
wire n_512;
wire n_685;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_2315;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_2272;
wire n_535;
wire n_1956;
wire n_681;
wire n_1718;
wire n_2225;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_505;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_1085;
wire n_2388;
wire n_2222;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_2135;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2232;
wire n_2121;
wire n_1893;
wire n_1570;
wire n_2231;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_1961;
wire n_1050;
wire n_2218;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_1632;
wire n_688;
wire n_1547;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1542;
wire n_1097;
wire n_1909;
wire n_2381;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_1940;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_1767;
wire n_1939;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_478;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2156;
wire n_753;
wire n_2126;
wire n_747;
wire n_645;
wire n_1147;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1518;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_682;
wire n_2061;
wire n_1373;
wire n_1686;
wire n_2131;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_755;
wire n_2091;
wire n_1029;
wire n_2394;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_2337;
wire n_854;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_2323;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_2371;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_569;
wire n_2305;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_2048;
wire n_987;
wire n_750;
wire n_1299;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_2227;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_1692;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_2291;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2303;
wire n_2357;
wire n_924;
wire n_2331;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2092;
wire n_566;
wire n_581;
wire n_1365;
wire n_1472;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_548;
wire n_1158;
wire n_1974;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_2168;
wire n_1948;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2378;
wire n_888;
wire n_1325;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2073;
wire n_952;
wire n_1947;
wire n_1675;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_1468;
wire n_2327;
wire n_913;
wire n_2353;
wire n_509;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_2321;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_519;
wire n_1843;
wire n_2186;
wire n_2030;
wire n_1665;
wire n_1091;
wire n_1780;
wire n_1678;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_2282;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;

INVx1_ASAP7_75t_SL g446 ( 
.A(n_177),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_274),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_170),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_119),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_84),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_297),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_408),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_175),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_231),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_254),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_386),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_161),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_334),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_442),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_193),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_419),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_285),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_266),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_392),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_444),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_196),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_396),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_435),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_389),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g470 ( 
.A(n_255),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_331),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_194),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_344),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_87),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_397),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_307),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_418),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_399),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_160),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_226),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_325),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_108),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_391),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_110),
.Y(n_484)
);

NOR2xp67_ASAP7_75t_L g485 ( 
.A(n_179),
.B(n_134),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_95),
.Y(n_486)
);

NOR2xp67_ASAP7_75t_L g487 ( 
.A(n_37),
.B(n_5),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_90),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_71),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_328),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_128),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_438),
.Y(n_492)
);

BUFx8_ASAP7_75t_SL g493 ( 
.A(n_421),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_113),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_401),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_45),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_343),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_254),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_62),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_336),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_409),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_443),
.B(n_199),
.Y(n_502)
);

NOR2xp67_ASAP7_75t_L g503 ( 
.A(n_413),
.B(n_102),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_317),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_259),
.Y(n_505)
);

CKINVDCx16_ASAP7_75t_R g506 ( 
.A(n_28),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_298),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_167),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_363),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_116),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_0),
.Y(n_511)
);

NOR2xp67_ASAP7_75t_L g512 ( 
.A(n_355),
.B(n_78),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_358),
.B(n_406),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_189),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_433),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_365),
.Y(n_516)
);

INVxp33_ASAP7_75t_SL g517 ( 
.A(n_427),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_128),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_200),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_102),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_415),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_122),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_318),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_405),
.Y(n_524)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_403),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_315),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_440),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_213),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_439),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_51),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_260),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_177),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_183),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_58),
.Y(n_534)
);

BUFx10_ASAP7_75t_L g535 ( 
.A(n_250),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_206),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_436),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_298),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_412),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_47),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_220),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_326),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_243),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_220),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_61),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_171),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_219),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_304),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_90),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_262),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_89),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_69),
.Y(n_552)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_360),
.Y(n_553)
);

NOR2xp67_ASAP7_75t_L g554 ( 
.A(n_313),
.B(n_267),
.Y(n_554)
);

INVx1_ASAP7_75t_SL g555 ( 
.A(n_96),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_19),
.Y(n_556)
);

NOR2xp67_ASAP7_75t_L g557 ( 
.A(n_1),
.B(n_236),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_278),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_300),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_398),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_341),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_285),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_245),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_84),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_387),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_366),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_420),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_44),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_106),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_445),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_99),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_273),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_422),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_191),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_290),
.Y(n_575)
);

BUFx10_ASAP7_75t_L g576 ( 
.A(n_156),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_49),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_100),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_372),
.Y(n_579)
);

BUFx2_ASAP7_75t_L g580 ( 
.A(n_100),
.Y(n_580)
);

BUFx5_ASAP7_75t_L g581 ( 
.A(n_306),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_346),
.Y(n_582)
);

INVxp67_ASAP7_75t_SL g583 ( 
.A(n_216),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_15),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_189),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_203),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_441),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_5),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_262),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_82),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_127),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_432),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_375),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_33),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_268),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_337),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_342),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_46),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_190),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_252),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_226),
.Y(n_601)
);

BUFx2_ASAP7_75t_L g602 ( 
.A(n_192),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_50),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_390),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_143),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_87),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_205),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_240),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_253),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_217),
.Y(n_610)
);

BUFx10_ASAP7_75t_L g611 ( 
.A(n_340),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_215),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_434),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_15),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_423),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_159),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_140),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_50),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_22),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_247),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_39),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_60),
.Y(n_622)
);

INVx4_ASAP7_75t_R g623 ( 
.A(n_275),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_74),
.B(n_71),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_271),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_253),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_49),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_170),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_368),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_255),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_97),
.Y(n_631)
);

INVxp67_ASAP7_75t_L g632 ( 
.A(n_36),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_184),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_73),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_240),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_286),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_176),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_350),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_301),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_335),
.Y(n_640)
);

NOR2xp67_ASAP7_75t_L g641 ( 
.A(n_188),
.B(n_277),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_144),
.Y(n_642)
);

INVxp67_ASAP7_75t_SL g643 ( 
.A(n_46),
.Y(n_643)
);

CKINVDCx14_ASAP7_75t_R g644 ( 
.A(n_53),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_296),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_17),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_227),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_349),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_426),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_376),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_224),
.B(n_113),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_195),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_22),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_293),
.B(n_385),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_430),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g656 ( 
.A(n_164),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_291),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_264),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_204),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_11),
.Y(n_660)
);

NOR2xp67_ASAP7_75t_L g661 ( 
.A(n_55),
.B(n_424),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_388),
.Y(n_662)
);

CKINVDCx16_ASAP7_75t_R g663 ( 
.A(n_206),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_17),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_214),
.Y(n_665)
);

BUFx2_ASAP7_75t_L g666 ( 
.A(n_4),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_261),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_41),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_154),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_251),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_43),
.Y(n_671)
);

CKINVDCx16_ASAP7_75t_R g672 ( 
.A(n_282),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_431),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_369),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_428),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_56),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_370),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_269),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_175),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_347),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_323),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_404),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_429),
.Y(n_683)
);

INVx1_ASAP7_75t_SL g684 ( 
.A(n_289),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_357),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_383),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_35),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_425),
.Y(n_688)
);

INVxp67_ASAP7_75t_SL g689 ( 
.A(n_402),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_288),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_166),
.Y(n_691)
);

BUFx10_ASAP7_75t_L g692 ( 
.A(n_382),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_299),
.Y(n_693)
);

INVx1_ASAP7_75t_SL g694 ( 
.A(n_89),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_284),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_131),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_171),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_322),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_242),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_407),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_211),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_192),
.B(n_359),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_292),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_384),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_381),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_356),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_394),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_345),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_211),
.Y(n_709)
);

CKINVDCx20_ASAP7_75t_R g710 ( 
.A(n_194),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_116),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_129),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_327),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_58),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_130),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_380),
.Y(n_716)
);

INVx1_ASAP7_75t_SL g717 ( 
.A(n_140),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_416),
.Y(n_718)
);

BUFx5_ASAP7_75t_L g719 ( 
.A(n_374),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_305),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_16),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_354),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_411),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_99),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_24),
.Y(n_725)
);

CKINVDCx16_ASAP7_75t_R g726 ( 
.A(n_4),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_52),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_437),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_400),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_51),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_414),
.Y(n_731)
);

CKINVDCx16_ASAP7_75t_R g732 ( 
.A(n_227),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_283),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_78),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_417),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_104),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_98),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_306),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_410),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_95),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_43),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_237),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_149),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_221),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_155),
.Y(n_745)
);

BUFx10_ASAP7_75t_L g746 ( 
.A(n_217),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_622),
.B(n_0),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_475),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_490),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_644),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_448),
.B(n_2),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_490),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_580),
.B(n_3),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_475),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_622),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_490),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_602),
.B(n_6),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_611),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_581),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_644),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_469),
.B(n_7),
.Y(n_761)
);

OAI22x1_ASAP7_75t_R g762 ( 
.A1(n_447),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_762)
);

INVx6_ASAP7_75t_L g763 ( 
.A(n_611),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_462),
.B(n_9),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_581),
.Y(n_765)
);

OAI21x1_ASAP7_75t_L g766 ( 
.A1(n_464),
.A2(n_310),
.B(n_309),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_470),
.A2(n_506),
.B1(n_672),
.B2(n_663),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_581),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_475),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_581),
.Y(n_770)
);

BUFx12f_ASAP7_75t_L g771 ( 
.A(n_611),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_634),
.B(n_10),
.Y(n_772)
);

INVxp67_ASAP7_75t_L g773 ( 
.A(n_666),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_614),
.B(n_12),
.Y(n_774)
);

OA21x2_ASAP7_75t_L g775 ( 
.A1(n_464),
.A2(n_312),
.B(n_311),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_504),
.Y(n_776)
);

OAI22x1_ASAP7_75t_L g777 ( 
.A1(n_690),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_462),
.Y(n_778)
);

BUFx8_ASAP7_75t_L g779 ( 
.A(n_581),
.Y(n_779)
);

INVxp67_ASAP7_75t_L g780 ( 
.A(n_636),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_504),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_549),
.A2(n_16),
.B1(n_13),
.B2(n_14),
.Y(n_782)
);

INVx5_ASAP7_75t_L g783 ( 
.A(n_504),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_549),
.B(n_714),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_714),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_581),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_569),
.B(n_18),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_527),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_SL g789 ( 
.A(n_493),
.B(n_314),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_719),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_656),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_660),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_727),
.Y(n_793)
);

BUFx2_ASAP7_75t_L g794 ( 
.A(n_733),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_726),
.B(n_18),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_727),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_719),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_719),
.Y(n_798)
);

BUFx2_ASAP7_75t_L g799 ( 
.A(n_733),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_719),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_690),
.Y(n_801)
);

AND2x4_ASAP7_75t_L g802 ( 
.A(n_463),
.B(n_19),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_719),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_732),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_577),
.B(n_20),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_472),
.B(n_20),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_529),
.B(n_21),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_527),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_527),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_632),
.B(n_21),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_719),
.Y(n_811)
);

CKINVDCx16_ASAP7_75t_R g812 ( 
.A(n_535),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_709),
.B(n_23),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_474),
.Y(n_814)
);

INVx4_ASAP7_75t_L g815 ( 
.A(n_692),
.Y(n_815)
);

BUFx2_ASAP7_75t_L g816 ( 
.A(n_493),
.Y(n_816)
);

BUFx2_ASAP7_75t_L g817 ( 
.A(n_709),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_517),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_474),
.Y(n_819)
);

INVx5_ASAP7_75t_L g820 ( 
.A(n_649),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_449),
.B(n_25),
.Y(n_821)
);

OA21x2_ASAP7_75t_L g822 ( 
.A1(n_497),
.A2(n_319),
.B(n_316),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_535),
.B(n_576),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_553),
.B(n_26),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_692),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_719),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_482),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_497),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_454),
.B(n_27),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_508),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_508),
.Y(n_831)
);

BUFx12f_ASAP7_75t_L g832 ( 
.A(n_692),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_501),
.Y(n_833)
);

OAI22xp5_ASAP7_75t_L g834 ( 
.A1(n_651),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_834)
);

INVx5_ASAP7_75t_L g835 ( 
.A(n_649),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_535),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_649),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_520),
.Y(n_838)
);

OA21x2_ASAP7_75t_L g839 ( 
.A1(n_501),
.A2(n_321),
.B(n_320),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_450),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_520),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_563),
.B(n_29),
.Y(n_842)
);

AND3x2_ASAP7_75t_L g843 ( 
.A(n_816),
.B(n_643),
.C(n_583),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_816),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_815),
.B(n_481),
.Y(n_845)
);

NAND2xp33_ASAP7_75t_SL g846 ( 
.A(n_807),
.B(n_468),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_779),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_759),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_817),
.Y(n_849)
);

OR2x2_ASAP7_75t_L g850 ( 
.A(n_817),
.B(n_446),
.Y(n_850)
);

OR2x6_ASAP7_75t_L g851 ( 
.A(n_771),
.B(n_485),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_765),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_765),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_768),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_779),
.Y(n_855)
);

BUFx2_ASAP7_75t_L g856 ( 
.A(n_823),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_768),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_770),
.Y(n_858)
);

OR2x2_ASAP7_75t_L g859 ( 
.A(n_812),
.B(n_466),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_770),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_784),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_747),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_786),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_784),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_786),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_790),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_758),
.B(n_680),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_823),
.B(n_680),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_794),
.B(n_763),
.Y(n_869)
);

INVx5_ASAP7_75t_L g870 ( 
.A(n_783),
.Y(n_870)
);

NAND2xp33_ASAP7_75t_L g871 ( 
.A(n_797),
.B(n_513),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_771),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_797),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_798),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_748),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_800),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_780),
.A2(n_517),
.B1(n_565),
.B2(n_468),
.Y(n_877)
);

AO21x2_ASAP7_75t_L g878 ( 
.A1(n_766),
.A2(n_456),
.B(n_452),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_758),
.B(n_682),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_779),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_803),
.Y(n_881)
);

AND3x2_ASAP7_75t_L g882 ( 
.A(n_789),
.B(n_624),
.C(n_689),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_803),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_801),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_811),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_802),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_811),
.Y(n_887)
);

BUFx6f_ASAP7_75t_SL g888 ( 
.A(n_764),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_826),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_802),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_756),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_773),
.A2(n_615),
.B1(n_629),
.B2(n_565),
.Y(n_892)
);

AO21x2_ASAP7_75t_L g893 ( 
.A1(n_766),
.A2(n_461),
.B(n_458),
.Y(n_893)
);

NAND2xp33_ASAP7_75t_L g894 ( 
.A(n_825),
.B(n_649),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_748),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_749),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_763),
.B(n_465),
.Y(n_897)
);

INVxp67_ASAP7_75t_SL g898 ( 
.A(n_791),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_748),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_763),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_748),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_754),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_764),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_778),
.B(n_785),
.Y(n_904)
);

NOR2x1p5_ASAP7_75t_L g905 ( 
.A(n_832),
.B(n_536),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_754),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_836),
.B(n_707),
.Y(n_907)
);

AOI21x1_ASAP7_75t_L g908 ( 
.A1(n_752),
.A2(n_686),
.B(n_638),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_754),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_754),
.Y(n_910)
);

AO21x2_ASAP7_75t_L g911 ( 
.A1(n_821),
.A2(n_477),
.B(n_473),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_769),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_752),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_793),
.B(n_478),
.Y(n_914)
);

AO21x2_ASAP7_75t_L g915 ( 
.A1(n_813),
.A2(n_495),
.B(n_483),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_769),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_802),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_828),
.Y(n_918)
);

OR2x2_ASAP7_75t_L g919 ( 
.A(n_792),
.B(n_555),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_806),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_828),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_799),
.B(n_746),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_806),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_832),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_784),
.B(n_681),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_796),
.B(n_681),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_840),
.B(n_683),
.Y(n_927)
);

INVx1_ASAP7_75t_SL g928 ( 
.A(n_807),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_833),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_833),
.Y(n_930)
);

INVx4_ASAP7_75t_L g931 ( 
.A(n_806),
.Y(n_931)
);

AO21x2_ASAP7_75t_L g932 ( 
.A1(n_805),
.A2(n_509),
.B(n_500),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_755),
.B(n_685),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_751),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_842),
.Y(n_935)
);

CKINVDCx20_ASAP7_75t_R g936 ( 
.A(n_804),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_751),
.B(n_685),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_776),
.Y(n_938)
);

BUFx10_ASAP7_75t_L g939 ( 
.A(n_842),
.Y(n_939)
);

INVx4_ASAP7_75t_L g940 ( 
.A(n_775),
.Y(n_940)
);

NAND2xp33_ASAP7_75t_L g941 ( 
.A(n_753),
.B(n_688),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_776),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_819),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_781),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_795),
.B(n_746),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_814),
.Y(n_946)
);

INVx5_ASAP7_75t_L g947 ( 
.A(n_783),
.Y(n_947)
);

NAND2xp33_ASAP7_75t_L g948 ( 
.A(n_829),
.B(n_688),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_788),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_841),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_795),
.Y(n_951)
);

AOI21x1_ASAP7_75t_L g952 ( 
.A1(n_775),
.A2(n_686),
.B(n_638),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_788),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_827),
.B(n_576),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_830),
.B(n_707),
.Y(n_955)
);

AO21x2_ASAP7_75t_L g956 ( 
.A1(n_774),
.A2(n_521),
.B(n_515),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_831),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_831),
.B(n_739),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_831),
.Y(n_959)
);

AOI21x1_ASAP7_75t_L g960 ( 
.A1(n_775),
.A2(n_722),
.B(n_704),
.Y(n_960)
);

AO21x2_ASAP7_75t_L g961 ( 
.A1(n_757),
.A2(n_524),
.B(n_523),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_829),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_838),
.Y(n_963)
);

BUFx10_ASAP7_75t_L g964 ( 
.A(n_824),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_808),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_808),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_767),
.B(n_526),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_809),
.Y(n_968)
);

AO21x2_ASAP7_75t_L g969 ( 
.A1(n_772),
.A2(n_539),
.B(n_537),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_824),
.B(n_542),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_783),
.Y(n_971)
);

AND3x2_ASAP7_75t_L g972 ( 
.A(n_762),
.B(n_476),
.C(n_457),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_809),
.Y(n_973)
);

INVx4_ASAP7_75t_L g974 ( 
.A(n_822),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_761),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_837),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_837),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_837),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_837),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_954),
.B(n_787),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_847),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_956),
.B(n_787),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_956),
.B(n_810),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_868),
.B(n_804),
.Y(n_984)
);

NAND3xp33_ASAP7_75t_L g985 ( 
.A(n_948),
.B(n_810),
.C(n_750),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_847),
.B(n_855),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_869),
.B(n_525),
.Y(n_987)
);

NOR3xp33_ASAP7_75t_L g988 ( 
.A(n_846),
.B(n_760),
.C(n_834),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_956),
.B(n_822),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_855),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_925),
.B(n_459),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_961),
.B(n_822),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_861),
.Y(n_993)
);

INVxp67_ASAP7_75t_L g994 ( 
.A(n_849),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_943),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_861),
.Y(n_996)
);

A2O1A1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_903),
.A2(n_480),
.B(n_498),
.C(n_484),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_898),
.B(n_451),
.Y(n_998)
);

OAI22xp33_ASAP7_75t_L g999 ( 
.A1(n_877),
.A2(n_928),
.B1(n_892),
.B2(n_919),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_961),
.B(n_839),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_880),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_969),
.B(n_839),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_975),
.B(n_937),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_969),
.B(n_560),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_969),
.B(n_566),
.Y(n_1005)
);

OR2x2_ASAP7_75t_L g1006 ( 
.A(n_919),
.B(n_684),
.Y(n_1006)
);

AOI221xp5_ASAP7_75t_L g1007 ( 
.A1(n_962),
.A2(n_777),
.B1(n_818),
.B2(n_507),
.C(n_514),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_943),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_867),
.B(n_467),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_880),
.B(n_471),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_943),
.Y(n_1011)
);

INVxp67_ASAP7_75t_SL g1012 ( 
.A(n_850),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_864),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_879),
.B(n_492),
.Y(n_1014)
);

NAND2x1_ASAP7_75t_L g1015 ( 
.A(n_931),
.B(n_623),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_934),
.B(n_782),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_964),
.B(n_845),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_856),
.B(n_516),
.Y(n_1018)
);

AOI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_948),
.A2(n_629),
.B1(n_706),
.B2(n_615),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_886),
.Y(n_1020)
);

BUFx5_ASAP7_75t_L g1021 ( 
.A(n_866),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_934),
.B(n_561),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_955),
.B(n_579),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_907),
.B(n_900),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_958),
.B(n_592),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_935),
.A2(n_723),
.B1(n_706),
.B2(n_455),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_939),
.B(n_593),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_945),
.B(n_613),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_940),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_939),
.B(n_640),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_939),
.B(n_648),
.Y(n_1031)
);

INVxp67_ASAP7_75t_L g1032 ( 
.A(n_859),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_922),
.B(n_655),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_922),
.B(n_675),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_967),
.A2(n_723),
.B1(n_738),
.B2(n_736),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_897),
.B(n_698),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_886),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_891),
.B(n_700),
.Y(n_1038)
);

NOR2xp67_ASAP7_75t_L g1039 ( 
.A(n_872),
.B(n_777),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_900),
.B(n_705),
.Y(n_1040)
);

NOR3xp33_ASAP7_75t_L g1041 ( 
.A(n_846),
.B(n_717),
.C(n_694),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_886),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_970),
.B(n_728),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_951),
.B(n_487),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_872),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_927),
.B(n_729),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_890),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_924),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_890),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_911),
.B(n_567),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_850),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_911),
.B(n_570),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_890),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_917),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_862),
.B(n_731),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_917),
.Y(n_1056)
);

OAI21xp33_ASAP7_75t_L g1057 ( 
.A1(n_935),
.A2(n_530),
.B(n_519),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_932),
.B(n_573),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_917),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_923),
.B(n_735),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_920),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_920),
.B(n_702),
.Y(n_1062)
);

AO221x1_ASAP7_75t_L g1063 ( 
.A1(n_972),
.A2(n_920),
.B1(n_844),
.B2(n_941),
.C(n_455),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_951),
.B(n_453),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_915),
.B(n_460),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_915),
.B(n_486),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_933),
.B(n_488),
.Y(n_1067)
);

NOR3xp33_ASAP7_75t_L g1068 ( 
.A(n_941),
.B(n_491),
.C(n_489),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_926),
.B(n_582),
.Y(n_1069)
);

OR2x2_ASAP7_75t_L g1070 ( 
.A(n_859),
.B(n_744),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_844),
.B(n_587),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_904),
.B(n_494),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_884),
.B(n_596),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_914),
.B(n_597),
.Y(n_1074)
);

NAND2xp33_ASAP7_75t_SL g1075 ( 
.A(n_888),
.B(n_502),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_871),
.B(n_950),
.Y(n_1076)
);

INVx2_ASAP7_75t_SL g1077 ( 
.A(n_905),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_851),
.B(n_496),
.Y(n_1078)
);

AO221x1_ASAP7_75t_L g1079 ( 
.A1(n_882),
.A2(n_505),
.B1(n_518),
.B2(n_479),
.C(n_447),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_871),
.B(n_950),
.Y(n_1080)
);

NAND3xp33_ASAP7_75t_L g1081 ( 
.A(n_940),
.B(n_510),
.C(n_499),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_946),
.B(n_511),
.Y(n_1082)
);

INVxp67_ASAP7_75t_L g1083 ( 
.A(n_918),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_851),
.B(n_604),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_921),
.B(n_929),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_957),
.Y(n_1086)
);

NAND2xp33_ASAP7_75t_SL g1087 ( 
.A(n_959),
.B(n_479),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_930),
.B(n_522),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_963),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_896),
.B(n_913),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_913),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_851),
.B(n_650),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_881),
.B(n_531),
.Y(n_1093)
);

INVx8_ASAP7_75t_L g1094 ( 
.A(n_851),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_843),
.B(n_532),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_857),
.B(n_534),
.Y(n_1096)
);

AOI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_894),
.A2(n_742),
.B1(n_734),
.B2(n_538),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_974),
.B(n_894),
.Y(n_1098)
);

OAI21xp33_ASAP7_75t_L g1099 ( 
.A1(n_858),
.A2(n_865),
.B(n_873),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_974),
.B(n_873),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_874),
.B(n_540),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_874),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_974),
.B(n_662),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_876),
.B(n_673),
.Y(n_1104)
);

NAND3xp33_ASAP7_75t_L g1105 ( 
.A(n_876),
.B(n_543),
.C(n_541),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_883),
.B(n_674),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_885),
.B(n_677),
.Y(n_1107)
);

AOI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_878),
.A2(n_548),
.B1(n_550),
.B2(n_545),
.Y(n_1108)
);

O2A1O1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_887),
.A2(n_547),
.B(n_552),
.C(n_546),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_889),
.B(n_551),
.Y(n_1110)
);

NOR2xp67_ASAP7_75t_L g1111 ( 
.A(n_908),
.B(n_30),
.Y(n_1111)
);

INVxp33_ASAP7_75t_L g1112 ( 
.A(n_936),
.Y(n_1112)
);

NOR3xp33_ASAP7_75t_L g1113 ( 
.A(n_936),
.B(n_564),
.C(n_558),
.Y(n_1113)
);

INVx2_ASAP7_75t_SL g1114 ( 
.A(n_878),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_848),
.B(n_568),
.Y(n_1115)
);

BUFx12f_ASAP7_75t_SL g1116 ( 
.A(n_875),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_848),
.B(n_572),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_878),
.B(n_578),
.Y(n_1118)
);

O2A1O1Ixp5_ASAP7_75t_L g1119 ( 
.A1(n_952),
.A2(n_708),
.B(n_716),
.C(n_713),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_852),
.B(n_586),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_853),
.B(n_589),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_853),
.B(n_590),
.Y(n_1122)
);

OR2x6_ASAP7_75t_L g1123 ( 
.A(n_960),
.B(n_557),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_854),
.B(n_718),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_893),
.B(n_641),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_893),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_854),
.B(n_860),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_893),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_863),
.B(n_591),
.Y(n_1129)
);

NAND2xp33_ASAP7_75t_L g1130 ( 
.A(n_971),
.B(n_528),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_971),
.B(n_563),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_870),
.B(n_659),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_870),
.B(n_659),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_SL g1134 ( 
.A(n_870),
.B(n_505),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_870),
.B(n_679),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_870),
.A2(n_544),
.B1(n_559),
.B2(n_518),
.Y(n_1136)
);

NAND2x1p5_ASAP7_75t_L g1137 ( 
.A(n_947),
.B(n_556),
.Y(n_1137)
);

INVx2_ASAP7_75t_SL g1138 ( 
.A(n_947),
.Y(n_1138)
);

O2A1O1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_968),
.A2(n_584),
.B(n_585),
.C(n_571),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_947),
.B(n_679),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_947),
.B(n_725),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_947),
.B(n_725),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_875),
.B(n_533),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_976),
.B(n_740),
.Y(n_1144)
);

NOR2x1p5_ASAP7_75t_L g1145 ( 
.A(n_895),
.B(n_598),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_899),
.B(n_740),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_875),
.B(n_533),
.Y(n_1147)
);

INVxp67_ASAP7_75t_L g1148 ( 
.A(n_899),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_SL g1149 ( 
.A(n_944),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_901),
.B(n_595),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_902),
.B(n_599),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_944),
.B(n_533),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_906),
.B(n_600),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_909),
.B(n_607),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_944),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_910),
.B(n_609),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_912),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_912),
.B(n_612),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_916),
.B(n_601),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1020),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1096),
.B(n_617),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1126),
.A2(n_654),
.B(n_512),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1037),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_981),
.B(n_603),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1076),
.A2(n_574),
.B1(n_594),
.B2(n_559),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_1032),
.B(n_574),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1080),
.A2(n_605),
.B1(n_695),
.B2(n_594),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_997),
.A2(n_618),
.B(n_625),
.C(n_621),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_994),
.B(n_605),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_999),
.A2(n_628),
.B(n_637),
.C(n_627),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1012),
.B(n_695),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_1029),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_1051),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_982),
.A2(n_642),
.B(n_647),
.C(n_639),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1070),
.B(n_696),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_989),
.A2(n_554),
.B(n_503),
.Y(n_1176)
);

INVx1_ASAP7_75t_SL g1177 ( 
.A(n_1021),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_1045),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1042),
.Y(n_1179)
);

OAI221xp5_ASAP7_75t_L g1180 ( 
.A1(n_1007),
.A2(n_610),
.B1(n_616),
.B2(n_608),
.C(n_606),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1047),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_982),
.B(n_983),
.Y(n_1182)
);

OAI22x1_ASAP7_75t_L g1183 ( 
.A1(n_1019),
.A2(n_697),
.B1(n_710),
.B2(n_696),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1026),
.Y(n_1184)
);

HB1xp67_ASAP7_75t_L g1185 ( 
.A(n_1026),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_989),
.A2(n_661),
.B(n_657),
.Y(n_1186)
);

INVx4_ASAP7_75t_L g1187 ( 
.A(n_990),
.Y(n_1187)
);

CKINVDCx10_ASAP7_75t_R g1188 ( 
.A(n_1112),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1110),
.B(n_619),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1129),
.B(n_620),
.Y(n_1190)
);

OAI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1000),
.A2(n_668),
.B(n_664),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1049),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1002),
.A2(n_1100),
.B(n_1103),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_983),
.A2(n_670),
.B(n_676),
.C(n_669),
.Y(n_1194)
);

INVx11_ASAP7_75t_L g1195 ( 
.A(n_1094),
.Y(n_1195)
);

INVxp67_ASAP7_75t_L g1196 ( 
.A(n_1134),
.Y(n_1196)
);

INVx1_ASAP7_75t_SL g1197 ( 
.A(n_1021),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_980),
.B(n_626),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_984),
.B(n_697),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_1136),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1083),
.B(n_630),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_998),
.B(n_631),
.Y(n_1202)
);

BUFx4f_ASAP7_75t_L g1203 ( 
.A(n_1094),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1098),
.A2(n_942),
.B(n_938),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_1094),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_988),
.A2(n_715),
.B1(n_724),
.B2(n_710),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_990),
.B(n_633),
.Y(n_1207)
);

INVxp67_ASAP7_75t_L g1208 ( 
.A(n_1006),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_1029),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1108),
.A2(n_985),
.B1(n_1052),
.B2(n_1050),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1053),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1114),
.A2(n_687),
.B(n_678),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1016),
.A2(n_645),
.B1(n_646),
.B2(n_635),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1102),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1119),
.A2(n_701),
.B(n_691),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_SL g1216 ( 
.A(n_990),
.B(n_652),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1054),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1016),
.A2(n_658),
.B1(n_665),
.B2(n_653),
.Y(n_1218)
);

AO21x1_ASAP7_75t_L g1219 ( 
.A1(n_1125),
.A2(n_712),
.B(n_711),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_987),
.B(n_667),
.Y(n_1220)
);

AO21x1_ASAP7_75t_L g1221 ( 
.A1(n_1058),
.A2(n_745),
.B(n_743),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1035),
.B(n_715),
.Y(n_1222)
);

AND2x2_ASAP7_75t_SL g1223 ( 
.A(n_1113),
.B(n_724),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1056),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_1136),
.B(n_671),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1087),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_1001),
.B(n_693),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_1048),
.Y(n_1228)
);

CKINVDCx6p67_ASAP7_75t_R g1229 ( 
.A(n_1071),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1127),
.A2(n_953),
.B(n_949),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1033),
.B(n_699),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1034),
.B(n_720),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_1116),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1028),
.B(n_730),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1059),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1075),
.Y(n_1236)
);

NAND3xp33_ASAP7_75t_L g1237 ( 
.A(n_1068),
.B(n_1041),
.C(n_1081),
.Y(n_1237)
);

BUFx4f_ASAP7_75t_L g1238 ( 
.A(n_1001),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1118),
.B(n_562),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1085),
.B(n_562),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1061),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1050),
.A2(n_588),
.B1(n_703),
.B2(n_575),
.Y(n_1242)
);

NAND2xp33_ASAP7_75t_L g1243 ( 
.A(n_1029),
.B(n_575),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1128),
.A2(n_966),
.B(n_965),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1018),
.B(n_575),
.Y(n_1245)
);

OR2x6_ASAP7_75t_L g1246 ( 
.A(n_1039),
.B(n_588),
.Y(n_1246)
);

AOI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1111),
.A2(n_977),
.B(n_973),
.Y(n_1247)
);

INVx4_ASAP7_75t_L g1248 ( 
.A(n_1137),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1131),
.Y(n_1249)
);

AOI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1052),
.A2(n_979),
.B(n_978),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1131),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1078),
.B(n_721),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1004),
.A2(n_1005),
.B(n_1017),
.Y(n_1253)
);

NOR2x1p5_ASAP7_75t_L g1254 ( 
.A(n_1015),
.B(n_737),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1064),
.B(n_1077),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1090),
.B(n_737),
.Y(n_1256)
);

AO21x1_ASAP7_75t_L g1257 ( 
.A1(n_1065),
.A2(n_835),
.B(n_820),
.Y(n_1257)
);

O2A1O1Ixp5_ASAP7_75t_L g1258 ( 
.A1(n_1074),
.A2(n_835),
.B(n_741),
.C(n_324),
.Y(n_1258)
);

O2A1O1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1109),
.A2(n_32),
.B(n_30),
.C(n_31),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1072),
.B(n_32),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1124),
.A2(n_1066),
.B1(n_1091),
.B2(n_1057),
.Y(n_1261)
);

INVxp67_ASAP7_75t_L g1262 ( 
.A(n_1022),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_993),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_996),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1073),
.B(n_33),
.Y(n_1265)
);

INVx3_ASAP7_75t_L g1266 ( 
.A(n_1137),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1038),
.A2(n_330),
.B(n_329),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1088),
.B(n_34),
.Y(n_1268)
);

BUFx8_ASAP7_75t_SL g1269 ( 
.A(n_1095),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1044),
.B(n_35),
.Y(n_1270)
);

INVx6_ASAP7_75t_L g1271 ( 
.A(n_1145),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1067),
.B(n_36),
.Y(n_1272)
);

INVxp67_ASAP7_75t_L g1273 ( 
.A(n_1082),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1084),
.B(n_38),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1093),
.B(n_38),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1092),
.B(n_40),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_SL g1277 ( 
.A(n_1149),
.B(n_1099),
.Y(n_1277)
);

BUFx12f_ASAP7_75t_L g1278 ( 
.A(n_1123),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1013),
.Y(n_1279)
);

O2A1O1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_1062),
.A2(n_45),
.B(n_42),
.C(n_44),
.Y(n_1280)
);

OAI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1086),
.A2(n_333),
.B(n_332),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1069),
.B(n_47),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1063),
.A2(n_53),
.B1(n_48),
.B2(n_52),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1132),
.Y(n_1284)
);

NAND3xp33_ASAP7_75t_SL g1285 ( 
.A(n_1139),
.B(n_48),
.C(n_54),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1079),
.B(n_54),
.Y(n_1286)
);

CKINVDCx11_ASAP7_75t_R g1287 ( 
.A(n_995),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1060),
.A2(n_339),
.B(n_338),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1101),
.B(n_57),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1138),
.Y(n_1290)
);

OR2x6_ASAP7_75t_L g1291 ( 
.A(n_986),
.B(n_57),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1132),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1133),
.Y(n_1293)
);

INVx2_ASAP7_75t_SL g1294 ( 
.A(n_1010),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1023),
.A2(n_1025),
.B(n_1055),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1027),
.Y(n_1296)
);

AO21x1_ASAP7_75t_L g1297 ( 
.A1(n_1124),
.A2(n_59),
.B(n_60),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1133),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1135),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_1155),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1046),
.B(n_63),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_991),
.B(n_63),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1089),
.B(n_64),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1115),
.A2(n_351),
.B(n_348),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1135),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1117),
.B(n_65),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1024),
.B(n_66),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1120),
.A2(n_353),
.B(n_352),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1121),
.B(n_1122),
.Y(n_1309)
);

INVx5_ASAP7_75t_L g1310 ( 
.A(n_1008),
.Y(n_1310)
);

OAI321xp33_ASAP7_75t_L g1311 ( 
.A1(n_1144),
.A2(n_67),
.A3(n_68),
.B1(n_70),
.B2(n_72),
.C(n_73),
.Y(n_1311)
);

BUFx4f_ASAP7_75t_L g1312 ( 
.A(n_1011),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1105),
.B(n_1097),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1150),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_1314)
);

INVx11_ASAP7_75t_L g1315 ( 
.A(n_1030),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1043),
.B(n_75),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1009),
.B(n_1014),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1031),
.A2(n_362),
.B(n_361),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1104),
.B(n_76),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1106),
.B(n_79),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1140),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1036),
.A2(n_367),
.B(n_364),
.Y(n_1322)
);

AND2x4_ASAP7_75t_L g1323 ( 
.A(n_1107),
.B(n_79),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1040),
.B(n_80),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1140),
.Y(n_1325)
);

AND2x4_ASAP7_75t_SL g1326 ( 
.A(n_1153),
.B(n_81),
.Y(n_1326)
);

INVxp67_ASAP7_75t_L g1327 ( 
.A(n_1141),
.Y(n_1327)
);

CKINVDCx10_ASAP7_75t_R g1328 ( 
.A(n_1149),
.Y(n_1328)
);

INVx4_ASAP7_75t_L g1329 ( 
.A(n_1155),
.Y(n_1329)
);

O2A1O1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1150),
.A2(n_86),
.B(n_83),
.C(n_85),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1142),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1148),
.A2(n_373),
.B(n_371),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1151),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1151),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1159),
.B(n_1158),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1154),
.A2(n_378),
.B(n_377),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_1155),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_SL g1338 ( 
.A(n_1158),
.B(n_379),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1154),
.B(n_88),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1156),
.B(n_91),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1146),
.Y(n_1341)
);

A2O1A1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1156),
.A2(n_93),
.B(n_91),
.C(n_92),
.Y(n_1342)
);

O2A1O1Ixp33_ASAP7_75t_L g1343 ( 
.A1(n_1146),
.A2(n_94),
.B(n_92),
.C(n_93),
.Y(n_1343)
);

INVx1_ASAP7_75t_SL g1344 ( 
.A(n_1130),
.Y(n_1344)
);

OAI21xp33_ASAP7_75t_L g1345 ( 
.A1(n_1157),
.A2(n_96),
.B(n_101),
.Y(n_1345)
);

AOI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1143),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1147),
.A2(n_1152),
.B1(n_107),
.B2(n_105),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1012),
.B(n_106),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1003),
.B(n_107),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1045),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1182),
.B(n_108),
.Y(n_1351)
);

INVx5_ASAP7_75t_L g1352 ( 
.A(n_1248),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1333),
.Y(n_1353)
);

OAI21xp33_ASAP7_75t_SL g1354 ( 
.A1(n_1212),
.A2(n_109),
.B(n_110),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1253),
.A2(n_109),
.B(n_111),
.Y(n_1355)
);

A2O1A1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1295),
.A2(n_114),
.B(n_111),
.C(n_112),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1193),
.A2(n_395),
.B(n_393),
.Y(n_1357)
);

A2O1A1Ixp33_ASAP7_75t_L g1358 ( 
.A1(n_1260),
.A2(n_117),
.B(n_114),
.C(n_115),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1249),
.B(n_115),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1251),
.B(n_117),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1321),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1210),
.B(n_118),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1210),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1199),
.B(n_120),
.Y(n_1364)
);

AND2x2_ASAP7_75t_SL g1365 ( 
.A(n_1203),
.B(n_121),
.Y(n_1365)
);

A2O1A1Ixp33_ASAP7_75t_L g1366 ( 
.A1(n_1170),
.A2(n_1302),
.B(n_1272),
.C(n_1309),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_1188),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1208),
.B(n_123),
.Y(n_1368)
);

NOR2xp67_ASAP7_75t_L g1369 ( 
.A(n_1183),
.B(n_124),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1331),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1165),
.B(n_124),
.Y(n_1371)
);

AO22x1_ASAP7_75t_L g1372 ( 
.A1(n_1165),
.A2(n_1167),
.B1(n_1175),
.B2(n_1166),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1174),
.B(n_1194),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1167),
.B(n_1171),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1212),
.B(n_125),
.Y(n_1375)
);

INVx5_ASAP7_75t_L g1376 ( 
.A(n_1248),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1263),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1300),
.Y(n_1378)
);

AOI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1169),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_SL g1380 ( 
.A(n_1203),
.B(n_126),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1200),
.B(n_129),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1296),
.B(n_131),
.Y(n_1382)
);

BUFx4f_ASAP7_75t_L g1383 ( 
.A(n_1246),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1191),
.B(n_132),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1184),
.B(n_132),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_SL g1386 ( 
.A1(n_1281),
.A2(n_133),
.B(n_134),
.Y(n_1386)
);

AOI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1173),
.A2(n_1222),
.B1(n_1185),
.B2(n_1273),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1334),
.B(n_1341),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1334),
.B(n_133),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1215),
.A2(n_1239),
.B(n_1261),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1264),
.Y(n_1391)
);

OAI22x1_ASAP7_75t_L g1392 ( 
.A1(n_1225),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_1392)
);

NAND2x1p5_ASAP7_75t_L g1393 ( 
.A(n_1177),
.B(n_136),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1279),
.Y(n_1394)
);

BUFx2_ASAP7_75t_L g1395 ( 
.A(n_1178),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1348),
.Y(n_1396)
);

BUFx6f_ASAP7_75t_L g1397 ( 
.A(n_1337),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1228),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1223),
.B(n_137),
.Y(n_1399)
);

NAND3xp33_ASAP7_75t_L g1400 ( 
.A(n_1237),
.B(n_138),
.C(n_139),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1160),
.B(n_139),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1262),
.B(n_141),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1161),
.B(n_141),
.Y(n_1403)
);

NAND3x1_ASAP7_75t_L g1404 ( 
.A(n_1286),
.B(n_142),
.C(n_143),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1197),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_1405)
);

INVx5_ASAP7_75t_L g1406 ( 
.A(n_1172),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_1337),
.Y(n_1407)
);

AOI21xp33_ASAP7_75t_L g1408 ( 
.A1(n_1242),
.A2(n_145),
.B(n_146),
.Y(n_1408)
);

AO31x2_ASAP7_75t_L g1409 ( 
.A1(n_1221),
.A2(n_146),
.A3(n_147),
.B(n_148),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1215),
.A2(n_147),
.B(n_148),
.Y(n_1410)
);

INVx4_ASAP7_75t_L g1411 ( 
.A(n_1195),
.Y(n_1411)
);

NAND3xp33_ASAP7_75t_SL g1412 ( 
.A(n_1283),
.B(n_149),
.C(n_150),
.Y(n_1412)
);

A2O1A1Ixp33_ASAP7_75t_L g1413 ( 
.A1(n_1349),
.A2(n_151),
.B(n_152),
.C(n_153),
.Y(n_1413)
);

INVx4_ASAP7_75t_SL g1414 ( 
.A(n_1172),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1261),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1163),
.B(n_157),
.Y(n_1416)
);

INVx6_ASAP7_75t_L g1417 ( 
.A(n_1350),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1233),
.Y(n_1418)
);

AO21x2_ASAP7_75t_L g1419 ( 
.A1(n_1176),
.A2(n_158),
.B(n_159),
.Y(n_1419)
);

OAI21xp33_ASAP7_75t_SL g1420 ( 
.A1(n_1246),
.A2(n_158),
.B(n_160),
.Y(n_1420)
);

A2O1A1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1259),
.A2(n_162),
.B(n_163),
.C(n_165),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_SL g1422 ( 
.A(n_1277),
.B(n_163),
.Y(n_1422)
);

CKINVDCx14_ASAP7_75t_R g1423 ( 
.A(n_1287),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1206),
.B(n_167),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1213),
.B(n_168),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1179),
.B(n_168),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1181),
.B(n_169),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1218),
.B(n_169),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1335),
.A2(n_172),
.B(n_173),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1192),
.B(n_174),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1339),
.A2(n_1303),
.B1(n_1327),
.B2(n_1268),
.Y(n_1431)
);

INVx3_ASAP7_75t_L g1432 ( 
.A(n_1266),
.Y(n_1432)
);

AO31x2_ASAP7_75t_L g1433 ( 
.A1(n_1297),
.A2(n_178),
.A3(n_179),
.B(n_180),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1211),
.B(n_180),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1217),
.B(n_181),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1224),
.B(n_182),
.Y(n_1436)
);

NAND3xp33_ASAP7_75t_SL g1437 ( 
.A(n_1219),
.B(n_182),
.C(n_183),
.Y(n_1437)
);

AOI221x1_ASAP7_75t_L g1438 ( 
.A1(n_1345),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.C(n_187),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1205),
.B(n_186),
.Y(n_1439)
);

INVx3_ASAP7_75t_L g1440 ( 
.A(n_1266),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1292),
.A2(n_195),
.B(n_197),
.Y(n_1441)
);

NOR2x1_ASAP7_75t_SL g1442 ( 
.A(n_1246),
.B(n_198),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1204),
.A2(n_200),
.B(n_201),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1235),
.B(n_201),
.Y(n_1444)
);

AOI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1274),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1317),
.A2(n_207),
.B(n_208),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1226),
.B(n_209),
.Y(n_1447)
);

CKINVDCx11_ASAP7_75t_R g1448 ( 
.A(n_1278),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1202),
.B(n_210),
.Y(n_1449)
);

AOI21xp33_ASAP7_75t_L g1450 ( 
.A1(n_1324),
.A2(n_212),
.B(n_213),
.Y(n_1450)
);

AO21x2_ASAP7_75t_L g1451 ( 
.A1(n_1162),
.A2(n_214),
.B(n_215),
.Y(n_1451)
);

AOI221x1_ASAP7_75t_L g1452 ( 
.A1(n_1162),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.C(n_221),
.Y(n_1452)
);

AO31x2_ASAP7_75t_L g1453 ( 
.A1(n_1240),
.A2(n_218),
.A3(n_222),
.B(n_223),
.Y(n_1453)
);

OAI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1293),
.A2(n_223),
.B(n_224),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1339),
.A2(n_225),
.B1(n_228),
.B2(n_229),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_1328),
.Y(n_1456)
);

A2O1A1Ixp33_ASAP7_75t_L g1457 ( 
.A1(n_1307),
.A2(n_225),
.B(n_228),
.C(n_229),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1241),
.B(n_230),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1256),
.A2(n_1313),
.B(n_1230),
.Y(n_1459)
);

INVx6_ASAP7_75t_L g1460 ( 
.A(n_1271),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1298),
.B(n_232),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1284),
.Y(n_1462)
);

A2O1A1Ixp33_ASAP7_75t_L g1463 ( 
.A1(n_1280),
.A2(n_232),
.B(n_233),
.C(n_234),
.Y(n_1463)
);

OAI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1299),
.A2(n_233),
.B(n_234),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1319),
.Y(n_1465)
);

BUFx12f_ASAP7_75t_L g1466 ( 
.A(n_1271),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1229),
.B(n_235),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1238),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1305),
.B(n_238),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1320),
.Y(n_1470)
);

BUFx2_ASAP7_75t_L g1471 ( 
.A(n_1291),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1325),
.B(n_239),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1198),
.B(n_241),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1320),
.Y(n_1474)
);

AO31x2_ASAP7_75t_L g1475 ( 
.A1(n_1342),
.A2(n_1314),
.A3(n_1322),
.B(n_1308),
.Y(n_1475)
);

AO31x2_ASAP7_75t_L g1476 ( 
.A1(n_1314),
.A2(n_241),
.A3(n_242),
.B(n_243),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1265),
.B(n_244),
.Y(n_1477)
);

A2O1A1Ixp33_ASAP7_75t_L g1478 ( 
.A1(n_1276),
.A2(n_246),
.B(n_248),
.C(n_249),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1238),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_1209),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1323),
.Y(n_1481)
);

BUFx6f_ASAP7_75t_L g1482 ( 
.A(n_1290),
.Y(n_1482)
);

OR2x6_ASAP7_75t_L g1483 ( 
.A(n_1291),
.B(n_308),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1301),
.B(n_256),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1340),
.B(n_257),
.Y(n_1485)
);

INVx6_ASAP7_75t_L g1486 ( 
.A(n_1291),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1270),
.B(n_258),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1275),
.B(n_260),
.Y(n_1488)
);

AO31x2_ASAP7_75t_L g1489 ( 
.A1(n_1304),
.A2(n_263),
.A3(n_264),
.B(n_265),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1168),
.B(n_265),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1189),
.B(n_266),
.Y(n_1491)
);

AO31x2_ASAP7_75t_L g1492 ( 
.A1(n_1267),
.A2(n_267),
.A3(n_268),
.B(n_269),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1231),
.B(n_270),
.Y(n_1493)
);

A2O1A1Ixp33_ASAP7_75t_L g1494 ( 
.A1(n_1330),
.A2(n_272),
.B(n_273),
.C(n_274),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1289),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1323),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_1269),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1232),
.B(n_1282),
.Y(n_1498)
);

NAND2x1p5_ASAP7_75t_L g1499 ( 
.A(n_1187),
.B(n_276),
.Y(n_1499)
);

A2O1A1Ixp33_ASAP7_75t_L g1500 ( 
.A1(n_1306),
.A2(n_279),
.B(n_280),
.C(n_281),
.Y(n_1500)
);

BUFx6f_ASAP7_75t_L g1501 ( 
.A(n_1290),
.Y(n_1501)
);

OR2x6_ASAP7_75t_L g1502 ( 
.A(n_1236),
.B(n_308),
.Y(n_1502)
);

AOI21xp33_ASAP7_75t_L g1503 ( 
.A1(n_1316),
.A2(n_283),
.B(n_284),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1190),
.B(n_286),
.Y(n_1504)
);

INVx1_ASAP7_75t_SL g1505 ( 
.A(n_1214),
.Y(n_1505)
);

OAI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1258),
.A2(n_287),
.B(n_288),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1180),
.A2(n_287),
.B1(n_289),
.B2(n_290),
.Y(n_1507)
);

BUFx6f_ASAP7_75t_L g1508 ( 
.A(n_1290),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_1315),
.Y(n_1509)
);

OAI21xp33_ASAP7_75t_L g1510 ( 
.A1(n_1220),
.A2(n_1234),
.B(n_1201),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1187),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1294),
.B(n_294),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1255),
.B(n_295),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1196),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1326),
.B(n_299),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_SL g1516 ( 
.A(n_1312),
.B(n_301),
.Y(n_1516)
);

OAI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1288),
.A2(n_302),
.B(n_303),
.Y(n_1517)
);

OAI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1336),
.A2(n_302),
.B(n_303),
.Y(n_1518)
);

AOI221xp5_ASAP7_75t_L g1519 ( 
.A1(n_1252),
.A2(n_304),
.B1(n_305),
.B2(n_307),
.C(n_1285),
.Y(n_1519)
);

BUFx6f_ASAP7_75t_L g1520 ( 
.A(n_1329),
.Y(n_1520)
);

OAI22x1_ASAP7_75t_L g1521 ( 
.A1(n_1254),
.A2(n_1346),
.B1(n_1164),
.B2(n_1207),
.Y(n_1521)
);

OAI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1318),
.A2(n_1332),
.B(n_1343),
.Y(n_1522)
);

AOI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1216),
.A2(n_1227),
.B(n_1338),
.Y(n_1523)
);

OAI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1245),
.A2(n_1311),
.B(n_1243),
.Y(n_1524)
);

AO31x2_ASAP7_75t_L g1525 ( 
.A1(n_1347),
.A2(n_1311),
.A3(n_1310),
.B(n_1344),
.Y(n_1525)
);

OAI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1182),
.A2(n_1253),
.B(n_1126),
.Y(n_1526)
);

AO31x2_ASAP7_75t_L g1527 ( 
.A1(n_1257),
.A2(n_1242),
.A3(n_1210),
.B(n_1126),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1250),
.A2(n_1247),
.B(n_1244),
.Y(n_1528)
);

AOI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1182),
.A2(n_989),
.B(n_992),
.Y(n_1529)
);

OAI21x1_ASAP7_75t_L g1530 ( 
.A1(n_1250),
.A2(n_1247),
.B(n_1244),
.Y(n_1530)
);

CKINVDCx20_ASAP7_75t_R g1531 ( 
.A(n_1287),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1182),
.B(n_1012),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1182),
.B(n_1012),
.Y(n_1533)
);

OAI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1250),
.A2(n_1247),
.B(n_1244),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1208),
.B(n_1012),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1182),
.A2(n_989),
.B(n_992),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1182),
.A2(n_1210),
.B1(n_1191),
.B2(n_1212),
.Y(n_1537)
);

AOI21xp5_ASAP7_75t_L g1538 ( 
.A1(n_1182),
.A2(n_989),
.B(n_992),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_SL g1539 ( 
.A(n_1203),
.B(n_847),
.Y(n_1539)
);

AOI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_1182),
.A2(n_989),
.B(n_992),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_SL g1541 ( 
.A(n_1203),
.B(n_847),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1208),
.B(n_1012),
.Y(n_1542)
);

BUFx12f_ASAP7_75t_L g1543 ( 
.A(n_1287),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1182),
.A2(n_989),
.B(n_992),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1182),
.B(n_1012),
.Y(n_1545)
);

AOI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1182),
.A2(n_989),
.B(n_992),
.Y(n_1546)
);

AOI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1182),
.A2(n_989),
.B(n_992),
.Y(n_1547)
);

NOR2x1_ASAP7_75t_SL g1548 ( 
.A(n_1246),
.B(n_1248),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1182),
.B(n_1012),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1182),
.A2(n_989),
.B(n_992),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1182),
.B(n_1012),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1182),
.B(n_1012),
.Y(n_1552)
);

OAI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1182),
.A2(n_1253),
.B(n_1126),
.Y(n_1553)
);

OAI22x1_ASAP7_75t_L g1554 ( 
.A1(n_1200),
.A2(n_892),
.B1(n_1019),
.B2(n_877),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1333),
.Y(n_1555)
);

AOI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1182),
.A2(n_989),
.B(n_992),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1182),
.B(n_1012),
.Y(n_1557)
);

O2A1O1Ixp5_ASAP7_75t_L g1558 ( 
.A1(n_1186),
.A2(n_1257),
.B(n_1176),
.C(n_1221),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1182),
.B(n_1012),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1182),
.B(n_1012),
.Y(n_1560)
);

OA22x2_ASAP7_75t_L g1561 ( 
.A1(n_1200),
.A2(n_1019),
.B1(n_892),
.B2(n_1026),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1182),
.B(n_1012),
.Y(n_1562)
);

A2O1A1Ixp33_ASAP7_75t_L g1563 ( 
.A1(n_1295),
.A2(n_1003),
.B(n_1260),
.C(n_1170),
.Y(n_1563)
);

AO31x2_ASAP7_75t_L g1564 ( 
.A1(n_1257),
.A2(n_1242),
.A3(n_1210),
.B(n_1126),
.Y(n_1564)
);

NAND3xp33_ASAP7_75t_L g1565 ( 
.A(n_1199),
.B(n_1186),
.C(n_1302),
.Y(n_1565)
);

AOI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1166),
.A2(n_1026),
.B1(n_1169),
.B2(n_846),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1199),
.B(n_1032),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1182),
.B(n_1012),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_L g1569 ( 
.A(n_1199),
.B(n_1032),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1333),
.Y(n_1570)
);

HB1xp67_ASAP7_75t_L g1571 ( 
.A(n_1173),
.Y(n_1571)
);

OAI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1182),
.A2(n_1253),
.B(n_1126),
.Y(n_1572)
);

BUFx12f_ASAP7_75t_L g1573 ( 
.A(n_1287),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1182),
.B(n_1012),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1321),
.Y(n_1575)
);

INVx4_ASAP7_75t_L g1576 ( 
.A(n_1195),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_1173),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1199),
.B(n_1032),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1208),
.B(n_1012),
.Y(n_1579)
);

BUFx2_ASAP7_75t_SL g1580 ( 
.A(n_1178),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1208),
.B(n_1012),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1333),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1182),
.B(n_1012),
.Y(n_1583)
);

OAI22x1_ASAP7_75t_L g1584 ( 
.A1(n_1200),
.A2(n_892),
.B1(n_1019),
.B2(n_877),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1182),
.B(n_1012),
.Y(n_1585)
);

BUFx2_ASAP7_75t_L g1586 ( 
.A(n_1173),
.Y(n_1586)
);

AO31x2_ASAP7_75t_L g1587 ( 
.A1(n_1257),
.A2(n_1242),
.A3(n_1210),
.B(n_1126),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1182),
.B(n_1012),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1182),
.A2(n_989),
.B(n_992),
.Y(n_1589)
);

BUFx2_ASAP7_75t_L g1590 ( 
.A(n_1173),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1387),
.B(n_1374),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_1586),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1388),
.Y(n_1593)
);

OAI21x1_ASAP7_75t_SL g1594 ( 
.A1(n_1548),
.A2(n_1442),
.B(n_1386),
.Y(n_1594)
);

BUFx3_ASAP7_75t_L g1595 ( 
.A(n_1352),
.Y(n_1595)
);

OR2x6_ASAP7_75t_L g1596 ( 
.A(n_1483),
.B(n_1486),
.Y(n_1596)
);

AOI22x1_ASAP7_75t_L g1597 ( 
.A1(n_1521),
.A2(n_1523),
.B1(n_1357),
.B2(n_1506),
.Y(n_1597)
);

AO21x2_ASAP7_75t_L g1598 ( 
.A1(n_1390),
.A2(n_1506),
.B(n_1362),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1462),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1353),
.Y(n_1600)
);

BUFx3_ASAP7_75t_L g1601 ( 
.A(n_1352),
.Y(n_1601)
);

OAI21x1_ASAP7_75t_L g1602 ( 
.A1(n_1526),
.A2(n_1572),
.B(n_1553),
.Y(n_1602)
);

BUFx2_ASAP7_75t_SL g1603 ( 
.A(n_1531),
.Y(n_1603)
);

AO21x2_ASAP7_75t_L g1604 ( 
.A1(n_1522),
.A2(n_1537),
.B(n_1518),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1532),
.B(n_1533),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1352),
.B(n_1376),
.Y(n_1606)
);

OAI21x1_ASAP7_75t_L g1607 ( 
.A1(n_1529),
.A2(n_1538),
.B(n_1536),
.Y(n_1607)
);

BUFx3_ASAP7_75t_L g1608 ( 
.A(n_1352),
.Y(n_1608)
);

OAI21x1_ASAP7_75t_L g1609 ( 
.A1(n_1540),
.A2(n_1546),
.B(n_1544),
.Y(n_1609)
);

BUFx2_ASAP7_75t_L g1610 ( 
.A(n_1590),
.Y(n_1610)
);

AO21x2_ASAP7_75t_L g1611 ( 
.A1(n_1537),
.A2(n_1518),
.B(n_1517),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1555),
.Y(n_1612)
);

OAI21x1_ASAP7_75t_L g1613 ( 
.A1(n_1547),
.A2(n_1556),
.B(n_1550),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1570),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1532),
.B(n_1533),
.Y(n_1615)
);

INVx6_ASAP7_75t_L g1616 ( 
.A(n_1376),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1577),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1456),
.Y(n_1618)
);

INVx3_ASAP7_75t_L g1619 ( 
.A(n_1376),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1577),
.B(n_1545),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1545),
.A2(n_1549),
.B1(n_1557),
.B2(n_1551),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1549),
.B(n_1551),
.Y(n_1622)
);

AO21x2_ASAP7_75t_L g1623 ( 
.A1(n_1517),
.A2(n_1355),
.B(n_1589),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1582),
.Y(n_1624)
);

OR2x6_ASAP7_75t_L g1625 ( 
.A(n_1483),
.B(n_1486),
.Y(n_1625)
);

INVx3_ASAP7_75t_L g1626 ( 
.A(n_1376),
.Y(n_1626)
);

INVx2_ASAP7_75t_SL g1627 ( 
.A(n_1383),
.Y(n_1627)
);

INVx3_ASAP7_75t_SL g1628 ( 
.A(n_1411),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1557),
.B(n_1560),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1377),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_1406),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_1367),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1391),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1561),
.A2(n_1483),
.B1(n_1424),
.B2(n_1365),
.Y(n_1634)
);

AO21x2_ASAP7_75t_L g1635 ( 
.A1(n_1355),
.A2(n_1524),
.B(n_1410),
.Y(n_1635)
);

BUFx2_ASAP7_75t_L g1636 ( 
.A(n_1571),
.Y(n_1636)
);

CKINVDCx11_ASAP7_75t_R g1637 ( 
.A(n_1543),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1431),
.A2(n_1562),
.B(n_1560),
.Y(n_1638)
);

OR2x6_ASAP7_75t_L g1639 ( 
.A(n_1502),
.B(n_1562),
.Y(n_1639)
);

OAI21x1_ASAP7_75t_SL g1640 ( 
.A1(n_1410),
.A2(n_1454),
.B(n_1441),
.Y(n_1640)
);

INVx2_ASAP7_75t_SL g1641 ( 
.A(n_1383),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1394),
.Y(n_1642)
);

INVx8_ASAP7_75t_L g1643 ( 
.A(n_1406),
.Y(n_1643)
);

BUFx3_ASAP7_75t_L g1644 ( 
.A(n_1406),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1361),
.Y(n_1645)
);

AO21x1_ASAP7_75t_L g1646 ( 
.A1(n_1415),
.A2(n_1363),
.B(n_1393),
.Y(n_1646)
);

OAI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1565),
.A2(n_1498),
.B(n_1568),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1568),
.B(n_1574),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1401),
.Y(n_1649)
);

AOI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1567),
.A2(n_1578),
.B1(n_1569),
.B2(n_1574),
.Y(n_1650)
);

OA21x2_ASAP7_75t_L g1651 ( 
.A1(n_1438),
.A2(n_1452),
.B(n_1441),
.Y(n_1651)
);

BUFx2_ASAP7_75t_SL g1652 ( 
.A(n_1411),
.Y(n_1652)
);

AO21x2_ASAP7_75t_L g1653 ( 
.A1(n_1454),
.A2(n_1464),
.B(n_1451),
.Y(n_1653)
);

INVx6_ASAP7_75t_L g1654 ( 
.A(n_1576),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1401),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1416),
.Y(n_1656)
);

AOI22xp33_ASAP7_75t_L g1657 ( 
.A1(n_1561),
.A2(n_1585),
.B1(n_1588),
.B2(n_1583),
.Y(n_1657)
);

BUFx3_ASAP7_75t_L g1658 ( 
.A(n_1406),
.Y(n_1658)
);

INVx2_ASAP7_75t_SL g1659 ( 
.A(n_1417),
.Y(n_1659)
);

NOR2xp67_ASAP7_75t_SL g1660 ( 
.A(n_1573),
.B(n_1576),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1583),
.B(n_1585),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1416),
.Y(n_1662)
);

AND2x6_ASAP7_75t_L g1663 ( 
.A(n_1482),
.B(n_1501),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1426),
.Y(n_1664)
);

INVx3_ASAP7_75t_L g1665 ( 
.A(n_1482),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1588),
.B(n_1552),
.Y(n_1666)
);

BUFx8_ASAP7_75t_SL g1667 ( 
.A(n_1497),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1559),
.B(n_1372),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1426),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1535),
.B(n_1542),
.Y(n_1670)
);

INVx1_ASAP7_75t_SL g1671 ( 
.A(n_1580),
.Y(n_1671)
);

INVx4_ASAP7_75t_L g1672 ( 
.A(n_1414),
.Y(n_1672)
);

OAI21x1_ASAP7_75t_L g1673 ( 
.A1(n_1351),
.A2(n_1389),
.B(n_1443),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1427),
.Y(n_1674)
);

INVx3_ASAP7_75t_L g1675 ( 
.A(n_1482),
.Y(n_1675)
);

INVx3_ASAP7_75t_SL g1676 ( 
.A(n_1509),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1430),
.Y(n_1677)
);

OAI21x1_ASAP7_75t_L g1678 ( 
.A1(n_1434),
.A2(n_1436),
.B(n_1435),
.Y(n_1678)
);

INVx3_ASAP7_75t_L g1679 ( 
.A(n_1501),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1566),
.B(n_1465),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1439),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1579),
.B(n_1581),
.Y(n_1682)
);

OAI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1498),
.A2(n_1510),
.B(n_1493),
.Y(n_1683)
);

OAI21x1_ASAP7_75t_L g1684 ( 
.A1(n_1444),
.A2(n_1458),
.B(n_1488),
.Y(n_1684)
);

AO31x2_ASAP7_75t_L g1685 ( 
.A1(n_1415),
.A2(n_1363),
.A3(n_1494),
.B(n_1356),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1370),
.Y(n_1686)
);

BUFx2_ASAP7_75t_L g1687 ( 
.A(n_1395),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1359),
.Y(n_1688)
);

BUFx2_ASAP7_75t_SL g1689 ( 
.A(n_1468),
.Y(n_1689)
);

BUFx3_ASAP7_75t_L g1690 ( 
.A(n_1417),
.Y(n_1690)
);

INVx6_ASAP7_75t_L g1691 ( 
.A(n_1511),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1359),
.Y(n_1692)
);

OA21x2_ASAP7_75t_L g1693 ( 
.A1(n_1408),
.A2(n_1463),
.B(n_1384),
.Y(n_1693)
);

BUFx3_ASAP7_75t_L g1694 ( 
.A(n_1501),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1470),
.B(n_1474),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1360),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1360),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1371),
.A2(n_1373),
.B1(n_1364),
.B2(n_1369),
.Y(n_1698)
);

OAI21x1_ASAP7_75t_L g1699 ( 
.A1(n_1499),
.A2(n_1469),
.B(n_1461),
.Y(n_1699)
);

OAI21x1_ASAP7_75t_L g1700 ( 
.A1(n_1499),
.A2(n_1469),
.B(n_1461),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1439),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1472),
.Y(n_1702)
);

NAND3xp33_ASAP7_75t_L g1703 ( 
.A(n_1400),
.B(n_1519),
.C(n_1420),
.Y(n_1703)
);

NOR2xp33_ASAP7_75t_L g1704 ( 
.A(n_1481),
.B(n_1496),
.Y(n_1704)
);

AOI22x1_ASAP7_75t_L g1705 ( 
.A1(n_1446),
.A2(n_1429),
.B1(n_1392),
.B2(n_1473),
.Y(n_1705)
);

BUFx3_ASAP7_75t_L g1706 ( 
.A(n_1508),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1554),
.B(n_1584),
.Y(n_1707)
);

AO21x2_ASAP7_75t_L g1708 ( 
.A1(n_1375),
.A2(n_1419),
.B(n_1484),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1396),
.B(n_1385),
.Y(n_1709)
);

AO21x2_ASAP7_75t_L g1710 ( 
.A1(n_1437),
.A2(n_1477),
.B(n_1485),
.Y(n_1710)
);

AND2x6_ASAP7_75t_L g1711 ( 
.A(n_1508),
.B(n_1378),
.Y(n_1711)
);

AO21x2_ASAP7_75t_L g1712 ( 
.A1(n_1477),
.A2(n_1421),
.B(n_1412),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1512),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1398),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1381),
.B(n_1425),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1512),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1382),
.Y(n_1717)
);

INVxp67_ASAP7_75t_L g1718 ( 
.A(n_1502),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1382),
.Y(n_1719)
);

INVx6_ASAP7_75t_L g1720 ( 
.A(n_1511),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1502),
.Y(n_1721)
);

AO31x2_ASAP7_75t_L g1722 ( 
.A1(n_1455),
.A2(n_1495),
.A3(n_1500),
.B(n_1413),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1432),
.B(n_1440),
.Y(n_1723)
);

OAI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1487),
.A2(n_1504),
.B(n_1491),
.Y(n_1724)
);

BUFx4_ASAP7_75t_SL g1725 ( 
.A(n_1418),
.Y(n_1725)
);

NAND2x1p5_ASAP7_75t_L g1726 ( 
.A(n_1479),
.B(n_1508),
.Y(n_1726)
);

OAI21x1_ASAP7_75t_SL g1727 ( 
.A1(n_1405),
.A2(n_1495),
.B(n_1490),
.Y(n_1727)
);

AND2x4_ASAP7_75t_L g1728 ( 
.A(n_1575),
.B(n_1414),
.Y(n_1728)
);

BUFx3_ASAP7_75t_L g1729 ( 
.A(n_1520),
.Y(n_1729)
);

OA21x2_ASAP7_75t_L g1730 ( 
.A1(n_1503),
.A2(n_1450),
.B(n_1358),
.Y(n_1730)
);

AO21x2_ASAP7_75t_L g1731 ( 
.A1(n_1503),
.A2(n_1450),
.B(n_1457),
.Y(n_1731)
);

OAI21x1_ASAP7_75t_L g1732 ( 
.A1(n_1516),
.A2(n_1405),
.B(n_1404),
.Y(n_1732)
);

AO21x2_ASAP7_75t_L g1733 ( 
.A1(n_1478),
.A2(n_1487),
.B(n_1527),
.Y(n_1733)
);

AO21x2_ASAP7_75t_L g1734 ( 
.A1(n_1527),
.A2(n_1564),
.B(n_1587),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1403),
.Y(n_1735)
);

OA21x2_ASAP7_75t_L g1736 ( 
.A1(n_1445),
.A2(n_1507),
.B(n_1379),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1428),
.B(n_1513),
.Y(n_1737)
);

NOR2x1_ASAP7_75t_R g1738 ( 
.A(n_1448),
.B(n_1466),
.Y(n_1738)
);

AND2x4_ASAP7_75t_L g1739 ( 
.A(n_1414),
.B(n_1471),
.Y(n_1739)
);

OAI21x1_ASAP7_75t_SL g1740 ( 
.A1(n_1402),
.A2(n_1422),
.B(n_1354),
.Y(n_1740)
);

OAI21x1_ASAP7_75t_L g1741 ( 
.A1(n_1380),
.A2(n_1449),
.B(n_1539),
.Y(n_1741)
);

OAI21x1_ASAP7_75t_L g1742 ( 
.A1(n_1541),
.A2(n_1475),
.B(n_1397),
.Y(n_1742)
);

INVx4_ASAP7_75t_L g1743 ( 
.A(n_1520),
.Y(n_1743)
);

NOR2xp33_ASAP7_75t_L g1744 ( 
.A(n_1514),
.B(n_1368),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1476),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1476),
.Y(n_1746)
);

OR2x6_ASAP7_75t_L g1747 ( 
.A(n_1520),
.B(n_1480),
.Y(n_1747)
);

OAI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1505),
.A2(n_1447),
.B(n_1422),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1399),
.B(n_1525),
.Y(n_1749)
);

OAI21x1_ASAP7_75t_L g1750 ( 
.A1(n_1407),
.A2(n_1492),
.B(n_1489),
.Y(n_1750)
);

OAI21x1_ASAP7_75t_L g1751 ( 
.A1(n_1492),
.A2(n_1489),
.B(n_1515),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_1467),
.B(n_1492),
.Y(n_1752)
);

BUFx3_ASAP7_75t_L g1753 ( 
.A(n_1460),
.Y(n_1753)
);

OA21x2_ASAP7_75t_L g1754 ( 
.A1(n_1433),
.A2(n_1409),
.B(n_1453),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1460),
.B(n_1423),
.Y(n_1755)
);

INVxp67_ASAP7_75t_L g1756 ( 
.A(n_1453),
.Y(n_1756)
);

NAND2x1p5_ASAP7_75t_L g1757 ( 
.A(n_1409),
.B(n_1352),
.Y(n_1757)
);

OR2x6_ASAP7_75t_L g1758 ( 
.A(n_1483),
.B(n_1486),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1353),
.Y(n_1759)
);

AOI21xp33_ASAP7_75t_L g1760 ( 
.A1(n_1498),
.A2(n_1565),
.B(n_1431),
.Y(n_1760)
);

NAND3xp33_ASAP7_75t_L g1761 ( 
.A(n_1400),
.B(n_1565),
.C(n_1452),
.Y(n_1761)
);

BUFx3_ASAP7_75t_L g1762 ( 
.A(n_1352),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1353),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1353),
.Y(n_1764)
);

OAI21x1_ASAP7_75t_SL g1765 ( 
.A1(n_1548),
.A2(n_1442),
.B(n_1386),
.Y(n_1765)
);

OA21x2_ASAP7_75t_L g1766 ( 
.A1(n_1528),
.A2(n_1534),
.B(n_1530),
.Y(n_1766)
);

BUFx3_ASAP7_75t_L g1767 ( 
.A(n_1352),
.Y(n_1767)
);

INVx2_ASAP7_75t_SL g1768 ( 
.A(n_1352),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1388),
.Y(n_1769)
);

AO222x2_ASAP7_75t_L g1770 ( 
.A1(n_1399),
.A2(n_1222),
.B1(n_1016),
.B2(n_1044),
.C1(n_1161),
.C2(n_945),
.Y(n_1770)
);

OR2x6_ASAP7_75t_L g1771 ( 
.A(n_1483),
.B(n_1486),
.Y(n_1771)
);

AO21x2_ASAP7_75t_L g1772 ( 
.A1(n_1390),
.A2(n_1386),
.B(n_1176),
.Y(n_1772)
);

AO21x2_ASAP7_75t_L g1773 ( 
.A1(n_1390),
.A2(n_1386),
.B(n_1176),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1532),
.B(n_1533),
.Y(n_1774)
);

INVx3_ASAP7_75t_L g1775 ( 
.A(n_1352),
.Y(n_1775)
);

BUFx2_ASAP7_75t_L g1776 ( 
.A(n_1586),
.Y(n_1776)
);

AO21x2_ASAP7_75t_L g1777 ( 
.A1(n_1390),
.A2(n_1386),
.B(n_1176),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1532),
.B(n_1533),
.Y(n_1778)
);

OAI21x1_ASAP7_75t_SL g1779 ( 
.A1(n_1548),
.A2(n_1442),
.B(n_1386),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1532),
.B(n_1533),
.Y(n_1780)
);

INVx6_ASAP7_75t_L g1781 ( 
.A(n_1352),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1353),
.Y(n_1782)
);

OAI21xp5_ASAP7_75t_L g1783 ( 
.A1(n_1366),
.A2(n_1558),
.B(n_1563),
.Y(n_1783)
);

INVxp67_ASAP7_75t_SL g1784 ( 
.A(n_1532),
.Y(n_1784)
);

AOI22x1_ASAP7_75t_L g1785 ( 
.A1(n_1521),
.A2(n_1254),
.B1(n_1459),
.B2(n_1523),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1353),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1532),
.A2(n_1545),
.B1(n_1549),
.B2(n_1533),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1353),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1532),
.B(n_1533),
.Y(n_1789)
);

OAI21x1_ASAP7_75t_SL g1790 ( 
.A1(n_1548),
.A2(n_1442),
.B(n_1386),
.Y(n_1790)
);

AOI22x1_ASAP7_75t_L g1791 ( 
.A1(n_1521),
.A2(n_1254),
.B1(n_1459),
.B2(n_1523),
.Y(n_1791)
);

OAI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1366),
.A2(n_1558),
.B(n_1563),
.Y(n_1792)
);

OAI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1366),
.A2(n_1558),
.B(n_1563),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1353),
.Y(n_1794)
);

INVx3_ASAP7_75t_L g1795 ( 
.A(n_1606),
.Y(n_1795)
);

BUFx2_ASAP7_75t_R g1796 ( 
.A(n_1618),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1600),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1612),
.Y(n_1798)
);

INVx5_ASAP7_75t_L g1799 ( 
.A(n_1643),
.Y(n_1799)
);

INVx4_ASAP7_75t_L g1800 ( 
.A(n_1643),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1593),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1614),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1624),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1759),
.Y(n_1804)
);

AOI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1621),
.A2(n_1787),
.B1(n_1661),
.B2(n_1774),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1763),
.Y(n_1806)
);

INVx3_ASAP7_75t_L g1807 ( 
.A(n_1606),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1764),
.Y(n_1808)
);

AOI22xp33_ASAP7_75t_SL g1809 ( 
.A1(n_1639),
.A2(n_1721),
.B1(n_1591),
.B2(n_1784),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1593),
.Y(n_1810)
);

INVx4_ASAP7_75t_L g1811 ( 
.A(n_1643),
.Y(n_1811)
);

AOI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1634),
.A2(n_1591),
.B1(n_1661),
.B2(n_1629),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1782),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1629),
.B(n_1774),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1786),
.Y(n_1815)
);

NAND2x1_ASAP7_75t_L g1816 ( 
.A(n_1594),
.B(n_1765),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1788),
.Y(n_1817)
);

INVx2_ASAP7_75t_SL g1818 ( 
.A(n_1654),
.Y(n_1818)
);

AOI22xp33_ASAP7_75t_L g1819 ( 
.A1(n_1634),
.A2(n_1778),
.B1(n_1780),
.B2(n_1760),
.Y(n_1819)
);

INVx3_ASAP7_75t_L g1820 ( 
.A(n_1643),
.Y(n_1820)
);

BUFx3_ASAP7_75t_L g1821 ( 
.A(n_1595),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1769),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1620),
.B(n_1682),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1778),
.A2(n_1780),
.B1(n_1646),
.B2(n_1639),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1794),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1630),
.Y(n_1826)
);

INVx3_ASAP7_75t_L g1827 ( 
.A(n_1619),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1633),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1607),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1609),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1650),
.B(n_1617),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1609),
.Y(n_1832)
);

INVx3_ASAP7_75t_L g1833 ( 
.A(n_1619),
.Y(n_1833)
);

AOI22xp33_ASAP7_75t_SL g1834 ( 
.A1(n_1639),
.A2(n_1727),
.B1(n_1640),
.B2(n_1596),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1642),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1670),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1645),
.Y(n_1837)
);

AOI22xp33_ASAP7_75t_L g1838 ( 
.A1(n_1646),
.A2(n_1639),
.B1(n_1657),
.B2(n_1680),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1613),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1599),
.B(n_1605),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1613),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1645),
.Y(n_1842)
);

OAI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1638),
.A2(n_1703),
.B(n_1761),
.Y(n_1843)
);

CKINVDCx20_ASAP7_75t_R g1844 ( 
.A(n_1637),
.Y(n_1844)
);

BUFx3_ASAP7_75t_L g1845 ( 
.A(n_1601),
.Y(n_1845)
);

BUFx3_ASAP7_75t_L g1846 ( 
.A(n_1608),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1686),
.Y(n_1847)
);

AOI222xp33_ASAP7_75t_L g1848 ( 
.A1(n_1718),
.A2(n_1715),
.B1(n_1737),
.B2(n_1657),
.C1(n_1770),
.C2(n_1680),
.Y(n_1848)
);

INVx4_ASAP7_75t_SL g1849 ( 
.A(n_1616),
.Y(n_1849)
);

INVx4_ASAP7_75t_L g1850 ( 
.A(n_1628),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1615),
.B(n_1622),
.Y(n_1851)
);

INVx6_ASAP7_75t_L g1852 ( 
.A(n_1616),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1648),
.B(n_1789),
.Y(n_1853)
);

INVx3_ASAP7_75t_L g1854 ( 
.A(n_1619),
.Y(n_1854)
);

INVx3_ASAP7_75t_L g1855 ( 
.A(n_1626),
.Y(n_1855)
);

AOI22xp33_ASAP7_75t_L g1856 ( 
.A1(n_1707),
.A2(n_1647),
.B1(n_1698),
.B2(n_1736),
.Y(n_1856)
);

AOI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1698),
.A2(n_1736),
.B1(n_1666),
.B2(n_1668),
.Y(n_1857)
);

OR2x6_ASAP7_75t_L g1858 ( 
.A(n_1596),
.B(n_1625),
.Y(n_1858)
);

INVx3_ASAP7_75t_L g1859 ( 
.A(n_1626),
.Y(n_1859)
);

OAI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1596),
.A2(n_1625),
.B1(n_1771),
.B2(n_1758),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1709),
.B(n_1649),
.Y(n_1861)
);

INVx2_ASAP7_75t_SL g1862 ( 
.A(n_1654),
.Y(n_1862)
);

AOI22xp33_ASAP7_75t_L g1863 ( 
.A1(n_1736),
.A2(n_1625),
.B1(n_1758),
.B2(n_1596),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1636),
.B(n_1592),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1695),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1655),
.B(n_1656),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1695),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1610),
.B(n_1776),
.Y(n_1868)
);

AOI22xp33_ASAP7_75t_L g1869 ( 
.A1(n_1625),
.A2(n_1758),
.B1(n_1771),
.B2(n_1683),
.Y(n_1869)
);

AO21x1_ASAP7_75t_L g1870 ( 
.A1(n_1745),
.A2(n_1746),
.B(n_1757),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1704),
.Y(n_1871)
);

INVx6_ASAP7_75t_L g1872 ( 
.A(n_1616),
.Y(n_1872)
);

AOI22xp33_ASAP7_75t_L g1873 ( 
.A1(n_1758),
.A2(n_1771),
.B1(n_1692),
.B2(n_1696),
.Y(n_1873)
);

BUFx3_ASAP7_75t_L g1874 ( 
.A(n_1608),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1701),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1713),
.Y(n_1876)
);

CKINVDCx8_ASAP7_75t_R g1877 ( 
.A(n_1652),
.Y(n_1877)
);

OAI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1771),
.A2(n_1681),
.B1(n_1724),
.B2(n_1748),
.Y(n_1878)
);

OR2x6_ASAP7_75t_L g1879 ( 
.A(n_1768),
.B(n_1781),
.Y(n_1879)
);

INVx2_ASAP7_75t_SL g1880 ( 
.A(n_1654),
.Y(n_1880)
);

INVx1_ASAP7_75t_SL g1881 ( 
.A(n_1725),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1602),
.Y(n_1882)
);

NOR2x1_ASAP7_75t_SL g1883 ( 
.A(n_1762),
.B(n_1767),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1744),
.B(n_1687),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1716),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1717),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1719),
.Y(n_1887)
);

CKINVDCx11_ASAP7_75t_R g1888 ( 
.A(n_1637),
.Y(n_1888)
);

AOI22xp33_ASAP7_75t_SL g1889 ( 
.A1(n_1732),
.A2(n_1740),
.B1(n_1749),
.B2(n_1705),
.Y(n_1889)
);

CKINVDCx20_ASAP7_75t_R g1890 ( 
.A(n_1618),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1768),
.Y(n_1891)
);

INVx6_ASAP7_75t_L g1892 ( 
.A(n_1781),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1662),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1664),
.B(n_1669),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1674),
.Y(n_1895)
);

INVx3_ASAP7_75t_L g1896 ( 
.A(n_1626),
.Y(n_1896)
);

AO21x1_ASAP7_75t_L g1897 ( 
.A1(n_1783),
.A2(n_1793),
.B(n_1792),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1677),
.Y(n_1898)
);

INVx3_ASAP7_75t_L g1899 ( 
.A(n_1775),
.Y(n_1899)
);

AOI22xp33_ASAP7_75t_L g1900 ( 
.A1(n_1688),
.A2(n_1702),
.B1(n_1697),
.B2(n_1752),
.Y(n_1900)
);

INVx6_ASAP7_75t_L g1901 ( 
.A(n_1781),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1762),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1744),
.B(n_1714),
.Y(n_1903)
);

BUFx2_ASAP7_75t_L g1904 ( 
.A(n_1743),
.Y(n_1904)
);

INVx3_ASAP7_75t_L g1905 ( 
.A(n_1672),
.Y(n_1905)
);

BUFx3_ASAP7_75t_L g1906 ( 
.A(n_1691),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1691),
.Y(n_1907)
);

AOI22xp33_ASAP7_75t_SL g1908 ( 
.A1(n_1732),
.A2(n_1749),
.B1(n_1611),
.B2(n_1752),
.Y(n_1908)
);

BUFx2_ASAP7_75t_L g1909 ( 
.A(n_1743),
.Y(n_1909)
);

AOI22xp33_ASAP7_75t_L g1910 ( 
.A1(n_1752),
.A2(n_1712),
.B1(n_1611),
.B2(n_1731),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1766),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1671),
.B(n_1735),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_SL g1913 ( 
.A(n_1779),
.B(n_1790),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1691),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1720),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1720),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1720),
.Y(n_1917)
);

AO21x1_ASAP7_75t_SL g1918 ( 
.A1(n_1672),
.A2(n_1663),
.B(n_1711),
.Y(n_1918)
);

NAND2x1p5_ASAP7_75t_L g1919 ( 
.A(n_1672),
.B(n_1631),
.Y(n_1919)
);

INVx2_ASAP7_75t_SL g1920 ( 
.A(n_1628),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1751),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1751),
.Y(n_1922)
);

BUFx2_ASAP7_75t_L g1923 ( 
.A(n_1743),
.Y(n_1923)
);

INVx3_ASAP7_75t_L g1924 ( 
.A(n_1631),
.Y(n_1924)
);

CKINVDCx20_ASAP7_75t_R g1925 ( 
.A(n_1632),
.Y(n_1925)
);

BUFx3_ASAP7_75t_L g1926 ( 
.A(n_1644),
.Y(n_1926)
);

INVx4_ASAP7_75t_L g1927 ( 
.A(n_1676),
.Y(n_1927)
);

OAI21xp5_ASAP7_75t_L g1928 ( 
.A1(n_1673),
.A2(n_1700),
.B(n_1699),
.Y(n_1928)
);

NAND2x1p5_ASAP7_75t_L g1929 ( 
.A(n_1658),
.B(n_1627),
.Y(n_1929)
);

OR2x2_ASAP7_75t_L g1930 ( 
.A(n_1627),
.B(n_1641),
.Y(n_1930)
);

BUFx2_ASAP7_75t_L g1931 ( 
.A(n_1729),
.Y(n_1931)
);

CKINVDCx20_ASAP7_75t_R g1932 ( 
.A(n_1632),
.Y(n_1932)
);

BUFx3_ASAP7_75t_L g1933 ( 
.A(n_1729),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1754),
.Y(n_1934)
);

OAI22xp33_ASAP7_75t_SL g1935 ( 
.A1(n_1641),
.A2(n_1739),
.B1(n_1770),
.B2(n_1756),
.Y(n_1935)
);

INVx3_ASAP7_75t_L g1936 ( 
.A(n_1728),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1754),
.Y(n_1937)
);

AOI22xp5_ASAP7_75t_SL g1938 ( 
.A1(n_1603),
.A2(n_1689),
.B1(n_1739),
.B2(n_1755),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1726),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1911),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1814),
.B(n_1659),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1840),
.B(n_1659),
.Y(n_1942)
);

BUFx2_ASAP7_75t_L g1943 ( 
.A(n_1821),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1797),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1798),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1831),
.B(n_1728),
.Y(n_1946)
);

INVx3_ASAP7_75t_L g1947 ( 
.A(n_1800),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1903),
.B(n_1728),
.Y(n_1948)
);

OR2x2_ASAP7_75t_L g1949 ( 
.A(n_1823),
.B(n_1733),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1802),
.Y(n_1950)
);

BUFx3_ASAP7_75t_L g1951 ( 
.A(n_1877),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1803),
.Y(n_1952)
);

BUFx2_ASAP7_75t_L g1953 ( 
.A(n_1821),
.Y(n_1953)
);

INVxp67_ASAP7_75t_L g1954 ( 
.A(n_1805),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1853),
.B(n_1836),
.Y(n_1955)
);

INVx2_ASAP7_75t_SL g1956 ( 
.A(n_1799),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1884),
.B(n_1690),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1804),
.Y(n_1958)
);

INVx4_ASAP7_75t_L g1959 ( 
.A(n_1799),
.Y(n_1959)
);

HB1xp67_ASAP7_75t_L g1960 ( 
.A(n_1801),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1848),
.B(n_1851),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1912),
.B(n_1690),
.Y(n_1962)
);

AOI22xp33_ASAP7_75t_L g1963 ( 
.A1(n_1812),
.A2(n_1712),
.B1(n_1731),
.B2(n_1710),
.Y(n_1963)
);

INVx3_ASAP7_75t_L g1964 ( 
.A(n_1800),
.Y(n_1964)
);

BUFx2_ASAP7_75t_L g1965 ( 
.A(n_1845),
.Y(n_1965)
);

AND2x4_ASAP7_75t_SL g1966 ( 
.A(n_1811),
.B(n_1747),
.Y(n_1966)
);

BUFx5_ASAP7_75t_L g1967 ( 
.A(n_1845),
.Y(n_1967)
);

HB1xp67_ASAP7_75t_L g1968 ( 
.A(n_1801),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1806),
.Y(n_1969)
);

OR2x2_ASAP7_75t_L g1970 ( 
.A(n_1864),
.B(n_1733),
.Y(n_1970)
);

OR2x2_ASAP7_75t_L g1971 ( 
.A(n_1868),
.B(n_1678),
.Y(n_1971)
);

HB1xp67_ASAP7_75t_L g1972 ( 
.A(n_1810),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1808),
.Y(n_1973)
);

INVx3_ASAP7_75t_L g1974 ( 
.A(n_1811),
.Y(n_1974)
);

AOI221xp5_ASAP7_75t_L g1975 ( 
.A1(n_1935),
.A2(n_1755),
.B1(n_1660),
.B2(n_1734),
.C(n_1723),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1813),
.Y(n_1976)
);

BUFx3_ASAP7_75t_L g1977 ( 
.A(n_1799),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1815),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1865),
.B(n_1867),
.Y(n_1979)
);

AOI22xp33_ASAP7_75t_L g1980 ( 
.A1(n_1812),
.A2(n_1710),
.B1(n_1730),
.B2(n_1635),
.Y(n_1980)
);

BUFx2_ASAP7_75t_L g1981 ( 
.A(n_1846),
.Y(n_1981)
);

AOI22xp33_ASAP7_75t_L g1982 ( 
.A1(n_1819),
.A2(n_1730),
.B1(n_1635),
.B2(n_1604),
.Y(n_1982)
);

BUFx2_ASAP7_75t_L g1983 ( 
.A(n_1846),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1817),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1825),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1826),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1828),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1835),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1893),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1926),
.B(n_1722),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1895),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1898),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1926),
.B(n_1722),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1866),
.Y(n_1994)
);

BUFx6f_ASAP7_75t_L g1995 ( 
.A(n_1918),
.Y(n_1995)
);

BUFx3_ASAP7_75t_L g1996 ( 
.A(n_1799),
.Y(n_1996)
);

AND2x4_ASAP7_75t_L g1997 ( 
.A(n_1858),
.B(n_1742),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1894),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1875),
.Y(n_1999)
);

NOR2xp67_ASAP7_75t_L g2000 ( 
.A(n_1850),
.B(n_1665),
.Y(n_2000)
);

BUFx3_ASAP7_75t_L g2001 ( 
.A(n_1820),
.Y(n_2001)
);

AO31x2_ASAP7_75t_L g2002 ( 
.A1(n_1897),
.A2(n_1870),
.A3(n_1829),
.B(n_1830),
.Y(n_2002)
);

NAND2x1p5_ASAP7_75t_L g2003 ( 
.A(n_1850),
.B(n_1694),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1876),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1871),
.B(n_1722),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1885),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1886),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1887),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1861),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1819),
.B(n_1685),
.Y(n_2010)
);

OAI22xp5_ASAP7_75t_L g2011 ( 
.A1(n_1824),
.A2(n_1597),
.B1(n_1747),
.B2(n_1651),
.Y(n_2011)
);

AND2x4_ASAP7_75t_L g2012 ( 
.A(n_1858),
.B(n_1742),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1837),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1842),
.Y(n_2014)
);

INVx4_ASAP7_75t_L g2015 ( 
.A(n_1820),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1847),
.Y(n_2016)
);

INVx3_ASAP7_75t_L g2017 ( 
.A(n_1919),
.Y(n_2017)
);

HB1xp67_ASAP7_75t_L g2018 ( 
.A(n_1822),
.Y(n_2018)
);

OAI21xp5_ASAP7_75t_SL g2019 ( 
.A1(n_1881),
.A2(n_1738),
.B(n_1679),
.Y(n_2019)
);

INVx2_ASAP7_75t_SL g2020 ( 
.A(n_1874),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1795),
.B(n_1741),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1795),
.B(n_1741),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1807),
.B(n_1685),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1807),
.B(n_1685),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1891),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1902),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1874),
.B(n_1685),
.Y(n_2027)
);

INVx4_ASAP7_75t_R g2028 ( 
.A(n_1920),
.Y(n_2028)
);

AOI22xp33_ASAP7_75t_L g2029 ( 
.A1(n_1824),
.A2(n_1604),
.B1(n_1772),
.B2(n_1777),
.Y(n_2029)
);

BUFx2_ASAP7_75t_L g2030 ( 
.A(n_1879),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1934),
.Y(n_2031)
);

OR2x2_ASAP7_75t_L g2032 ( 
.A(n_1904),
.B(n_1684),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1909),
.B(n_1694),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1937),
.Y(n_2034)
);

AND2x4_ASAP7_75t_L g2035 ( 
.A(n_1913),
.B(n_1750),
.Y(n_2035)
);

INVxp67_ASAP7_75t_L g2036 ( 
.A(n_1923),
.Y(n_2036)
);

NOR2x1_ASAP7_75t_L g2037 ( 
.A(n_1927),
.B(n_1706),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1906),
.B(n_1706),
.Y(n_2038)
);

AOI22xp33_ASAP7_75t_L g2039 ( 
.A1(n_1838),
.A2(n_1777),
.B1(n_1773),
.B2(n_1772),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1856),
.B(n_1684),
.Y(n_2040)
);

AND2x4_ASAP7_75t_SL g2041 ( 
.A(n_1927),
.B(n_1665),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1883),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1906),
.B(n_1753),
.Y(n_2043)
);

AOI22xp33_ASAP7_75t_L g2044 ( 
.A1(n_1838),
.A2(n_1773),
.B1(n_1623),
.B2(n_1693),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1930),
.Y(n_2045)
);

BUFx3_ASAP7_75t_L g2046 ( 
.A(n_1879),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1856),
.B(n_1734),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1924),
.B(n_1753),
.Y(n_2048)
);

AOI22xp33_ASAP7_75t_L g2049 ( 
.A1(n_1860),
.A2(n_1623),
.B1(n_1693),
.B2(n_1653),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1907),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1857),
.B(n_1598),
.Y(n_2051)
);

AND2x4_ASAP7_75t_L g2052 ( 
.A(n_1913),
.B(n_1750),
.Y(n_2052)
);

AOI22xp33_ASAP7_75t_L g2053 ( 
.A1(n_1860),
.A2(n_1693),
.B1(n_1653),
.B2(n_1651),
.Y(n_2053)
);

INVx2_ASAP7_75t_SL g2054 ( 
.A(n_1995),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_2005),
.B(n_1908),
.Y(n_2055)
);

BUFx3_ASAP7_75t_L g2056 ( 
.A(n_1943),
.Y(n_2056)
);

AND2x2_ASAP7_75t_SL g2057 ( 
.A(n_1995),
.B(n_1863),
.Y(n_2057)
);

INVx2_ASAP7_75t_SL g2058 ( 
.A(n_1995),
.Y(n_2058)
);

BUFx3_ASAP7_75t_L g2059 ( 
.A(n_1953),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1944),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_2023),
.B(n_1908),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1940),
.Y(n_2062)
);

OR2x2_ASAP7_75t_L g2063 ( 
.A(n_1955),
.B(n_1900),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_2024),
.B(n_1910),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1945),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_2027),
.B(n_1910),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1990),
.B(n_1921),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_1993),
.B(n_1922),
.Y(n_2068)
);

OR2x2_ASAP7_75t_L g2069 ( 
.A(n_1949),
.B(n_1857),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1950),
.Y(n_2070)
);

OR2x2_ASAP7_75t_L g2071 ( 
.A(n_1971),
.B(n_1900),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_2031),
.B(n_2034),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1954),
.B(n_1863),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1952),
.Y(n_2074)
);

OAI222xp33_ASAP7_75t_L g2075 ( 
.A1(n_1954),
.A2(n_1809),
.B1(n_1834),
.B2(n_1878),
.C1(n_1869),
.C2(n_1873),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1958),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1969),
.Y(n_2077)
);

INVx1_ASAP7_75t_SL g2078 ( 
.A(n_1951),
.Y(n_2078)
);

OR2x2_ASAP7_75t_L g2079 ( 
.A(n_2036),
.B(n_1931),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_1960),
.B(n_1889),
.Y(n_2080)
);

INVx2_ASAP7_75t_SL g2081 ( 
.A(n_1995),
.Y(n_2081)
);

BUFx2_ASAP7_75t_L g2082 ( 
.A(n_2042),
.Y(n_2082)
);

INVx3_ASAP7_75t_L g2083 ( 
.A(n_2035),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_1968),
.B(n_1889),
.Y(n_2084)
);

NOR2xp67_ASAP7_75t_L g2085 ( 
.A(n_1959),
.B(n_1905),
.Y(n_2085)
);

AND2x4_ASAP7_75t_SL g2086 ( 
.A(n_1959),
.B(n_1905),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1973),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1976),
.Y(n_2088)
);

INVx2_ASAP7_75t_SL g2089 ( 
.A(n_1965),
.Y(n_2089)
);

OR2x2_ASAP7_75t_L g2090 ( 
.A(n_1970),
.B(n_1882),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_1968),
.B(n_1972),
.Y(n_2091)
);

NAND3x1_ASAP7_75t_L g2092 ( 
.A(n_1947),
.B(n_1938),
.C(n_1924),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_SL g2093 ( 
.A(n_1967),
.B(n_1809),
.Y(n_2093)
);

HB1xp67_ASAP7_75t_L g2094 ( 
.A(n_2036),
.Y(n_2094)
);

NAND2xp33_ASAP7_75t_SL g2095 ( 
.A(n_2015),
.B(n_1816),
.Y(n_2095)
);

HB1xp67_ASAP7_75t_L g2096 ( 
.A(n_1981),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1978),
.Y(n_2097)
);

BUFx2_ASAP7_75t_L g2098 ( 
.A(n_1983),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1984),
.Y(n_2099)
);

BUFx2_ASAP7_75t_L g2100 ( 
.A(n_2020),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1985),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1986),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1987),
.Y(n_2103)
);

OAI222xp33_ASAP7_75t_L g2104 ( 
.A1(n_2015),
.A2(n_1834),
.B1(n_1869),
.B2(n_1873),
.C1(n_1929),
.C2(n_1919),
.Y(n_2104)
);

NOR2xp33_ASAP7_75t_L g2105 ( 
.A(n_1961),
.B(n_1914),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1988),
.Y(n_2106)
);

NOR2xp33_ASAP7_75t_L g2107 ( 
.A(n_2009),
.B(n_1915),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1989),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1991),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_1994),
.B(n_1843),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_1998),
.B(n_1936),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1992),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1999),
.Y(n_2113)
);

AOI22xp5_ASAP7_75t_L g2114 ( 
.A1(n_1975),
.A2(n_1818),
.B1(n_1862),
.B2(n_1880),
.Y(n_2114)
);

INVx1_ASAP7_75t_SL g2115 ( 
.A(n_1951),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2004),
.Y(n_2116)
);

HB1xp67_ASAP7_75t_L g2117 ( 
.A(n_2020),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_1979),
.B(n_1936),
.Y(n_2118)
);

OR2x2_ASAP7_75t_L g2119 ( 
.A(n_2010),
.B(n_2018),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2006),
.Y(n_2120)
);

AOI22xp33_ASAP7_75t_L g2121 ( 
.A1(n_1946),
.A2(n_1708),
.B1(n_1785),
.B2(n_1791),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2007),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_2029),
.B(n_1832),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_2029),
.B(n_1832),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_2045),
.B(n_1827),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_2008),
.B(n_1827),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_2044),
.B(n_1839),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2044),
.B(n_1839),
.Y(n_2128)
);

OR2x2_ASAP7_75t_L g2129 ( 
.A(n_1941),
.B(n_1933),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2021),
.B(n_1841),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2026),
.Y(n_2131)
);

INVx4_ASAP7_75t_L g2132 ( 
.A(n_1977),
.Y(n_2132)
);

INVx2_ASAP7_75t_SL g2133 ( 
.A(n_1967),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_2022),
.B(n_2049),
.Y(n_2134)
);

AND2x4_ASAP7_75t_L g2135 ( 
.A(n_1997),
.B(n_1928),
.Y(n_2135)
);

OR2x2_ASAP7_75t_SL g2136 ( 
.A(n_2028),
.B(n_1888),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2064),
.B(n_2049),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_2062),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2064),
.B(n_2035),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2055),
.B(n_2035),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_2110),
.B(n_2025),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_2105),
.B(n_2013),
.Y(n_2142)
);

OR2x2_ASAP7_75t_L g2143 ( 
.A(n_2119),
.B(n_2069),
.Y(n_2143)
);

CKINVDCx5p33_ASAP7_75t_R g2144 ( 
.A(n_2078),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2072),
.Y(n_2145)
);

NOR2xp67_ASAP7_75t_L g2146 ( 
.A(n_2132),
.B(n_1956),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_SL g2147 ( 
.A(n_2132),
.B(n_2000),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2105),
.B(n_2014),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2055),
.B(n_1980),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_2066),
.B(n_2052),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2066),
.B(n_2052),
.Y(n_2151)
);

AND2x4_ASAP7_75t_L g2152 ( 
.A(n_2135),
.B(n_2052),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2061),
.B(n_1997),
.Y(n_2153)
);

INVx3_ASAP7_75t_L g2154 ( 
.A(n_2083),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_2072),
.B(n_1980),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_2069),
.B(n_1963),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2060),
.Y(n_2157)
);

OR2x2_ASAP7_75t_L g2158 ( 
.A(n_2119),
.B(n_2047),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2061),
.B(n_1997),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_2065),
.B(n_1963),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2070),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_2082),
.B(n_2016),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_2067),
.B(n_2012),
.Y(n_2163)
);

AND2x4_ASAP7_75t_L g2164 ( 
.A(n_2135),
.B(n_2012),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2067),
.B(n_2012),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2074),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2076),
.Y(n_2167)
);

INVx1_ASAP7_75t_SL g2168 ( 
.A(n_2056),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2077),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_2068),
.B(n_2053),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_2068),
.B(n_2053),
.Y(n_2171)
);

OR2x2_ASAP7_75t_L g2172 ( 
.A(n_2071),
.B(n_2051),
.Y(n_2172)
);

HB1xp67_ASAP7_75t_L g2173 ( 
.A(n_2096),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_2134),
.B(n_2039),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_2134),
.B(n_2130),
.Y(n_2175)
);

OR2x2_ASAP7_75t_L g2176 ( 
.A(n_2091),
.B(n_2040),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_2130),
.B(n_2039),
.Y(n_2177)
);

AND2x4_ASAP7_75t_L g2178 ( 
.A(n_2135),
.B(n_2002),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2087),
.Y(n_2179)
);

INVx1_ASAP7_75t_SL g2180 ( 
.A(n_2056),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2088),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_2097),
.B(n_1982),
.Y(n_2182)
);

NOR2xp33_ASAP7_75t_L g2183 ( 
.A(n_2115),
.B(n_2019),
.Y(n_2183)
);

OR2x2_ASAP7_75t_L g2184 ( 
.A(n_2091),
.B(n_2032),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_2123),
.B(n_1982),
.Y(n_2185)
);

OR2x2_ASAP7_75t_L g2186 ( 
.A(n_2143),
.B(n_2090),
.Y(n_2186)
);

INVxp67_ASAP7_75t_L g2187 ( 
.A(n_2173),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2157),
.Y(n_2188)
);

NAND3xp33_ASAP7_75t_L g2189 ( 
.A(n_2156),
.B(n_2094),
.C(n_2114),
.Y(n_2189)
);

OAI211xp5_ASAP7_75t_L g2190 ( 
.A1(n_2183),
.A2(n_2098),
.B(n_1888),
.C(n_2095),
.Y(n_2190)
);

OAI21xp33_ASAP7_75t_L g2191 ( 
.A1(n_2153),
.A2(n_2057),
.B(n_2080),
.Y(n_2191)
);

OR2x2_ASAP7_75t_L g2192 ( 
.A(n_2143),
.B(n_2158),
.Y(n_2192)
);

AND2x2_ASAP7_75t_L g2193 ( 
.A(n_2175),
.B(n_2080),
.Y(n_2193)
);

NAND2x1_ASAP7_75t_L g2194 ( 
.A(n_2146),
.B(n_2132),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_2137),
.B(n_2089),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2157),
.Y(n_2196)
);

HB1xp67_ASAP7_75t_L g2197 ( 
.A(n_2168),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_2175),
.B(n_2084),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2139),
.B(n_2084),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2161),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2161),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_2139),
.B(n_2123),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2166),
.Y(n_2203)
);

HB1xp67_ASAP7_75t_L g2204 ( 
.A(n_2168),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_2140),
.B(n_2124),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2166),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_2140),
.B(n_2124),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2167),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_2138),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2137),
.B(n_2149),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2167),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2169),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2169),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2179),
.Y(n_2214)
);

OR2x2_ASAP7_75t_L g2215 ( 
.A(n_2158),
.B(n_2176),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_2150),
.B(n_2127),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_2150),
.B(n_2127),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_2149),
.B(n_2089),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_2151),
.B(n_2128),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2179),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2181),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2181),
.Y(n_2222)
);

BUFx2_ASAP7_75t_L g2223 ( 
.A(n_2180),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_2151),
.B(n_2153),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_2159),
.B(n_2128),
.Y(n_2225)
);

AOI221xp5_ASAP7_75t_L g2226 ( 
.A1(n_2187),
.A2(n_2148),
.B1(n_2142),
.B2(n_2174),
.C(n_2075),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_SL g2227 ( 
.A(n_2223),
.B(n_2146),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2193),
.B(n_2198),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2192),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2192),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_2193),
.B(n_2159),
.Y(n_2231)
);

INVx1_ASAP7_75t_SL g2232 ( 
.A(n_2223),
.Y(n_2232)
);

AND2x4_ASAP7_75t_L g2233 ( 
.A(n_2194),
.B(n_2164),
.Y(n_2233)
);

AOI22xp5_ASAP7_75t_L g2234 ( 
.A1(n_2191),
.A2(n_2057),
.B1(n_2174),
.B2(n_2185),
.Y(n_2234)
);

AND2x2_ASAP7_75t_L g2235 ( 
.A(n_2198),
.B(n_2163),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2215),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2224),
.B(n_2163),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_2209),
.Y(n_2238)
);

AOI22xp5_ASAP7_75t_L g2239 ( 
.A1(n_2190),
.A2(n_2185),
.B1(n_2156),
.B2(n_2171),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2215),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2186),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_2209),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2186),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2210),
.B(n_2170),
.Y(n_2244)
);

AND2x2_ASAP7_75t_L g2245 ( 
.A(n_2224),
.B(n_2165),
.Y(n_2245)
);

OAI22xp33_ASAP7_75t_L g2246 ( 
.A1(n_2194),
.A2(n_2180),
.B1(n_2059),
.B2(n_2100),
.Y(n_2246)
);

OR2x2_ASAP7_75t_L g2247 ( 
.A(n_2218),
.B(n_2176),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2196),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_2196),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_2200),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2199),
.B(n_2170),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2200),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_SL g2253 ( 
.A(n_2197),
.B(n_2144),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_2199),
.B(n_2171),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_2189),
.B(n_2172),
.Y(n_2255)
);

OAI22xp5_ASAP7_75t_L g2256 ( 
.A1(n_2204),
.A2(n_2092),
.B1(n_2136),
.B2(n_2162),
.Y(n_2256)
);

OAI21xp33_ASAP7_75t_L g2257 ( 
.A1(n_2195),
.A2(n_2172),
.B(n_2165),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2201),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2225),
.B(n_2177),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2201),
.Y(n_2260)
);

OR2x2_ASAP7_75t_L g2261 ( 
.A(n_2216),
.B(n_2184),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_2225),
.B(n_2178),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2203),
.Y(n_2263)
);

AOI21xp5_ASAP7_75t_L g2264 ( 
.A1(n_2227),
.A2(n_2095),
.B(n_2147),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2248),
.Y(n_2265)
);

OAI22xp5_ASAP7_75t_L g2266 ( 
.A1(n_2256),
.A2(n_2092),
.B1(n_2059),
.B2(n_2164),
.Y(n_2266)
);

HB1xp67_ASAP7_75t_L g2267 ( 
.A(n_2232),
.Y(n_2267)
);

OAI22xp5_ASAP7_75t_L g2268 ( 
.A1(n_2239),
.A2(n_2164),
.B1(n_2184),
.B2(n_2205),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2252),
.Y(n_2269)
);

OAI22xp5_ASAP7_75t_L g2270 ( 
.A1(n_2227),
.A2(n_2164),
.B1(n_2207),
.B2(n_2205),
.Y(n_2270)
);

BUFx3_ASAP7_75t_L g2271 ( 
.A(n_2233),
.Y(n_2271)
);

INVxp67_ASAP7_75t_L g2272 ( 
.A(n_2253),
.Y(n_2272)
);

OAI22xp33_ASAP7_75t_L g2273 ( 
.A1(n_2234),
.A2(n_2058),
.B1(n_2081),
.B2(n_2054),
.Y(n_2273)
);

AOI21xp5_ASAP7_75t_L g2274 ( 
.A1(n_2246),
.A2(n_2093),
.B(n_2104),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2258),
.Y(n_2275)
);

AOI22xp33_ASAP7_75t_L g2276 ( 
.A1(n_2226),
.A2(n_2229),
.B1(n_2230),
.B2(n_2255),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_2262),
.B(n_2216),
.Y(n_2277)
);

OAI22xp33_ASAP7_75t_L g2278 ( 
.A1(n_2261),
.A2(n_2058),
.B1(n_2081),
.B2(n_2054),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2260),
.Y(n_2279)
);

OAI22xp5_ASAP7_75t_L g2280 ( 
.A1(n_2253),
.A2(n_2093),
.B1(n_2129),
.B2(n_2117),
.Y(n_2280)
);

AND3x1_ASAP7_75t_L g2281 ( 
.A(n_2257),
.B(n_1964),
.C(n_1947),
.Y(n_2281)
);

OAI22xp33_ASAP7_75t_L g2282 ( 
.A1(n_2261),
.A2(n_2154),
.B1(n_2085),
.B2(n_2133),
.Y(n_2282)
);

AOI22xp5_ASAP7_75t_L g2283 ( 
.A1(n_2236),
.A2(n_2207),
.B1(n_2202),
.B2(n_2177),
.Y(n_2283)
);

OAI21xp33_ASAP7_75t_L g2284 ( 
.A1(n_2262),
.A2(n_2240),
.B(n_2241),
.Y(n_2284)
);

AOI22xp5_ASAP7_75t_L g2285 ( 
.A1(n_2243),
.A2(n_2202),
.B1(n_2219),
.B2(n_2217),
.Y(n_2285)
);

OA22x2_ASAP7_75t_L g2286 ( 
.A1(n_2233),
.A2(n_2086),
.B1(n_2152),
.B2(n_1974),
.Y(n_2286)
);

AOI21xp33_ASAP7_75t_SL g2287 ( 
.A1(n_2233),
.A2(n_1956),
.B(n_1964),
.Y(n_2287)
);

AOI22xp5_ASAP7_75t_SL g2288 ( 
.A1(n_2266),
.A2(n_1844),
.B1(n_1925),
.B2(n_1890),
.Y(n_2288)
);

AOI211xp5_ASAP7_75t_L g2289 ( 
.A1(n_2274),
.A2(n_2073),
.B(n_2178),
.C(n_2247),
.Y(n_2289)
);

OAI211xp5_ASAP7_75t_SL g2290 ( 
.A1(n_2276),
.A2(n_2247),
.B(n_2244),
.C(n_2259),
.Y(n_2290)
);

NAND3xp33_ASAP7_75t_L g2291 ( 
.A(n_2267),
.B(n_2263),
.C(n_2206),
.Y(n_2291)
);

XNOR2xp5_ASAP7_75t_L g2292 ( 
.A(n_2281),
.B(n_1844),
.Y(n_2292)
);

NOR2x1_ASAP7_75t_L g2293 ( 
.A(n_2264),
.B(n_2280),
.Y(n_2293)
);

AOI21xp5_ASAP7_75t_L g2294 ( 
.A1(n_2280),
.A2(n_2086),
.B(n_2182),
.Y(n_2294)
);

O2A1O1Ixp33_ASAP7_75t_L g2295 ( 
.A1(n_2272),
.A2(n_2141),
.B(n_2254),
.C(n_2251),
.Y(n_2295)
);

OAI21xp33_ASAP7_75t_L g2296 ( 
.A1(n_2268),
.A2(n_2228),
.B(n_2237),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2283),
.B(n_2228),
.Y(n_2297)
);

OAI21xp5_ASAP7_75t_L g2298 ( 
.A1(n_2286),
.A2(n_2287),
.B(n_2270),
.Y(n_2298)
);

NOR2xp33_ASAP7_75t_L g2299 ( 
.A(n_2271),
.B(n_2284),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2265),
.Y(n_2300)
);

AOI21xp5_ASAP7_75t_L g2301 ( 
.A1(n_2286),
.A2(n_2182),
.B(n_2160),
.Y(n_2301)
);

NOR2xp33_ASAP7_75t_L g2302 ( 
.A(n_2285),
.B(n_1796),
.Y(n_2302)
);

AOI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_2273),
.A2(n_2178),
.B1(n_2245),
.B2(n_2237),
.Y(n_2303)
);

AOI32xp33_ASAP7_75t_L g2304 ( 
.A1(n_2282),
.A2(n_2245),
.A3(n_2235),
.B1(n_2231),
.B2(n_2219),
.Y(n_2304)
);

OAI221xp5_ASAP7_75t_SL g2305 ( 
.A1(n_2278),
.A2(n_2063),
.B1(n_2155),
.B2(n_2231),
.C(n_2235),
.Y(n_2305)
);

OAI22xp5_ASAP7_75t_L g2306 ( 
.A1(n_2277),
.A2(n_2217),
.B1(n_2152),
.B2(n_2249),
.Y(n_2306)
);

O2A1O1Ixp33_ASAP7_75t_L g2307 ( 
.A1(n_2269),
.A2(n_1925),
.B(n_1932),
.C(n_1890),
.Y(n_2307)
);

AND2x4_ASAP7_75t_L g2308 ( 
.A(n_2275),
.B(n_2188),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_2279),
.B(n_2211),
.Y(n_2309)
);

OAI211xp5_ASAP7_75t_L g2310 ( 
.A1(n_2276),
.A2(n_1974),
.B(n_1932),
.C(n_2037),
.Y(n_2310)
);

CKINVDCx14_ASAP7_75t_R g2311 ( 
.A(n_2267),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2267),
.Y(n_2312)
);

NAND4xp25_ASAP7_75t_L g2313 ( 
.A(n_2276),
.B(n_2121),
.C(n_2107),
.D(n_1977),
.Y(n_2313)
);

OAI21xp33_ASAP7_75t_L g2314 ( 
.A1(n_2276),
.A2(n_2178),
.B(n_2155),
.Y(n_2314)
);

NOR2xp33_ASAP7_75t_L g2315 ( 
.A(n_2311),
.B(n_1667),
.Y(n_2315)
);

AOI21xp5_ASAP7_75t_SL g2316 ( 
.A1(n_2292),
.A2(n_1996),
.B(n_2003),
.Y(n_2316)
);

OAI21xp5_ASAP7_75t_SL g2317 ( 
.A1(n_2293),
.A2(n_2041),
.B(n_1966),
.Y(n_2317)
);

AOI222xp33_ASAP7_75t_L g2318 ( 
.A1(n_2314),
.A2(n_2120),
.B1(n_2109),
.B2(n_2099),
.C1(n_2101),
.C2(n_2122),
.Y(n_2318)
);

AOI221xp5_ASAP7_75t_L g2319 ( 
.A1(n_2289),
.A2(n_2214),
.B1(n_2220),
.B2(n_2213),
.C(n_2212),
.Y(n_2319)
);

NOR3xp33_ASAP7_75t_L g2320 ( 
.A(n_2310),
.B(n_1667),
.C(n_1916),
.Y(n_2320)
);

AND4x1_ASAP7_75t_L g2321 ( 
.A(n_2302),
.B(n_1676),
.C(n_2043),
.D(n_1962),
.Y(n_2321)
);

NOR4xp25_ASAP7_75t_L g2322 ( 
.A(n_2307),
.B(n_1942),
.C(n_1957),
.D(n_2102),
.Y(n_2322)
);

NAND4xp25_ASAP7_75t_SL g2323 ( 
.A(n_2298),
.B(n_2160),
.C(n_2079),
.D(n_2249),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2312),
.Y(n_2324)
);

A2O1A1Ixp33_ASAP7_75t_L g2325 ( 
.A1(n_2288),
.A2(n_1996),
.B(n_2041),
.C(n_1966),
.Y(n_2325)
);

OAI21xp33_ASAP7_75t_SL g2326 ( 
.A1(n_2304),
.A2(n_2133),
.B(n_2238),
.Y(n_2326)
);

NOR4xp25_ASAP7_75t_L g2327 ( 
.A(n_2305),
.B(n_2103),
.C(n_2108),
.D(n_2106),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2309),
.Y(n_2328)
);

AOI22xp5_ASAP7_75t_L g2329 ( 
.A1(n_2313),
.A2(n_2221),
.B1(n_2206),
.B2(n_2208),
.Y(n_2329)
);

AOI21xp5_ASAP7_75t_L g2330 ( 
.A1(n_2294),
.A2(n_2299),
.B(n_2296),
.Y(n_2330)
);

NAND4xp75_ASAP7_75t_L g2331 ( 
.A(n_2303),
.B(n_2048),
.C(n_2038),
.D(n_2107),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_2295),
.B(n_2203),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2301),
.B(n_2208),
.Y(n_2333)
);

OAI211xp5_ASAP7_75t_L g2334 ( 
.A1(n_2317),
.A2(n_2290),
.B(n_2297),
.C(n_2291),
.Y(n_2334)
);

NAND4xp25_ASAP7_75t_L g2335 ( 
.A(n_2330),
.B(n_2306),
.C(n_2300),
.D(n_2001),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_2322),
.B(n_2308),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2324),
.Y(n_2337)
);

NOR3x1_ASAP7_75t_L g2338 ( 
.A(n_2331),
.B(n_2030),
.C(n_2011),
.Y(n_2338)
);

AOI22xp5_ASAP7_75t_L g2339 ( 
.A1(n_2320),
.A2(n_2308),
.B1(n_2250),
.B2(n_2152),
.Y(n_2339)
);

NOR2x1_ASAP7_75t_L g2340 ( 
.A(n_2315),
.B(n_2001),
.Y(n_2340)
);

NOR3xp33_ASAP7_75t_L g2341 ( 
.A(n_2323),
.B(n_1917),
.C(n_2017),
.Y(n_2341)
);

NOR3xp33_ASAP7_75t_L g2342 ( 
.A(n_2320),
.B(n_2017),
.C(n_1854),
.Y(n_2342)
);

NAND4xp25_ASAP7_75t_L g2343 ( 
.A(n_2325),
.B(n_2316),
.C(n_2318),
.D(n_2329),
.Y(n_2343)
);

NAND4xp25_ASAP7_75t_SL g2344 ( 
.A(n_2326),
.B(n_2238),
.C(n_2242),
.D(n_2250),
.Y(n_2344)
);

NOR2x1_ASAP7_75t_L g2345 ( 
.A(n_2328),
.B(n_2046),
.Y(n_2345)
);

NOR3x1_ASAP7_75t_L g2346 ( 
.A(n_2332),
.B(n_2333),
.C(n_2321),
.Y(n_2346)
);

INVx1_ASAP7_75t_SL g2347 ( 
.A(n_2327),
.Y(n_2347)
);

OAI221xp5_ASAP7_75t_L g2348 ( 
.A1(n_2319),
.A2(n_2003),
.B1(n_2154),
.B2(n_2222),
.C(n_2242),
.Y(n_2348)
);

NOR3xp33_ASAP7_75t_L g2349 ( 
.A(n_2317),
.B(n_1854),
.C(n_1833),
.Y(n_2349)
);

NOR3xp33_ASAP7_75t_L g2350 ( 
.A(n_2343),
.B(n_1859),
.C(n_1855),
.Y(n_2350)
);

AND2x2_ASAP7_75t_SL g2351 ( 
.A(n_2338),
.B(n_1849),
.Y(n_2351)
);

NOR2xp33_ASAP7_75t_L g2352 ( 
.A(n_2347),
.B(n_2112),
.Y(n_2352)
);

NAND4xp75_ASAP7_75t_L g2353 ( 
.A(n_2346),
.B(n_2033),
.C(n_2111),
.D(n_2050),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2337),
.Y(n_2354)
);

INVx2_ASAP7_75t_SL g2355 ( 
.A(n_2340),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2336),
.Y(n_2356)
);

NOR2xp33_ASAP7_75t_L g2357 ( 
.A(n_2335),
.B(n_2113),
.Y(n_2357)
);

NOR3xp33_ASAP7_75t_L g2358 ( 
.A(n_2334),
.B(n_1859),
.C(n_1855),
.Y(n_2358)
);

INVx5_ASAP7_75t_L g2359 ( 
.A(n_2345),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2341),
.Y(n_2360)
);

AOI21xp5_ASAP7_75t_L g2361 ( 
.A1(n_2344),
.A2(n_2222),
.B(n_2126),
.Y(n_2361)
);

NOR3xp33_ASAP7_75t_L g2362 ( 
.A(n_2342),
.B(n_1899),
.C(n_1896),
.Y(n_2362)
);

AND3x4_ASAP7_75t_L g2363 ( 
.A(n_2350),
.B(n_2349),
.C(n_2348),
.Y(n_2363)
);

AND2x2_ASAP7_75t_L g2364 ( 
.A(n_2355),
.B(n_2339),
.Y(n_2364)
);

NOR3xp33_ASAP7_75t_L g2365 ( 
.A(n_2356),
.B(n_2116),
.C(n_1675),
.Y(n_2365)
);

BUFx3_ASAP7_75t_L g2366 ( 
.A(n_2354),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2359),
.Y(n_2367)
);

NAND4xp75_ASAP7_75t_L g2368 ( 
.A(n_2360),
.B(n_2125),
.C(n_1939),
.D(n_2118),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_2359),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2352),
.Y(n_2370)
);

NAND3x1_ASAP7_75t_L g2371 ( 
.A(n_2357),
.B(n_2154),
.C(n_1899),
.Y(n_2371)
);

XOR2xp5_ASAP7_75t_L g2372 ( 
.A(n_2353),
.B(n_1929),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_2351),
.B(n_2145),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_2367),
.B(n_2369),
.Y(n_2374)
);

AND2x4_ASAP7_75t_L g2375 ( 
.A(n_2366),
.B(n_2359),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_2364),
.B(n_2358),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2370),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_2368),
.Y(n_2378)
);

NOR2xp33_ASAP7_75t_L g2379 ( 
.A(n_2370),
.B(n_2361),
.Y(n_2379)
);

AOI22xp5_ASAP7_75t_L g2380 ( 
.A1(n_2363),
.A2(n_2362),
.B1(n_1852),
.B2(n_1892),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2372),
.Y(n_2381)
);

AND2x4_ASAP7_75t_L g2382 ( 
.A(n_2365),
.B(n_2131),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_2373),
.Y(n_2383)
);

AND2x2_ASAP7_75t_L g2384 ( 
.A(n_2365),
.B(n_2363),
.Y(n_2384)
);

INVx1_ASAP7_75t_SL g2385 ( 
.A(n_2374),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2377),
.Y(n_2386)
);

OAI22xp33_ASAP7_75t_L g2387 ( 
.A1(n_2380),
.A2(n_2371),
.B1(n_1852),
.B2(n_1892),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2375),
.B(n_1948),
.Y(n_2388)
);

NOR2xp33_ASAP7_75t_L g2389 ( 
.A(n_2375),
.B(n_1852),
.Y(n_2389)
);

AOI22x1_ASAP7_75t_L g2390 ( 
.A1(n_2381),
.A2(n_1896),
.B1(n_2154),
.B2(n_1675),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2385),
.Y(n_2391)
);

AO22x1_ASAP7_75t_L g2392 ( 
.A1(n_2389),
.A2(n_2384),
.B1(n_2377),
.B2(n_2378),
.Y(n_2392)
);

INVx1_ASAP7_75t_SL g2393 ( 
.A(n_2386),
.Y(n_2393)
);

OAI31xp33_ASAP7_75t_SL g2394 ( 
.A1(n_2390),
.A2(n_2379),
.A3(n_2376),
.B(n_2383),
.Y(n_2394)
);

XNOR2xp5_ASAP7_75t_L g2395 ( 
.A(n_2388),
.B(n_2382),
.Y(n_2395)
);

INVx2_ASAP7_75t_SL g2396 ( 
.A(n_2387),
.Y(n_2396)
);

INVxp67_ASAP7_75t_L g2397 ( 
.A(n_2391),
.Y(n_2397)
);

INVxp67_ASAP7_75t_L g2398 ( 
.A(n_2396),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2395),
.Y(n_2399)
);

OAI22x1_ASAP7_75t_SL g2400 ( 
.A1(n_2399),
.A2(n_2393),
.B1(n_2392),
.B2(n_2394),
.Y(n_2400)
);

OAI22xp5_ASAP7_75t_L g2401 ( 
.A1(n_2398),
.A2(n_2382),
.B1(n_1872),
.B2(n_1901),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2400),
.Y(n_2402)
);

AOI21xp5_ASAP7_75t_L g2403 ( 
.A1(n_2402),
.A2(n_2397),
.B(n_2401),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2403),
.Y(n_2404)
);

AOI22xp33_ASAP7_75t_L g2405 ( 
.A1(n_2404),
.A2(n_1872),
.B1(n_1901),
.B2(n_1892),
.Y(n_2405)
);


endmodule