module fake_jpeg_17813_n_250 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_250);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_7),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_40),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_14),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_25),
.B1(n_19),
.B2(n_18),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_41),
.A2(n_15),
.B1(n_17),
.B2(n_24),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_25),
.Y(n_48)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_18),
.B1(n_27),
.B2(n_26),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_35),
.B1(n_33),
.B2(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_23),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_53),
.B(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_23),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_35),
.A2(n_18),
.B1(n_27),
.B2(n_26),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_23),
.B1(n_17),
.B2(n_15),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_38),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_33),
.B1(n_17),
.B2(n_15),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_31),
.C(n_32),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_82),
.C(n_54),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_35),
.B1(n_39),
.B2(n_36),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_63),
.A2(n_66),
.B1(n_44),
.B2(n_39),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_64),
.A2(n_76),
.B1(n_85),
.B2(n_49),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

AO22x2_ASAP7_75t_L g66 ( 
.A1(n_41),
.A2(n_26),
.B1(n_36),
.B2(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_53),
.B1(n_22),
.B2(n_20),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_78),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_42),
.B1(n_58),
.B2(n_57),
.Y(n_86)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_69),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_51),
.A2(n_24),
.B1(n_16),
.B2(n_29),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_42),
.A2(n_28),
.B(n_29),
.C(n_24),
.Y(n_80)
);

NAND3xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_13),
.C(n_12),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_45),
.A2(n_31),
.B(n_32),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_60),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_16),
.B1(n_28),
.B2(n_22),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_86),
.A2(n_88),
.B1(n_90),
.B2(n_95),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_87),
.A2(n_89),
.B1(n_91),
.B2(n_93),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_55),
.B1(n_49),
.B2(n_44),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_61),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_68),
.A2(n_13),
.B1(n_11),
.B2(n_9),
.Y(n_95)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_97),
.B(n_104),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_66),
.A2(n_60),
.B1(n_56),
.B2(n_52),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_98),
.A2(n_105),
.B1(n_106),
.B2(n_65),
.Y(n_127)
);

AOI32xp33_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_54),
.A3(n_31),
.B1(n_32),
.B2(n_46),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_101),
.Y(n_116)
);

BUFx4f_ASAP7_75t_SL g103 ( 
.A(n_70),
.Y(n_103)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_68),
.B(n_20),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_66),
.A2(n_9),
.B1(n_6),
.B2(n_12),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_66),
.A2(n_8),
.B1(n_6),
.B2(n_30),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_84),
.Y(n_107)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_62),
.A2(n_56),
.B1(n_52),
.B2(n_20),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_108),
.A2(n_77),
.B1(n_79),
.B2(n_71),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_109),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_56),
.B1(n_52),
.B2(n_30),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_54),
.B1(n_8),
.B2(n_2),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_108),
.C(n_104),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_93),
.C(n_103),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_80),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_115),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_75),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_73),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_128),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_121),
.B(n_0),
.Y(n_155)
);

OR2x2_ASAP7_75t_SL g122 ( 
.A(n_100),
.B(n_72),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_122),
.A2(n_127),
.B1(n_109),
.B2(n_1),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_70),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_98),
.A2(n_71),
.B1(n_67),
.B2(n_74),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_132),
.B1(n_117),
.B2(n_126),
.Y(n_139)
);

OAI32xp33_ASAP7_75t_L g128 ( 
.A1(n_87),
.A2(n_63),
.A3(n_30),
.B1(n_65),
.B2(n_78),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_77),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_130),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_87),
.A2(n_54),
.B(n_21),
.C(n_2),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_131),
.A2(n_21),
.B1(n_103),
.B2(n_2),
.Y(n_148)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_86),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_144),
.C(n_116),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_91),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_141),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_140),
.B1(n_149),
.B2(n_0),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_126),
.A2(n_110),
.B1(n_92),
.B2(n_99),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_103),
.Y(n_141)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_114),
.B(n_102),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_111),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_148),
.A2(n_153),
.B(n_155),
.Y(n_158)
);

OA22x2_ASAP7_75t_L g149 ( 
.A1(n_128),
.A2(n_109),
.B1(n_21),
.B2(n_2),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_151),
.A2(n_132),
.B1(n_131),
.B2(n_127),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_115),
.B(n_0),
.Y(n_152)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

NOR2x1_ASAP7_75t_R g153 ( 
.A(n_122),
.B(n_0),
.Y(n_153)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_154),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_159),
.B(n_163),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_113),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_162),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_123),
.C(n_121),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_123),
.C(n_129),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_1),
.B(n_4),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_165),
.A2(n_167),
.B1(n_169),
.B2(n_170),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_153),
.A2(n_120),
.B1(n_125),
.B2(n_119),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_119),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_175),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_135),
.A2(n_137),
.B1(n_151),
.B2(n_139),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_134),
.A2(n_112),
.B1(n_3),
.B2(n_4),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_171),
.A2(n_172),
.B1(n_154),
.B2(n_148),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_134),
.A2(n_112),
.B1(n_3),
.B2(n_4),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_145),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_173),
.B(n_145),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_112),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_176),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_170),
.A2(n_155),
.B1(n_141),
.B2(n_138),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_179),
.A2(n_181),
.B1(n_182),
.B2(n_188),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_180),
.B(n_189),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_161),
.A2(n_138),
.B1(n_149),
.B2(n_150),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_147),
.B1(n_153),
.B2(n_149),
.Y(n_182)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_161),
.A2(n_142),
.B1(n_143),
.B2(n_146),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_186),
.Y(n_198)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_187),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_163),
.A2(n_149),
.B1(n_142),
.B2(n_154),
.Y(n_188)
);

AO22x2_ASAP7_75t_L g190 ( 
.A1(n_164),
.A2(n_149),
.B1(n_152),
.B2(n_5),
.Y(n_190)
);

AOI21x1_ASAP7_75t_SL g196 ( 
.A1(n_190),
.A2(n_158),
.B(n_172),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_171),
.Y(n_203)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_192),
.Y(n_194)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_190),
.Y(n_197)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_197),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_178),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_201),
.C(n_205),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_160),
.Y(n_201)
);

AOI21x1_ASAP7_75t_SL g202 ( 
.A1(n_190),
.A2(n_175),
.B(n_165),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_202),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_177),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_159),
.C(n_168),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_202),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_216),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_209),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_206),
.B(n_184),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_214),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_205),
.B(n_184),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_217),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_201),
.C(n_199),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_188),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_207),
.A2(n_180),
.B(n_198),
.Y(n_218)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_218),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_195),
.C(n_181),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_179),
.C(n_182),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_212),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_226),
.Y(n_228)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_211),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_222),
.A2(n_194),
.B1(n_196),
.B2(n_190),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_204),
.Y(n_226)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_227),
.Y(n_237)
);

OAI21x1_ASAP7_75t_L g229 ( 
.A1(n_219),
.A2(n_210),
.B(n_203),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_223),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_209),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_232),
.C(n_233),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_157),
.C(n_194),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_221),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_235),
.B(n_236),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_231),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_238),
.A2(n_224),
.B(n_232),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_239),
.A2(n_240),
.B(n_241),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_236),
.A2(n_233),
.B1(n_225),
.B2(n_191),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_167),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_L g243 ( 
.A(n_242),
.B(n_237),
.C(n_174),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_243),
.A2(n_245),
.B(n_1),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_239),
.A2(n_158),
.B(n_4),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_1),
.C(n_5),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_247),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_5),
.Y(n_249)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_249),
.Y(n_250)
);


endmodule