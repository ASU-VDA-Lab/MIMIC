module fake_netlist_1_4158_n_559 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_559);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_559;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_357;
wire n_90;
wire n_245;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_445;
wire n_398;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_15), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_21), .Y(n_80) );
BUFx6f_ASAP7_75t_L g81 ( .A(n_23), .Y(n_81) );
BUFx10_ASAP7_75t_L g82 ( .A(n_70), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_19), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_78), .Y(n_84) );
BUFx2_ASAP7_75t_L g85 ( .A(n_18), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_25), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_29), .Y(n_87) );
NOR2xp33_ASAP7_75t_L g88 ( .A(n_35), .B(n_48), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_54), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_56), .Y(n_90) );
BUFx2_ASAP7_75t_L g91 ( .A(n_30), .Y(n_91) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_6), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_67), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_27), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_1), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_57), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_77), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_72), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_41), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_17), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_6), .Y(n_101) );
BUFx3_ASAP7_75t_L g102 ( .A(n_58), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_52), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_16), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_38), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_24), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_37), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_71), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g109 ( .A(n_33), .B(n_5), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_53), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_13), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_46), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_59), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_17), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_9), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_75), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_4), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_85), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_94), .Y(n_120) );
INVx6_ASAP7_75t_L g121 ( .A(n_82), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_85), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_94), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_81), .Y(n_124) );
NAND2xp33_ASAP7_75t_L g125 ( .A(n_86), .B(n_76), .Y(n_125) );
INVx4_ASAP7_75t_L g126 ( .A(n_91), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_103), .Y(n_127) );
AND2x6_ASAP7_75t_L g128 ( .A(n_102), .B(n_36), .Y(n_128) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_79), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_81), .Y(n_130) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_79), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_87), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_87), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_81), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_91), .B(n_0), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_103), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_101), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_81), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_95), .B(n_3), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_95), .B(n_3), .Y(n_140) );
OAI22x1_ASAP7_75t_R g141 ( .A1(n_118), .A2(n_4), .B1(n_5), .B2(n_7), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_120), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_124), .Y(n_143) );
NAND3xp33_ASAP7_75t_L g144 ( .A(n_126), .B(n_111), .C(n_100), .Y(n_144) );
NOR3xp33_ASAP7_75t_L g145 ( .A(n_129), .B(n_104), .C(n_116), .Y(n_145) );
NAND3xp33_ASAP7_75t_L g146 ( .A(n_126), .B(n_112), .C(n_115), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_126), .B(n_82), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_126), .B(n_80), .Y(n_148) );
AOI22xp33_ASAP7_75t_L g149 ( .A1(n_132), .A2(n_118), .B1(n_101), .B2(n_92), .Y(n_149) );
OAI21xp33_ASAP7_75t_SL g150 ( .A1(n_132), .A2(n_99), .B(n_90), .Y(n_150) );
OR2x6_ASAP7_75t_L g151 ( .A(n_129), .B(n_92), .Y(n_151) );
AOI22xp33_ASAP7_75t_L g152 ( .A1(n_133), .A2(n_92), .B1(n_99), .B2(n_90), .Y(n_152) );
NAND2xp33_ASAP7_75t_L g153 ( .A(n_128), .B(n_97), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_119), .B(n_82), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_124), .Y(n_155) );
BUFx3_ASAP7_75t_L g156 ( .A(n_128), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_120), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_123), .Y(n_158) );
INVx4_ASAP7_75t_L g159 ( .A(n_128), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_124), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_121), .B(n_98), .Y(n_161) );
OAI22xp5_ASAP7_75t_L g162 ( .A1(n_119), .A2(n_98), .B1(n_89), .B2(n_97), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_124), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_124), .Y(n_164) );
INVx1_ASAP7_75t_SL g165 ( .A(n_131), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_130), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_122), .Y(n_167) );
AOI22xp33_ASAP7_75t_L g168 ( .A1(n_144), .A2(n_128), .B1(n_133), .B2(n_135), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_142), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_142), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_153), .A2(n_125), .B(n_123), .Y(n_171) );
NOR2xp33_ASAP7_75t_SL g172 ( .A(n_159), .B(n_128), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_159), .B(n_122), .Y(n_173) );
BUFx3_ASAP7_75t_L g174 ( .A(n_156), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_159), .A2(n_127), .B(n_136), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_157), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_157), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_L g178 ( .A1(n_150), .A2(n_140), .B(n_139), .C(n_127), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_158), .Y(n_179) );
INVxp67_ASAP7_75t_SL g180 ( .A(n_156), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_147), .B(n_121), .Y(n_181) );
BUFx12f_ASAP7_75t_L g182 ( .A(n_167), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_147), .B(n_121), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_150), .A2(n_128), .B1(n_121), .B2(n_136), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_154), .B(n_86), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_159), .B(n_106), .Y(n_186) );
INVxp67_ASAP7_75t_SL g187 ( .A(n_156), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_161), .B(n_110), .Y(n_188) );
AND2x2_ASAP7_75t_SL g189 ( .A(n_145), .B(n_117), .Y(n_189) );
INVx2_ASAP7_75t_SL g190 ( .A(n_161), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_148), .B(n_110), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_146), .B(n_106), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_165), .B(n_89), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_162), .B(n_152), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_158), .B(n_128), .Y(n_195) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_149), .A2(n_137), .B(n_83), .C(n_107), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_143), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_143), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_151), .B(n_137), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_143), .Y(n_200) );
NOR2xp33_ASAP7_75t_R g201 ( .A(n_151), .B(n_137), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_184), .A2(n_151), .B1(n_92), .B2(n_84), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_193), .B(n_190), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_190), .B(n_151), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_170), .Y(n_205) );
OAI22xp5_ASAP7_75t_L g206 ( .A1(n_184), .A2(n_151), .B1(n_92), .B2(n_93), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_170), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_170), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_172), .A2(n_114), .B(n_96), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_172), .B(n_108), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_188), .B(n_113), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g212 ( .A1(n_189), .A2(n_109), .B1(n_105), .B2(n_117), .Y(n_212) );
OAI21xp33_ASAP7_75t_L g213 ( .A1(n_201), .A2(n_102), .B(n_88), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_199), .B(n_7), .Y(n_214) );
INVx4_ASAP7_75t_L g215 ( .A(n_179), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_195), .A2(n_166), .B(n_164), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_175), .A2(n_166), .B(n_164), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_181), .A2(n_166), .B(n_164), .Y(n_218) );
INVx3_ASAP7_75t_L g219 ( .A(n_179), .Y(n_219) );
OAI22xp5_ASAP7_75t_SL g220 ( .A1(n_182), .A2(n_141), .B1(n_81), .B2(n_10), .Y(n_220) );
OAI21xp33_ASAP7_75t_L g221 ( .A1(n_191), .A2(n_141), .B(n_138), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_179), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_183), .A2(n_163), .B(n_160), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_174), .B(n_138), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_174), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_171), .A2(n_173), .B(n_186), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_169), .B(n_8), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_169), .B(n_8), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_176), .B(n_9), .Y(n_229) );
INVx2_ASAP7_75t_SL g230 ( .A(n_182), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_174), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_189), .A2(n_138), .B1(n_134), .B2(n_130), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_178), .A2(n_163), .B(n_160), .C(n_155), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g234 ( .A1(n_176), .A2(n_138), .B1(n_134), .B2(n_130), .Y(n_234) );
AO22x1_ASAP7_75t_L g235 ( .A1(n_185), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_226), .A2(n_194), .B(n_187), .Y(n_236) );
OAI21xp5_ASAP7_75t_L g237 ( .A1(n_233), .A2(n_177), .B(n_168), .Y(n_237) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_215), .Y(n_238) );
CKINVDCx6p67_ASAP7_75t_R g239 ( .A(n_215), .Y(n_239) );
OAI21x1_ASAP7_75t_L g240 ( .A1(n_216), .A2(n_177), .B(n_198), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_217), .A2(n_180), .B(n_196), .Y(n_241) );
AO31x2_ASAP7_75t_L g242 ( .A1(n_202), .A2(n_200), .A3(n_197), .B(n_198), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_207), .B(n_222), .Y(n_243) );
OA21x2_ASAP7_75t_L g244 ( .A1(n_218), .A2(n_200), .B(n_197), .Y(n_244) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_225), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_204), .B(n_189), .Y(n_246) );
BUFx2_ASAP7_75t_L g247 ( .A(n_230), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_221), .B(n_192), .Y(n_248) );
OAI21x1_ASAP7_75t_L g249 ( .A1(n_223), .A2(n_198), .B(n_163), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_227), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_203), .B(n_11), .Y(n_251) );
OAI21xp5_ASAP7_75t_L g252 ( .A1(n_205), .A2(n_160), .B(n_155), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_219), .B(n_12), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_211), .A2(n_155), .B(n_138), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_209), .A2(n_134), .B(n_130), .Y(n_255) );
AOI221xp5_ASAP7_75t_L g256 ( .A1(n_220), .A2(n_134), .B1(n_130), .B2(n_15), .C(n_16), .Y(n_256) );
AO31x2_ASAP7_75t_L g257 ( .A1(n_202), .A2(n_134), .A3(n_14), .B(n_13), .Y(n_257) );
OAI21x1_ASAP7_75t_L g258 ( .A1(n_219), .A2(n_49), .B(n_20), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_210), .A2(n_50), .B(n_22), .Y(n_259) );
OR2x2_ASAP7_75t_L g260 ( .A(n_227), .B(n_14), .Y(n_260) );
AO31x2_ASAP7_75t_L g261 ( .A1(n_206), .A2(n_26), .A3(n_28), .B(n_31), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_208), .A2(n_32), .B(n_34), .Y(n_262) );
OAI21xp33_ASAP7_75t_L g263 ( .A1(n_206), .A2(n_39), .B(n_40), .Y(n_263) );
AOI21xp33_ASAP7_75t_L g264 ( .A1(n_260), .A2(n_228), .B(n_229), .Y(n_264) );
AO31x2_ASAP7_75t_L g265 ( .A1(n_236), .A2(n_234), .A3(n_214), .B(n_235), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_247), .B(n_212), .Y(n_266) );
OA21x2_ASAP7_75t_L g267 ( .A1(n_249), .A2(n_232), .B(n_213), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_250), .B(n_231), .Y(n_268) );
INVx2_ASAP7_75t_SL g269 ( .A(n_239), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_243), .A2(n_224), .B(n_234), .Y(n_270) );
AOI21xp33_ASAP7_75t_L g271 ( .A1(n_248), .A2(n_231), .B(n_225), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_243), .A2(n_231), .B1(n_225), .B2(n_44), .Y(n_272) );
INVx3_ASAP7_75t_L g273 ( .A(n_238), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_238), .B(n_42), .Y(n_274) );
OAI21xp5_ASAP7_75t_L g275 ( .A1(n_237), .A2(n_43), .B(n_45), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_244), .Y(n_276) );
AOI22x1_ASAP7_75t_L g277 ( .A1(n_255), .A2(n_47), .B1(n_51), .B2(n_55), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_244), .Y(n_278) );
OAI21x1_ASAP7_75t_SL g279 ( .A1(n_253), .A2(n_60), .B(n_61), .Y(n_279) );
OAI21x1_ASAP7_75t_L g280 ( .A1(n_258), .A2(n_62), .B(n_63), .Y(n_280) );
OR2x6_ASAP7_75t_L g281 ( .A(n_238), .B(n_64), .Y(n_281) );
AO21x2_ASAP7_75t_L g282 ( .A1(n_237), .A2(n_65), .B(n_66), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_254), .A2(n_68), .B(n_69), .Y(n_283) );
AO21x2_ASAP7_75t_L g284 ( .A1(n_241), .A2(n_73), .B(n_74), .Y(n_284) );
AO21x2_ASAP7_75t_L g285 ( .A1(n_241), .A2(n_254), .B(n_263), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_246), .B(n_251), .Y(n_286) );
AO31x2_ASAP7_75t_L g287 ( .A1(n_253), .A2(n_246), .A3(n_255), .B(n_262), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_276), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_276), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_286), .B(n_242), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_276), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_286), .B(n_257), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_278), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_278), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_278), .Y(n_295) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_269), .Y(n_296) );
BUFx3_ASAP7_75t_L g297 ( .A(n_269), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_273), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_285), .Y(n_299) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_273), .Y(n_300) );
INVx2_ASAP7_75t_SL g301 ( .A(n_273), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_268), .B(n_242), .Y(n_302) );
BUFx2_ASAP7_75t_L g303 ( .A(n_281), .Y(n_303) );
AO21x1_ASAP7_75t_SL g304 ( .A1(n_275), .A2(n_252), .B(n_261), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_268), .Y(n_305) );
INVx2_ASAP7_75t_SL g306 ( .A(n_273), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_274), .B(n_257), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_279), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_266), .B(n_242), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_279), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_292), .B(n_257), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_292), .B(n_271), .Y(n_312) );
BUFx2_ASAP7_75t_L g313 ( .A(n_303), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_289), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_307), .B(n_261), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_288), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_288), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_289), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_288), .Y(n_319) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_291), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_307), .B(n_261), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_293), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_291), .B(n_284), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_294), .B(n_284), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_294), .B(n_284), .Y(n_325) );
AO21x2_ASAP7_75t_L g326 ( .A1(n_299), .A2(n_285), .B(n_275), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_309), .B(n_284), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_309), .B(n_274), .Y(n_328) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_297), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_293), .Y(n_330) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_293), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_296), .B(n_256), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_295), .B(n_285), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_295), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_295), .B(n_285), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_290), .B(n_305), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_290), .B(n_271), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_299), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_303), .B(n_281), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_302), .Y(n_340) );
NOR2xp67_ASAP7_75t_L g341 ( .A(n_320), .B(n_310), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_314), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_311), .B(n_302), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_340), .B(n_305), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_338), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_311), .B(n_299), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_331), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_340), .B(n_297), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_315), .B(n_310), .Y(n_349) );
INVxp67_ASAP7_75t_L g350 ( .A(n_329), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_315), .B(n_308), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_314), .Y(n_352) );
INVx2_ASAP7_75t_SL g353 ( .A(n_320), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_336), .B(n_297), .Y(n_354) );
AND2x4_ASAP7_75t_L g355 ( .A(n_339), .B(n_308), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_318), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_318), .Y(n_357) );
AND2x4_ASAP7_75t_L g358 ( .A(n_339), .B(n_306), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_312), .B(n_300), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_336), .B(n_332), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_330), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_321), .B(n_304), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_339), .B(n_321), .Y(n_363) );
AND2x4_ASAP7_75t_L g364 ( .A(n_339), .B(n_306), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_331), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_328), .B(n_304), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_328), .B(n_306), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_333), .B(n_301), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_338), .Y(n_369) );
BUFx2_ASAP7_75t_SL g370 ( .A(n_316), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_312), .B(n_298), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_330), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_337), .B(n_301), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_316), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_337), .B(n_301), .Y(n_375) );
BUFx3_ASAP7_75t_L g376 ( .A(n_316), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_327), .A2(n_256), .B1(n_264), .B2(n_281), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_327), .B(n_287), .Y(n_378) );
AND2x4_ASAP7_75t_L g379 ( .A(n_333), .B(n_281), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_317), .B(n_287), .Y(n_380) );
INVx2_ASAP7_75t_SL g381 ( .A(n_317), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_317), .B(n_264), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_338), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_319), .B(n_265), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_342), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_343), .B(n_324), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_343), .B(n_324), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_342), .Y(n_388) );
NAND3xp33_ASAP7_75t_L g389 ( .A(n_350), .B(n_313), .C(n_323), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_360), .B(n_323), .Y(n_390) );
INVx1_ASAP7_75t_SL g391 ( .A(n_354), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_378), .B(n_325), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_352), .B(n_325), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_366), .A2(n_313), .B1(n_281), .B2(n_282), .Y(n_394) );
AOI21xp33_ASAP7_75t_L g395 ( .A1(n_382), .A2(n_335), .B(n_326), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_352), .B(n_334), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_378), .B(n_335), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_346), .B(n_334), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_356), .B(n_322), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_346), .B(n_334), .Y(n_400) );
OR2x6_ASAP7_75t_L g401 ( .A(n_370), .B(n_322), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_356), .B(n_322), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_349), .B(n_319), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_357), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_357), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_349), .B(n_351), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_359), .B(n_319), .Y(n_407) );
OAI21xp33_ASAP7_75t_L g408 ( .A1(n_362), .A2(n_272), .B(n_283), .Y(n_408) );
INVx3_ASAP7_75t_L g409 ( .A(n_376), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_345), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_351), .B(n_326), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_345), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_361), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_362), .B(n_326), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_359), .B(n_326), .Y(n_415) );
INVxp67_ASAP7_75t_SL g416 ( .A(n_353), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_344), .B(n_265), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_361), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_372), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_371), .B(n_353), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_363), .B(n_265), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_371), .B(n_265), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_363), .B(n_265), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_372), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_383), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_383), .Y(n_426) );
NOR2xp67_ASAP7_75t_L g427 ( .A(n_341), .B(n_272), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_373), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_363), .B(n_265), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_373), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_363), .B(n_287), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_366), .B(n_287), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_347), .Y(n_433) );
AND2x4_ASAP7_75t_L g434 ( .A(n_355), .B(n_282), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_345), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_375), .B(n_287), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_367), .B(n_287), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_428), .B(n_380), .Y(n_438) );
BUFx2_ASAP7_75t_L g439 ( .A(n_416), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_406), .B(n_368), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_397), .B(n_347), .Y(n_441) );
BUFx2_ASAP7_75t_L g442 ( .A(n_401), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_420), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_430), .B(n_380), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_420), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_406), .B(n_368), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_404), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_414), .B(n_368), .Y(n_448) );
INVxp67_ASAP7_75t_L g449 ( .A(n_433), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_410), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_390), .B(n_367), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_404), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_397), .B(n_365), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_392), .B(n_365), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_405), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_414), .B(n_368), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_392), .B(n_379), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_405), .Y(n_458) );
NAND4xp25_ASAP7_75t_L g459 ( .A(n_394), .B(n_377), .C(n_348), .D(n_341), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_410), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_419), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_391), .B(n_355), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_431), .B(n_411), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_419), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_424), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_424), .Y(n_466) );
INVx1_ASAP7_75t_SL g467 ( .A(n_407), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_385), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_388), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_413), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_386), .B(n_355), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_386), .B(n_381), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_387), .B(n_381), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_418), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_403), .Y(n_475) );
AO21x1_ASAP7_75t_SL g476 ( .A1(n_407), .A2(n_370), .B(n_384), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_387), .B(n_355), .Y(n_477) );
NAND4xp25_ASAP7_75t_L g478 ( .A(n_408), .B(n_379), .C(n_358), .D(n_364), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_431), .B(n_379), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_393), .B(n_364), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_403), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_412), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_437), .B(n_376), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_463), .B(n_411), .Y(n_484) );
AOI221xp5_ASAP7_75t_L g485 ( .A1(n_478), .A2(n_395), .B1(n_432), .B2(n_421), .C(n_423), .Y(n_485) );
AOI222xp33_ASAP7_75t_L g486 ( .A1(n_443), .A2(n_432), .B1(n_421), .B2(n_423), .C1(n_429), .C2(n_437), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_442), .A2(n_401), .B(n_389), .Y(n_487) );
NOR4xp25_ASAP7_75t_SL g488 ( .A(n_439), .B(n_426), .C(n_425), .D(n_435), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_447), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_463), .B(n_436), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_449), .B(n_409), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_445), .B(n_415), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_SL g493 ( .A1(n_467), .A2(n_422), .B(n_409), .C(n_415), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_471), .B(n_409), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_462), .B(n_427), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_475), .B(n_481), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_480), .B(n_429), .Y(n_497) );
INVx1_ASAP7_75t_SL g498 ( .A(n_473), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_480), .B(n_398), .Y(n_499) );
NOR3xp33_ASAP7_75t_L g500 ( .A(n_459), .B(n_417), .C(n_422), .Y(n_500) );
INVxp67_ASAP7_75t_L g501 ( .A(n_462), .Y(n_501) );
AOI221xp5_ASAP7_75t_L g502 ( .A1(n_471), .A2(n_426), .B1(n_425), .B2(n_398), .C(n_400), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_451), .B(n_400), .Y(n_503) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_440), .A2(n_401), .B(n_434), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_452), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_441), .B(n_435), .Y(n_506) );
NOR3xp33_ASAP7_75t_L g507 ( .A(n_468), .B(n_469), .C(n_470), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_441), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_455), .Y(n_509) );
INVxp67_ASAP7_75t_L g510 ( .A(n_476), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_453), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_438), .B(n_412), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_458), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_477), .B(n_396), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_501), .B(n_446), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_489), .Y(n_516) );
OAI31xp33_ASAP7_75t_L g517 ( .A1(n_493), .A2(n_440), .A3(n_446), .B(n_479), .Y(n_517) );
OAI22xp5_ASAP7_75t_SL g518 ( .A1(n_510), .A2(n_401), .B1(n_472), .B2(n_453), .Y(n_518) );
NAND2xp33_ASAP7_75t_L g519 ( .A(n_500), .B(n_457), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_490), .B(n_454), .Y(n_520) );
OAI322xp33_ASAP7_75t_L g521 ( .A1(n_487), .A2(n_483), .A3(n_444), .B1(n_474), .B2(n_461), .C1(n_466), .C2(n_465), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_492), .B(n_448), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_488), .A2(n_448), .B(n_456), .Y(n_523) );
AOI221xp5_ASAP7_75t_L g524 ( .A1(n_485), .A2(n_457), .B1(n_456), .B2(n_479), .C(n_464), .Y(n_524) );
INVx1_ASAP7_75t_SL g525 ( .A(n_498), .Y(n_525) );
AOI221xp5_ASAP7_75t_L g526 ( .A1(n_502), .A2(n_482), .B1(n_460), .B2(n_450), .C(n_434), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_494), .A2(n_434), .B1(n_364), .B2(n_358), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_505), .Y(n_528) );
AOI31xp33_ASAP7_75t_L g529 ( .A1(n_495), .A2(n_379), .A3(n_358), .B(n_364), .Y(n_529) );
OA33x2_ASAP7_75t_L g530 ( .A1(n_496), .A2(n_402), .A3(n_399), .B1(n_450), .B2(n_482), .B3(n_460), .Y(n_530) );
AO221x1_ASAP7_75t_L g531 ( .A1(n_508), .A2(n_369), .B1(n_374), .B2(n_358), .C(n_376), .Y(n_531) );
AOI21xp33_ASAP7_75t_L g532 ( .A1(n_495), .A2(n_369), .B(n_374), .Y(n_532) );
NAND4xp75_ASAP7_75t_L g533 ( .A(n_504), .B(n_283), .C(n_369), .D(n_267), .Y(n_533) );
NOR3xp33_ASAP7_75t_L g534 ( .A(n_491), .B(n_280), .C(n_259), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_497), .B(n_282), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_494), .B(n_282), .Y(n_536) );
OAI21xp33_ASAP7_75t_L g537 ( .A1(n_486), .A2(n_277), .B(n_280), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_491), .B(n_245), .Y(n_538) );
NAND4xp75_ASAP7_75t_L g539 ( .A(n_514), .B(n_267), .C(n_270), .D(n_252), .Y(n_539) );
AOI311xp33_ASAP7_75t_L g540 ( .A1(n_507), .A2(n_277), .A3(n_280), .B(n_267), .C(n_240), .Y(n_540) );
AOI221xp5_ASAP7_75t_L g541 ( .A1(n_514), .A2(n_245), .B1(n_267), .B2(n_509), .C(n_513), .Y(n_541) );
NAND4xp75_ASAP7_75t_L g542 ( .A(n_484), .B(n_245), .C(n_499), .D(n_512), .Y(n_542) );
AOI221xp5_ASAP7_75t_L g543 ( .A1(n_521), .A2(n_519), .B1(n_524), .B2(n_537), .C(n_525), .Y(n_543) );
OAI21xp5_ASAP7_75t_L g544 ( .A1(n_517), .A2(n_523), .B(n_525), .Y(n_544) );
NAND4xp75_ASAP7_75t_L g545 ( .A(n_526), .B(n_527), .C(n_532), .D(n_541), .Y(n_545) );
NAND4xp75_ASAP7_75t_L g546 ( .A(n_536), .B(n_538), .C(n_515), .D(n_535), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_528), .Y(n_547) );
NAND4xp75_ASAP7_75t_L g548 ( .A(n_544), .B(n_516), .C(n_518), .D(n_529), .Y(n_548) );
NOR3xp33_ASAP7_75t_L g549 ( .A(n_543), .B(n_542), .C(n_533), .Y(n_549) );
NAND3xp33_ASAP7_75t_SL g550 ( .A(n_547), .B(n_534), .C(n_531), .Y(n_550) );
NOR2xp67_ASAP7_75t_L g551 ( .A(n_550), .B(n_520), .Y(n_551) );
OR2x6_ASAP7_75t_L g552 ( .A(n_548), .B(n_545), .Y(n_552) );
INVx4_ASAP7_75t_L g553 ( .A(n_552), .Y(n_553) );
INVx3_ASAP7_75t_SL g554 ( .A(n_553), .Y(n_554) );
XNOR2xp5_ASAP7_75t_L g555 ( .A(n_554), .B(n_551), .Y(n_555) );
OA21x2_ASAP7_75t_L g556 ( .A1(n_555), .A2(n_549), .B(n_546), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_556), .A2(n_522), .B(n_503), .Y(n_557) );
OAI21xp5_ASAP7_75t_L g558 ( .A1(n_557), .A2(n_539), .B(n_511), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_558), .A2(n_506), .B1(n_530), .B2(n_540), .Y(n_559) );
endmodule