module fake_netlist_5_2055_n_2895 (n_137, n_676, n_294, n_431, n_318, n_380, n_419, n_653, n_611, n_444, n_642, n_469, n_615, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_619, n_408, n_61, n_664, n_376, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_667, n_515, n_57, n_353, n_351, n_367, n_620, n_643, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_649, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_590, n_629, n_672, n_4, n_378, n_551, n_17, n_581, n_382, n_554, n_254, n_33, n_23, n_583, n_671, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_625, n_621, n_100, n_455, n_674, n_417, n_612, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_606, n_559, n_275, n_640, n_252, n_624, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_610, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_668, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_659, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_650, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_658, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_654, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_636, n_600, n_660, n_223, n_392, n_158, n_655, n_138, n_264, n_109, n_669, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_635, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_662, n_459, n_646, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_622, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_661, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_670, n_15, n_336, n_584, n_591, n_145, n_48, n_521, n_614, n_663, n_50, n_337, n_430, n_313, n_631, n_673, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_675, n_296, n_613, n_241, n_637, n_357, n_598, n_608, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_638, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_652, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_595, n_502, n_239, n_466, n_420, n_630, n_489, n_632, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_627, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_648, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_641, n_628, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_647, n_237, n_425, n_513, n_407, n_527, n_180, n_560, n_656, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_665, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_623, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_572, n_113, n_246, n_596, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_657, n_126, n_644, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_651, n_435, n_159, n_334, n_599, n_541, n_391, n_434, n_645, n_539, n_175, n_538, n_666, n_262, n_238, n_639, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_634, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_2895);

input n_137;
input n_676;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_653;
input n_611;
input n_444;
input n_642;
input n_469;
input n_615;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_619;
input n_408;
input n_61;
input n_664;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_667;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_643;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_649;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_629;
input n_672;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_583;
input n_671;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_625;
input n_621;
input n_100;
input n_455;
input n_674;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_606;
input n_559;
input n_275;
input n_640;
input n_252;
input n_624;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_610;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_668;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_659;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_650;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_658;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_654;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_636;
input n_600;
input n_660;
input n_223;
input n_392;
input n_158;
input n_655;
input n_138;
input n_264;
input n_109;
input n_669;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_635;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_662;
input n_459;
input n_646;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_661;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_670;
input n_15;
input n_336;
input n_584;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_663;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_673;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_675;
input n_296;
input n_613;
input n_241;
input n_637;
input n_357;
input n_598;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_638;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_652;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_502;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_627;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_648;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_641;
input n_628;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_647;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_560;
input n_656;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_665;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_623;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_657;
input n_126;
input n_644;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_651;
input n_435;
input n_159;
input n_334;
input n_599;
input n_541;
input n_391;
input n_434;
input n_645;
input n_539;
input n_175;
input n_538;
input n_666;
input n_262;
input n_238;
input n_639;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_634;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2895;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2417;
wire n_2253;
wire n_2756;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_785;
wire n_2617;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_1007;
wire n_2369;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_2143;
wire n_2853;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1107;
wire n_1728;
wire n_2031;
wire n_2076;
wire n_2482;
wire n_2677;
wire n_1230;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_2770;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1243;
wire n_1016;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_2761;
wire n_731;
wire n_1483;
wire n_2888;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2635;
wire n_2652;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_2651;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_696;
wire n_897;
wire n_798;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_1414;
wire n_1216;
wire n_2693;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_926;
wire n_2249;
wire n_2180;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_1070;
wire n_777;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_1513;
wire n_1600;
wire n_845;
wire n_2235;
wire n_1862;
wire n_837;
wire n_1239;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_1587;
wire n_680;
wire n_1473;
wire n_2682;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_1672;
wire n_2506;
wire n_2699;
wire n_888;
wire n_1880;
wire n_2769;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_2753;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_1836;
wire n_2868;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_2833;
wire n_1585;
wire n_2684;
wire n_2712;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_2855;
wire n_2713;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_2100;
wire n_2258;
wire n_748;
wire n_1058;
wire n_1667;
wire n_838;
wire n_2784;
wire n_1053;
wire n_1224;
wire n_2865;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2757;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_1385;
wire n_793;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2862;
wire n_2175;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_1565;
wire n_2828;
wire n_1809;
wire n_1856;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_857;
wire n_832;
wire n_2305;
wire n_2636;
wire n_2450;
wire n_1319;
wire n_2379;
wire n_2616;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2798;
wire n_2331;
wire n_2293;
wire n_686;
wire n_2837;
wire n_847;
wire n_1393;
wire n_2319;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_2762;
wire n_2808;
wire n_702;
wire n_1276;
wire n_2548;
wire n_822;
wire n_1412;
wire n_2679;
wire n_1709;
wire n_2676;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_1038;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_2698;
wire n_809;
wire n_870;
wire n_931;
wire n_1891;
wire n_1662;
wire n_1711;
wire n_1481;
wire n_2626;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_868;
wire n_2454;
wire n_2804;
wire n_914;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_2009;
wire n_1888;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_1189;
wire n_2690;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_2621;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2491;
wire n_2177;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_2671;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_2022;
wire n_1798;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_2007;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_1510;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_2718;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_2577;
wire n_1760;
wire n_2875;
wire n_936;
wire n_1500;
wire n_1090;
wire n_2796;
wire n_757;
wire n_2342;
wire n_2856;
wire n_1832;
wire n_1851;
wire n_999;
wire n_758;
wire n_2046;
wire n_2848;
wire n_2741;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_2787;
wire n_1964;
wire n_2869;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_2846;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_2061;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_2857;
wire n_1586;
wire n_959;
wire n_2459;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_1017;
wire n_2481;
wire n_2171;
wire n_978;
wire n_2768;
wire n_2314;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2320;
wire n_2339;
wire n_2473;
wire n_2137;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_2882;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_2812;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_2565;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_2418;
wire n_829;
wire n_2519;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_700;
wire n_1237;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_2681;
wire n_1562;
wire n_834;
wire n_765;
wire n_2424;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_2878;
wire n_1823;
wire n_874;
wire n_2464;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_860;
wire n_2849;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_1849;
wire n_2410;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_2645;
wire n_2467;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_1205;
wire n_1044;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_2508;
wire n_2593;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_2088;
wire n_824;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_2658;
wire n_1717;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_1821;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2890;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_716;
wire n_1630;
wire n_2512;
wire n_2122;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_2647;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_2824;
wire n_2650;
wire n_968;
wire n_912;
wire n_2440;
wire n_1699;
wire n_1386;
wire n_967;
wire n_1442;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_2333;
wire n_885;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_2870;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_2637;
wire n_690;
wire n_1974;
wire n_2463;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_2881;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_753;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_2415;
wire n_2309;
wire n_2646;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_1312;
wire n_1439;
wire n_804;
wire n_2827;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_2755;
wire n_842;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_2153;
wire n_1977;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_2533;
wire n_896;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2860;
wire n_2291;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_2318;
wire n_833;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2749;
wire n_2043;
wire n_1940;
wire n_814;
wire n_2707;
wire n_2751;
wire n_2793;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_2758;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_2559;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_2295;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_2840;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_2893;
wire n_1188;
wire n_2588;
wire n_1722;
wire n_2441;
wire n_1802;
wire n_2600;
wire n_849;
wire n_2795;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_2800;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_749;
wire n_1895;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_2653;
wire n_836;
wire n_990;
wire n_2867;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_1465;
wire n_778;
wire n_1122;
wire n_2608;
wire n_2657;
wire n_770;
wire n_1375;
wire n_2494;
wire n_2649;
wire n_1102;
wire n_2852;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_2633;
wire n_1441;
wire n_2522;
wire n_2435;
wire n_1597;
wire n_1392;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2542;
wire n_2313;
wire n_2097;
wire n_1174;
wire n_2431;
wire n_2835;
wire n_2558;
wire n_1371;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_726;
wire n_982;
wire n_2575;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2722;
wire n_2117;
wire n_2745;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1345;
wire n_1059;
wire n_1133;
wire n_1912;
wire n_1771;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_2877;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_1584;
wire n_1835;
wire n_1726;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_2634;
wire n_910;
wire n_2232;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_2811;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_708;
wire n_1812;
wire n_735;
wire n_2501;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_2665;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_1067;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_2003;
wire n_766;
wire n_1457;
wire n_2692;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_872;
wire n_2012;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_2103;
wire n_2160;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_1178;
wire n_855;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_2421;
wire n_2286;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_2430;
wire n_2363;
wire n_916;
wire n_1081;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_1235;
wire n_980;
wire n_698;
wire n_703;
wire n_1115;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2601;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_2686;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_2316;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2817;
wire n_2773;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_2687;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_2850;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_2654;
wire n_997;
wire n_932;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_2884;
wire n_1268;
wire n_825;
wire n_2819;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_812;
wire n_2104;
wire n_2748;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_2717;
wire n_2818;
wire n_1100;
wire n_2129;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_2889;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_1675;
wire n_1924;
wire n_2573;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_1745;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2447;
wire n_1813;
wire n_2343;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_2726;
wire n_2774;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_786;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_930;
wire n_1873;
wire n_1411;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_2854;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_682;
wire n_1567;
wire n_2567;
wire n_1247;
wire n_2709;
wire n_922;
wire n_816;
wire n_1648;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_685;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_2834;
wire n_2531;
wire n_1589;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2883;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_2809;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2591;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_1546;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_699;
wire n_979;
wire n_1515;
wire n_2841;
wire n_1627;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2505;
wire n_2438;
wire n_1673;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_2112;
wire n_1739;
wire n_2278;
wire n_2594;
wire n_2394;
wire n_1914;
wire n_2335;
wire n_2135;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2569;
wire n_2349;
wire n_1103;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_2655;
wire n_2027;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_2513;
wire n_2525;
wire n_2695;
wire n_1764;
wire n_2892;
wire n_712;
wire n_2414;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2044;
wire n_1990;
wire n_2013;
wire n_2689;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_1693;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_2839;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_2802;
wire n_1542;
wire n_1251;
wire n_2728;
wire n_2268;

INVx1_ASAP7_75t_L g677 ( 
.A(n_494),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_674),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_613),
.Y(n_679)
);

CKINVDCx14_ASAP7_75t_R g680 ( 
.A(n_136),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_490),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_617),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_63),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_514),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_648),
.Y(n_685)
);

BUFx10_ASAP7_75t_L g686 ( 
.A(n_621),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_176),
.Y(n_687)
);

CKINVDCx20_ASAP7_75t_R g688 ( 
.A(n_663),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_47),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_148),
.Y(n_690)
);

BUFx10_ASAP7_75t_L g691 ( 
.A(n_630),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_587),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_81),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_645),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_631),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_276),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_27),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_166),
.Y(n_698)
);

BUFx10_ASAP7_75t_L g699 ( 
.A(n_622),
.Y(n_699)
);

CKINVDCx20_ASAP7_75t_R g700 ( 
.A(n_605),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_658),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_336),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_477),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_665),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_655),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_309),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_242),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_217),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_51),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_157),
.Y(n_710)
);

BUFx10_ASAP7_75t_L g711 ( 
.A(n_316),
.Y(n_711)
);

CKINVDCx20_ASAP7_75t_R g712 ( 
.A(n_480),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_390),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_337),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_666),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_517),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_75),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_236),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_582),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_24),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_588),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_602),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_29),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_110),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_129),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_453),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_63),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_590),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_533),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_511),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_319),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_563),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_600),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_81),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_281),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_132),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_541),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_654),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_549),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_378),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_669),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_271),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_596),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_670),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_33),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_157),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_429),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_552),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_664),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_323),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_660),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_564),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_651),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_623),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_653),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_609),
.Y(n_756)
);

INVxp67_ASAP7_75t_L g757 ( 
.A(n_329),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_339),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_124),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_649),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_521),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_554),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_539),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_235),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_296),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_579),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_475),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_461),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_393),
.Y(n_769)
);

CKINVDCx16_ASAP7_75t_R g770 ( 
.A(n_297),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_601),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_634),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_200),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_149),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_467),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_370),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_525),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_280),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_312),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_637),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_94),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_620),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_628),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_0),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_567),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_69),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_279),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_108),
.Y(n_788)
);

BUFx2_ASAP7_75t_L g789 ( 
.A(n_497),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_591),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_27),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_127),
.Y(n_792)
);

CKINVDCx14_ASAP7_75t_R g793 ( 
.A(n_133),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_124),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_360),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_603),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_186),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_228),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_254),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_189),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_95),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_173),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_126),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_200),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_614),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_440),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_446),
.Y(n_807)
);

BUFx10_ASAP7_75t_L g808 ( 
.A(n_300),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_586),
.Y(n_809)
);

CKINVDCx20_ASAP7_75t_R g810 ( 
.A(n_185),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_661),
.Y(n_811)
);

INVx1_ASAP7_75t_SL g812 ( 
.A(n_499),
.Y(n_812)
);

BUFx10_ASAP7_75t_L g813 ( 
.A(n_404),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_400),
.Y(n_814)
);

CKINVDCx16_ASAP7_75t_R g815 ( 
.A(n_589),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_284),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_188),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_322),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_120),
.Y(n_819)
);

CKINVDCx16_ASAP7_75t_R g820 ( 
.A(n_565),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_451),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_426),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_223),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_468),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_485),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_150),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_387),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_54),
.Y(n_828)
);

INVx1_ASAP7_75t_SL g829 ( 
.A(n_391),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_574),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_182),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_39),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_438),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_282),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_518),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_325),
.Y(n_836)
);

INVxp67_ASAP7_75t_L g837 ( 
.A(n_434),
.Y(n_837)
);

CKINVDCx20_ASAP7_75t_R g838 ( 
.A(n_313),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_334),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_572),
.Y(n_840)
);

BUFx2_ASAP7_75t_L g841 ( 
.A(n_366),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_435),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_538),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_15),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_147),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_382),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_225),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_328),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_553),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_243),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_667),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_65),
.Y(n_852)
);

INVx1_ASAP7_75t_SL g853 ( 
.A(n_551),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_626),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_397),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_220),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_70),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_240),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_329),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_263),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_189),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_166),
.Y(n_862)
);

CKINVDCx16_ASAP7_75t_R g863 ( 
.A(n_624),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_305),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_584),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_284),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_546),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_278),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_544),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_51),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_126),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_50),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_526),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_668),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_310),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_616),
.Y(n_876)
);

CKINVDCx16_ASAP7_75t_R g877 ( 
.A(n_267),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_594),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_633),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_328),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_615),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_636),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_123),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_127),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_547),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_372),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_618),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_578),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_611),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_320),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_13),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_144),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_642),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_437),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_560),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_386),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_97),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_52),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_534),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_415),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_671),
.Y(n_901)
);

CKINVDCx20_ASAP7_75t_R g902 ( 
.A(n_556),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_492),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_465),
.Y(n_904)
);

CKINVDCx20_ASAP7_75t_R g905 ( 
.A(n_285),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_137),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_137),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_568),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_199),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_454),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_495),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_108),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_128),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_643),
.Y(n_914)
);

CKINVDCx20_ASAP7_75t_R g915 ( 
.A(n_673),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_304),
.Y(n_916)
);

CKINVDCx20_ASAP7_75t_R g917 ( 
.A(n_241),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_431),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_656),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_581),
.Y(n_920)
);

CKINVDCx20_ASAP7_75t_R g921 ( 
.A(n_88),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_675),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_273),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_91),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_639),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_510),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_7),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_606),
.Y(n_928)
);

BUFx2_ASAP7_75t_L g929 ( 
.A(n_66),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_522),
.Y(n_930)
);

CKINVDCx20_ASAP7_75t_R g931 ( 
.A(n_330),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_248),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_395),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_266),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_430),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_272),
.Y(n_936)
);

BUFx5_ASAP7_75t_L g937 ( 
.A(n_376),
.Y(n_937)
);

INVx1_ASAP7_75t_SL g938 ( 
.A(n_8),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_158),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_411),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_175),
.Y(n_941)
);

CKINVDCx20_ASAP7_75t_R g942 ( 
.A(n_350),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_26),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_30),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_632),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_566),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_472),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_333),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_128),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_417),
.Y(n_950)
);

BUFx2_ASAP7_75t_L g951 ( 
.A(n_321),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_18),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_571),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_263),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_326),
.Y(n_955)
);

BUFx8_ASAP7_75t_SL g956 ( 
.A(n_121),
.Y(n_956)
);

CKINVDCx20_ASAP7_75t_R g957 ( 
.A(n_550),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_161),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_65),
.Y(n_959)
);

BUFx10_ASAP7_75t_L g960 ( 
.A(n_629),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_249),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_250),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_151),
.Y(n_963)
);

BUFx8_ASAP7_75t_SL g964 ( 
.A(n_368),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_44),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_471),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_290),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_319),
.Y(n_968)
);

BUFx2_ASAP7_75t_L g969 ( 
.A(n_413),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_569),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_181),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_48),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_223),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_132),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_294),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_57),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_540),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_233),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_595),
.Y(n_979)
);

BUFx10_ASAP7_75t_L g980 ( 
.A(n_268),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_191),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_39),
.Y(n_982)
);

BUFx10_ASAP7_75t_L g983 ( 
.A(n_317),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_257),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_32),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_364),
.Y(n_986)
);

BUFx10_ASAP7_75t_L g987 ( 
.A(n_308),
.Y(n_987)
);

CKINVDCx16_ASAP7_75t_R g988 ( 
.A(n_190),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_185),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_168),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_249),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_593),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_300),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_327),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_165),
.Y(n_995)
);

BUFx5_ASAP7_75t_L g996 ( 
.A(n_118),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_6),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_362),
.Y(n_998)
);

BUFx3_ASAP7_75t_L g999 ( 
.A(n_394),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_318),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_237),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_198),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_55),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_462),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_529),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_389),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_10),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_242),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_555),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_117),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_190),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_577),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_187),
.Y(n_1013)
);

CKINVDCx16_ASAP7_75t_R g1014 ( 
.A(n_307),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_96),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_652),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_343),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_352),
.Y(n_1018)
);

BUFx3_ASAP7_75t_L g1019 ( 
.A(n_123),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_314),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_302),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_576),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_501),
.Y(n_1023)
);

INVx1_ASAP7_75t_SL g1024 ( 
.A(n_575),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_1),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_452),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_598),
.Y(n_1027)
);

BUFx10_ASAP7_75t_L g1028 ( 
.A(n_342),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_62),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_379),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_82),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_619),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_516),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_479),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_608),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_445),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_299),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_152),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_160),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_646),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_17),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_73),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_28),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_418),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_449),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_558),
.Y(n_1046)
);

CKINVDCx20_ASAP7_75t_R g1047 ( 
.A(n_464),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_341),
.Y(n_1048)
);

BUFx5_ASAP7_75t_L g1049 ( 
.A(n_97),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_78),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_47),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_196),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_531),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_498),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_457),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_315),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_562),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_543),
.Y(n_1058)
);

CKINVDCx20_ASAP7_75t_R g1059 ( 
.A(n_676),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_573),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_316),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_218),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_599),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_71),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_217),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_385),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_322),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_612),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_357),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_176),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_198),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_231),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_476),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_10),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_133),
.Y(n_1075)
);

INVx1_ASAP7_75t_SL g1076 ( 
.A(n_650),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_580),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_657),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_308),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_155),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_261),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_459),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_44),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_659),
.Y(n_1084)
);

BUFx8_ASAP7_75t_SL g1085 ( 
.A(n_56),
.Y(n_1085)
);

CKINVDCx20_ASAP7_75t_R g1086 ( 
.A(n_583),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_305),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_496),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_272),
.Y(n_1089)
);

CKINVDCx20_ASAP7_75t_R g1090 ( 
.A(n_380),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_76),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_635),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_256),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_469),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_98),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_428),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_203),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_235),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_135),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_56),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_203),
.Y(n_1101)
);

BUFx5_ASAP7_75t_L g1102 ( 
.A(n_513),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_115),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_306),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_148),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_151),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_561),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_597),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_307),
.Y(n_1109)
);

CKINVDCx16_ASAP7_75t_R g1110 ( 
.A(n_16),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_545),
.Y(n_1111)
);

CKINVDCx20_ASAP7_75t_R g1112 ( 
.A(n_196),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_142),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_354),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_559),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_265),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_192),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_261),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_647),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_274),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_52),
.Y(n_1121)
);

INVx2_ASAP7_75t_SL g1122 ( 
.A(n_425),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_36),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_180),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_32),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_201),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_331),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_625),
.Y(n_1128)
);

CKINVDCx14_ASAP7_75t_R g1129 ( 
.A(n_335),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_229),
.Y(n_1130)
);

CKINVDCx20_ASAP7_75t_R g1131 ( 
.A(n_570),
.Y(n_1131)
);

INVx1_ASAP7_75t_SL g1132 ( 
.A(n_592),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_191),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_142),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_324),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_672),
.Y(n_1136)
);

CKINVDCx14_ASAP7_75t_R g1137 ( 
.A(n_160),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_304),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_240),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_318),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_254),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_173),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_74),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_75),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_92),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_121),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_427),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_9),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_408),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_347),
.Y(n_1150)
);

INVx1_ASAP7_75t_SL g1151 ( 
.A(n_264),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_401),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_78),
.Y(n_1153)
);

INVx1_ASAP7_75t_SL g1154 ( 
.A(n_607),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_460),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_644),
.Y(n_1156)
);

INVx2_ASAP7_75t_SL g1157 ( 
.A(n_62),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_299),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_147),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_610),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_112),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_520),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_134),
.Y(n_1163)
);

BUFx10_ASAP7_75t_L g1164 ( 
.A(n_585),
.Y(n_1164)
);

CKINVDCx16_ASAP7_75t_R g1165 ( 
.A(n_627),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_114),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_548),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_283),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_29),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_106),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_532),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_99),
.Y(n_1172)
);

BUFx3_ASAP7_75t_L g1173 ( 
.A(n_15),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_207),
.Y(n_1174)
);

CKINVDCx16_ASAP7_75t_R g1175 ( 
.A(n_311),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_638),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_96),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_662),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_523),
.Y(n_1179)
);

CKINVDCx16_ASAP7_75t_R g1180 ( 
.A(n_218),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_303),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_138),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_491),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_49),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_641),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_25),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_239),
.Y(n_1187)
);

INVxp67_ASAP7_75t_L g1188 ( 
.A(n_268),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_604),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_232),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_557),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_640),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_834),
.Y(n_1193)
);

BUFx3_ASAP7_75t_L g1194 ( 
.A(n_681),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_789),
.B(n_0),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_834),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_996),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_680),
.B(n_1),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_996),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_841),
.B(n_2),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_680),
.B(n_2),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_834),
.Y(n_1202)
);

INVx5_ASAP7_75t_L g1203 ( 
.A(n_753),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_996),
.Y(n_1204)
);

BUFx8_ASAP7_75t_SL g1205 ( 
.A(n_956),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_969),
.B(n_3),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_996),
.Y(n_1207)
);

CKINVDCx16_ASAP7_75t_R g1208 ( 
.A(n_770),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_793),
.B(n_3),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_SL g1210 ( 
.A(n_815),
.B(n_4),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_731),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1178),
.B(n_4),
.Y(n_1212)
);

INVx5_ASAP7_75t_L g1213 ( 
.A(n_753),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_996),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_681),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_999),
.B(n_5),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_956),
.Y(n_1217)
);

BUFx8_ASAP7_75t_L g1218 ( 
.A(n_929),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_834),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_996),
.Y(n_1220)
);

INVx5_ASAP7_75t_L g1221 ( 
.A(n_753),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_886),
.B(n_5),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_996),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_1085),
.Y(n_1224)
);

NOR2x1_ASAP7_75t_L g1225 ( 
.A(n_999),
.B(n_332),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_793),
.B(n_6),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1137),
.B(n_7),
.Y(n_1227)
);

INVx3_ASAP7_75t_L g1228 ( 
.A(n_731),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_1114),
.B(n_8),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_966),
.B(n_9),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1137),
.B(n_11),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1114),
.B(n_11),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1049),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_951),
.B(n_12),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1143),
.B(n_12),
.Y(n_1235)
);

INVx4_ASAP7_75t_L g1236 ( 
.A(n_753),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_826),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1129),
.B(n_13),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1129),
.B(n_14),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_826),
.B(n_14),
.Y(n_1240)
);

INVx5_ASAP7_75t_L g1241 ( 
.A(n_833),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1049),
.Y(n_1242)
);

AND2x6_ASAP7_75t_L g1243 ( 
.A(n_833),
.B(n_338),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1049),
.B(n_16),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_856),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_856),
.Y(n_1246)
);

CKINVDCx6p67_ASAP7_75t_R g1247 ( 
.A(n_820),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_722),
.B(n_17),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1049),
.B(n_18),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1049),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1049),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1049),
.B(n_19),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_856),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_782),
.B(n_19),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_856),
.Y(n_1255)
);

BUFx12f_ASAP7_75t_L g1256 ( 
.A(n_711),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_975),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_865),
.B(n_20),
.Y(n_1258)
);

BUFx2_ASAP7_75t_L g1259 ( 
.A(n_1085),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_975),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1122),
.B(n_20),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_882),
.B(n_21),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_949),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_949),
.B(n_21),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_677),
.B(n_22),
.Y(n_1265)
);

AND2x4_ASAP7_75t_L g1266 ( 
.A(n_679),
.B(n_22),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_684),
.B(n_23),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_882),
.B(n_23),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_928),
.B(n_24),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_686),
.Y(n_1270)
);

INVxp67_ASAP7_75t_L g1271 ( 
.A(n_1079),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_975),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_837),
.B(n_25),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1019),
.B(n_26),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_928),
.B(n_28),
.Y(n_1275)
);

BUFx8_ASAP7_75t_SL g1276 ( 
.A(n_964),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1096),
.B(n_30),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_975),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_692),
.B(n_31),
.Y(n_1279)
);

BUFx12f_ASAP7_75t_L g1280 ( 
.A(n_711),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1096),
.B(n_31),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_994),
.Y(n_1282)
);

INVx5_ASAP7_75t_L g1283 ( 
.A(n_833),
.Y(n_1283)
);

INVx5_ASAP7_75t_L g1284 ( 
.A(n_833),
.Y(n_1284)
);

INVx3_ASAP7_75t_L g1285 ( 
.A(n_1019),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1176),
.B(n_33),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_702),
.B(n_34),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_994),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1176),
.B(n_34),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_994),
.Y(n_1290)
);

BUFx8_ASAP7_75t_L g1291 ( 
.A(n_994),
.Y(n_1291)
);

AND2x6_ASAP7_75t_L g1292 ( 
.A(n_1150),
.B(n_340),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1083),
.B(n_35),
.Y(n_1293)
);

INVx5_ASAP7_75t_L g1294 ( 
.A(n_1150),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_812),
.B(n_35),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1083),
.B(n_36),
.Y(n_1296)
);

BUFx12f_ASAP7_75t_L g1297 ( 
.A(n_711),
.Y(n_1297)
);

BUFx6f_ASAP7_75t_L g1298 ( 
.A(n_1169),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1169),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1146),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1169),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_705),
.B(n_37),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1169),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1146),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_L g1305 ( 
.A(n_1173),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_L g1306 ( 
.A(n_829),
.B(n_37),
.Y(n_1306)
);

INVx3_ASAP7_75t_L g1307 ( 
.A(n_1173),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_877),
.B(n_38),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1150),
.Y(n_1309)
);

INVx5_ASAP7_75t_L g1310 ( 
.A(n_1150),
.Y(n_1310)
);

INVx5_ASAP7_75t_L g1311 ( 
.A(n_686),
.Y(n_1311)
);

INVx5_ASAP7_75t_L g1312 ( 
.A(n_686),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_698),
.Y(n_1313)
);

BUFx6f_ASAP7_75t_L g1314 ( 
.A(n_696),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_937),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_937),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_988),
.Y(n_1317)
);

INVx5_ASAP7_75t_L g1318 ( 
.A(n_691),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_719),
.B(n_38),
.Y(n_1319)
);

INVxp67_ASAP7_75t_L g1320 ( 
.A(n_808),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_696),
.Y(n_1321)
);

BUFx12f_ASAP7_75t_L g1322 ( 
.A(n_808),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_764),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_853),
.B(n_40),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_1024),
.B(n_40),
.Y(n_1325)
);

AND2x4_ASAP7_75t_L g1326 ( 
.A(n_729),
.B(n_41),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1076),
.B(n_41),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_SL g1328 ( 
.A(n_863),
.B(n_42),
.Y(n_1328)
);

BUFx6f_ASAP7_75t_L g1329 ( 
.A(n_764),
.Y(n_1329)
);

INVx5_ASAP7_75t_L g1330 ( 
.A(n_691),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_732),
.B(n_42),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_725),
.Y(n_1332)
);

BUFx6f_ASAP7_75t_L g1333 ( 
.A(n_864),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1014),
.B(n_43),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1110),
.B(n_43),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_864),
.Y(n_1336)
);

BUFx12f_ASAP7_75t_L g1337 ( 
.A(n_808),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_875),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_875),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_927),
.Y(n_1340)
);

BUFx12f_ASAP7_75t_L g1341 ( 
.A(n_980),
.Y(n_1341)
);

INVx5_ASAP7_75t_L g1342 ( 
.A(n_691),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_736),
.Y(n_1343)
);

INVx5_ASAP7_75t_L g1344 ( 
.A(n_699),
.Y(n_1344)
);

INVx2_ASAP7_75t_SL g1345 ( 
.A(n_980),
.Y(n_1345)
);

INVxp67_ASAP7_75t_L g1346 ( 
.A(n_980),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1175),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_927),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_954),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_937),
.B(n_45),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_738),
.B(n_45),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_937),
.Y(n_1352)
);

INVx5_ASAP7_75t_L g1353 ( 
.A(n_699),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_954),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1180),
.Y(n_1355)
);

INVx5_ASAP7_75t_L g1356 ( 
.A(n_699),
.Y(n_1356)
);

AND2x6_ASAP7_75t_L g1357 ( 
.A(n_1132),
.B(n_344),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_742),
.Y(n_1358)
);

INVx5_ASAP7_75t_L g1359 ( 
.A(n_813),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_937),
.B(n_46),
.Y(n_1360)
);

INVx2_ASAP7_75t_SL g1361 ( 
.A(n_983),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_740),
.B(n_46),
.Y(n_1362)
);

NAND3xp33_ASAP7_75t_L g1363 ( 
.A(n_757),
.B(n_48),
.C(n_49),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1154),
.B(n_50),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_937),
.B(n_53),
.Y(n_1365)
);

AOI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1238),
.A2(n_1165),
.B1(n_688),
.B2(n_712),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1270),
.B(n_741),
.Y(n_1367)
);

OAI22xp33_ASAP7_75t_SL g1368 ( 
.A1(n_1210),
.A2(n_1188),
.B1(n_687),
.B2(n_745),
.Y(n_1368)
);

AO22x2_ASAP7_75t_L g1369 ( 
.A1(n_1234),
.A2(n_847),
.B1(n_870),
.B2(n_709),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_SL g1370 ( 
.A1(n_1208),
.A2(n_921),
.B1(n_931),
.B2(n_917),
.Y(n_1370)
);

AOI22xp5_ASAP7_75t_SL g1371 ( 
.A1(n_1308),
.A2(n_921),
.B1(n_931),
.B2(n_917),
.Y(n_1371)
);

OR2x6_ASAP7_75t_L g1372 ( 
.A(n_1259),
.B(n_968),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1239),
.A2(n_754),
.B1(n_762),
.B2(n_700),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_1276),
.Y(n_1374)
);

AND2x2_ASAP7_75t_SL g1375 ( 
.A(n_1328),
.B(n_972),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1193),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1311),
.B(n_743),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1253),
.Y(n_1378)
);

AOI22x1_ASAP7_75t_SL g1379 ( 
.A1(n_1224),
.A2(n_720),
.B1(n_727),
.B2(n_708),
.Y(n_1379)
);

AO22x2_ASAP7_75t_L g1380 ( 
.A1(n_1235),
.A2(n_1157),
.B1(n_1020),
.B2(n_1031),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1193),
.Y(n_1381)
);

AOI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1231),
.A2(n_915),
.B1(n_942),
.B2(n_902),
.Y(n_1382)
);

AO22x2_ASAP7_75t_L g1383 ( 
.A1(n_1226),
.A2(n_1020),
.B1(n_1031),
.B2(n_972),
.Y(n_1383)
);

OA22x2_ASAP7_75t_L g1384 ( 
.A1(n_1271),
.A2(n_765),
.B1(n_773),
.B2(n_746),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1311),
.B(n_813),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1317),
.B(n_860),
.Y(n_1386)
);

OAI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1198),
.A2(n_1151),
.B1(n_938),
.B2(n_689),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1312),
.B(n_813),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1196),
.Y(n_1389)
);

OR2x6_ASAP7_75t_L g1390 ( 
.A(n_1217),
.B(n_1148),
.Y(n_1390)
);

OAI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1201),
.A2(n_690),
.B1(n_693),
.B2(n_683),
.Y(n_1391)
);

INVx2_ASAP7_75t_SL g1392 ( 
.A(n_1312),
.Y(n_1392)
);

AOI22x1_ASAP7_75t_L g1393 ( 
.A1(n_1248),
.A2(n_1148),
.B1(n_786),
.B2(n_799),
.Y(n_1393)
);

OAI22xp33_ASAP7_75t_SL g1394 ( 
.A1(n_1209),
.A2(n_706),
.B1(n_707),
.B2(n_697),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1318),
.B(n_960),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1196),
.Y(n_1396)
);

AND2x2_ASAP7_75t_SL g1397 ( 
.A(n_1334),
.B(n_749),
.Y(n_1397)
);

AO22x2_ASAP7_75t_L g1398 ( 
.A1(n_1335),
.A2(n_801),
.B1(n_802),
.B2(n_781),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1255),
.Y(n_1399)
);

AO22x2_ASAP7_75t_L g1400 ( 
.A1(n_1216),
.A2(n_818),
.B1(n_823),
.B2(n_804),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1318),
.B(n_960),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1330),
.B(n_960),
.Y(n_1402)
);

OAI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1227),
.A2(n_717),
.B1(n_718),
.B2(n_710),
.Y(n_1403)
);

OAI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1347),
.A2(n_724),
.B1(n_734),
.B2(n_723),
.Y(n_1404)
);

XNOR2xp5_ASAP7_75t_L g1405 ( 
.A(n_1355),
.B(n_759),
.Y(n_1405)
);

OA22x2_ASAP7_75t_L g1406 ( 
.A1(n_1320),
.A2(n_845),
.B1(n_857),
.B2(n_844),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1260),
.Y(n_1407)
);

OAI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1345),
.A2(n_774),
.B1(n_778),
.B2(n_735),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1299),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1330),
.B(n_1028),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1202),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1303),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1342),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1342),
.B(n_761),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1202),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1219),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1344),
.B(n_1028),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1344),
.B(n_1028),
.Y(n_1418)
);

AO22x2_ASAP7_75t_L g1419 ( 
.A1(n_1229),
.A2(n_871),
.B1(n_880),
.B2(n_859),
.Y(n_1419)
);

OR2x6_ASAP7_75t_L g1420 ( 
.A(n_1345),
.B(n_883),
.Y(n_1420)
);

AOI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1195),
.A2(n_1023),
.B1(n_1047),
.B2(n_957),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1353),
.B(n_1164),
.Y(n_1422)
);

OA22x2_ASAP7_75t_L g1423 ( 
.A1(n_1346),
.A2(n_906),
.B1(n_913),
.B2(n_892),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1353),
.B(n_1164),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_SL g1425 ( 
.A1(n_1200),
.A2(n_810),
.B1(n_828),
.B2(n_750),
.Y(n_1425)
);

AO22x2_ASAP7_75t_L g1426 ( 
.A1(n_1232),
.A2(n_932),
.B1(n_943),
.B2(n_923),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1219),
.Y(n_1427)
);

AOI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1206),
.A2(n_1086),
.B1(n_1090),
.B2(n_1059),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1245),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_SL g1430 ( 
.A(n_1356),
.B(n_1164),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1245),
.Y(n_1431)
);

OAI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1361),
.A2(n_784),
.B1(n_787),
.B2(n_779),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1246),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1246),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1257),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1356),
.B(n_983),
.Y(n_1436)
);

AO22x2_ASAP7_75t_L g1437 ( 
.A1(n_1363),
.A2(n_958),
.B1(n_959),
.B2(n_944),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1257),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1212),
.A2(n_791),
.B1(n_792),
.B2(n_788),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_SL g1440 ( 
.A1(n_1222),
.A2(n_905),
.B1(n_939),
.B2(n_838),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1247),
.A2(n_797),
.B1(n_798),
.B2(n_794),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_SL g1442 ( 
.A1(n_1230),
.A2(n_1112),
.B1(n_1021),
.B2(n_803),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1359),
.B(n_983),
.Y(n_1443)
);

OAI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1361),
.A2(n_816),
.B1(n_817),
.B2(n_800),
.Y(n_1444)
);

AO22x2_ASAP7_75t_L g1445 ( 
.A1(n_1240),
.A2(n_967),
.B1(n_971),
.B2(n_962),
.Y(n_1445)
);

AO22x2_ASAP7_75t_L g1446 ( 
.A1(n_1240),
.A2(n_978),
.B1(n_982),
.B2(n_973),
.Y(n_1446)
);

INVx1_ASAP7_75t_SL g1447 ( 
.A(n_1205),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1359),
.B(n_987),
.Y(n_1448)
);

AOI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1295),
.A2(n_1131),
.B1(n_1189),
.B2(n_1108),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1237),
.B(n_819),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1194),
.B(n_987),
.Y(n_1451)
);

AOI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1306),
.A2(n_832),
.B1(n_836),
.B2(n_831),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1272),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1272),
.Y(n_1454)
);

AOI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1324),
.A2(n_850),
.B1(n_852),
.B2(n_848),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1325),
.A2(n_861),
.B1(n_862),
.B2(n_858),
.Y(n_1456)
);

OAI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1247),
.A2(n_866),
.B1(n_872),
.B2(n_868),
.Y(n_1457)
);

AOI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1327),
.A2(n_890),
.B1(n_891),
.B2(n_884),
.Y(n_1458)
);

XOR2xp5_ASAP7_75t_L g1459 ( 
.A(n_1225),
.B(n_678),
.Y(n_1459)
);

OAI22xp33_ASAP7_75t_SL g1460 ( 
.A1(n_1254),
.A2(n_898),
.B1(n_907),
.B2(n_897),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1215),
.B(n_771),
.Y(n_1461)
);

AOI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1364),
.A2(n_912),
.B1(n_916),
.B2(n_909),
.Y(n_1462)
);

AOI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1273),
.A2(n_934),
.B1(n_936),
.B2(n_924),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1291),
.B(n_772),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1237),
.B(n_987),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1211),
.B(n_682),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1278),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1278),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1282),
.Y(n_1469)
);

OAI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1261),
.A2(n_952),
.B1(n_955),
.B2(n_941),
.Y(n_1470)
);

OA22x2_ASAP7_75t_L g1471 ( 
.A1(n_1263),
.A2(n_1003),
.B1(n_1039),
.B2(n_991),
.Y(n_1471)
);

AND2x4_ASAP7_75t_L g1472 ( 
.A(n_1274),
.B(n_783),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_SL g1473 ( 
.A(n_1258),
.B(n_961),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1228),
.B(n_685),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1285),
.B(n_694),
.Y(n_1475)
);

AOI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1256),
.A2(n_965),
.B1(n_974),
.B2(n_963),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1282),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1288),
.Y(n_1478)
);

AO22x2_ASAP7_75t_L g1479 ( 
.A1(n_1264),
.A2(n_1296),
.B1(n_1293),
.B2(n_1266),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1288),
.Y(n_1480)
);

AOI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1280),
.A2(n_981),
.B1(n_984),
.B2(n_976),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1290),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1297),
.A2(n_989),
.B1(n_990),
.B2(n_985),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1290),
.Y(n_1484)
);

AOI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1322),
.A2(n_995),
.B1(n_997),
.B2(n_993),
.Y(n_1485)
);

OAI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1262),
.A2(n_1000),
.B1(n_1002),
.B2(n_1001),
.Y(n_1486)
);

AO22x2_ASAP7_75t_L g1487 ( 
.A1(n_1264),
.A2(n_1267),
.B1(n_1279),
.B2(n_1265),
.Y(n_1487)
);

AND2x2_ASAP7_75t_SL g1488 ( 
.A(n_1287),
.B(n_785),
.Y(n_1488)
);

AOI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1337),
.A2(n_1341),
.B1(n_1357),
.B2(n_1275),
.Y(n_1489)
);

BUFx10_ASAP7_75t_L g1490 ( 
.A(n_1300),
.Y(n_1490)
);

OAI22xp33_ASAP7_75t_SL g1491 ( 
.A1(n_1350),
.A2(n_1008),
.B1(n_1010),
.B2(n_1007),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_SL g1492 ( 
.A1(n_1289),
.A2(n_1013),
.B1(n_1015),
.B2(n_1011),
.Y(n_1492)
);

OR2x6_ASAP7_75t_L g1493 ( 
.A(n_1304),
.B(n_1050),
.Y(n_1493)
);

AO22x2_ASAP7_75t_L g1494 ( 
.A1(n_1302),
.A2(n_1061),
.B1(n_1065),
.B2(n_1052),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1298),
.Y(n_1495)
);

BUFx2_ASAP7_75t_L g1496 ( 
.A(n_1218),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1203),
.B(n_796),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1304),
.Y(n_1498)
);

AO22x2_ASAP7_75t_L g1499 ( 
.A1(n_1319),
.A2(n_1075),
.B1(n_1091),
.B2(n_1074),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1307),
.B(n_1025),
.Y(n_1500)
);

AO22x2_ASAP7_75t_L g1501 ( 
.A1(n_1326),
.A2(n_1105),
.B1(n_1109),
.B2(n_1097),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1298),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_SL g1503 ( 
.A1(n_1268),
.A2(n_1037),
.B1(n_1038),
.B2(n_1029),
.Y(n_1503)
);

AOI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1357),
.A2(n_1042),
.B1(n_1043),
.B2(n_1041),
.Y(n_1504)
);

OAI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1269),
.A2(n_1056),
.B1(n_1062),
.B2(n_1051),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_SL g1506 ( 
.A1(n_1277),
.A2(n_1067),
.B1(n_1070),
.B2(n_1064),
.Y(n_1506)
);

OR2x6_ASAP7_75t_L g1507 ( 
.A(n_1305),
.B(n_1313),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1301),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1301),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1281),
.B(n_805),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1305),
.Y(n_1511)
);

AO22x2_ASAP7_75t_L g1512 ( 
.A1(n_1331),
.A2(n_1121),
.B1(n_1123),
.B2(n_1118),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1203),
.B(n_1213),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1309),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1286),
.B(n_807),
.Y(n_1515)
);

AO22x2_ASAP7_75t_L g1516 ( 
.A1(n_1351),
.A2(n_1126),
.B1(n_1127),
.B2(n_1124),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1309),
.Y(n_1517)
);

AO22x2_ASAP7_75t_L g1518 ( 
.A1(n_1362),
.A2(n_1139),
.B1(n_1141),
.B2(n_1130),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_1314),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_R g1520 ( 
.A(n_1357),
.B(n_695),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1213),
.B(n_701),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_SL g1522 ( 
.A1(n_1360),
.A2(n_1072),
.B1(n_1080),
.B2(n_1071),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1221),
.B(n_1241),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1199),
.Y(n_1524)
);

AOI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1365),
.A2(n_1087),
.B1(n_1089),
.B2(n_1081),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1221),
.B(n_703),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1244),
.B(n_835),
.Y(n_1527)
);

OAI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1249),
.A2(n_1095),
.B1(n_1098),
.B2(n_1093),
.Y(n_1528)
);

OAI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1252),
.A2(n_1100),
.B1(n_1101),
.B2(n_1099),
.Y(n_1529)
);

AOI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1243),
.A2(n_1104),
.B1(n_1106),
.B2(n_1103),
.Y(n_1530)
);

OAI22xp33_ASAP7_75t_SL g1531 ( 
.A1(n_1332),
.A2(n_1116),
.B1(n_1117),
.B2(n_1113),
.Y(n_1531)
);

OA22x2_ASAP7_75t_L g1532 ( 
.A1(n_1358),
.A2(n_1343),
.B1(n_1177),
.B2(n_1187),
.Y(n_1532)
);

OR2x6_ASAP7_75t_L g1533 ( 
.A(n_1314),
.B(n_1158),
.Y(n_1533)
);

AO22x2_ASAP7_75t_L g1534 ( 
.A1(n_1197),
.A2(n_846),
.B1(n_854),
.B2(n_840),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1241),
.B(n_704),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1204),
.Y(n_1536)
);

OA22x2_ASAP7_75t_L g1537 ( 
.A1(n_1207),
.A2(n_1125),
.B1(n_1133),
.B2(n_1120),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1214),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1233),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1220),
.Y(n_1540)
);

OR2x6_ASAP7_75t_L g1541 ( 
.A(n_1321),
.B(n_867),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1283),
.B(n_713),
.Y(n_1542)
);

OAI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1321),
.A2(n_1135),
.B1(n_1138),
.B2(n_1134),
.Y(n_1543)
);

AO22x2_ASAP7_75t_L g1544 ( 
.A1(n_1242),
.A2(n_900),
.B1(n_903),
.B2(n_887),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1323),
.Y(n_1545)
);

OAI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1323),
.A2(n_1142),
.B1(n_1144),
.B2(n_1140),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1223),
.Y(n_1547)
);

AO22x2_ASAP7_75t_L g1548 ( 
.A1(n_1315),
.A2(n_922),
.B1(n_925),
.B2(n_918),
.Y(n_1548)
);

AOI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1243),
.A2(n_1153),
.B1(n_1159),
.B2(n_1145),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1329),
.Y(n_1550)
);

NAND2x1p5_ASAP7_75t_L g1551 ( 
.A(n_1283),
.B(n_1192),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1284),
.B(n_714),
.Y(n_1552)
);

AO22x2_ASAP7_75t_L g1553 ( 
.A1(n_1316),
.A2(n_946),
.B1(n_950),
.B2(n_926),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1284),
.B(n_715),
.Y(n_1554)
);

AOI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1243),
.A2(n_1163),
.B1(n_1166),
.B2(n_1161),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1294),
.B(n_716),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1294),
.B(n_1005),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1250),
.Y(n_1558)
);

OAI22xp33_ASAP7_75t_SL g1559 ( 
.A1(n_1352),
.A2(n_1170),
.B1(n_1172),
.B2(n_1168),
.Y(n_1559)
);

AOI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1292),
.A2(n_1181),
.B1(n_1182),
.B2(n_1174),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1329),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1251),
.A2(n_1186),
.B1(n_1190),
.B2(n_1184),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1333),
.Y(n_1563)
);

AO22x2_ASAP7_75t_L g1564 ( 
.A1(n_1236),
.A2(n_1030),
.B1(n_1033),
.B2(n_1009),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1333),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1336),
.Y(n_1566)
);

OAI22xp33_ASAP7_75t_SL g1567 ( 
.A1(n_1310),
.A2(n_1036),
.B1(n_1040),
.B2(n_1034),
.Y(n_1567)
);

AOI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1292),
.A2(n_726),
.B1(n_728),
.B2(n_721),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1310),
.B(n_730),
.Y(n_1569)
);

AOI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1292),
.A2(n_737),
.B1(n_739),
.B2(n_733),
.Y(n_1570)
);

NAND3x1_ASAP7_75t_L g1571 ( 
.A(n_1336),
.B(n_1046),
.C(n_1044),
.Y(n_1571)
);

OR2x6_ASAP7_75t_L g1572 ( 
.A(n_1338),
.B(n_1048),
.Y(n_1572)
);

AOI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1338),
.A2(n_747),
.B1(n_748),
.B2(n_744),
.Y(n_1573)
);

OAI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1339),
.A2(n_1054),
.B1(n_1066),
.B2(n_1053),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1339),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1340),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1340),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1354),
.Y(n_1578)
);

AOI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1354),
.A2(n_752),
.B1(n_755),
.B2(n_751),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1348),
.B(n_756),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1348),
.Y(n_1581)
);

AND2x4_ASAP7_75t_L g1582 ( 
.A(n_1349),
.B(n_1078),
.Y(n_1582)
);

AO22x2_ASAP7_75t_L g1583 ( 
.A1(n_1349),
.A2(n_1088),
.B1(n_1162),
.B2(n_1084),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_SL g1584 ( 
.A1(n_1208),
.A2(n_1183),
.B1(n_1191),
.B2(n_1185),
.Y(n_1584)
);

AOI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1238),
.A2(n_760),
.B1(n_763),
.B2(n_758),
.Y(n_1585)
);

AOI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1238),
.A2(n_767),
.B1(n_768),
.B2(n_766),
.Y(n_1586)
);

OAI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1210),
.A2(n_775),
.B1(n_776),
.B2(n_769),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1193),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1193),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1193),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1253),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1311),
.B(n_777),
.Y(n_1592)
);

INVx3_ASAP7_75t_L g1593 ( 
.A(n_1304),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1253),
.Y(n_1594)
);

NAND3xp33_ASAP7_75t_L g1595 ( 
.A(n_1210),
.B(n_1160),
.C(n_1156),
.Y(n_1595)
);

AOI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1238),
.A2(n_790),
.B1(n_795),
.B2(n_780),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1193),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1253),
.Y(n_1598)
);

BUFx10_ASAP7_75t_L g1599 ( 
.A(n_1224),
.Y(n_1599)
);

AOI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1238),
.A2(n_809),
.B1(n_811),
.B2(n_806),
.Y(n_1600)
);

OAI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1198),
.A2(n_821),
.B1(n_822),
.B2(n_814),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1253),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1317),
.B(n_53),
.Y(n_1603)
);

OAI22xp33_ASAP7_75t_SL g1604 ( 
.A1(n_1210),
.A2(n_825),
.B1(n_827),
.B2(n_824),
.Y(n_1604)
);

AOI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1238),
.A2(n_839),
.B1(n_842),
.B2(n_830),
.Y(n_1605)
);

AOI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1238),
.A2(n_849),
.B1(n_851),
.B2(n_843),
.Y(n_1606)
);

NAND3x1_ASAP7_75t_L g1607 ( 
.A(n_1308),
.B(n_54),
.C(n_55),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1193),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1311),
.B(n_855),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1254),
.B(n_869),
.Y(n_1610)
);

NAND3x1_ASAP7_75t_L g1611 ( 
.A(n_1308),
.B(n_57),
.C(n_58),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_SL g1612 ( 
.A1(n_1208),
.A2(n_874),
.B1(n_876),
.B2(n_873),
.Y(n_1612)
);

AO22x2_ASAP7_75t_L g1613 ( 
.A1(n_1234),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_1613)
);

AOI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1238),
.A2(n_879),
.B1(n_881),
.B2(n_878),
.Y(n_1614)
);

CKINVDCx6p67_ASAP7_75t_R g1615 ( 
.A(n_1247),
.Y(n_1615)
);

OAI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1210),
.A2(n_888),
.B1(n_889),
.B2(n_885),
.Y(n_1616)
);

AO22x2_ASAP7_75t_L g1617 ( 
.A1(n_1234),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1193),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1193),
.Y(n_1619)
);

OAI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1210),
.A2(n_894),
.B1(n_895),
.B2(n_893),
.Y(n_1620)
);

OAI22xp33_ASAP7_75t_SL g1621 ( 
.A1(n_1210),
.A2(n_899),
.B1(n_901),
.B2(n_896),
.Y(n_1621)
);

AOI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1238),
.A2(n_908),
.B1(n_910),
.B2(n_904),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1193),
.Y(n_1623)
);

INVx8_ASAP7_75t_L g1624 ( 
.A(n_1276),
.Y(n_1624)
);

AOI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1238),
.A2(n_914),
.B1(n_919),
.B2(n_911),
.Y(n_1625)
);

AO22x2_ASAP7_75t_L g1626 ( 
.A1(n_1234),
.A2(n_66),
.B1(n_61),
.B2(n_64),
.Y(n_1626)
);

OAI22xp33_ASAP7_75t_R g1627 ( 
.A1(n_1345),
.A2(n_68),
.B1(n_64),
.B2(n_67),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_1254),
.B(n_920),
.Y(n_1628)
);

OAI22xp33_ASAP7_75t_SL g1629 ( 
.A1(n_1210),
.A2(n_933),
.B1(n_935),
.B2(n_930),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1193),
.Y(n_1630)
);

AO22x2_ASAP7_75t_L g1631 ( 
.A1(n_1234),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1311),
.B(n_940),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1193),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1254),
.B(n_945),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1253),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1253),
.Y(n_1636)
);

OAI22xp33_ASAP7_75t_SL g1637 ( 
.A1(n_1210),
.A2(n_947),
.B1(n_953),
.B2(n_948),
.Y(n_1637)
);

AOI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1238),
.A2(n_970),
.B1(n_979),
.B2(n_977),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1311),
.B(n_986),
.Y(n_1639)
);

INVx3_ASAP7_75t_L g1640 ( 
.A(n_1304),
.Y(n_1640)
);

AOI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1238),
.A2(n_992),
.B1(n_1004),
.B2(n_998),
.Y(n_1641)
);

AO22x2_ASAP7_75t_L g1642 ( 
.A1(n_1234),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_1642)
);

AO22x2_ASAP7_75t_L g1643 ( 
.A1(n_1234),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_1643)
);

AOI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1238),
.A2(n_1006),
.B1(n_1016),
.B2(n_1012),
.Y(n_1644)
);

OR2x6_ASAP7_75t_L g1645 ( 
.A(n_1259),
.B(n_964),
.Y(n_1645)
);

AND2x2_ASAP7_75t_SL g1646 ( 
.A(n_1210),
.B(n_76),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1253),
.Y(n_1647)
);

OAI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1210),
.A2(n_1018),
.B1(n_1022),
.B2(n_1017),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1193),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1253),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1311),
.B(n_1026),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1198),
.A2(n_1027),
.B1(n_1035),
.B2(n_1032),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_L g1653 ( 
.A(n_1254),
.B(n_1045),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1311),
.B(n_1055),
.Y(n_1654)
);

OA22x2_ASAP7_75t_L g1655 ( 
.A1(n_1271),
.A2(n_1057),
.B1(n_1060),
.B2(n_1058),
.Y(n_1655)
);

AO22x2_ASAP7_75t_L g1656 ( 
.A1(n_1234),
.A2(n_80),
.B1(n_77),
.B2(n_79),
.Y(n_1656)
);

AOI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1238),
.A2(n_1063),
.B1(n_1069),
.B2(n_1068),
.Y(n_1657)
);

OR2x6_ASAP7_75t_L g1658 ( 
.A(n_1259),
.B(n_77),
.Y(n_1658)
);

OA22x2_ASAP7_75t_L g1659 ( 
.A1(n_1271),
.A2(n_1073),
.B1(n_1082),
.B2(n_1077),
.Y(n_1659)
);

OA22x2_ASAP7_75t_L g1660 ( 
.A1(n_1271),
.A2(n_1092),
.B1(n_1107),
.B2(n_1094),
.Y(n_1660)
);

BUFx6f_ASAP7_75t_SL g1661 ( 
.A(n_1345),
.Y(n_1661)
);

AO22x2_ASAP7_75t_L g1662 ( 
.A1(n_1234),
.A2(n_82),
.B1(n_79),
.B2(n_80),
.Y(n_1662)
);

INVx3_ASAP7_75t_L g1663 ( 
.A(n_1304),
.Y(n_1663)
);

OR2x6_ASAP7_75t_L g1664 ( 
.A(n_1259),
.B(n_83),
.Y(n_1664)
);

OAI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1198),
.A2(n_1115),
.B1(n_1119),
.B2(n_1111),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1311),
.B(n_1128),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1253),
.Y(n_1667)
);

OAI22xp33_ASAP7_75t_SL g1668 ( 
.A1(n_1210),
.A2(n_1147),
.B1(n_1149),
.B2(n_1136),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1317),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1311),
.B(n_1152),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1253),
.Y(n_1671)
);

AOI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1238),
.A2(n_1167),
.B1(n_1171),
.B2(n_1155),
.Y(n_1672)
);

AOI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1238),
.A2(n_1179),
.B1(n_1102),
.B2(n_937),
.Y(n_1673)
);

AO22x2_ASAP7_75t_L g1674 ( 
.A1(n_1234),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_SL g1675 ( 
.A1(n_1208),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1675)
);

BUFx6f_ASAP7_75t_L g1676 ( 
.A(n_1193),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1193),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1253),
.Y(n_1678)
);

AOI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1238),
.A2(n_1102),
.B1(n_88),
.B2(n_86),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1193),
.Y(n_1680)
);

INVx2_ASAP7_75t_SL g1681 ( 
.A(n_1311),
.Y(n_1681)
);

BUFx6f_ASAP7_75t_L g1682 ( 
.A(n_1193),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1311),
.B(n_1102),
.Y(n_1683)
);

AO22x2_ASAP7_75t_L g1684 ( 
.A1(n_1234),
.A2(n_90),
.B1(n_87),
.B2(n_89),
.Y(n_1684)
);

AOI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1238),
.A2(n_1102),
.B1(n_90),
.B2(n_87),
.Y(n_1685)
);

OAI22xp33_ASAP7_75t_SL g1686 ( 
.A1(n_1210),
.A2(n_1102),
.B1(n_92),
.B2(n_89),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1311),
.B(n_1102),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1253),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_1276),
.Y(n_1689)
);

OAI22xp33_ASAP7_75t_L g1690 ( 
.A1(n_1210),
.A2(n_94),
.B1(n_91),
.B2(n_93),
.Y(n_1690)
);

INVx1_ASAP7_75t_SL g1691 ( 
.A(n_1276),
.Y(n_1691)
);

AOI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1238),
.A2(n_1102),
.B1(n_98),
.B2(n_93),
.Y(n_1692)
);

AO22x2_ASAP7_75t_L g1693 ( 
.A1(n_1234),
.A2(n_100),
.B1(n_95),
.B2(n_99),
.Y(n_1693)
);

AOI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1238),
.A2(n_102),
.B1(n_100),
.B2(n_101),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1311),
.B(n_345),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1311),
.B(n_346),
.Y(n_1696)
);

OA22x2_ASAP7_75t_L g1697 ( 
.A1(n_1271),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1193),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_1276),
.Y(n_1699)
);

BUFx2_ASAP7_75t_L g1700 ( 
.A(n_1276),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1311),
.B(n_348),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1610),
.B(n_1628),
.Y(n_1702)
);

XOR2xp5_ASAP7_75t_L g1703 ( 
.A(n_1405),
.B(n_349),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1536),
.Y(n_1704)
);

NAND2x1p5_ASAP7_75t_L g1705 ( 
.A(n_1593),
.B(n_351),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1587),
.B(n_103),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1465),
.B(n_104),
.Y(n_1707)
);

CKINVDCx20_ASAP7_75t_R g1708 ( 
.A(n_1615),
.Y(n_1708)
);

BUFx5_ASAP7_75t_L g1709 ( 
.A(n_1538),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1539),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1616),
.B(n_104),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1524),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1540),
.Y(n_1713)
);

CKINVDCx20_ASAP7_75t_R g1714 ( 
.A(n_1373),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1545),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_L g1716 ( 
.A(n_1620),
.B(n_105),
.Y(n_1716)
);

CKINVDCx6p67_ASAP7_75t_R g1717 ( 
.A(n_1624),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1550),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1634),
.B(n_353),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1436),
.B(n_105),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1443),
.B(n_106),
.Y(n_1721)
);

OR2x6_ASAP7_75t_L g1722 ( 
.A(n_1624),
.B(n_107),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1561),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1563),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1565),
.Y(n_1725)
);

OR2x6_ASAP7_75t_L g1726 ( 
.A(n_1645),
.B(n_107),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1577),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1566),
.Y(n_1728)
);

XOR2xp5_ASAP7_75t_L g1729 ( 
.A(n_1382),
.B(n_355),
.Y(n_1729)
);

XNOR2xp5_ASAP7_75t_L g1730 ( 
.A(n_1371),
.B(n_109),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1575),
.Y(n_1731)
);

INVxp67_ASAP7_75t_SL g1732 ( 
.A(n_1519),
.Y(n_1732)
);

INVxp67_ASAP7_75t_L g1733 ( 
.A(n_1448),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1576),
.Y(n_1734)
);

INVx2_ASAP7_75t_SL g1735 ( 
.A(n_1385),
.Y(n_1735)
);

BUFx6f_ASAP7_75t_L g1736 ( 
.A(n_1519),
.Y(n_1736)
);

INVx2_ASAP7_75t_SL g1737 ( 
.A(n_1388),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1578),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1581),
.Y(n_1739)
);

NOR2xp67_ASAP7_75t_L g1740 ( 
.A(n_1449),
.B(n_356),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1653),
.B(n_358),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1514),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1547),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1558),
.Y(n_1744)
);

NAND2xp33_ASAP7_75t_R g1745 ( 
.A(n_1520),
.B(n_109),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1517),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1648),
.B(n_110),
.Y(n_1747)
);

BUFx3_ASAP7_75t_L g1748 ( 
.A(n_1580),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1416),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1427),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1429),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1378),
.Y(n_1752)
);

AOI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1487),
.A2(n_361),
.B(n_359),
.Y(n_1753)
);

CKINVDCx20_ASAP7_75t_R g1754 ( 
.A(n_1421),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_1374),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1431),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1434),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1435),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1453),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1477),
.Y(n_1760)
);

CKINVDCx20_ASAP7_75t_R g1761 ( 
.A(n_1428),
.Y(n_1761)
);

AOI21xp5_ASAP7_75t_L g1762 ( 
.A1(n_1487),
.A2(n_365),
.B(n_363),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_L g1763 ( 
.A(n_1595),
.B(n_111),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1399),
.Y(n_1764)
);

AND2x2_ASAP7_75t_SL g1765 ( 
.A(n_1646),
.B(n_111),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_1689),
.Y(n_1766)
);

INVx2_ASAP7_75t_SL g1767 ( 
.A(n_1395),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1407),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1482),
.Y(n_1769)
);

CKINVDCx20_ASAP7_75t_R g1770 ( 
.A(n_1366),
.Y(n_1770)
);

XOR2xp5_ASAP7_75t_L g1771 ( 
.A(n_1699),
.B(n_367),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1409),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1451),
.B(n_1401),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1502),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1509),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1412),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_1599),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1510),
.B(n_1515),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1381),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1389),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1396),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1411),
.Y(n_1782)
);

BUFx3_ASAP7_75t_L g1783 ( 
.A(n_1640),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1415),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1433),
.Y(n_1785)
);

OAI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1527),
.A2(n_371),
.B(n_369),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1438),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1521),
.B(n_373),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1604),
.B(n_1621),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1591),
.Y(n_1790)
);

XOR2xp5_ASAP7_75t_L g1791 ( 
.A(n_1379),
.B(n_374),
.Y(n_1791)
);

INVx2_ASAP7_75t_SL g1792 ( 
.A(n_1402),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1454),
.Y(n_1793)
);

CKINVDCx20_ASAP7_75t_R g1794 ( 
.A(n_1669),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_1700),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1410),
.B(n_112),
.Y(n_1796)
);

XNOR2x1_ASAP7_75t_L g1797 ( 
.A(n_1613),
.B(n_113),
.Y(n_1797)
);

XOR2xp5_ASAP7_75t_L g1798 ( 
.A(n_1459),
.B(n_375),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1467),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1417),
.B(n_113),
.Y(n_1800)
);

NOR2xp33_ASAP7_75t_L g1801 ( 
.A(n_1629),
.B(n_114),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1468),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1418),
.B(n_115),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1469),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1478),
.Y(n_1805)
);

NAND2xp33_ASAP7_75t_R g1806 ( 
.A(n_1386),
.B(n_1603),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1480),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1484),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1422),
.B(n_116),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1495),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1450),
.B(n_116),
.Y(n_1811)
);

AND2x4_ASAP7_75t_L g1812 ( 
.A(n_1461),
.B(n_377),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_SL g1813 ( 
.A(n_1375),
.B(n_117),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1526),
.B(n_381),
.Y(n_1814)
);

INVxp67_ASAP7_75t_SL g1815 ( 
.A(n_1513),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1508),
.Y(n_1816)
);

AND2x4_ASAP7_75t_L g1817 ( 
.A(n_1367),
.B(n_383),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_1661),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1588),
.Y(n_1819)
);

XNOR2xp5_ASAP7_75t_L g1820 ( 
.A(n_1425),
.B(n_118),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1589),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1594),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1590),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1597),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1608),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1618),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1598),
.Y(n_1827)
);

CKINVDCx20_ASAP7_75t_R g1828 ( 
.A(n_1612),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1619),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1623),
.Y(n_1830)
);

AND2x2_ASAP7_75t_SL g1831 ( 
.A(n_1397),
.B(n_119),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1630),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1633),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1649),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1677),
.Y(n_1835)
);

INVx3_ASAP7_75t_R g1836 ( 
.A(n_1496),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1535),
.B(n_384),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1680),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1424),
.B(n_119),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1542),
.B(n_1552),
.Y(n_1840)
);

NAND2xp33_ASAP7_75t_R g1841 ( 
.A(n_1390),
.B(n_120),
.Y(n_1841)
);

INVx2_ASAP7_75t_SL g1842 ( 
.A(n_1500),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1698),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1602),
.Y(n_1844)
);

CKINVDCx20_ASAP7_75t_R g1845 ( 
.A(n_1584),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1635),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1554),
.B(n_388),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1466),
.B(n_122),
.Y(n_1848)
);

INVxp33_ASAP7_75t_L g1849 ( 
.A(n_1370),
.Y(n_1849)
);

INVxp33_ASAP7_75t_L g1850 ( 
.A(n_1492),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1636),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1647),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1650),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1637),
.B(n_122),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1474),
.B(n_125),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1667),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1671),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1678),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_SL g1859 ( 
.A(n_1504),
.B(n_125),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1475),
.B(n_129),
.Y(n_1860)
);

NAND2xp33_ASAP7_75t_SL g1861 ( 
.A(n_1442),
.B(n_130),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1592),
.B(n_130),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1688),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1498),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1511),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1663),
.Y(n_1866)
);

CKINVDCx20_ASAP7_75t_R g1867 ( 
.A(n_1585),
.Y(n_1867)
);

XOR2xp5_ASAP7_75t_L g1868 ( 
.A(n_1440),
.B(n_392),
.Y(n_1868)
);

AND2x4_ASAP7_75t_L g1869 ( 
.A(n_1582),
.B(n_396),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1376),
.Y(n_1870)
);

CKINVDCx20_ASAP7_75t_R g1871 ( 
.A(n_1586),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1609),
.B(n_131),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1376),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1676),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1676),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1668),
.B(n_131),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1488),
.B(n_134),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1682),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1682),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1632),
.B(n_135),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1532),
.Y(n_1881)
);

NOR2xp33_ASAP7_75t_L g1882 ( 
.A(n_1596),
.B(n_136),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1533),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1533),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1471),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1651),
.B(n_138),
.Y(n_1886)
);

AND2x4_ASAP7_75t_L g1887 ( 
.A(n_1507),
.B(n_1541),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1493),
.Y(n_1888)
);

AND2x4_ASAP7_75t_L g1889 ( 
.A(n_1507),
.B(n_398),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1493),
.Y(n_1890)
);

INVx4_ASAP7_75t_L g1891 ( 
.A(n_1523),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1490),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1654),
.B(n_139),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1497),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1557),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1541),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1572),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1572),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1393),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1548),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1548),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1553),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1553),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1383),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1666),
.B(n_139),
.Y(n_1905)
);

CKINVDCx20_ASAP7_75t_R g1906 ( 
.A(n_1600),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1406),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1383),
.Y(n_1908)
);

AOI21x1_ASAP7_75t_L g1909 ( 
.A1(n_1683),
.A2(n_402),
.B(n_399),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1423),
.Y(n_1910)
);

XOR2xp5_ASAP7_75t_L g1911 ( 
.A(n_1655),
.B(n_403),
.Y(n_1911)
);

CKINVDCx16_ASAP7_75t_R g1912 ( 
.A(n_1372),
.Y(n_1912)
);

XOR2xp5_ASAP7_75t_L g1913 ( 
.A(n_1659),
.B(n_405),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1670),
.B(n_140),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1384),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1556),
.B(n_406),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1569),
.B(n_407),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1392),
.B(n_140),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_L g1919 ( 
.A(n_1605),
.B(n_1606),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1681),
.B(n_141),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1687),
.Y(n_1921)
);

INVx2_ASAP7_75t_SL g1922 ( 
.A(n_1660),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1583),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1583),
.Y(n_1924)
);

BUFx3_ASAP7_75t_L g1925 ( 
.A(n_1695),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1534),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1534),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1544),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1544),
.Y(n_1929)
);

INVx1_ASAP7_75t_SL g1930 ( 
.A(n_1413),
.Y(n_1930)
);

INVxp33_ASAP7_75t_L g1931 ( 
.A(n_1439),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1472),
.Y(n_1932)
);

NOR2xp33_ASAP7_75t_L g1933 ( 
.A(n_1614),
.B(n_1622),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1377),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1673),
.B(n_409),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1400),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_SL g1937 ( 
.A(n_1368),
.B(n_141),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1414),
.Y(n_1938)
);

NOR2xp33_ASAP7_75t_L g1939 ( 
.A(n_1625),
.B(n_143),
.Y(n_1939)
);

AND2x2_ASAP7_75t_SL g1940 ( 
.A(n_1679),
.B(n_143),
.Y(n_1940)
);

INVx1_ASAP7_75t_SL g1941 ( 
.A(n_1522),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1420),
.B(n_144),
.Y(n_1942)
);

NAND2x1p5_ASAP7_75t_L g1943 ( 
.A(n_1696),
.B(n_1701),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1400),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1419),
.Y(n_1945)
);

XOR2x2_ASAP7_75t_L g1946 ( 
.A(n_1607),
.B(n_145),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1419),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1420),
.B(n_145),
.Y(n_1948)
);

CKINVDCx20_ASAP7_75t_R g1949 ( 
.A(n_1638),
.Y(n_1949)
);

INVx2_ASAP7_75t_SL g1950 ( 
.A(n_1537),
.Y(n_1950)
);

INVx2_ASAP7_75t_SL g1951 ( 
.A(n_1390),
.Y(n_1951)
);

BUFx8_ASAP7_75t_L g1952 ( 
.A(n_1447),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1426),
.Y(n_1953)
);

AOI21xp5_ASAP7_75t_L g1954 ( 
.A1(n_1479),
.A2(n_412),
.B(n_410),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1530),
.B(n_1549),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1426),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1479),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1494),
.Y(n_1958)
);

NOR2xp33_ASAP7_75t_L g1959 ( 
.A(n_1641),
.B(n_146),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1452),
.B(n_146),
.Y(n_1960)
);

NOR2x1p5_ASAP7_75t_L g1961 ( 
.A(n_1464),
.B(n_149),
.Y(n_1961)
);

INVx5_ASAP7_75t_L g1962 ( 
.A(n_1372),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1494),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1499),
.Y(n_1964)
);

INVx2_ASAP7_75t_SL g1965 ( 
.A(n_1499),
.Y(n_1965)
);

BUFx8_ASAP7_75t_L g1966 ( 
.A(n_1691),
.Y(n_1966)
);

BUFx3_ASAP7_75t_L g1967 ( 
.A(n_1573),
.Y(n_1967)
);

XOR2x2_ASAP7_75t_L g1968 ( 
.A(n_1611),
.B(n_150),
.Y(n_1968)
);

BUFx6f_ASAP7_75t_L g1969 ( 
.A(n_1658),
.Y(n_1969)
);

XOR2xp5_ASAP7_75t_L g1970 ( 
.A(n_1476),
.B(n_414),
.Y(n_1970)
);

NOR2xp33_ASAP7_75t_L g1971 ( 
.A(n_1644),
.B(n_152),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1501),
.Y(n_1972)
);

OR2x2_ASAP7_75t_SL g1973 ( 
.A(n_1627),
.B(n_153),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1501),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1512),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1512),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1516),
.Y(n_1977)
);

INVxp33_ASAP7_75t_L g1978 ( 
.A(n_1503),
.Y(n_1978)
);

NOR2xp33_ASAP7_75t_L g1979 ( 
.A(n_1657),
.B(n_153),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1516),
.Y(n_1980)
);

XOR2xp5_ASAP7_75t_L g1981 ( 
.A(n_1481),
.B(n_416),
.Y(n_1981)
);

CKINVDCx20_ASAP7_75t_R g1982 ( 
.A(n_1672),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_SL g1983 ( 
.A(n_1489),
.B(n_154),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1518),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1555),
.B(n_419),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1455),
.B(n_154),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1518),
.Y(n_1987)
);

INVx2_ASAP7_75t_SL g1988 ( 
.A(n_1398),
.Y(n_1988)
);

AOI21xp5_ASAP7_75t_L g1989 ( 
.A1(n_1473),
.A2(n_421),
.B(n_420),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1456),
.B(n_155),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1437),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1437),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1445),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1445),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1458),
.B(n_156),
.Y(n_1995)
);

XOR2xp5_ASAP7_75t_L g1996 ( 
.A(n_1483),
.B(n_422),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1446),
.Y(n_1997)
);

NOR2xp33_ASAP7_75t_L g1998 ( 
.A(n_1579),
.B(n_1601),
.Y(n_1998)
);

INVx2_ASAP7_75t_SL g1999 ( 
.A(n_1398),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1462),
.B(n_156),
.Y(n_2000)
);

OAI21xp5_ASAP7_75t_L g2001 ( 
.A1(n_1568),
.A2(n_424),
.B(n_423),
.Y(n_2001)
);

NOR2xp33_ASAP7_75t_L g2002 ( 
.A(n_1652),
.B(n_158),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1446),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1380),
.Y(n_2004)
);

OR2x2_ASAP7_75t_L g2005 ( 
.A(n_1441),
.B(n_159),
.Y(n_2005)
);

BUFx3_ASAP7_75t_L g2006 ( 
.A(n_1551),
.Y(n_2006)
);

CKINVDCx5p33_ASAP7_75t_R g2007 ( 
.A(n_1645),
.Y(n_2007)
);

AND2x6_ASAP7_75t_L g2008 ( 
.A(n_1570),
.B(n_432),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1380),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1685),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1692),
.Y(n_2011)
);

XOR2xp5_ASAP7_75t_L g2012 ( 
.A(n_1485),
.B(n_433),
.Y(n_2012)
);

NOR2xp33_ASAP7_75t_L g2013 ( 
.A(n_1665),
.B(n_159),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1463),
.B(n_161),
.Y(n_2014)
);

OR2x6_ASAP7_75t_L g2015 ( 
.A(n_1658),
.B(n_162),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1525),
.B(n_162),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1564),
.Y(n_2017)
);

CKINVDCx20_ASAP7_75t_R g2018 ( 
.A(n_1506),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1560),
.B(n_436),
.Y(n_2019)
);

INVxp67_ASAP7_75t_SL g2020 ( 
.A(n_1571),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1564),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1697),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1694),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1369),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1752),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1778),
.B(n_1528),
.Y(n_2026)
);

AND2x4_ASAP7_75t_L g2027 ( 
.A(n_1881),
.B(n_1639),
.Y(n_2027)
);

CKINVDCx5p33_ASAP7_75t_R g2028 ( 
.A(n_1755),
.Y(n_2028)
);

NOR2xp33_ASAP7_75t_L g2029 ( 
.A(n_1702),
.B(n_1408),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1764),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1921),
.B(n_1529),
.Y(n_2031)
);

NAND2x1p5_ASAP7_75t_L g2032 ( 
.A(n_1748),
.B(n_1430),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1863),
.Y(n_2033)
);

AND2x4_ASAP7_75t_L g2034 ( 
.A(n_1885),
.B(n_1664),
.Y(n_2034)
);

INVxp67_ASAP7_75t_L g2035 ( 
.A(n_1806),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1768),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1863),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1772),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1704),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1704),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1776),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1925),
.B(n_1391),
.Y(n_2042)
);

BUFx6f_ASAP7_75t_L g2043 ( 
.A(n_1736),
.Y(n_2043)
);

INVx2_ASAP7_75t_SL g2044 ( 
.A(n_1842),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1773),
.B(n_1369),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1710),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1710),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1840),
.B(n_1403),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1790),
.Y(n_2049)
);

BUFx3_ASAP7_75t_L g2050 ( 
.A(n_1783),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1735),
.B(n_1664),
.Y(n_2051)
);

AND2x2_ASAP7_75t_SL g2052 ( 
.A(n_1765),
.B(n_1613),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1846),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1943),
.B(n_1486),
.Y(n_2054)
);

AND2x4_ASAP7_75t_L g2055 ( 
.A(n_1932),
.B(n_439),
.Y(n_2055)
);

BUFx3_ASAP7_75t_L g2056 ( 
.A(n_1736),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1851),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1852),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_1737),
.B(n_1562),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_SL g2060 ( 
.A(n_1767),
.B(n_1491),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1853),
.Y(n_2061)
);

NOR2xp67_ASAP7_75t_L g2062 ( 
.A(n_1777),
.B(n_441),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_SL g2063 ( 
.A(n_1792),
.B(n_1869),
.Y(n_2063)
);

AND2x2_ASAP7_75t_SL g2064 ( 
.A(n_1831),
.B(n_1813),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1856),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1822),
.Y(n_2066)
);

OAI21xp5_ASAP7_75t_L g2067 ( 
.A1(n_1998),
.A2(n_1505),
.B(n_1470),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1899),
.B(n_1432),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1827),
.Y(n_2069)
);

OAI21xp5_ASAP7_75t_L g2070 ( 
.A1(n_1919),
.A2(n_1444),
.B(n_1559),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1844),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1857),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1858),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_1733),
.B(n_1617),
.Y(n_2074)
);

INVx1_ASAP7_75t_SL g2075 ( 
.A(n_1794),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1869),
.B(n_1394),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_1815),
.B(n_1617),
.Y(n_2077)
);

INVx3_ASAP7_75t_L g2078 ( 
.A(n_1725),
.Y(n_2078)
);

OAI21xp5_ASAP7_75t_L g2079 ( 
.A1(n_1933),
.A2(n_1460),
.B(n_1686),
.Y(n_2079)
);

NOR2xp33_ASAP7_75t_L g2080 ( 
.A(n_1931),
.B(n_1404),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1712),
.Y(n_2081)
);

AND2x4_ASAP7_75t_L g2082 ( 
.A(n_1907),
.B(n_442),
.Y(n_2082)
);

AND2x2_ASAP7_75t_SL g2083 ( 
.A(n_1940),
.B(n_1626),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_1934),
.B(n_1626),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_1938),
.B(n_1631),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1712),
.Y(n_2086)
);

AND2x6_ASAP7_75t_L g2087 ( 
.A(n_1904),
.B(n_1631),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1713),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1713),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_1894),
.B(n_1567),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_1887),
.B(n_1642),
.Y(n_2091)
);

AND2x4_ASAP7_75t_L g2092 ( 
.A(n_1910),
.B(n_443),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_SL g2093 ( 
.A(n_1740),
.B(n_1955),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_1887),
.B(n_1642),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1743),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1744),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1728),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1731),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1742),
.Y(n_2099)
);

INVx4_ASAP7_75t_L g2100 ( 
.A(n_1736),
.Y(n_2100)
);

AND2x4_ASAP7_75t_L g2101 ( 
.A(n_1902),
.B(n_444),
.Y(n_2101)
);

HB1xp67_ASAP7_75t_L g2102 ( 
.A(n_1915),
.Y(n_2102)
);

NOR2xp33_ASAP7_75t_L g2103 ( 
.A(n_1895),
.B(n_1457),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1734),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_1930),
.B(n_1643),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_1891),
.B(n_1643),
.Y(n_2106)
);

INVxp67_ASAP7_75t_SL g2107 ( 
.A(n_1715),
.Y(n_2107)
);

INVx1_ASAP7_75t_SL g2108 ( 
.A(n_1811),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_1891),
.B(n_1656),
.Y(n_2109)
);

NOR2xp33_ASAP7_75t_SL g2110 ( 
.A(n_1818),
.B(n_1690),
.Y(n_2110)
);

BUFx6f_ASAP7_75t_L g2111 ( 
.A(n_1879),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1738),
.Y(n_2112)
);

AND2x2_ASAP7_75t_SL g2113 ( 
.A(n_1706),
.B(n_1656),
.Y(n_2113)
);

INVx4_ASAP7_75t_L g2114 ( 
.A(n_1812),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_1848),
.B(n_1531),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_1855),
.B(n_1543),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1739),
.Y(n_2117)
);

NOR2xp33_ASAP7_75t_L g2118 ( 
.A(n_1941),
.B(n_1387),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1749),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1750),
.Y(n_2120)
);

BUFx6f_ASAP7_75t_L g2121 ( 
.A(n_1812),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1751),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_1892),
.B(n_1662),
.Y(n_2123)
);

INVx3_ASAP7_75t_L g2124 ( 
.A(n_1817),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_1707),
.B(n_1662),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_1756),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_1960),
.B(n_1674),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1860),
.B(n_1546),
.Y(n_2128)
);

HB1xp67_ASAP7_75t_L g2129 ( 
.A(n_1965),
.Y(n_2129)
);

INVx3_ASAP7_75t_L g2130 ( 
.A(n_1817),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1757),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1758),
.Y(n_2132)
);

INVx4_ASAP7_75t_L g2133 ( 
.A(n_1889),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1709),
.B(n_1574),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1759),
.Y(n_2135)
);

INVx1_ASAP7_75t_SL g2136 ( 
.A(n_1795),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_1760),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_1986),
.B(n_1674),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1769),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1774),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1775),
.Y(n_2141)
);

AND2x4_ASAP7_75t_L g2142 ( 
.A(n_1732),
.B(n_447),
.Y(n_2142)
);

CKINVDCx5p33_ASAP7_75t_R g2143 ( 
.A(n_1766),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1718),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_1990),
.B(n_1684),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_1995),
.B(n_1684),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_1723),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_1724),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1709),
.B(n_1693),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_2000),
.B(n_1693),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_1727),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_2014),
.B(n_163),
.Y(n_2152)
);

INVx4_ASAP7_75t_L g2153 ( 
.A(n_1889),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_1709),
.B(n_448),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1709),
.B(n_450),
.Y(n_2155)
);

OR2x2_ASAP7_75t_L g2156 ( 
.A(n_1991),
.B(n_1675),
.Y(n_2156)
);

AND2x4_ASAP7_75t_L g2157 ( 
.A(n_1957),
.B(n_455),
.Y(n_2157)
);

HB1xp67_ASAP7_75t_L g2158 ( 
.A(n_1908),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_1942),
.B(n_163),
.Y(n_2159)
);

HB1xp67_ASAP7_75t_L g2160 ( 
.A(n_2004),
.Y(n_2160)
);

AND2x4_ASAP7_75t_L g2161 ( 
.A(n_1900),
.B(n_456),
.Y(n_2161)
);

HB1xp67_ASAP7_75t_L g2162 ( 
.A(n_2004),
.Y(n_2162)
);

HB1xp67_ASAP7_75t_L g2163 ( 
.A(n_2009),
.Y(n_2163)
);

AND2x4_ASAP7_75t_L g2164 ( 
.A(n_1901),
.B(n_458),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_1948),
.B(n_2016),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_1709),
.B(n_463),
.Y(n_2166)
);

INVx4_ASAP7_75t_L g2167 ( 
.A(n_1705),
.Y(n_2167)
);

AND2x6_ASAP7_75t_L g2168 ( 
.A(n_1926),
.B(n_466),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_1796),
.B(n_1800),
.Y(n_2169)
);

INVx3_ASAP7_75t_SL g2170 ( 
.A(n_1717),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_1746),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2006),
.B(n_1888),
.Y(n_2172)
);

INVx2_ASAP7_75t_SL g2173 ( 
.A(n_1720),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_1890),
.B(n_164),
.Y(n_2174)
);

INVxp67_ASAP7_75t_L g2175 ( 
.A(n_1789),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_1896),
.B(n_164),
.Y(n_2176)
);

OAI21xp5_ASAP7_75t_L g2177 ( 
.A1(n_2009),
.A2(n_473),
.B(n_470),
.Y(n_2177)
);

INVx3_ASAP7_75t_L g2178 ( 
.A(n_1779),
.Y(n_2178)
);

OAI21xp5_ASAP7_75t_L g2179 ( 
.A1(n_1903),
.A2(n_478),
.B(n_474),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_1780),
.Y(n_2180)
);

INVx3_ASAP7_75t_L g2181 ( 
.A(n_1781),
.Y(n_2181)
);

INVx3_ASAP7_75t_L g2182 ( 
.A(n_1782),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_1721),
.B(n_165),
.Y(n_2183)
);

BUFx4f_ASAP7_75t_L g2184 ( 
.A(n_1969),
.Y(n_2184)
);

AND2x4_ASAP7_75t_L g2185 ( 
.A(n_1972),
.B(n_481),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1784),
.Y(n_2186)
);

INVxp67_ASAP7_75t_L g2187 ( 
.A(n_1841),
.Y(n_2187)
);

INVx8_ASAP7_75t_L g2188 ( 
.A(n_1962),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_SL g2189 ( 
.A(n_1877),
.B(n_167),
.Y(n_2189)
);

INVx1_ASAP7_75t_SL g2190 ( 
.A(n_2005),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_1803),
.B(n_482),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1785),
.Y(n_2192)
);

AND2x2_ASAP7_75t_L g2193 ( 
.A(n_2022),
.B(n_167),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_2022),
.B(n_2024),
.Y(n_2194)
);

INVxp67_ASAP7_75t_L g2195 ( 
.A(n_1801),
.Y(n_2195)
);

BUFx3_ASAP7_75t_L g2196 ( 
.A(n_1870),
.Y(n_2196)
);

AND2x4_ASAP7_75t_L g2197 ( 
.A(n_1936),
.B(n_483),
.Y(n_2197)
);

INVx3_ASAP7_75t_L g2198 ( 
.A(n_1787),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_1988),
.B(n_168),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_1809),
.B(n_484),
.Y(n_2200)
);

BUFx6f_ASAP7_75t_L g2201 ( 
.A(n_1873),
.Y(n_2201)
);

INVxp67_ASAP7_75t_L g2202 ( 
.A(n_1854),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_1999),
.B(n_169),
.Y(n_2203)
);

NOR2xp33_ASAP7_75t_R g2204 ( 
.A(n_1708),
.B(n_486),
.Y(n_2204)
);

AND2x4_ASAP7_75t_L g2205 ( 
.A(n_1865),
.B(n_487),
.Y(n_2205)
);

NOR2xp33_ASAP7_75t_L g2206 ( 
.A(n_1850),
.B(n_169),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_1793),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_1799),
.Y(n_2208)
);

AND2x2_ASAP7_75t_L g2209 ( 
.A(n_2010),
.B(n_170),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_1839),
.B(n_488),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_1802),
.Y(n_2211)
);

NOR2xp33_ASAP7_75t_L g2212 ( 
.A(n_1978),
.B(n_170),
.Y(n_2212)
);

AND2x4_ASAP7_75t_L g2213 ( 
.A(n_1950),
.B(n_489),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1804),
.Y(n_2214)
);

AND2x2_ASAP7_75t_SL g2215 ( 
.A(n_1711),
.B(n_171),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_2010),
.B(n_171),
.Y(n_2216)
);

OAI21xp5_ASAP7_75t_L g2217 ( 
.A1(n_1786),
.A2(n_500),
.B(n_493),
.Y(n_2217)
);

INVx4_ASAP7_75t_L g2218 ( 
.A(n_2008),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1805),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_2011),
.B(n_172),
.Y(n_2220)
);

INVx4_ASAP7_75t_L g2221 ( 
.A(n_2008),
.Y(n_2221)
);

HB1xp67_ASAP7_75t_L g2222 ( 
.A(n_1922),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1807),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_2011),
.B(n_172),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1808),
.Y(n_2225)
);

OAI21xp5_ASAP7_75t_L g2226 ( 
.A1(n_1927),
.A2(n_503),
.B(n_502),
.Y(n_2226)
);

AND2x4_ASAP7_75t_L g2227 ( 
.A(n_1864),
.B(n_504),
.Y(n_2227)
);

NOR2xp67_ASAP7_75t_L g2228 ( 
.A(n_1985),
.B(n_505),
.Y(n_2228)
);

INVxp67_ASAP7_75t_L g2229 ( 
.A(n_1876),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1810),
.Y(n_2230)
);

BUFx6f_ASAP7_75t_L g2231 ( 
.A(n_1874),
.Y(n_2231)
);

INVx4_ASAP7_75t_L g2232 ( 
.A(n_2008),
.Y(n_2232)
);

BUFx6f_ASAP7_75t_L g2233 ( 
.A(n_1875),
.Y(n_2233)
);

CKINVDCx5p33_ASAP7_75t_R g2234 ( 
.A(n_1952),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_1862),
.B(n_506),
.Y(n_2235)
);

OR2x6_ASAP7_75t_L g2236 ( 
.A(n_1722),
.B(n_174),
.Y(n_2236)
);

AND2x4_ASAP7_75t_L g2237 ( 
.A(n_1866),
.B(n_507),
.Y(n_2237)
);

AND2x4_ASAP7_75t_L g2238 ( 
.A(n_1928),
.B(n_508),
.Y(n_2238)
);

NOR2xp33_ASAP7_75t_L g2239 ( 
.A(n_1967),
.B(n_2017),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1816),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1819),
.Y(n_2241)
);

INVx3_ASAP7_75t_L g2242 ( 
.A(n_1821),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_1993),
.B(n_174),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_1823),
.Y(n_2244)
);

HB1xp67_ASAP7_75t_L g2245 ( 
.A(n_1992),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_1872),
.B(n_509),
.Y(n_2246)
);

INVx3_ASAP7_75t_L g2247 ( 
.A(n_1824),
.Y(n_2247)
);

INVx3_ASAP7_75t_L g2248 ( 
.A(n_1825),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_1994),
.B(n_175),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_1880),
.B(n_512),
.Y(n_2250)
);

BUFx8_ASAP7_75t_L g2251 ( 
.A(n_1969),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_1886),
.B(n_515),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_1997),
.B(n_177),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_1893),
.B(n_519),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1826),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_1905),
.B(n_524),
.Y(n_2256)
);

HB1xp67_ASAP7_75t_L g2257 ( 
.A(n_2021),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_2003),
.B(n_2023),
.Y(n_2258)
);

NOR2xp33_ASAP7_75t_L g2259 ( 
.A(n_2017),
.B(n_177),
.Y(n_2259)
);

AND2x2_ASAP7_75t_SL g2260 ( 
.A(n_1716),
.B(n_178),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_1914),
.B(n_527),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_1929),
.B(n_528),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_SL g2263 ( 
.A(n_1882),
.B(n_178),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1829),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2023),
.B(n_179),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1830),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_SL g2267 ( 
.A(n_1939),
.B(n_179),
.Y(n_2267)
);

AND2x6_ASAP7_75t_L g2268 ( 
.A(n_1923),
.B(n_530),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_SL g2269 ( 
.A(n_1959),
.B(n_180),
.Y(n_2269)
);

BUFx6f_ASAP7_75t_L g2270 ( 
.A(n_1878),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_2081),
.Y(n_2271)
);

OR2x2_ASAP7_75t_L g2272 ( 
.A(n_2190),
.B(n_1944),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2257),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2129),
.Y(n_2274)
);

OR2x6_ASAP7_75t_L g2275 ( 
.A(n_2188),
.B(n_1951),
.Y(n_2275)
);

INVxp67_ASAP7_75t_L g2276 ( 
.A(n_2222),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2029),
.B(n_1747),
.Y(n_2277)
);

NOR2xp33_ASAP7_75t_SL g2278 ( 
.A(n_2028),
.B(n_2143),
.Y(n_2278)
);

AND2x6_ASAP7_75t_L g2279 ( 
.A(n_2082),
.B(n_1924),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2102),
.Y(n_2280)
);

OR2x2_ASAP7_75t_L g2281 ( 
.A(n_2035),
.B(n_1945),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_2165),
.B(n_1971),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2039),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2124),
.B(n_1979),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_2025),
.Y(n_2285)
);

AND2x2_ASAP7_75t_L g2286 ( 
.A(n_2108),
.B(n_1947),
.Y(n_2286)
);

INVx5_ASAP7_75t_L g2287 ( 
.A(n_2188),
.Y(n_2287)
);

BUFx6f_ASAP7_75t_L g2288 ( 
.A(n_2043),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_2030),
.Y(n_2289)
);

AND2x4_ASAP7_75t_L g2290 ( 
.A(n_2050),
.B(n_1883),
.Y(n_2290)
);

INVx4_ASAP7_75t_L g2291 ( 
.A(n_2121),
.Y(n_2291)
);

INVx5_ASAP7_75t_L g2292 ( 
.A(n_2043),
.Y(n_2292)
);

BUFx8_ASAP7_75t_SL g2293 ( 
.A(n_2234),
.Y(n_2293)
);

NAND2x1p5_ASAP7_75t_L g2294 ( 
.A(n_2133),
.B(n_1962),
.Y(n_2294)
);

NOR2xp33_ASAP7_75t_SL g2295 ( 
.A(n_2136),
.B(n_1828),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2124),
.B(n_1953),
.Y(n_2296)
);

INVx2_ASAP7_75t_SL g2297 ( 
.A(n_2172),
.Y(n_2297)
);

INVx4_ASAP7_75t_L g2298 ( 
.A(n_2121),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2040),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2046),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2187),
.B(n_1956),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2047),
.Y(n_2302)
);

NAND2x1p5_ASAP7_75t_L g2303 ( 
.A(n_2133),
.B(n_1962),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_2036),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_2044),
.B(n_1958),
.Y(n_2305)
);

AND2x4_ASAP7_75t_L g2306 ( 
.A(n_2194),
.B(n_1884),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2130),
.B(n_1963),
.Y(n_2307)
);

BUFx6f_ASAP7_75t_L g2308 ( 
.A(n_2043),
.Y(n_2308)
);

NAND2x1p5_ASAP7_75t_L g2309 ( 
.A(n_2153),
.B(n_1964),
.Y(n_2309)
);

INVx4_ASAP7_75t_L g2310 ( 
.A(n_2121),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2038),
.Y(n_2311)
);

AND2x4_ASAP7_75t_L g2312 ( 
.A(n_2196),
.B(n_1897),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2033),
.Y(n_2313)
);

CKINVDCx14_ASAP7_75t_R g2314 ( 
.A(n_2204),
.Y(n_2314)
);

NAND2x1p5_ASAP7_75t_L g2315 ( 
.A(n_2153),
.B(n_1974),
.Y(n_2315)
);

NOR2xp33_ASAP7_75t_L g2316 ( 
.A(n_2026),
.B(n_1849),
.Y(n_2316)
);

NOR2x1p5_ASAP7_75t_SL g2317 ( 
.A(n_2041),
.B(n_1909),
.Y(n_2317)
);

AND2x4_ASAP7_75t_L g2318 ( 
.A(n_2213),
.B(n_1898),
.Y(n_2318)
);

NAND2x1p5_ASAP7_75t_L g2319 ( 
.A(n_2114),
.B(n_1975),
.Y(n_2319)
);

AND2x6_ASAP7_75t_L g2320 ( 
.A(n_2082),
.B(n_1976),
.Y(n_2320)
);

AND2x4_ASAP7_75t_L g2321 ( 
.A(n_2213),
.B(n_1977),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2037),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2086),
.Y(n_2323)
);

NAND2x1_ASAP7_75t_L g2324 ( 
.A(n_2114),
.B(n_1832),
.Y(n_2324)
);

AND2x4_ASAP7_75t_L g2325 ( 
.A(n_2056),
.B(n_1980),
.Y(n_2325)
);

INVxp67_ASAP7_75t_L g2326 ( 
.A(n_2239),
.Y(n_2326)
);

NOR2xp33_ASAP7_75t_SL g2327 ( 
.A(n_2064),
.B(n_1912),
.Y(n_2327)
);

BUFx4f_ASAP7_75t_L g2328 ( 
.A(n_2170),
.Y(n_2328)
);

BUFx2_ASAP7_75t_L g2329 ( 
.A(n_2175),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2130),
.B(n_1984),
.Y(n_2330)
);

INVx8_ASAP7_75t_L g2331 ( 
.A(n_2268),
.Y(n_2331)
);

BUFx6f_ASAP7_75t_L g2332 ( 
.A(n_2184),
.Y(n_2332)
);

NOR2xp33_ASAP7_75t_SL g2333 ( 
.A(n_2083),
.B(n_2052),
.Y(n_2333)
);

BUFx4f_ASAP7_75t_L g2334 ( 
.A(n_2238),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2088),
.Y(n_2335)
);

NOR2xp33_ASAP7_75t_L g2336 ( 
.A(n_2080),
.B(n_1754),
.Y(n_2336)
);

AND2x4_ASAP7_75t_L g2337 ( 
.A(n_2055),
.B(n_1987),
.Y(n_2337)
);

NOR2xp33_ASAP7_75t_L g2338 ( 
.A(n_2195),
.B(n_1761),
.Y(n_2338)
);

NOR2xp33_ASAP7_75t_L g2339 ( 
.A(n_2202),
.B(n_1714),
.Y(n_2339)
);

BUFx6f_ASAP7_75t_L g2340 ( 
.A(n_2100),
.Y(n_2340)
);

BUFx8_ASAP7_75t_L g2341 ( 
.A(n_2091),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2118),
.B(n_1969),
.Y(n_2342)
);

AO21x2_ASAP7_75t_L g2343 ( 
.A1(n_2217),
.A2(n_2001),
.B(n_1814),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2169),
.B(n_2002),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_2049),
.Y(n_2345)
);

AND2x2_ASAP7_75t_SL g2346 ( 
.A(n_2215),
.B(n_2013),
.Y(n_2346)
);

INVx4_ASAP7_75t_L g2347 ( 
.A(n_2100),
.Y(n_2347)
);

AND2x4_ASAP7_75t_L g2348 ( 
.A(n_2055),
.B(n_1833),
.Y(n_2348)
);

BUFx8_ASAP7_75t_L g2349 ( 
.A(n_2094),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2068),
.B(n_1763),
.Y(n_2350)
);

INVxp67_ASAP7_75t_L g2351 ( 
.A(n_2212),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2092),
.B(n_2019),
.Y(n_2352)
);

BUFx6f_ASAP7_75t_L g2353 ( 
.A(n_2111),
.Y(n_2353)
);

AND2x4_ASAP7_75t_L g2354 ( 
.A(n_2174),
.B(n_1834),
.Y(n_2354)
);

INVx3_ASAP7_75t_L g2355 ( 
.A(n_2111),
.Y(n_2355)
);

BUFx12f_ASAP7_75t_L g2356 ( 
.A(n_2251),
.Y(n_2356)
);

INVx3_ASAP7_75t_L g2357 ( 
.A(n_2111),
.Y(n_2357)
);

INVx6_ASAP7_75t_L g2358 ( 
.A(n_2251),
.Y(n_2358)
);

INVx1_ASAP7_75t_SL g2359 ( 
.A(n_2075),
.Y(n_2359)
);

INVx3_ASAP7_75t_L g2360 ( 
.A(n_2201),
.Y(n_2360)
);

BUFx12f_ASAP7_75t_L g2361 ( 
.A(n_2236),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_2066),
.Y(n_2362)
);

NAND2x1p5_ASAP7_75t_L g2363 ( 
.A(n_2092),
.B(n_1835),
.Y(n_2363)
);

INVx2_ASAP7_75t_SL g2364 ( 
.A(n_2258),
.Y(n_2364)
);

CKINVDCx8_ASAP7_75t_R g2365 ( 
.A(n_2034),
.Y(n_2365)
);

BUFx5_ASAP7_75t_L g2366 ( 
.A(n_2168),
.Y(n_2366)
);

OR2x2_ASAP7_75t_L g2367 ( 
.A(n_2229),
.B(n_1973),
.Y(n_2367)
);

BUFx6f_ASAP7_75t_L g2368 ( 
.A(n_2201),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2048),
.B(n_2020),
.Y(n_2369)
);

NOR2xp33_ASAP7_75t_SL g2370 ( 
.A(n_2260),
.B(n_1845),
.Y(n_2370)
);

BUFx6f_ASAP7_75t_L g2371 ( 
.A(n_2201),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_2173),
.B(n_1859),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_2152),
.B(n_1983),
.Y(n_2373)
);

AND2x4_ASAP7_75t_L g2374 ( 
.A(n_2176),
.B(n_1838),
.Y(n_2374)
);

INVx1_ASAP7_75t_SL g2375 ( 
.A(n_2265),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2067),
.B(n_1719),
.Y(n_2376)
);

AND2x4_ASAP7_75t_L g2377 ( 
.A(n_2144),
.B(n_1843),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_2069),
.Y(n_2378)
);

BUFx2_ASAP7_75t_L g2379 ( 
.A(n_2087),
.Y(n_2379)
);

INVx6_ASAP7_75t_L g2380 ( 
.A(n_2034),
.Y(n_2380)
);

BUFx5_ASAP7_75t_L g2381 ( 
.A(n_2168),
.Y(n_2381)
);

NAND2x1_ASAP7_75t_L g2382 ( 
.A(n_2218),
.B(n_2008),
.Y(n_2382)
);

AND2x4_ASAP7_75t_L g2383 ( 
.A(n_2147),
.B(n_1961),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2101),
.B(n_1741),
.Y(n_2384)
);

OR2x6_ASAP7_75t_L g2385 ( 
.A(n_2236),
.B(n_1722),
.Y(n_2385)
);

AND2x2_ASAP7_75t_L g2386 ( 
.A(n_2059),
.B(n_2015),
.Y(n_2386)
);

BUFx6f_ASAP7_75t_L g2387 ( 
.A(n_2231),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2089),
.Y(n_2388)
);

AND2x2_ASAP7_75t_L g2389 ( 
.A(n_2209),
.B(n_2015),
.Y(n_2389)
);

INVx6_ASAP7_75t_L g2390 ( 
.A(n_2231),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2158),
.Y(n_2391)
);

HB1xp67_ASAP7_75t_L g2392 ( 
.A(n_2245),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_2216),
.B(n_1729),
.Y(n_2393)
);

INVx8_ASAP7_75t_L g2394 ( 
.A(n_2268),
.Y(n_2394)
);

AND2x4_ASAP7_75t_L g2395 ( 
.A(n_2148),
.B(n_2007),
.Y(n_2395)
);

BUFx6f_ASAP7_75t_L g2396 ( 
.A(n_2231),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2186),
.Y(n_2397)
);

OR2x4_ASAP7_75t_L g2398 ( 
.A(n_2206),
.B(n_1797),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_SL g2399 ( 
.A(n_2185),
.B(n_2197),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2192),
.Y(n_2400)
);

BUFx6f_ASAP7_75t_L g2401 ( 
.A(n_2233),
.Y(n_2401)
);

INVx4_ASAP7_75t_L g2402 ( 
.A(n_2142),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2101),
.B(n_1935),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_2185),
.B(n_1788),
.Y(n_2404)
);

CKINVDCx8_ASAP7_75t_R g2405 ( 
.A(n_2087),
.Y(n_2405)
);

NOR2xp33_ASAP7_75t_SL g2406 ( 
.A(n_2218),
.B(n_1952),
.Y(n_2406)
);

INVxp67_ASAP7_75t_L g2407 ( 
.A(n_2103),
.Y(n_2407)
);

NAND2x1p5_ASAP7_75t_L g2408 ( 
.A(n_2197),
.B(n_1937),
.Y(n_2408)
);

INVxp67_ASAP7_75t_SL g2409 ( 
.A(n_2178),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2214),
.Y(n_2410)
);

CKINVDCx5p33_ASAP7_75t_R g2411 ( 
.A(n_2070),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2219),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_2031),
.B(n_2183),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2223),
.Y(n_2414)
);

AND2x2_ASAP7_75t_SL g2415 ( 
.A(n_2113),
.B(n_1868),
.Y(n_2415)
);

AND2x4_ASAP7_75t_L g2416 ( 
.A(n_2151),
.B(n_1918),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2225),
.Y(n_2417)
);

NAND2x1p5_ASAP7_75t_L g2418 ( 
.A(n_2221),
.B(n_1954),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_2071),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2095),
.Y(n_2420)
);

OR2x6_ASAP7_75t_L g2421 ( 
.A(n_2157),
.B(n_1726),
.Y(n_2421)
);

NOR2xp33_ASAP7_75t_L g2422 ( 
.A(n_2110),
.B(n_1770),
.Y(n_2422)
);

INVx2_ASAP7_75t_L g2423 ( 
.A(n_2099),
.Y(n_2423)
);

BUFx2_ASAP7_75t_SL g2424 ( 
.A(n_2062),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2053),
.Y(n_2425)
);

AND2x2_ASAP7_75t_L g2426 ( 
.A(n_2220),
.B(n_1867),
.Y(n_2426)
);

OR2x2_ASAP7_75t_L g2427 ( 
.A(n_2156),
.B(n_1703),
.Y(n_2427)
);

AND2x2_ASAP7_75t_L g2428 ( 
.A(n_2224),
.B(n_1871),
.Y(n_2428)
);

BUFx6f_ASAP7_75t_L g2429 ( 
.A(n_2233),
.Y(n_2429)
);

AOI22xp5_ASAP7_75t_L g2430 ( 
.A1(n_2411),
.A2(n_2093),
.B1(n_1949),
.B2(n_1982),
.Y(n_2430)
);

INVx6_ASAP7_75t_SL g2431 ( 
.A(n_2385),
.Y(n_2431)
);

BUFx12f_ASAP7_75t_L g2432 ( 
.A(n_2356),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2277),
.B(n_2079),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2283),
.Y(n_2434)
);

BUFx4f_ASAP7_75t_L g2435 ( 
.A(n_2332),
.Y(n_2435)
);

INVx1_ASAP7_75t_SL g2436 ( 
.A(n_2359),
.Y(n_2436)
);

INVx2_ASAP7_75t_SL g2437 ( 
.A(n_2332),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2299),
.Y(n_2438)
);

INVxp67_ASAP7_75t_SL g2439 ( 
.A(n_2399),
.Y(n_2439)
);

INVx1_ASAP7_75t_SL g2440 ( 
.A(n_2329),
.Y(n_2440)
);

INVx3_ASAP7_75t_L g2441 ( 
.A(n_2340),
.Y(n_2441)
);

NOR2xp33_ASAP7_75t_L g2442 ( 
.A(n_2407),
.B(n_1906),
.Y(n_2442)
);

BUFx2_ASAP7_75t_L g2443 ( 
.A(n_2342),
.Y(n_2443)
);

CKINVDCx20_ASAP7_75t_R g2444 ( 
.A(n_2293),
.Y(n_2444)
);

BUFx6f_ASAP7_75t_L g2445 ( 
.A(n_2288),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2300),
.Y(n_2446)
);

AND2x2_ASAP7_75t_L g2447 ( 
.A(n_2282),
.B(n_2127),
.Y(n_2447)
);

BUFx6f_ASAP7_75t_L g2448 ( 
.A(n_2288),
.Y(n_2448)
);

CKINVDCx6p67_ASAP7_75t_R g2449 ( 
.A(n_2287),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_2425),
.Y(n_2450)
);

INVxp67_ASAP7_75t_SL g2451 ( 
.A(n_2340),
.Y(n_2451)
);

INVx2_ASAP7_75t_SL g2452 ( 
.A(n_2380),
.Y(n_2452)
);

AOI22xp33_ASAP7_75t_L g2453 ( 
.A1(n_2346),
.A2(n_2263),
.B1(n_2269),
.B2(n_2267),
.Y(n_2453)
);

BUFx12f_ASAP7_75t_L g2454 ( 
.A(n_2358),
.Y(n_2454)
);

NAND2x1p5_ASAP7_75t_L g2455 ( 
.A(n_2292),
.B(n_2221),
.Y(n_2455)
);

INVx3_ASAP7_75t_L g2456 ( 
.A(n_2292),
.Y(n_2456)
);

OR2x6_ASAP7_75t_L g2457 ( 
.A(n_2331),
.B(n_2394),
.Y(n_2457)
);

CKINVDCx11_ASAP7_75t_R g2458 ( 
.A(n_2365),
.Y(n_2458)
);

INVxp67_ASAP7_75t_SL g2459 ( 
.A(n_2368),
.Y(n_2459)
);

BUFx6f_ASAP7_75t_L g2460 ( 
.A(n_2308),
.Y(n_2460)
);

CKINVDCx20_ASAP7_75t_R g2461 ( 
.A(n_2314),
.Y(n_2461)
);

BUFx3_ASAP7_75t_L g2462 ( 
.A(n_2290),
.Y(n_2462)
);

NAND2x1p5_ASAP7_75t_L g2463 ( 
.A(n_2291),
.B(n_2232),
.Y(n_2463)
);

CKINVDCx5p33_ASAP7_75t_R g2464 ( 
.A(n_2328),
.Y(n_2464)
);

INVx1_ASAP7_75t_SL g2465 ( 
.A(n_2272),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_SL g2466 ( 
.A(n_2316),
.B(n_2054),
.Y(n_2466)
);

INVx3_ASAP7_75t_L g2467 ( 
.A(n_2368),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2413),
.B(n_2138),
.Y(n_2468)
);

NOR2x1_ASAP7_75t_R g2469 ( 
.A(n_2287),
.B(n_2105),
.Y(n_2469)
);

CKINVDCx16_ASAP7_75t_R g2470 ( 
.A(n_2278),
.Y(n_2470)
);

NAND2x1p5_ASAP7_75t_L g2471 ( 
.A(n_2298),
.B(n_2232),
.Y(n_2471)
);

CKINVDCx8_ASAP7_75t_R g2472 ( 
.A(n_2395),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2302),
.Y(n_2473)
);

INVx3_ASAP7_75t_L g2474 ( 
.A(n_2371),
.Y(n_2474)
);

NAND2x1p5_ASAP7_75t_L g2475 ( 
.A(n_2310),
.B(n_2178),
.Y(n_2475)
);

BUFx3_ASAP7_75t_L g2476 ( 
.A(n_2341),
.Y(n_2476)
);

INVx8_ASAP7_75t_L g2477 ( 
.A(n_2275),
.Y(n_2477)
);

INVx1_ASAP7_75t_SL g2478 ( 
.A(n_2367),
.Y(n_2478)
);

INVx1_ASAP7_75t_SL g2479 ( 
.A(n_2286),
.Y(n_2479)
);

BUFx5_ASAP7_75t_L g2480 ( 
.A(n_2320),
.Y(n_2480)
);

INVx1_ASAP7_75t_SL g2481 ( 
.A(n_2392),
.Y(n_2481)
);

INVx2_ASAP7_75t_SL g2482 ( 
.A(n_2312),
.Y(n_2482)
);

INVx2_ASAP7_75t_L g2483 ( 
.A(n_2271),
.Y(n_2483)
);

NOR2xp33_ASAP7_75t_L g2484 ( 
.A(n_2351),
.B(n_2145),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2397),
.Y(n_2485)
);

BUFx6f_ASAP7_75t_L g2486 ( 
.A(n_2308),
.Y(n_2486)
);

BUFx12f_ASAP7_75t_L g2487 ( 
.A(n_2361),
.Y(n_2487)
);

CKINVDCx5p33_ASAP7_75t_R g2488 ( 
.A(n_2349),
.Y(n_2488)
);

INVx5_ASAP7_75t_L g2489 ( 
.A(n_2421),
.Y(n_2489)
);

CKINVDCx5p33_ASAP7_75t_R g2490 ( 
.A(n_2339),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2400),
.Y(n_2491)
);

BUFx2_ASAP7_75t_SL g2492 ( 
.A(n_2366),
.Y(n_2492)
);

INVx3_ASAP7_75t_L g2493 ( 
.A(n_2371),
.Y(n_2493)
);

BUFx4f_ASAP7_75t_L g2494 ( 
.A(n_2294),
.Y(n_2494)
);

BUFx6f_ASAP7_75t_L g2495 ( 
.A(n_2306),
.Y(n_2495)
);

BUFx3_ASAP7_75t_L g2496 ( 
.A(n_2391),
.Y(n_2496)
);

BUFx3_ASAP7_75t_L g2497 ( 
.A(n_2274),
.Y(n_2497)
);

INVx3_ASAP7_75t_L g2498 ( 
.A(n_2387),
.Y(n_2498)
);

INVxp67_ASAP7_75t_SL g2499 ( 
.A(n_2387),
.Y(n_2499)
);

BUFx12f_ASAP7_75t_L g2500 ( 
.A(n_2383),
.Y(n_2500)
);

NAND2x1p5_ASAP7_75t_L g2501 ( 
.A(n_2347),
.B(n_2181),
.Y(n_2501)
);

CKINVDCx5p33_ASAP7_75t_R g2502 ( 
.A(n_2338),
.Y(n_2502)
);

INVx3_ASAP7_75t_L g2503 ( 
.A(n_2396),
.Y(n_2503)
);

BUFx8_ASAP7_75t_L g2504 ( 
.A(n_2389),
.Y(n_2504)
);

OR2x2_ASAP7_75t_L g2505 ( 
.A(n_2427),
.B(n_2042),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2410),
.Y(n_2506)
);

BUFx6f_ASAP7_75t_L g2507 ( 
.A(n_2325),
.Y(n_2507)
);

INVx5_ASAP7_75t_L g2508 ( 
.A(n_2301),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2412),
.Y(n_2509)
);

BUFx6f_ASAP7_75t_L g2510 ( 
.A(n_2353),
.Y(n_2510)
);

BUFx6f_ASAP7_75t_L g2511 ( 
.A(n_2353),
.Y(n_2511)
);

BUFx3_ASAP7_75t_L g2512 ( 
.A(n_2280),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2313),
.Y(n_2513)
);

BUFx6f_ASAP7_75t_L g2514 ( 
.A(n_2318),
.Y(n_2514)
);

BUFx6f_ASAP7_75t_L g2515 ( 
.A(n_2396),
.Y(n_2515)
);

BUFx2_ASAP7_75t_SL g2516 ( 
.A(n_2366),
.Y(n_2516)
);

INVx2_ASAP7_75t_L g2517 ( 
.A(n_2322),
.Y(n_2517)
);

AND2x2_ASAP7_75t_L g2518 ( 
.A(n_2350),
.B(n_2344),
.Y(n_2518)
);

BUFx2_ASAP7_75t_L g2519 ( 
.A(n_2279),
.Y(n_2519)
);

INVx3_ASAP7_75t_L g2520 ( 
.A(n_2401),
.Y(n_2520)
);

BUFx3_ASAP7_75t_L g2521 ( 
.A(n_2273),
.Y(n_2521)
);

BUFx2_ASAP7_75t_SL g2522 ( 
.A(n_2366),
.Y(n_2522)
);

BUFx5_ASAP7_75t_L g2523 ( 
.A(n_2320),
.Y(n_2523)
);

BUFx3_ASAP7_75t_L g2524 ( 
.A(n_2305),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2414),
.Y(n_2525)
);

BUFx6f_ASAP7_75t_L g2526 ( 
.A(n_2401),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2417),
.Y(n_2527)
);

AND2x4_ASAP7_75t_L g2528 ( 
.A(n_2297),
.B(n_2051),
.Y(n_2528)
);

AOI22xp33_ASAP7_75t_L g2529 ( 
.A1(n_2453),
.A2(n_2370),
.B1(n_2336),
.B2(n_2422),
.Y(n_2529)
);

AOI22xp33_ASAP7_75t_L g2530 ( 
.A1(n_2443),
.A2(n_2189),
.B1(n_2415),
.B2(n_2386),
.Y(n_2530)
);

INVx6_ASAP7_75t_L g2531 ( 
.A(n_2454),
.Y(n_2531)
);

BUFx10_ASAP7_75t_L g2532 ( 
.A(n_2464),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2485),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2513),
.Y(n_2534)
);

AOI22xp33_ASAP7_75t_L g2535 ( 
.A1(n_2443),
.A2(n_2447),
.B1(n_2505),
.B2(n_2518),
.Y(n_2535)
);

AOI22xp33_ASAP7_75t_SL g2536 ( 
.A1(n_2470),
.A2(n_2393),
.B1(n_2428),
.B2(n_2426),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2491),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2506),
.Y(n_2538)
);

HB1xp67_ASAP7_75t_L g2539 ( 
.A(n_2440),
.Y(n_2539)
);

OAI22xp5_ASAP7_75t_L g2540 ( 
.A1(n_2433),
.A2(n_2334),
.B1(n_2352),
.B2(n_2403),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2509),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2517),
.Y(n_2542)
);

AOI22xp33_ASAP7_75t_L g2543 ( 
.A1(n_2447),
.A2(n_2505),
.B1(n_2518),
.B2(n_2376),
.Y(n_2543)
);

BUFx4f_ASAP7_75t_L g2544 ( 
.A(n_2449),
.Y(n_2544)
);

INVx4_ASAP7_75t_L g2545 ( 
.A(n_2435),
.Y(n_2545)
);

INVx2_ASAP7_75t_SL g2546 ( 
.A(n_2437),
.Y(n_2546)
);

BUFx10_ASAP7_75t_L g2547 ( 
.A(n_2528),
.Y(n_2547)
);

OAI22xp5_ASAP7_75t_L g2548 ( 
.A1(n_2430),
.A2(n_2284),
.B1(n_2402),
.B2(n_2384),
.Y(n_2548)
);

AOI22xp33_ASAP7_75t_L g2549 ( 
.A1(n_2468),
.A2(n_2373),
.B1(n_2018),
.B2(n_2279),
.Y(n_2549)
);

BUFx6f_ASAP7_75t_SL g2550 ( 
.A(n_2476),
.Y(n_2550)
);

AOI22xp33_ASAP7_75t_SL g2551 ( 
.A1(n_2490),
.A2(n_2333),
.B1(n_2327),
.B2(n_2406),
.Y(n_2551)
);

CKINVDCx20_ASAP7_75t_R g2552 ( 
.A(n_2444),
.Y(n_2552)
);

INVx6_ASAP7_75t_L g2553 ( 
.A(n_2504),
.Y(n_2553)
);

AOI22xp33_ASAP7_75t_SL g2554 ( 
.A1(n_2502),
.A2(n_2295),
.B1(n_2150),
.B2(n_2146),
.Y(n_2554)
);

OAI21xp33_ASAP7_75t_L g2555 ( 
.A1(n_2479),
.A2(n_2369),
.B(n_2375),
.Y(n_2555)
);

INVx4_ASAP7_75t_L g2556 ( 
.A(n_2515),
.Y(n_2556)
);

OAI22xp33_ASAP7_75t_L g2557 ( 
.A1(n_2508),
.A2(n_2398),
.B1(n_2326),
.B2(n_1745),
.Y(n_2557)
);

INVx2_ASAP7_75t_SL g2558 ( 
.A(n_2462),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_2525),
.Y(n_2559)
);

INVx6_ASAP7_75t_L g2560 ( 
.A(n_2477),
.Y(n_2560)
);

OAI22xp5_ASAP7_75t_L g2561 ( 
.A1(n_2466),
.A2(n_2404),
.B1(n_2363),
.B2(n_2408),
.Y(n_2561)
);

AOI22xp33_ASAP7_75t_L g2562 ( 
.A1(n_2468),
.A2(n_2279),
.B1(n_2320),
.B2(n_1861),
.Y(n_2562)
);

BUFx4_ASAP7_75t_R g2563 ( 
.A(n_2480),
.Y(n_2563)
);

AOI22xp33_ASAP7_75t_L g2564 ( 
.A1(n_2442),
.A2(n_2343),
.B1(n_1820),
.B2(n_2045),
.Y(n_2564)
);

OAI22xp5_ASAP7_75t_L g2565 ( 
.A1(n_2439),
.A2(n_2405),
.B1(n_2409),
.B2(n_2484),
.Y(n_2565)
);

OAI22xp5_ASAP7_75t_L g2566 ( 
.A1(n_2508),
.A2(n_2116),
.B1(n_2128),
.B2(n_2379),
.Y(n_2566)
);

BUFx6f_ASAP7_75t_L g2567 ( 
.A(n_2445),
.Y(n_2567)
);

CKINVDCx5p33_ASAP7_75t_R g2568 ( 
.A(n_2432),
.Y(n_2568)
);

OAI22xp33_ASAP7_75t_L g2569 ( 
.A1(n_2465),
.A2(n_2364),
.B1(n_2076),
.B2(n_2372),
.Y(n_2569)
);

CKINVDCx20_ASAP7_75t_R g2570 ( 
.A(n_2461),
.Y(n_2570)
);

BUFx6f_ASAP7_75t_L g2571 ( 
.A(n_2445),
.Y(n_2571)
);

INVx6_ASAP7_75t_L g2572 ( 
.A(n_2477),
.Y(n_2572)
);

AOI22xp33_ASAP7_75t_L g2573 ( 
.A1(n_2478),
.A2(n_1968),
.B1(n_1946),
.B2(n_1970),
.Y(n_2573)
);

AOI22xp33_ASAP7_75t_SL g2574 ( 
.A1(n_2496),
.A2(n_2159),
.B1(n_2268),
.B2(n_2168),
.Y(n_2574)
);

AOI22xp33_ASAP7_75t_SL g2575 ( 
.A1(n_2512),
.A2(n_2268),
.B1(n_2168),
.B2(n_2177),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_2527),
.Y(n_2576)
);

BUFx3_ASAP7_75t_L g2577 ( 
.A(n_2472),
.Y(n_2577)
);

INVx6_ASAP7_75t_L g2578 ( 
.A(n_2489),
.Y(n_2578)
);

AOI22xp33_ASAP7_75t_L g2579 ( 
.A1(n_2524),
.A2(n_1996),
.B1(n_2012),
.B2(n_1981),
.Y(n_2579)
);

AOI22xp33_ASAP7_75t_SL g2580 ( 
.A1(n_2521),
.A2(n_2331),
.B1(n_2394),
.B2(n_2226),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2434),
.Y(n_2581)
);

BUFx12f_ASAP7_75t_L g2582 ( 
.A(n_2458),
.Y(n_2582)
);

AOI22xp33_ASAP7_75t_L g2583 ( 
.A1(n_2450),
.A2(n_2179),
.B1(n_2027),
.B2(n_2109),
.Y(n_2583)
);

HB1xp67_ASAP7_75t_L g2584 ( 
.A(n_2481),
.Y(n_2584)
);

INVx3_ASAP7_75t_L g2585 ( 
.A(n_2497),
.Y(n_2585)
);

AOI22xp33_ASAP7_75t_L g2586 ( 
.A1(n_2483),
.A2(n_2027),
.B1(n_2106),
.B2(n_2157),
.Y(n_2586)
);

AOI22xp5_ASAP7_75t_L g2587 ( 
.A1(n_2436),
.A2(n_2354),
.B1(n_2374),
.B2(n_2348),
.Y(n_2587)
);

AOI22xp33_ASAP7_75t_L g2588 ( 
.A1(n_2438),
.A2(n_2074),
.B1(n_2123),
.B2(n_2161),
.Y(n_2588)
);

AOI22xp33_ASAP7_75t_L g2589 ( 
.A1(n_2446),
.A2(n_2164),
.B1(n_2161),
.B2(n_2337),
.Y(n_2589)
);

INVx1_ASAP7_75t_SL g2590 ( 
.A(n_2482),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2473),
.Y(n_2591)
);

BUFx3_ASAP7_75t_L g2592 ( 
.A(n_2495),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2459),
.Y(n_2593)
);

OAI22xp5_ASAP7_75t_L g2594 ( 
.A1(n_2519),
.A2(n_2424),
.B1(n_2382),
.B2(n_2296),
.Y(n_2594)
);

CKINVDCx6p67_ASAP7_75t_R g2595 ( 
.A(n_2489),
.Y(n_2595)
);

CKINVDCx11_ASAP7_75t_R g2596 ( 
.A(n_2487),
.Y(n_2596)
);

OAI21xp5_ASAP7_75t_SL g2597 ( 
.A1(n_2495),
.A2(n_1730),
.B(n_1798),
.Y(n_2597)
);

INVx1_ASAP7_75t_SL g2598 ( 
.A(n_2507),
.Y(n_2598)
);

OAI22xp5_ASAP7_75t_L g2599 ( 
.A1(n_2519),
.A2(n_2307),
.B1(n_2330),
.B2(n_2063),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2499),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2467),
.Y(n_2601)
);

CKINVDCx5p33_ASAP7_75t_R g2602 ( 
.A(n_2488),
.Y(n_2602)
);

AOI22xp33_ASAP7_75t_L g2603 ( 
.A1(n_2507),
.A2(n_2164),
.B1(n_2238),
.B2(n_2077),
.Y(n_2603)
);

INVx1_ASAP7_75t_SL g2604 ( 
.A(n_2448),
.Y(n_2604)
);

CKINVDCx20_ASAP7_75t_R g2605 ( 
.A(n_2500),
.Y(n_2605)
);

INVx1_ASAP7_75t_SL g2606 ( 
.A(n_2448),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2474),
.Y(n_2607)
);

CKINVDCx5p33_ASAP7_75t_R g2608 ( 
.A(n_2431),
.Y(n_2608)
);

INVx6_ASAP7_75t_L g2609 ( 
.A(n_2514),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2559),
.Y(n_2610)
);

AOI22xp33_ASAP7_75t_L g2611 ( 
.A1(n_2529),
.A2(n_2060),
.B1(n_2115),
.B2(n_2205),
.Y(n_2611)
);

OAI21xp5_ASAP7_75t_SL g2612 ( 
.A1(n_2579),
.A2(n_2573),
.B(n_1791),
.Y(n_2612)
);

INVx3_ASAP7_75t_L g2613 ( 
.A(n_2576),
.Y(n_2613)
);

OAI211xp5_ASAP7_75t_L g2614 ( 
.A1(n_2564),
.A2(n_1911),
.B(n_1913),
.C(n_2259),
.Y(n_2614)
);

BUFx12f_ASAP7_75t_SL g2615 ( 
.A(n_2545),
.Y(n_2615)
);

BUFx4f_ASAP7_75t_SL g2616 ( 
.A(n_2582),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2533),
.Y(n_2617)
);

AOI21xp33_ASAP7_75t_L g2618 ( 
.A1(n_2540),
.A2(n_2246),
.B(n_2235),
.Y(n_2618)
);

OAI22xp5_ASAP7_75t_L g2619 ( 
.A1(n_2589),
.A2(n_2494),
.B1(n_2319),
.B2(n_2309),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_2543),
.B(n_2281),
.Y(n_2620)
);

INVx2_ASAP7_75t_L g2621 ( 
.A(n_2534),
.Y(n_2621)
);

AOI22xp33_ASAP7_75t_L g2622 ( 
.A1(n_2548),
.A2(n_2205),
.B1(n_2377),
.B2(n_2228),
.Y(n_2622)
);

AOI22xp33_ASAP7_75t_L g2623 ( 
.A1(n_2536),
.A2(n_2252),
.B1(n_2254),
.B2(n_2250),
.Y(n_2623)
);

BUFx2_ASAP7_75t_L g2624 ( 
.A(n_2539),
.Y(n_2624)
);

AND2x2_ASAP7_75t_L g2625 ( 
.A(n_2535),
.B(n_2084),
.Y(n_2625)
);

OAI22xp5_ASAP7_75t_L g2626 ( 
.A1(n_2549),
.A2(n_2315),
.B1(n_2390),
.B2(n_2335),
.Y(n_2626)
);

INVx4_ASAP7_75t_L g2627 ( 
.A(n_2567),
.Y(n_2627)
);

AOI22xp33_ASAP7_75t_L g2628 ( 
.A1(n_2554),
.A2(n_2261),
.B1(n_2256),
.B2(n_2420),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2537),
.Y(n_2629)
);

AOI22xp33_ASAP7_75t_L g2630 ( 
.A1(n_2530),
.A2(n_2182),
.B1(n_2198),
.B2(n_2181),
.Y(n_2630)
);

AOI22xp33_ASAP7_75t_L g2631 ( 
.A1(n_2566),
.A2(n_2198),
.B1(n_2242),
.B2(n_2182),
.Y(n_2631)
);

INVx3_ASAP7_75t_SL g2632 ( 
.A(n_2608),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_2555),
.B(n_2321),
.Y(n_2633)
);

AOI22xp33_ASAP7_75t_SL g2634 ( 
.A1(n_2553),
.A2(n_1726),
.B1(n_2381),
.B2(n_2125),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_2542),
.Y(n_2635)
);

OAI22xp33_ASAP7_75t_L g2636 ( 
.A1(n_2557),
.A2(n_2323),
.B1(n_2388),
.B2(n_2032),
.Y(n_2636)
);

AOI22xp5_ASAP7_75t_L g2637 ( 
.A1(n_2569),
.A2(n_2599),
.B1(n_2588),
.B2(n_2586),
.Y(n_2637)
);

OAI22xp5_ASAP7_75t_L g2638 ( 
.A1(n_2551),
.A2(n_2575),
.B1(n_2603),
.B2(n_2562),
.Y(n_2638)
);

OAI22xp33_ASAP7_75t_L g2639 ( 
.A1(n_2587),
.A2(n_2167),
.B1(n_2149),
.B2(n_2262),
.Y(n_2639)
);

AOI22xp33_ASAP7_75t_L g2640 ( 
.A1(n_2561),
.A2(n_2242),
.B1(n_2248),
.B2(n_2247),
.Y(n_2640)
);

INVx6_ASAP7_75t_L g2641 ( 
.A(n_2531),
.Y(n_2641)
);

AOI22xp33_ASAP7_75t_L g2642 ( 
.A1(n_2583),
.A2(n_2247),
.B1(n_2248),
.B2(n_2227),
.Y(n_2642)
);

AND2x2_ASAP7_75t_L g2643 ( 
.A(n_2584),
.B(n_2085),
.Y(n_2643)
);

AOI22xp5_ASAP7_75t_L g2644 ( 
.A1(n_2565),
.A2(n_2416),
.B1(n_2227),
.B2(n_2107),
.Y(n_2644)
);

BUFx4f_ASAP7_75t_SL g2645 ( 
.A(n_2552),
.Y(n_2645)
);

HB1xp67_ASAP7_75t_L g2646 ( 
.A(n_2585),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2538),
.Y(n_2647)
);

AOI22xp33_ASAP7_75t_L g2648 ( 
.A1(n_2580),
.A2(n_2574),
.B1(n_2577),
.B2(n_2237),
.Y(n_2648)
);

AOI22xp33_ASAP7_75t_L g2649 ( 
.A1(n_2578),
.A2(n_2237),
.B1(n_2200),
.B2(n_2210),
.Y(n_2649)
);

INVx5_ASAP7_75t_SL g2650 ( 
.A(n_2595),
.Y(n_2650)
);

AND2x2_ASAP7_75t_L g2651 ( 
.A(n_2541),
.B(n_2193),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2581),
.Y(n_2652)
);

OAI21xp5_ASAP7_75t_SL g2653 ( 
.A1(n_2597),
.A2(n_1771),
.B(n_1762),
.Y(n_2653)
);

AOI22xp33_ASAP7_75t_SL g2654 ( 
.A1(n_2553),
.A2(n_2381),
.B1(n_1966),
.B2(n_2492),
.Y(n_2654)
);

AOI22xp33_ASAP7_75t_SL g2655 ( 
.A1(n_2578),
.A2(n_2381),
.B1(n_1966),
.B2(n_2492),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2591),
.Y(n_2656)
);

INVx2_ASAP7_75t_SL g2657 ( 
.A(n_2560),
.Y(n_2657)
);

OAI21xp33_ASAP7_75t_L g2658 ( 
.A1(n_2590),
.A2(n_2090),
.B(n_2058),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2593),
.B(n_2600),
.Y(n_2659)
);

AOI22xp33_ASAP7_75t_L g2660 ( 
.A1(n_2594),
.A2(n_2191),
.B1(n_2057),
.B2(n_2065),
.Y(n_2660)
);

AOI22xp33_ASAP7_75t_L g2661 ( 
.A1(n_2531),
.A2(n_2061),
.B1(n_2073),
.B2(n_2072),
.Y(n_2661)
);

NOR2xp33_ASAP7_75t_L g2662 ( 
.A(n_2570),
.B(n_2276),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_2598),
.B(n_2087),
.Y(n_2663)
);

AOI22xp5_ASAP7_75t_L g2664 ( 
.A1(n_2605),
.A2(n_2514),
.B1(n_2167),
.B2(n_2451),
.Y(n_2664)
);

AOI22xp33_ASAP7_75t_L g2665 ( 
.A1(n_2558),
.A2(n_2096),
.B1(n_2240),
.B2(n_2230),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2601),
.Y(n_2666)
);

NAND3xp33_ASAP7_75t_L g2667 ( 
.A(n_2607),
.B(n_1989),
.C(n_2241),
.Y(n_2667)
);

OAI22xp5_ASAP7_75t_L g2668 ( 
.A1(n_2560),
.A2(n_2457),
.B1(n_2475),
.B2(n_2471),
.Y(n_2668)
);

AND2x2_ASAP7_75t_L g2669 ( 
.A(n_2547),
.B(n_2199),
.Y(n_2669)
);

OAI21xp5_ASAP7_75t_SL g2670 ( 
.A1(n_2604),
.A2(n_1753),
.B(n_2243),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2563),
.Y(n_2671)
);

AND2x2_ASAP7_75t_L g2672 ( 
.A(n_2606),
.B(n_2203),
.Y(n_2672)
);

OAI222xp33_ASAP7_75t_L g2673 ( 
.A1(n_2568),
.A2(n_2457),
.B1(n_2253),
.B2(n_2249),
.C1(n_2134),
.C2(n_2501),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_2546),
.Y(n_2674)
);

AOI22xp33_ASAP7_75t_L g2675 ( 
.A1(n_2572),
.A2(n_2255),
.B1(n_2264),
.B2(n_2244),
.Y(n_2675)
);

INVx3_ASAP7_75t_L g2676 ( 
.A(n_2556),
.Y(n_2676)
);

AOI22xp5_ASAP7_75t_L g2677 ( 
.A1(n_2550),
.A2(n_2266),
.B1(n_2180),
.B2(n_2207),
.Y(n_2677)
);

OAI22xp5_ASAP7_75t_L g2678 ( 
.A1(n_2572),
.A2(n_2463),
.B1(n_2303),
.B2(n_2429),
.Y(n_2678)
);

BUFx2_ASAP7_75t_L g2679 ( 
.A(n_2592),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2567),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2567),
.Y(n_2681)
);

HB1xp67_ASAP7_75t_L g2682 ( 
.A(n_2571),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2571),
.Y(n_2683)
);

AOI22xp33_ASAP7_75t_L g2684 ( 
.A1(n_2609),
.A2(n_2171),
.B1(n_2211),
.B2(n_2208),
.Y(n_2684)
);

AOI22xp33_ASAP7_75t_L g2685 ( 
.A1(n_2638),
.A2(n_2097),
.B1(n_2119),
.B2(n_2098),
.Y(n_2685)
);

NAND4xp25_ASAP7_75t_L g2686 ( 
.A(n_2614),
.B(n_2122),
.C(n_2132),
.D(n_2120),
.Y(n_2686)
);

OAI22xp33_ASAP7_75t_L g2687 ( 
.A1(n_2637),
.A2(n_2544),
.B1(n_2441),
.B2(n_2609),
.Y(n_2687)
);

OAI22xp5_ASAP7_75t_L g2688 ( 
.A1(n_2677),
.A2(n_2360),
.B1(n_2429),
.B2(n_2456),
.Y(n_2688)
);

AOI22xp33_ASAP7_75t_L g2689 ( 
.A1(n_2637),
.A2(n_2625),
.B1(n_2658),
.B2(n_2611),
.Y(n_2689)
);

AOI22xp33_ASAP7_75t_L g2690 ( 
.A1(n_2648),
.A2(n_2142),
.B1(n_2140),
.B2(n_2141),
.Y(n_2690)
);

OAI22xp5_ASAP7_75t_L g2691 ( 
.A1(n_2677),
.A2(n_2455),
.B1(n_2498),
.B2(n_2493),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2620),
.B(n_2285),
.Y(n_2692)
);

AND2x2_ASAP7_75t_L g2693 ( 
.A(n_2643),
.B(n_2503),
.Y(n_2693)
);

AOI22xp33_ASAP7_75t_L g2694 ( 
.A1(n_2671),
.A2(n_2135),
.B1(n_2112),
.B2(n_2117),
.Y(n_2694)
);

OAI22xp5_ASAP7_75t_L g2695 ( 
.A1(n_2634),
.A2(n_2520),
.B1(n_2418),
.B2(n_2357),
.Y(n_2695)
);

NAND2xp33_ASAP7_75t_SL g2696 ( 
.A(n_2632),
.B(n_1836),
.Y(n_2696)
);

NAND3xp33_ASAP7_75t_L g2697 ( 
.A(n_2612),
.B(n_2126),
.C(n_2104),
.Y(n_2697)
);

AOI221xp5_ASAP7_75t_L g2698 ( 
.A1(n_2636),
.A2(n_1920),
.B1(n_2162),
.B2(n_2163),
.C(n_2160),
.Y(n_2698)
);

OAI22xp5_ASAP7_75t_L g2699 ( 
.A1(n_2644),
.A2(n_2355),
.B1(n_2526),
.B2(n_2515),
.Y(n_2699)
);

AOI22xp33_ASAP7_75t_L g2700 ( 
.A1(n_2639),
.A2(n_2137),
.B1(n_2139),
.B2(n_2131),
.Y(n_2700)
);

AOI22xp33_ASAP7_75t_L g2701 ( 
.A1(n_2623),
.A2(n_2270),
.B1(n_2233),
.B2(n_2480),
.Y(n_2701)
);

AOI22xp33_ASAP7_75t_L g2702 ( 
.A1(n_2622),
.A2(n_2270),
.B1(n_2523),
.B2(n_2480),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_L g2703 ( 
.A(n_2624),
.B(n_2289),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2621),
.B(n_2304),
.Y(n_2704)
);

AOI22xp5_ASAP7_75t_L g2705 ( 
.A1(n_2653),
.A2(n_2602),
.B1(n_2596),
.B2(n_2532),
.Y(n_2705)
);

OAI21xp5_ASAP7_75t_L g2706 ( 
.A1(n_2618),
.A2(n_1847),
.B(n_1837),
.Y(n_2706)
);

AOI22xp33_ASAP7_75t_L g2707 ( 
.A1(n_2628),
.A2(n_2270),
.B1(n_2523),
.B2(n_2480),
.Y(n_2707)
);

CKINVDCx20_ASAP7_75t_R g2708 ( 
.A(n_2645),
.Y(n_2708)
);

AOI22xp33_ASAP7_75t_SL g2709 ( 
.A1(n_2626),
.A2(n_2619),
.B1(n_2633),
.B2(n_2646),
.Y(n_2709)
);

AOI22xp5_ASAP7_75t_L g2710 ( 
.A1(n_2662),
.A2(n_2523),
.B1(n_2452),
.B2(n_2324),
.Y(n_2710)
);

AOI221xp5_ASAP7_75t_L g2711 ( 
.A1(n_2673),
.A2(n_2419),
.B1(n_2311),
.B2(n_2345),
.C(n_2362),
.Y(n_2711)
);

AND2x2_ASAP7_75t_L g2712 ( 
.A(n_2613),
.B(n_2526),
.Y(n_2712)
);

AOI22xp33_ASAP7_75t_L g2713 ( 
.A1(n_2649),
.A2(n_2523),
.B1(n_2423),
.B2(n_2378),
.Y(n_2713)
);

AOI22xp33_ASAP7_75t_L g2714 ( 
.A1(n_2644),
.A2(n_1917),
.B1(n_1916),
.B2(n_2078),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_SL g2715 ( 
.A(n_2655),
.B(n_2510),
.Y(n_2715)
);

INVx2_ASAP7_75t_L g2716 ( 
.A(n_2613),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2635),
.B(n_2087),
.Y(n_2717)
);

AOI22xp33_ASAP7_75t_L g2718 ( 
.A1(n_2642),
.A2(n_2078),
.B1(n_2522),
.B2(n_2516),
.Y(n_2718)
);

AOI22xp33_ASAP7_75t_L g2719 ( 
.A1(n_2669),
.A2(n_2522),
.B1(n_2516),
.B2(n_2155),
.Y(n_2719)
);

AOI22xp33_ASAP7_75t_L g2720 ( 
.A1(n_2630),
.A2(n_2166),
.B1(n_2154),
.B2(n_2510),
.Y(n_2720)
);

OAI22xp5_ASAP7_75t_L g2721 ( 
.A1(n_2675),
.A2(n_2511),
.B1(n_2571),
.B2(n_2460),
.Y(n_2721)
);

NAND3xp33_ASAP7_75t_L g2722 ( 
.A(n_2670),
.B(n_2511),
.C(n_2486),
.Y(n_2722)
);

AND2x2_ASAP7_75t_L g2723 ( 
.A(n_2651),
.B(n_2460),
.Y(n_2723)
);

AOI22xp33_ASAP7_75t_SL g2724 ( 
.A1(n_2641),
.A2(n_2486),
.B1(n_2469),
.B2(n_183),
.Y(n_2724)
);

AOI22xp33_ASAP7_75t_L g2725 ( 
.A1(n_2667),
.A2(n_2317),
.B1(n_183),
.B2(n_181),
.Y(n_2725)
);

BUFx3_ASAP7_75t_L g2726 ( 
.A(n_2641),
.Y(n_2726)
);

AOI22xp33_ASAP7_75t_L g2727 ( 
.A1(n_2661),
.A2(n_186),
.B1(n_182),
.B2(n_184),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2610),
.B(n_184),
.Y(n_2728)
);

AOI22xp33_ASAP7_75t_L g2729 ( 
.A1(n_2660),
.A2(n_192),
.B1(n_187),
.B2(n_188),
.Y(n_2729)
);

AOI22xp33_ASAP7_75t_L g2730 ( 
.A1(n_2665),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.Y(n_2730)
);

AND2x2_ASAP7_75t_L g2731 ( 
.A(n_2672),
.B(n_535),
.Y(n_2731)
);

AOI22xp33_ASAP7_75t_L g2732 ( 
.A1(n_2654),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.Y(n_2732)
);

AOI221xp5_ASAP7_75t_L g2733 ( 
.A1(n_2666),
.A2(n_197),
.B1(n_199),
.B2(n_201),
.C(n_202),
.Y(n_2733)
);

AOI22xp33_ASAP7_75t_L g2734 ( 
.A1(n_2631),
.A2(n_204),
.B1(n_197),
.B2(n_202),
.Y(n_2734)
);

AOI22xp33_ASAP7_75t_L g2735 ( 
.A1(n_2617),
.A2(n_206),
.B1(n_204),
.B2(n_205),
.Y(n_2735)
);

AOI22xp33_ASAP7_75t_L g2736 ( 
.A1(n_2629),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_2736)
);

OAI221xp5_ASAP7_75t_L g2737 ( 
.A1(n_2664),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.C(n_211),
.Y(n_2737)
);

AOI222xp33_ASAP7_75t_L g2738 ( 
.A1(n_2616),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.C1(n_211),
.C2(n_212),
.Y(n_2738)
);

OAI222xp33_ASAP7_75t_L g2739 ( 
.A1(n_2659),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.C1(n_215),
.C2(n_216),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2689),
.B(n_2647),
.Y(n_2740)
);

NOR2xp33_ASAP7_75t_L g2741 ( 
.A(n_2687),
.B(n_2652),
.Y(n_2741)
);

AND2x2_ASAP7_75t_L g2742 ( 
.A(n_2723),
.B(n_2693),
.Y(n_2742)
);

NAND3xp33_ASAP7_75t_L g2743 ( 
.A(n_2738),
.B(n_2684),
.C(n_2640),
.Y(n_2743)
);

AND2x2_ASAP7_75t_L g2744 ( 
.A(n_2712),
.B(n_2656),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_SL g2745 ( 
.A(n_2687),
.B(n_2668),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2689),
.B(n_2692),
.Y(n_2746)
);

NAND4xp25_ASAP7_75t_L g2747 ( 
.A(n_2735),
.B(n_2674),
.C(n_2679),
.D(n_2663),
.Y(n_2747)
);

NAND3xp33_ASAP7_75t_SL g2748 ( 
.A(n_2737),
.B(n_2678),
.C(n_2681),
.Y(n_2748)
);

OA211x2_ASAP7_75t_L g2749 ( 
.A1(n_2733),
.A2(n_2650),
.B(n_2615),
.C(n_2682),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_SL g2750 ( 
.A(n_2709),
.B(n_2676),
.Y(n_2750)
);

AOI22xp33_ASAP7_75t_L g2751 ( 
.A1(n_2735),
.A2(n_2683),
.B1(n_2680),
.B2(n_2657),
.Y(n_2751)
);

OAI21xp33_ASAP7_75t_SL g2752 ( 
.A1(n_2736),
.A2(n_2627),
.B(n_2676),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2703),
.B(n_2627),
.Y(n_2753)
);

AND2x2_ASAP7_75t_L g2754 ( 
.A(n_2731),
.B(n_2650),
.Y(n_2754)
);

NAND3xp33_ASAP7_75t_L g2755 ( 
.A(n_2736),
.B(n_213),
.C(n_214),
.Y(n_2755)
);

NOR3xp33_ASAP7_75t_L g2756 ( 
.A(n_2686),
.B(n_215),
.C(n_216),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2716),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2728),
.B(n_219),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_SL g2759 ( 
.A(n_2705),
.B(n_536),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2685),
.B(n_219),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2685),
.B(n_220),
.Y(n_2761)
);

AND2x2_ASAP7_75t_L g2762 ( 
.A(n_2710),
.B(n_221),
.Y(n_2762)
);

OAI21xp33_ASAP7_75t_L g2763 ( 
.A1(n_2732),
.A2(n_221),
.B(n_222),
.Y(n_2763)
);

OAI221xp5_ASAP7_75t_L g2764 ( 
.A1(n_2724),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.C(n_226),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_2704),
.B(n_224),
.Y(n_2765)
);

AND2x2_ASAP7_75t_L g2766 ( 
.A(n_2715),
.B(n_226),
.Y(n_2766)
);

NAND3xp33_ASAP7_75t_L g2767 ( 
.A(n_2697),
.B(n_2729),
.C(n_2722),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_2719),
.B(n_227),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2717),
.B(n_227),
.Y(n_2769)
);

NAND2xp33_ASAP7_75t_SL g2770 ( 
.A(n_2708),
.B(n_228),
.Y(n_2770)
);

AOI221xp5_ASAP7_75t_L g2771 ( 
.A1(n_2739),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.C(n_232),
.Y(n_2771)
);

AND2x2_ASAP7_75t_L g2772 ( 
.A(n_2726),
.B(n_230),
.Y(n_2772)
);

AND2x2_ASAP7_75t_L g2773 ( 
.A(n_2707),
.B(n_233),
.Y(n_2773)
);

AOI21xp5_ASAP7_75t_SL g2774 ( 
.A1(n_2706),
.A2(n_542),
.B(n_537),
.Y(n_2774)
);

NAND3xp33_ASAP7_75t_SL g2775 ( 
.A(n_2756),
.B(n_2730),
.C(n_2725),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2757),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2744),
.Y(n_2777)
);

NAND4xp75_ASAP7_75t_L g2778 ( 
.A(n_2749),
.B(n_2711),
.C(n_2698),
.D(n_2696),
.Y(n_2778)
);

NOR3xp33_ASAP7_75t_L g2779 ( 
.A(n_2767),
.B(n_2755),
.C(n_2764),
.Y(n_2779)
);

AOI22xp33_ASAP7_75t_L g2780 ( 
.A1(n_2756),
.A2(n_2727),
.B1(n_2690),
.B2(n_2702),
.Y(n_2780)
);

NAND2xp33_ASAP7_75t_SL g2781 ( 
.A(n_2750),
.B(n_2721),
.Y(n_2781)
);

HB1xp67_ASAP7_75t_L g2782 ( 
.A(n_2741),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2740),
.Y(n_2783)
);

NAND4xp25_ASAP7_75t_L g2784 ( 
.A(n_2771),
.B(n_2734),
.C(n_2694),
.D(n_2701),
.Y(n_2784)
);

OR2x2_ASAP7_75t_L g2785 ( 
.A(n_2753),
.B(n_2695),
.Y(n_2785)
);

AND2x2_ASAP7_75t_L g2786 ( 
.A(n_2742),
.B(n_2699),
.Y(n_2786)
);

AND2x2_ASAP7_75t_L g2787 ( 
.A(n_2754),
.B(n_2713),
.Y(n_2787)
);

NOR3xp33_ASAP7_75t_L g2788 ( 
.A(n_2763),
.B(n_2691),
.C(n_2688),
.Y(n_2788)
);

BUFx3_ASAP7_75t_L g2789 ( 
.A(n_2772),
.Y(n_2789)
);

OAI211xp5_ASAP7_75t_L g2790 ( 
.A1(n_2751),
.A2(n_2714),
.B(n_2700),
.C(n_2718),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2741),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_2746),
.B(n_2720),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2758),
.B(n_234),
.Y(n_2793)
);

OR2x2_ASAP7_75t_L g2794 ( 
.A(n_2765),
.B(n_234),
.Y(n_2794)
);

AOI22xp5_ASAP7_75t_L g2795 ( 
.A1(n_2745),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_2795)
);

INVx1_ASAP7_75t_SL g2796 ( 
.A(n_2789),
.Y(n_2796)
);

NOR4xp25_ASAP7_75t_L g2797 ( 
.A(n_2775),
.B(n_2766),
.C(n_2762),
.D(n_2750),
.Y(n_2797)
);

XNOR2xp5_ASAP7_75t_L g2798 ( 
.A(n_2787),
.B(n_2770),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2776),
.Y(n_2799)
);

NAND4xp75_ASAP7_75t_SL g2800 ( 
.A(n_2778),
.B(n_2773),
.C(n_2781),
.D(n_2779),
.Y(n_2800)
);

AND2x2_ASAP7_75t_L g2801 ( 
.A(n_2777),
.B(n_2752),
.Y(n_2801)
);

NAND4xp75_ASAP7_75t_L g2802 ( 
.A(n_2795),
.B(n_2759),
.C(n_2761),
.D(n_2760),
.Y(n_2802)
);

OR2x2_ASAP7_75t_L g2803 ( 
.A(n_2783),
.B(n_2769),
.Y(n_2803)
);

XOR2xp5_ASAP7_75t_L g2804 ( 
.A(n_2792),
.B(n_2747),
.Y(n_2804)
);

NAND4xp75_ASAP7_75t_SL g2805 ( 
.A(n_2786),
.B(n_2774),
.C(n_2748),
.D(n_2751),
.Y(n_2805)
);

NAND4xp75_ASAP7_75t_SL g2806 ( 
.A(n_2788),
.B(n_2743),
.C(n_2768),
.D(n_241),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2782),
.Y(n_2807)
);

NAND4xp25_ASAP7_75t_L g2808 ( 
.A(n_2793),
.B(n_238),
.C(n_239),
.D(n_243),
.Y(n_2808)
);

INVx2_ASAP7_75t_L g2809 ( 
.A(n_2799),
.Y(n_2809)
);

XNOR2x1_ASAP7_75t_L g2810 ( 
.A(n_2798),
.B(n_2794),
.Y(n_2810)
);

OA22x2_ASAP7_75t_L g2811 ( 
.A1(n_2804),
.A2(n_2791),
.B1(n_2793),
.B2(n_2790),
.Y(n_2811)
);

XNOR2x1_ASAP7_75t_L g2812 ( 
.A(n_2800),
.B(n_2785),
.Y(n_2812)
);

XOR2x2_ASAP7_75t_L g2813 ( 
.A(n_2806),
.B(n_2805),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_2807),
.Y(n_2814)
);

XOR2x2_ASAP7_75t_L g2815 ( 
.A(n_2796),
.B(n_2780),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2809),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2814),
.Y(n_2817)
);

AO22x2_ASAP7_75t_L g2818 ( 
.A1(n_2812),
.A2(n_2803),
.B1(n_2802),
.B2(n_2801),
.Y(n_2818)
);

OA22x2_ASAP7_75t_L g2819 ( 
.A1(n_2811),
.A2(n_2813),
.B1(n_2797),
.B2(n_2815),
.Y(n_2819)
);

AOI22xp5_ASAP7_75t_L g2820 ( 
.A1(n_2811),
.A2(n_2808),
.B1(n_2784),
.B2(n_246),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2810),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2809),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2816),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2822),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2817),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2818),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2818),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2820),
.B(n_2808),
.Y(n_2828)
);

OAI22xp5_ASAP7_75t_L g2829 ( 
.A1(n_2826),
.A2(n_2819),
.B1(n_2821),
.B2(n_2784),
.Y(n_2829)
);

AO22x2_ASAP7_75t_L g2830 ( 
.A1(n_2827),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_2830)
);

OAI22xp5_ASAP7_75t_L g2831 ( 
.A1(n_2828),
.A2(n_244),
.B1(n_245),
.B2(n_247),
.Y(n_2831)
);

NAND4xp25_ASAP7_75t_SL g2832 ( 
.A(n_2823),
.B(n_247),
.C(n_248),
.D(n_250),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2824),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2833),
.Y(n_2834)
);

OA22x2_ASAP7_75t_L g2835 ( 
.A1(n_2829),
.A2(n_2825),
.B1(n_252),
.B2(n_253),
.Y(n_2835)
);

AOI22xp5_ASAP7_75t_L g2836 ( 
.A1(n_2832),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_2836)
);

AOI22xp5_ASAP7_75t_L g2837 ( 
.A1(n_2831),
.A2(n_251),
.B1(n_255),
.B2(n_256),
.Y(n_2837)
);

INVx2_ASAP7_75t_SL g2838 ( 
.A(n_2830),
.Y(n_2838)
);

NOR4xp25_ASAP7_75t_L g2839 ( 
.A(n_2838),
.B(n_255),
.C(n_257),
.D(n_258),
.Y(n_2839)
);

NOR2xp33_ASAP7_75t_L g2840 ( 
.A(n_2835),
.B(n_2836),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2834),
.Y(n_2841)
);

NOR2x1_ASAP7_75t_L g2842 ( 
.A(n_2837),
.B(n_258),
.Y(n_2842)
);

NOR2x1_ASAP7_75t_L g2843 ( 
.A(n_2834),
.B(n_259),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_2838),
.Y(n_2844)
);

INVxp67_ASAP7_75t_SL g2845 ( 
.A(n_2838),
.Y(n_2845)
);

NOR4xp25_ASAP7_75t_L g2846 ( 
.A(n_2838),
.B(n_259),
.C(n_260),
.D(n_262),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2845),
.B(n_260),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2844),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2843),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2841),
.Y(n_2850)
);

INVxp67_ASAP7_75t_SL g2851 ( 
.A(n_2842),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2840),
.Y(n_2852)
);

AOI22xp5_ASAP7_75t_L g2853 ( 
.A1(n_2839),
.A2(n_262),
.B1(n_264),
.B2(n_265),
.Y(n_2853)
);

AOI22xp5_ASAP7_75t_L g2854 ( 
.A1(n_2846),
.A2(n_266),
.B1(n_267),
.B2(n_269),
.Y(n_2854)
);

AOI22xp5_ASAP7_75t_L g2855 ( 
.A1(n_2852),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.Y(n_2855)
);

HB1xp67_ASAP7_75t_L g2856 ( 
.A(n_2849),
.Y(n_2856)
);

INVx2_ASAP7_75t_L g2857 ( 
.A(n_2848),
.Y(n_2857)
);

INVx2_ASAP7_75t_L g2858 ( 
.A(n_2847),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2851),
.Y(n_2859)
);

AOI22xp5_ASAP7_75t_L g2860 ( 
.A1(n_2853),
.A2(n_270),
.B1(n_273),
.B2(n_274),
.Y(n_2860)
);

OR3x2_ASAP7_75t_L g2861 ( 
.A(n_2850),
.B(n_275),
.C(n_276),
.Y(n_2861)
);

AOI22xp5_ASAP7_75t_L g2862 ( 
.A1(n_2854),
.A2(n_275),
.B1(n_277),
.B2(n_278),
.Y(n_2862)
);

INVx2_ASAP7_75t_L g2863 ( 
.A(n_2849),
.Y(n_2863)
);

OAI22xp5_ASAP7_75t_L g2864 ( 
.A1(n_2861),
.A2(n_277),
.B1(n_279),
.B2(n_280),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2856),
.Y(n_2865)
);

BUFx2_ASAP7_75t_L g2866 ( 
.A(n_2859),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2863),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2857),
.Y(n_2868)
);

OR2x2_ASAP7_75t_L g2869 ( 
.A(n_2858),
.B(n_281),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2855),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2860),
.Y(n_2871)
);

HB1xp67_ASAP7_75t_L g2872 ( 
.A(n_2862),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2866),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2865),
.Y(n_2874)
);

AO22x2_ASAP7_75t_L g2875 ( 
.A1(n_2864),
.A2(n_282),
.B1(n_283),
.B2(n_285),
.Y(n_2875)
);

AOI22xp33_ASAP7_75t_L g2876 ( 
.A1(n_2871),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2869),
.Y(n_2877)
);

OAI22x1_ASAP7_75t_L g2878 ( 
.A1(n_2872),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_2878)
);

OAI22x1_ASAP7_75t_L g2879 ( 
.A1(n_2870),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2875),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2875),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2873),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2878),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2879),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2874),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2877),
.Y(n_2886)
);

AOI22xp5_ASAP7_75t_L g2887 ( 
.A1(n_2883),
.A2(n_2867),
.B1(n_2868),
.B2(n_2876),
.Y(n_2887)
);

NAND4xp25_ASAP7_75t_L g2888 ( 
.A(n_2884),
.B(n_289),
.C(n_291),
.D(n_292),
.Y(n_2888)
);

AOI22xp5_ASAP7_75t_L g2889 ( 
.A1(n_2882),
.A2(n_2886),
.B1(n_2881),
.B2(n_2880),
.Y(n_2889)
);

AOI221xp5_ASAP7_75t_SL g2890 ( 
.A1(n_2885),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.C(n_295),
.Y(n_2890)
);

INVx3_ASAP7_75t_L g2891 ( 
.A(n_2890),
.Y(n_2891)
);

AOI22xp5_ASAP7_75t_L g2892 ( 
.A1(n_2891),
.A2(n_2887),
.B1(n_2889),
.B2(n_2888),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2892),
.Y(n_2893)
);

AOI221xp5_ASAP7_75t_L g2894 ( 
.A1(n_2893),
.A2(n_293),
.B1(n_295),
.B2(n_296),
.C(n_297),
.Y(n_2894)
);

AOI211xp5_ASAP7_75t_L g2895 ( 
.A1(n_2894),
.A2(n_298),
.B(n_301),
.C(n_302),
.Y(n_2895)
);


endmodule