module fake_netlist_1_5913_n_448 (n_53, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_448);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_448;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_137;
wire n_277;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_67;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_203;
wire n_102;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_68;
wire n_123;
wire n_223;
wire n_372;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g66 ( .A(n_22), .Y(n_66) );
INVx1_ASAP7_75t_L g67 ( .A(n_36), .Y(n_67) );
INVx1_ASAP7_75t_L g68 ( .A(n_50), .Y(n_68) );
INVxp67_ASAP7_75t_L g69 ( .A(n_51), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_43), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_57), .Y(n_71) );
BUFx2_ASAP7_75t_L g72 ( .A(n_31), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_17), .Y(n_73) );
INVxp67_ASAP7_75t_SL g74 ( .A(n_63), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_42), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_55), .Y(n_76) );
INVxp67_ASAP7_75t_SL g77 ( .A(n_32), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_5), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_5), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_64), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_14), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_14), .Y(n_82) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_20), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_30), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_41), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_62), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_0), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_23), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_8), .Y(n_89) );
INVxp67_ASAP7_75t_L g90 ( .A(n_19), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_54), .Y(n_91) );
INVx1_ASAP7_75t_SL g92 ( .A(n_56), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_45), .Y(n_93) );
AND2x2_ASAP7_75t_L g94 ( .A(n_35), .B(n_37), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_4), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_65), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_46), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_7), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_72), .Y(n_99) );
NAND2xp5_ASAP7_75t_SL g100 ( .A(n_72), .B(n_0), .Y(n_100) );
BUFx6f_ASAP7_75t_L g101 ( .A(n_91), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_87), .B(n_1), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_79), .Y(n_103) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_91), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_66), .Y(n_105) );
INVxp67_ASAP7_75t_SL g106 ( .A(n_79), .Y(n_106) );
AND2x6_ASAP7_75t_L g107 ( .A(n_94), .B(n_33), .Y(n_107) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_70), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_84), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_81), .Y(n_110) );
BUFx3_ASAP7_75t_L g111 ( .A(n_70), .Y(n_111) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_78), .Y(n_112) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_78), .Y(n_113) );
AND2x4_ASAP7_75t_L g114 ( .A(n_82), .B(n_1), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_84), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_81), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_96), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_96), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_71), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_83), .Y(n_120) );
NOR2x1_ASAP7_75t_L g121 ( .A(n_95), .B(n_34), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_109), .Y(n_122) );
AOI22xp5_ASAP7_75t_L g123 ( .A1(n_109), .A2(n_82), .B1(n_89), .B2(n_98), .Y(n_123) );
OAI22xp5_ASAP7_75t_L g124 ( .A1(n_99), .A2(n_89), .B1(n_69), .B2(n_90), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_101), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_101), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_101), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_101), .Y(n_128) );
INVx4_ASAP7_75t_L g129 ( .A(n_107), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_108), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_115), .B(n_97), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_101), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_108), .Y(n_133) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_115), .Y(n_134) );
BUFx4f_ASAP7_75t_L g135 ( .A(n_107), .Y(n_135) );
BUFx2_ASAP7_75t_L g136 ( .A(n_117), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_108), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_111), .B(n_67), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_111), .B(n_68), .Y(n_139) );
AND2x4_ASAP7_75t_L g140 ( .A(n_106), .B(n_71), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_104), .Y(n_141) );
BUFx4_ASAP7_75t_L g142 ( .A(n_102), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_117), .B(n_80), .Y(n_143) );
OAI21xp33_ASAP7_75t_L g144 ( .A1(n_114), .A2(n_73), .B(n_93), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_108), .Y(n_145) );
BUFx3_ASAP7_75t_L g146 ( .A(n_107), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_104), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_130), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_129), .B(n_118), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_140), .B(n_118), .Y(n_150) );
NAND3xp33_ASAP7_75t_SL g151 ( .A(n_122), .B(n_120), .C(n_105), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_140), .B(n_114), .Y(n_152) );
BUFx2_ASAP7_75t_L g153 ( .A(n_136), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_146), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_130), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_140), .B(n_112), .Y(n_156) );
CKINVDCx16_ASAP7_75t_R g157 ( .A(n_136), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_146), .Y(n_158) );
INVx1_ASAP7_75t_SL g159 ( .A(n_142), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_122), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_143), .B(n_113), .Y(n_161) );
BUFx3_ASAP7_75t_L g162 ( .A(n_135), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_133), .Y(n_163) );
BUFx3_ASAP7_75t_L g164 ( .A(n_135), .Y(n_164) );
BUFx2_ASAP7_75t_L g165 ( .A(n_134), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_133), .Y(n_166) );
INVx3_ASAP7_75t_L g167 ( .A(n_129), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_137), .Y(n_168) );
AND2x4_ASAP7_75t_L g169 ( .A(n_129), .B(n_114), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_131), .B(n_100), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_135), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_138), .B(n_107), .Y(n_172) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_127), .Y(n_173) );
OR2x2_ASAP7_75t_L g174 ( .A(n_123), .B(n_120), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_137), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_139), .B(n_107), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_145), .Y(n_177) );
BUFx2_ASAP7_75t_L g178 ( .A(n_124), .Y(n_178) );
OR2x2_ASAP7_75t_L g179 ( .A(n_144), .B(n_110), .Y(n_179) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_145), .A2(n_107), .B1(n_119), .B2(n_108), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_142), .B(n_116), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_152), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_153), .B(n_103), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_152), .Y(n_184) );
BUFx2_ASAP7_75t_L g185 ( .A(n_153), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_152), .B(n_119), .Y(n_186) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_171), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_157), .Y(n_188) );
BUFx2_ASAP7_75t_L g189 ( .A(n_165), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_169), .Y(n_190) );
BUFx12f_ASAP7_75t_L g191 ( .A(n_165), .Y(n_191) );
OAI221xp5_ASAP7_75t_L g192 ( .A1(n_156), .A2(n_161), .B1(n_178), .B2(n_150), .C(n_179), .Y(n_192) );
BUFx2_ASAP7_75t_L g193 ( .A(n_157), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_154), .Y(n_194) );
INVx5_ASAP7_75t_L g195 ( .A(n_154), .Y(n_195) );
AOI221xp5_ASAP7_75t_L g196 ( .A1(n_178), .A2(n_119), .B1(n_93), .B2(n_75), .C(n_76), .Y(n_196) );
BUFx3_ASAP7_75t_L g197 ( .A(n_171), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_171), .Y(n_198) );
INVx4_ASAP7_75t_L g199 ( .A(n_169), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_170), .A2(n_119), .B1(n_121), .B2(n_74), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_171), .Y(n_201) );
OR2x6_ASAP7_75t_L g202 ( .A(n_169), .B(n_73), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_148), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_181), .B(n_119), .Y(n_204) );
INVx3_ASAP7_75t_L g205 ( .A(n_154), .Y(n_205) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_159), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_181), .B(n_75), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_170), .B(n_76), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_171), .B(n_94), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_179), .Y(n_210) );
BUFx3_ASAP7_75t_L g211 ( .A(n_154), .Y(n_211) );
INVx4_ASAP7_75t_L g212 ( .A(n_154), .Y(n_212) );
BUFx3_ASAP7_75t_L g213 ( .A(n_158), .Y(n_213) );
OR2x2_ASAP7_75t_L g214 ( .A(n_174), .B(n_2), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g215 ( .A1(n_192), .A2(n_170), .B1(n_174), .B2(n_176), .Y(n_215) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_189), .Y(n_216) );
AOI21xp5_ASAP7_75t_SL g217 ( .A1(n_202), .A2(n_180), .B(n_162), .Y(n_217) );
OR2x2_ASAP7_75t_L g218 ( .A(n_189), .B(n_151), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_185), .A2(n_160), .B1(n_172), .B2(n_149), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_203), .Y(n_220) );
OAI22xp33_ASAP7_75t_L g221 ( .A1(n_191), .A2(n_180), .B1(n_167), .B2(n_164), .Y(n_221) );
BUFx4f_ASAP7_75t_SL g222 ( .A(n_191), .Y(n_222) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_187), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_199), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_192), .B(n_167), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_187), .Y(n_226) );
OR2x2_ASAP7_75t_L g227 ( .A(n_193), .B(n_2), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g228 ( .A1(n_202), .A2(n_162), .B1(n_164), .B2(n_167), .Y(n_228) );
OAI21x1_ASAP7_75t_L g229 ( .A1(n_194), .A2(n_88), .B(n_85), .Y(n_229) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_200), .A2(n_88), .B(n_86), .Y(n_230) );
OAI22xp33_ASAP7_75t_L g231 ( .A1(n_191), .A2(n_158), .B1(n_77), .B2(n_92), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_203), .Y(n_232) );
OAI21x1_ASAP7_75t_L g233 ( .A1(n_194), .A2(n_141), .B(n_125), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_207), .B(n_158), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_188), .Y(n_235) );
NAND2x1_ASAP7_75t_L g236 ( .A(n_203), .B(n_158), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_190), .Y(n_237) );
BUFx2_ASAP7_75t_L g238 ( .A(n_185), .Y(n_238) );
OAI22xp33_ASAP7_75t_L g239 ( .A1(n_214), .A2(n_158), .B1(n_104), .B2(n_168), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_220), .Y(n_240) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_229), .A2(n_196), .B(n_200), .Y(n_241) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_220), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_220), .B(n_207), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_232), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_215), .A2(n_193), .B1(n_214), .B2(n_202), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_232), .Y(n_246) );
INVx3_ASAP7_75t_L g247 ( .A(n_232), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_215), .A2(n_202), .B1(n_207), .B2(n_208), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_234), .B(n_183), .Y(n_249) );
OAI22xp33_ASAP7_75t_L g250 ( .A1(n_227), .A2(n_202), .B1(n_210), .B2(n_196), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_238), .A2(n_202), .B1(n_208), .B2(n_204), .Y(n_251) );
OAI221xp5_ASAP7_75t_L g252 ( .A1(n_218), .A2(n_182), .B1(n_184), .B2(n_183), .C(n_206), .Y(n_252) );
BUFx8_ASAP7_75t_SL g253 ( .A(n_235), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_238), .A2(n_204), .B1(n_206), .B2(n_184), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_218), .A2(n_182), .B1(n_190), .B2(n_199), .Y(n_255) );
AOI22xp33_ASAP7_75t_SL g256 ( .A1(n_222), .A2(n_199), .B1(n_195), .B2(n_201), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_216), .B(n_199), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_237), .Y(n_258) );
AOI221xp5_ASAP7_75t_SL g259 ( .A1(n_239), .A2(n_209), .B1(n_186), .B2(n_104), .C(n_201), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_242), .A2(n_217), .B(n_250), .Y(n_260) );
OR2x2_ASAP7_75t_L g261 ( .A(n_242), .B(n_227), .Y(n_261) );
INVx3_ASAP7_75t_L g262 ( .A(n_247), .Y(n_262) );
INVx3_ASAP7_75t_L g263 ( .A(n_247), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_246), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_240), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_249), .B(n_219), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_240), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_240), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_244), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_245), .B(n_224), .Y(n_270) );
NOR3xp33_ASAP7_75t_SL g271 ( .A(n_252), .B(n_231), .C(n_221), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_243), .B(n_230), .Y(n_272) );
AOI221xp5_ASAP7_75t_L g273 ( .A1(n_250), .A2(n_225), .B1(n_186), .B2(n_224), .C(n_217), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_247), .Y(n_274) );
AO21x2_ASAP7_75t_L g275 ( .A1(n_246), .A2(n_229), .B(n_230), .Y(n_275) );
AOI221xp5_ASAP7_75t_L g276 ( .A1(n_252), .A2(n_224), .B1(n_104), .B2(n_228), .C(n_148), .Y(n_276) );
AOI221xp5_ASAP7_75t_L g277 ( .A1(n_248), .A2(n_224), .B1(n_155), .B2(n_163), .C(n_166), .Y(n_277) );
AOI222xp33_ASAP7_75t_L g278 ( .A1(n_258), .A2(n_212), .B1(n_211), .B2(n_213), .C1(n_197), .C2(n_205), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_244), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_265), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_265), .Y(n_281) );
NAND3xp33_ASAP7_75t_L g282 ( .A(n_271), .B(n_259), .C(n_254), .Y(n_282) );
NOR3xp33_ASAP7_75t_L g283 ( .A(n_266), .B(n_257), .C(n_256), .Y(n_283) );
INVx1_ASAP7_75t_SL g284 ( .A(n_265), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_264), .Y(n_285) );
BUFx2_ASAP7_75t_L g286 ( .A(n_267), .Y(n_286) );
OAI221xp5_ASAP7_75t_SL g287 ( .A1(n_260), .A2(n_251), .B1(n_255), .B2(n_259), .C(n_256), .Y(n_287) );
INVxp67_ASAP7_75t_L g288 ( .A(n_261), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_267), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_279), .B(n_244), .Y(n_290) );
AND2x4_ASAP7_75t_L g291 ( .A(n_267), .B(n_247), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_268), .B(n_241), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_276), .A2(n_241), .B1(n_212), .B2(n_197), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_272), .B(n_241), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_268), .Y(n_295) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_261), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_268), .Y(n_297) );
AOI221xp5_ASAP7_75t_L g298 ( .A1(n_270), .A2(n_125), .B1(n_126), .B2(n_141), .C(n_128), .Y(n_298) );
INVxp67_ASAP7_75t_SL g299 ( .A(n_269), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_272), .B(n_253), .Y(n_300) );
OAI33xp33_ASAP7_75t_L g301 ( .A1(n_269), .A2(n_126), .A3(n_128), .B1(n_6), .B2(n_7), .B3(n_8), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_279), .B(n_241), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_279), .B(n_241), .Y(n_303) );
INVx3_ASAP7_75t_L g304 ( .A(n_262), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_269), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_275), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_262), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_286), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_296), .B(n_273), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_288), .B(n_275), .Y(n_310) );
NOR2x1_ASAP7_75t_L g311 ( .A(n_282), .B(n_275), .Y(n_311) );
NAND2x1p5_ASAP7_75t_L g312 ( .A(n_286), .B(n_263), .Y(n_312) );
AOI211xp5_ASAP7_75t_L g313 ( .A1(n_287), .A2(n_277), .B(n_263), .C(n_274), .Y(n_313) );
INVx2_ASAP7_75t_SL g314 ( .A(n_290), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_294), .B(n_274), .Y(n_315) );
INVx2_ASAP7_75t_SL g316 ( .A(n_290), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_285), .B(n_274), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_281), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_300), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_283), .B(n_274), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_291), .B(n_278), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_282), .B(n_3), .Y(n_322) );
AOI211xp5_ASAP7_75t_L g323 ( .A1(n_306), .A2(n_127), .B(n_132), .C(n_147), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_295), .B(n_3), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_292), .B(n_4), .Y(n_325) );
OAI32xp33_ASAP7_75t_L g326 ( .A1(n_284), .A2(n_297), .A3(n_305), .B1(n_295), .B2(n_306), .Y(n_326) );
INVx2_ASAP7_75t_SL g327 ( .A(n_291), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_292), .B(n_6), .Y(n_328) );
NAND2x1p5_ASAP7_75t_L g329 ( .A(n_291), .B(n_304), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_305), .Y(n_330) );
NOR3xp33_ASAP7_75t_L g331 ( .A(n_301), .B(n_236), .C(n_212), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_299), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_291), .B(n_9), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_280), .B(n_9), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_281), .Y(n_335) );
INVxp67_ASAP7_75t_L g336 ( .A(n_289), .Y(n_336) );
AND2x2_ASAP7_75t_SL g337 ( .A(n_281), .B(n_223), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_289), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_293), .A2(n_236), .B1(n_212), .B2(n_226), .Y(n_339) );
INVx1_ASAP7_75t_SL g340 ( .A(n_303), .Y(n_340) );
INVx2_ASAP7_75t_SL g341 ( .A(n_304), .Y(n_341) );
AND2x4_ASAP7_75t_L g342 ( .A(n_304), .B(n_223), .Y(n_342) );
INVx4_ASAP7_75t_L g343 ( .A(n_304), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g344 ( .A1(n_322), .A2(n_307), .B1(n_302), .B2(n_298), .Y(n_344) );
AOI222xp33_ASAP7_75t_L g345 ( .A1(n_322), .A2(n_307), .B1(n_11), .B2(n_12), .C1(n_13), .C2(n_15), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_323), .A2(n_226), .B(n_223), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_325), .B(n_10), .Y(n_347) );
AOI21xp33_ASAP7_75t_L g348 ( .A1(n_320), .A2(n_10), .B(n_11), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_325), .B(n_12), .Y(n_349) );
OAI21xp5_ASAP7_75t_L g350 ( .A1(n_328), .A2(n_233), .B(n_195), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_314), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_314), .B(n_13), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_319), .B(n_15), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_319), .B(n_16), .Y(n_354) );
OAI221xp5_ASAP7_75t_SL g355 ( .A1(n_309), .A2(n_213), .B1(n_211), .B2(n_197), .C(n_205), .Y(n_355) );
AOI22xp5_ASAP7_75t_SL g356 ( .A1(n_328), .A2(n_226), .B1(n_223), .B2(n_213), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_316), .B(n_226), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_321), .A2(n_226), .B1(n_223), .B2(n_211), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_313), .A2(n_226), .B1(n_223), .B2(n_195), .Y(n_359) );
INVx1_ASAP7_75t_SL g360 ( .A(n_340), .Y(n_360) );
OAI21xp5_ASAP7_75t_L g361 ( .A1(n_333), .A2(n_233), .B(n_195), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_334), .Y(n_362) );
OAI21xp33_ASAP7_75t_L g363 ( .A1(n_311), .A2(n_127), .B(n_132), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_315), .B(n_18), .Y(n_364) );
NAND2x1_ASAP7_75t_L g365 ( .A(n_343), .B(n_205), .Y(n_365) );
OAI321xp33_ASAP7_75t_L g366 ( .A1(n_310), .A2(n_147), .A3(n_132), .B1(n_127), .B2(n_201), .C(n_198), .Y(n_366) );
OAI21xp33_ASAP7_75t_L g367 ( .A1(n_315), .A2(n_127), .B(n_132), .Y(n_367) );
AOI321xp33_ASAP7_75t_L g368 ( .A1(n_326), .A2(n_205), .A3(n_194), .B1(n_168), .B2(n_166), .C(n_163), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_331), .A2(n_194), .B1(n_195), .B2(n_198), .Y(n_369) );
O2A1O1Ixp33_ASAP7_75t_L g370 ( .A1(n_324), .A2(n_155), .B(n_177), .C(n_175), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_327), .B(n_21), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_330), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_332), .Y(n_373) );
OAI221xp5_ASAP7_75t_SL g374 ( .A1(n_308), .A2(n_24), .B1(n_25), .B2(n_26), .C(n_27), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_336), .B(n_28), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_327), .B(n_29), .Y(n_376) );
NAND2xp33_ASAP7_75t_L g377 ( .A(n_312), .B(n_329), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_317), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_317), .B(n_38), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_338), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_373), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_360), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_351), .B(n_329), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_362), .B(n_308), .Y(n_384) );
NAND2x1_ASAP7_75t_L g385 ( .A(n_346), .B(n_343), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_354), .B(n_341), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_345), .A2(n_337), .B1(n_335), .B2(n_318), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_378), .B(n_312), .Y(n_388) );
NAND2xp33_ASAP7_75t_SL g389 ( .A(n_352), .B(n_339), .Y(n_389) );
OAI21xp33_ASAP7_75t_L g390 ( .A1(n_347), .A2(n_349), .B(n_369), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_372), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_380), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_344), .B(n_318), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_356), .B(n_337), .Y(n_394) );
INVx1_ASAP7_75t_SL g395 ( .A(n_377), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_374), .A2(n_339), .B1(n_342), .B2(n_195), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_348), .B(n_342), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_359), .B(n_342), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_358), .B(n_39), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_364), .B(n_350), .Y(n_400) );
NOR3xp33_ASAP7_75t_SL g401 ( .A(n_374), .B(n_40), .C(n_44), .Y(n_401) );
INVxp33_ASAP7_75t_L g402 ( .A(n_365), .Y(n_402) );
XOR2xp5_ASAP7_75t_L g403 ( .A(n_357), .B(n_47), .Y(n_403) );
NOR3xp33_ASAP7_75t_L g404 ( .A(n_375), .B(n_48), .C(n_49), .Y(n_404) );
INVxp67_ASAP7_75t_L g405 ( .A(n_368), .Y(n_405) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_346), .A2(n_195), .B1(n_198), .B2(n_201), .Y(n_406) );
NOR2x1_ASAP7_75t_L g407 ( .A(n_395), .B(n_370), .Y(n_407) );
INVx2_ASAP7_75t_SL g408 ( .A(n_382), .Y(n_408) );
AOI22xp33_ASAP7_75t_SL g409 ( .A1(n_405), .A2(n_361), .B1(n_371), .B2(n_376), .Y(n_409) );
NOR2xp33_ASAP7_75t_R g410 ( .A(n_389), .B(n_379), .Y(n_410) );
NAND3xp33_ASAP7_75t_L g411 ( .A(n_405), .B(n_355), .C(n_370), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_393), .B(n_367), .Y(n_412) );
AOI21xp5_ASAP7_75t_L g413 ( .A1(n_385), .A2(n_355), .B(n_366), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_387), .A2(n_363), .B1(n_201), .B2(n_198), .Y(n_414) );
AOI221xp5_ASAP7_75t_L g415 ( .A1(n_387), .A2(n_201), .B1(n_198), .B2(n_187), .C(n_177), .Y(n_415) );
INVxp67_ASAP7_75t_L g416 ( .A(n_384), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_390), .B(n_52), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_391), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_401), .A2(n_198), .B1(n_187), .B2(n_53), .Y(n_419) );
OAI32xp33_ASAP7_75t_L g420 ( .A1(n_402), .A2(n_58), .A3(n_59), .B1(n_60), .B2(n_61), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_392), .Y(n_421) );
OAI21xp5_ASAP7_75t_SL g422 ( .A1(n_394), .A2(n_403), .B(n_396), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_422), .A2(n_400), .B1(n_398), .B2(n_386), .Y(n_423) );
BUFx2_ASAP7_75t_L g424 ( .A(n_408), .Y(n_424) );
NOR2x1_ASAP7_75t_L g425 ( .A(n_407), .B(n_406), .Y(n_425) );
INVxp33_ASAP7_75t_L g426 ( .A(n_410), .Y(n_426) );
O2A1O1Ixp33_ASAP7_75t_L g427 ( .A1(n_419), .A2(n_404), .B(n_406), .C(n_381), .Y(n_427) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_411), .B(n_397), .C(n_404), .Y(n_428) );
OAI221xp5_ASAP7_75t_L g429 ( .A1(n_409), .A2(n_388), .B1(n_399), .B2(n_383), .C(n_187), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_418), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_416), .B(n_173), .Y(n_431) );
AOI221xp5_ASAP7_75t_L g432 ( .A1(n_421), .A2(n_173), .B1(n_415), .B2(n_412), .C(n_417), .Y(n_432) );
OAI211xp5_ASAP7_75t_SL g433 ( .A1(n_409), .A2(n_173), .B(n_414), .C(n_413), .Y(n_433) );
NAND3xp33_ASAP7_75t_L g434 ( .A(n_420), .B(n_407), .C(n_411), .Y(n_434) );
AOI222xp33_ASAP7_75t_L g435 ( .A1(n_411), .A2(n_405), .B1(n_389), .B2(n_407), .C1(n_422), .C2(n_353), .Y(n_435) );
OAI211xp5_ASAP7_75t_SL g436 ( .A1(n_407), .A2(n_405), .B(n_422), .C(n_387), .Y(n_436) );
INVx6_ASAP7_75t_L g437 ( .A(n_431), .Y(n_437) );
INVxp67_ASAP7_75t_L g438 ( .A(n_434), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_430), .Y(n_439) );
OAI221xp5_ASAP7_75t_L g440 ( .A1(n_436), .A2(n_435), .B1(n_425), .B2(n_428), .C(n_423), .Y(n_440) );
NAND3xp33_ASAP7_75t_L g441 ( .A(n_438), .B(n_433), .C(n_432), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_439), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_437), .Y(n_443) );
INVxp33_ASAP7_75t_L g444 ( .A(n_443), .Y(n_444) );
BUFx2_ASAP7_75t_L g445 ( .A(n_442), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_445), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_446), .A2(n_440), .B1(n_444), .B2(n_441), .Y(n_447) );
AOI221xp5_ASAP7_75t_L g448 ( .A1(n_447), .A2(n_426), .B1(n_429), .B2(n_424), .C(n_427), .Y(n_448) );
endmodule