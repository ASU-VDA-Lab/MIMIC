module fake_netlist_6_3091_n_4331 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_442, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_67, n_15, n_443, n_246, n_38, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_466, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_397, n_155, n_109, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_414, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_363, n_395, n_323, n_393, n_411, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_102, n_204, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_433, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_464, n_33, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_328, n_429, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_64, n_288, n_427, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_4331);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_466;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_397;
input n_155;
input n_109;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_102;
input n_204;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_433;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_464;
input n_33;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_328;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_64;
input n_288;
input n_427;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_4331;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_801;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_2576;
wire n_1234;
wire n_3254;
wire n_3684;
wire n_1199;
wire n_1674;
wire n_3392;
wire n_741;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_625;
wire n_1189;
wire n_3152;
wire n_4154;
wire n_3579;
wire n_1212;
wire n_4251;
wire n_726;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3783;
wire n_700;
wire n_3773;
wire n_4177;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_4127;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_3844;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3301;
wire n_3089;
wire n_4099;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_3741;
wire n_4168;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_509;
wire n_1342;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_1708;
wire n_677;
wire n_805;
wire n_1151;
wire n_2977;
wire n_3952;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_3911;
wire n_2359;
wire n_480;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_3332;
wire n_4134;
wire n_4285;
wire n_3465;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_3706;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2997;
wire n_2179;
wire n_2386;
wire n_2570;
wire n_4092;
wire n_1724;
wire n_1032;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_4078;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_4249;
wire n_1264;
wire n_1192;
wire n_471;
wire n_3564;
wire n_1844;
wire n_3619;
wire n_4087;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_4302;
wire n_2291;
wire n_830;
wire n_2299;
wire n_3340;
wire n_4179;
wire n_873;
wire n_1285;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_3946;
wire n_4213;
wire n_1985;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_852;
wire n_2509;
wire n_4065;
wire n_4026;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_3904;
wire n_4178;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_4273;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_4029;
wire n_836;
wire n_3345;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2919;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_3879;
wire n_4010;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_3979;
wire n_616;
wire n_658;
wire n_4308;
wire n_1874;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2739;
wire n_3023;
wire n_822;
wire n_3232;
wire n_693;
wire n_1313;
wire n_2791;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_1056;
wire n_3877;
wire n_3316;
wire n_4325;
wire n_2212;
wire n_3929;
wire n_758;
wire n_516;
wire n_3494;
wire n_3048;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3063;
wire n_4311;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_4060;
wire n_1550;
wire n_2703;
wire n_491;
wire n_3998;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_772;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_666;
wire n_4187;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_538;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_4164;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3624;
wire n_3077;
wire n_3737;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3655;
wire n_494;
wire n_539;
wire n_493;
wire n_3107;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_4117;
wire n_3948;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_4327;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_3765;
wire n_713;
wire n_2655;
wire n_4125;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_4221;
wire n_1467;
wire n_3297;
wire n_4250;
wire n_976;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_3906;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_4262;
wire n_1894;
wire n_2996;
wire n_1231;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3963;
wire n_3368;
wire n_917;
wire n_574;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_907;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_2591;
wire n_3507;
wire n_659;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_4253;
wire n_913;
wire n_4110;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_4071;
wire n_4255;
wire n_3506;
wire n_4268;
wire n_3568;
wire n_3269;
wire n_4047;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_473;
wire n_1193;
wire n_1967;
wire n_3999;
wire n_1054;
wire n_3928;
wire n_559;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_4139;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_551;
wire n_1986;
wire n_699;
wire n_2300;
wire n_3943;
wire n_4320;
wire n_4305;
wire n_564;
wire n_2397;
wire n_3884;
wire n_3931;
wire n_824;
wire n_686;
wire n_4102;
wire n_4297;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_3871;
wire n_2907;
wire n_577;
wire n_3438;
wire n_2735;
wire n_4141;
wire n_1843;
wire n_619;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_2778;
wire n_4227;
wire n_2850;
wire n_572;
wire n_4314;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_3822;
wire n_4163;
wire n_606;
wire n_1441;
wire n_818;
wire n_3373;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_1699;
wire n_3910;
wire n_916;
wire n_3934;
wire n_2093;
wire n_4033;
wire n_4296;
wire n_4009;
wire n_2633;
wire n_483;
wire n_3883;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_630;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_541;
wire n_512;
wire n_2669;
wire n_2925;
wire n_3728;
wire n_4094;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_792;
wire n_2522;
wire n_476;
wire n_3949;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_3912;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_3923;
wire n_2529;
wire n_3900;
wire n_1162;
wire n_860;
wire n_1530;
wire n_3798;
wire n_788;
wire n_939;
wire n_3488;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_3732;
wire n_982;
wire n_4257;
wire n_2674;
wire n_2832;
wire n_4226;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_932;
wire n_2831;
wire n_2998;
wire n_4318;
wire n_3446;
wire n_4158;
wire n_3857;
wire n_3978;
wire n_3317;
wire n_1876;
wire n_4107;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_4074;
wire n_3716;
wire n_1873;
wire n_4294;
wire n_905;
wire n_3630;
wire n_3518;
wire n_3824;
wire n_3859;
wire n_1866;
wire n_4013;
wire n_1680;
wire n_2692;
wire n_993;
wire n_3842;
wire n_689;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1413;
wire n_1605;
wire n_1330;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3914;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_547;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_558;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_4032;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_634;
wire n_2355;
wire n_3927;
wire n_4147;
wire n_966;
wire n_3888;
wire n_2908;
wire n_3168;
wire n_764;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_4161;
wire n_4130;
wire n_2895;
wire n_2009;
wire n_4172;
wire n_692;
wire n_3403;
wire n_733;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_3882;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_487;
wire n_3055;
wire n_3092;
wire n_3492;
wire n_3895;
wire n_3966;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_1014;
wire n_3734;
wire n_3686;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_4118;
wire n_882;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_586;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_2459;
wire n_3746;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_715;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3935;
wire n_3384;
wire n_1265;
wire n_4277;
wire n_2711;
wire n_3490;
wire n_4291;
wire n_4199;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_4319;
wire n_3369;
wire n_3419;
wire n_1982;
wire n_3872;
wire n_2878;
wire n_618;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_3875;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_3794;
wire n_674;
wire n_3247;
wire n_871;
wire n_3069;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_1722;
wire n_1664;
wire n_612;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_3933;
wire n_702;
wire n_2008;
wire n_2749;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_2254;
wire n_3346;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_3691;
wire n_780;
wire n_3861;
wire n_675;
wire n_2624;
wire n_4066;
wire n_903;
wire n_4146;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_3891;
wire n_2193;
wire n_3961;
wire n_2676;
wire n_1655;
wire n_3940;
wire n_4072;
wire n_4220;
wire n_835;
wire n_928;
wire n_1801;
wire n_850;
wire n_690;
wire n_1214;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3410;
wire n_3153;
wire n_3428;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_604;
wire n_4004;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_4043;
wire n_825;
wire n_4313;
wire n_728;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_4292;
wire n_1588;
wire n_3785;
wire n_3942;
wire n_3997;
wire n_2963;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_1124;
wire n_1624;
wire n_3873;
wire n_3983;
wire n_515;
wire n_2096;
wire n_2980;
wire n_3968;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_598;
wire n_3434;
wire n_696;
wire n_1515;
wire n_961;
wire n_3510;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_593;
wire n_4169;
wire n_514;
wire n_4055;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_3271;
wire n_950;
wire n_4248;
wire n_2812;
wire n_484;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_3889;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_3707;
wire n_2075;
wire n_4045;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_4070;
wire n_1987;
wire n_3545;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_3578;
wire n_3885;
wire n_881;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_760;
wire n_3993;
wire n_1546;
wire n_2583;
wire n_590;
wire n_4116;
wire n_2606;
wire n_4031;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_2431;
wire n_3073;
wire n_4018;
wire n_2987;
wire n_694;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_3696;
wire n_3780;
wire n_4082;
wire n_1634;
wire n_2078;
wire n_3252;
wire n_2932;
wire n_595;
wire n_1767;
wire n_627;
wire n_3253;
wire n_1779;
wire n_524;
wire n_1465;
wire n_3337;
wire n_3431;
wire n_3450;
wire n_3209;
wire n_4002;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_4329;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_2893;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_3477;
wire n_4288;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_4289;
wire n_2712;
wire n_2684;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_495;
wire n_815;
wire n_3953;
wire n_1100;
wire n_585;
wire n_1487;
wire n_2691;
wire n_3614;
wire n_840;
wire n_2913;
wire n_3421;
wire n_874;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_4019;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_3616;
wire n_4228;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_4044;
wire n_3436;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_4191;
wire n_1364;
wire n_4322;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_3937;
wire n_615;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_4287;
wire n_1293;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_3941;
wire n_963;
wire n_639;
wire n_794;
wire n_2767;
wire n_3793;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_3385;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_1139;
wire n_1714;
wire n_872;
wire n_3922;
wire n_3179;
wire n_718;
wire n_1018;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_4330;
wire n_542;
wire n_847;
wire n_851;
wire n_644;
wire n_682;
wire n_2897;
wire n_2537;
wire n_3970;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_1513;
wire n_2747;
wire n_3924;
wire n_3171;
wire n_791;
wire n_1913;
wire n_4216;
wire n_3608;
wire n_510;
wire n_837;
wire n_4315;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_4156;
wire n_3491;
wire n_4240;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_704;
wire n_2148;
wire n_4284;
wire n_4162;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_536;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2590;
wire n_2643;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_3782;
wire n_3975;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_4011;
wire n_1835;
wire n_3470;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_4098;
wire n_4021;
wire n_765;
wire n_1492;
wire n_987;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_4058;
wire n_4103;
wire n_3104;
wire n_631;
wire n_720;
wire n_3435;
wire n_842;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_4022;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_4310;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_499;
wire n_2675;
wire n_1426;
wire n_3580;
wire n_705;
wire n_3418;
wire n_3775;
wire n_3537;
wire n_2134;
wire n_1176;
wire n_1004;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_3887;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_684;
wire n_2667;
wire n_2698;
wire n_2539;
wire n_4096;
wire n_1431;
wire n_4123;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_3835;
wire n_1571;
wire n_3312;
wire n_4286;
wire n_1809;
wire n_3119;
wire n_4280;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_3731;
wire n_1822;
wire n_486;
wire n_947;
wire n_2936;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_648;
wire n_657;
wire n_1049;
wire n_3223;
wire n_3996;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_4097;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_4218;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_3880;
wire n_1849;
wire n_2848;
wire n_919;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_478;
wire n_4100;
wire n_2231;
wire n_3609;
wire n_929;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_4264;
wire n_2857;
wire n_3693;
wire n_3788;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_2896;
wire n_526;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_4079;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_4175;
wire n_998;
wire n_717;
wire n_3200;
wire n_1665;
wire n_4306;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_4224;
wire n_3390;
wire n_3656;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_3593;
wire n_3867;
wire n_3341;
wire n_3324;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_3559;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_4005;
wire n_1507;
wire n_2482;
wire n_552;
wire n_3810;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_912;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_1284;
wire n_745;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_3201;
wire n_3633;
wire n_3447;
wire n_3971;
wire n_1142;
wire n_2849;
wire n_716;
wire n_1475;
wire n_1774;
wire n_1048;
wire n_1398;
wire n_623;
wire n_884;
wire n_1201;
wire n_2682;
wire n_2354;
wire n_3103;
wire n_3032;
wire n_3638;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_3393;
wire n_474;
wire n_683;
wire n_811;
wire n_527;
wire n_1207;
wire n_2442;
wire n_3627;
wire n_1791;
wire n_1368;
wire n_3480;
wire n_3451;
wire n_1418;
wire n_958;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_4222;
wire n_2545;
wire n_3540;
wire n_3577;
wire n_889;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_589;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_819;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_3591;
wire n_767;
wire n_3641;
wire n_1314;
wire n_600;
wire n_1837;
wire n_831;
wire n_2218;
wire n_2788;
wire n_964;
wire n_477;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_4120;
wire n_1382;
wire n_1534;
wire n_3892;
wire n_1736;
wire n_1564;
wire n_4069;
wire n_4053;
wire n_2748;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_505;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2511;
wire n_537;
wire n_2475;
wire n_3964;
wire n_1993;
wire n_2281;
wire n_4167;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_596;
wire n_3944;
wire n_3909;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2301;
wire n_2209;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_4223;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_970;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_642;
wire n_3481;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_4299;
wire n_3724;
wire n_3033;
wire n_1252;
wire n_1784;
wire n_3913;
wire n_3571;
wire n_1223;
wire n_3311;
wire n_4276;
wire n_511;
wire n_2990;
wire n_3847;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_520;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3323;
wire n_3226;
wire n_4020;
wire n_3364;
wire n_4176;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_3407;
wire n_518;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_2384;
wire n_3894;
wire n_4204;
wire n_4261;
wire n_1745;
wire n_914;
wire n_759;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_4063;
wire n_1625;
wire n_3986;
wire n_4237;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_1453;
wire n_2146;
wire n_4006;
wire n_2226;
wire n_2131;
wire n_488;
wire n_2502;
wire n_2801;
wire n_3646;
wire n_497;
wire n_2920;
wire n_4015;
wire n_773;
wire n_3547;
wire n_1901;
wire n_3869;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_3188;
wire n_3742;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_4034;
wire n_4056;
wire n_1617;
wire n_3260;
wire n_3816;
wire n_3386;
wire n_3370;
wire n_3960;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_3175;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_848;
wire n_2732;
wire n_2928;
wire n_4206;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_1580;
wire n_2227;
wire n_4247;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_4180;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_3284;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_1390;
wire n_906;
wire n_688;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2289;
wire n_1419;
wire n_2863;
wire n_3299;
wire n_3663;
wire n_4132;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_3360;
wire n_2135;
wire n_3956;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_4001;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_4149;
wire n_1331;
wire n_613;
wire n_736;
wire n_2627;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_3234;
wire n_3917;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_3016;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_2993;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_4003;
wire n_1129;
wire n_3870;
wire n_4030;
wire n_4126;
wire n_554;
wire n_602;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_3845;
wire n_664;
wire n_1869;
wire n_2911;
wire n_3625;
wire n_3751;
wire n_3804;
wire n_1764;
wire n_4207;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_4113;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_793;
wire n_587;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_4014;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_4067;
wire n_4252;
wire n_607;
wire n_1551;
wire n_4028;
wire n_4054;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_3907;
wire n_2555;
wire n_4048;
wire n_3338;
wire n_4217;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_3919;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_2984;
wire n_575;
wire n_994;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_2304;
wire n_4024;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3276;
wire n_3250;
wire n_1934;
wire n_3194;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_4214;
wire n_1728;
wire n_3973;
wire n_557;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_617;
wire n_3886;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_485;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_3637;
wire n_3120;
wire n_1468;
wire n_3991;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3797;
wire n_3926;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_4234;
wire n_4304;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_4101;
wire n_3548;
wire n_3767;
wire n_1024;
wire n_3864;
wire n_4036;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_3974;
wire n_1847;
wire n_2052;
wire n_3634;
wire n_2302;
wire n_517;
wire n_4211;
wire n_4182;
wire n_1667;
wire n_667;
wire n_1206;
wire n_3230;
wire n_4016;
wire n_1037;
wire n_1397;
wire n_621;
wire n_3268;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_3592;
wire n_468;
wire n_2755;
wire n_3141;
wire n_923;
wire n_504;
wire n_1409;
wire n_4230;
wire n_1841;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_3967;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_4328;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_4274;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_4189;
wire n_4270;
wire n_4151;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_1818;
wire n_1108;
wire n_710;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3730;
wire n_1298;
wire n_4124;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_785;
wire n_4155;
wire n_2740;
wire n_746;
wire n_4238;
wire n_609;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2401;
wire n_2337;
wire n_1356;
wire n_1589;
wire n_3213;
wire n_3042;
wire n_3820;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_4152;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_4219;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_3529;
wire n_4193;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_4109;
wire n_4192;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_3424;
wire n_3957;
wire n_4038;
wire n_2790;
wire n_4131;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_4159;
wire n_4195;
wire n_3784;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_3594;
wire n_809;
wire n_1043;
wire n_3819;
wire n_4090;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_4165;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_4144;
wire n_1870;
wire n_2964;
wire n_4174;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3475;
wire n_662;
wire n_3501;
wire n_1840;
wire n_1152;
wire n_1705;
wire n_3905;
wire n_3262;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_4008;
wire n_2244;
wire n_4290;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_3692;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_4258;
wire n_650;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_1405;
wire n_972;
wire n_2376;
wire n_3826;
wire n_1406;
wire n_3790;
wire n_3878;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_4323;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_4300;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_2882;
wire n_3675;
wire n_3666;
wire n_4017;
wire n_4260;
wire n_3320;
wire n_2541;
wire n_654;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_1974;
wire n_3988;
wire n_4122;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_934;
wire n_482;
wire n_1637;
wire n_2635;
wire n_3307;
wire n_3439;
wire n_3588;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_4135;
wire n_4209;
wire n_2871;
wire n_4279;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_3858;
wire n_4183;
wire n_1489;
wire n_4321;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_4128;
wire n_543;
wire n_2229;
wire n_1964;
wire n_4133;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_4145;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_4271;
wire n_1946;
wire n_1355;
wire n_4181;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_4040;
wire n_804;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_4111;
wire n_533;
wire n_2390;
wire n_4007;
wire n_806;
wire n_3712;
wire n_959;
wire n_879;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_4239;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_4184;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_4037;
wire n_523;
wire n_1319;
wire n_707;
wire n_2986;
wire n_1900;
wire n_3930;
wire n_3246;
wire n_799;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_3915;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_787;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_4215;
wire n_1282;
wire n_2561;
wire n_550;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_3377;
wire n_2939;
wire n_560;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_4185;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_1914;
wire n_1318;
wire n_737;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_3893;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_3762;
wire n_3469;
wire n_3932;
wire n_2266;
wire n_2960;
wire n_3958;
wire n_3005;
wire n_3985;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1029;
wire n_4196;
wire n_3779;
wire n_1447;
wire n_2388;
wire n_3984;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_1706;
wire n_4242;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_4232;
wire n_4190;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_4052;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_3899;
wire n_4084;
wire n_3558;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_4326;
wire n_3156;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_502;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_3939;
wire n_1375;
wire n_1941;
wire n_3483;
wire n_3613;
wire n_3972;
wire n_4153;
wire n_2128;
wire n_655;
wire n_1045;
wire n_1650;
wire n_1794;
wire n_786;
wire n_1962;
wire n_1236;
wire n_706;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_3855;
wire n_3743;
wire n_1872;
wire n_3091;
wire n_4317;
wire n_834;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_4269;
wire n_743;
wire n_766;
wire n_3124;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_4088;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_545;
wire n_3524;
wire n_2671;
wire n_489;
wire n_2761;
wire n_2923;
wire n_2793;
wire n_2715;
wire n_2885;
wire n_1804;
wire n_2888;
wire n_3711;
wire n_3776;
wire n_4235;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_4301;
wire n_3511;
wire n_2054;
wire n_4143;
wire n_4170;
wire n_729;
wire n_876;
wire n_774;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_2062;
wire n_660;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_479;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_869;
wire n_1154;
wire n_3308;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_897;
wire n_846;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_841;
wire n_1476;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_3515;
wire n_1150;
wire n_4203;
wire n_3808;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1076;
wire n_1118;
wire n_2949;
wire n_3726;
wire n_1807;
wire n_1007;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_3758;
wire n_1879;
wire n_853;
wire n_695;
wire n_3806;
wire n_4081;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_875;
wire n_680;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_3866;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_671;
wire n_3565;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_3343;
wire n_3303;
wire n_978;
wire n_4157;
wire n_2752;
wire n_4173;
wire n_3135;
wire n_4324;
wire n_1976;
wire n_4229;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_3990;
wire n_751;
wire n_749;
wire n_3865;
wire n_1824;
wire n_3954;
wire n_1628;
wire n_4073;
wire n_1324;
wire n_3890;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_988;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_3658;
wire n_1516;
wire n_1536;
wire n_3846;
wire n_2163;
wire n_2186;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3951;
wire n_3034;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_3874;
wire n_1379;
wire n_2814;
wire n_2528;
wire n_2787;
wire n_2969;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_3027;
wire n_781;
wire n_789;
wire n_1554;
wire n_3231;
wire n_4083;
wire n_1130;
wire n_3083;
wire n_4212;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_4295;
wire n_1120;
wire n_1583;
wire n_832;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_4225;
wire n_4171;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_747;
wire n_3541;
wire n_2565;
wire n_4023;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_721;
wire n_1461;
wire n_742;
wire n_3432;
wire n_535;
wire n_691;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_3860;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_4282;
wire n_1598;
wire n_3493;
wire n_2935;
wire n_4046;
wire n_3807;
wire n_863;
wire n_3015;
wire n_2175;
wire n_601;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3701;
wire n_3154;
wire n_4027;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_3473;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_3739;
wire n_2284;
wire n_3898;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_744;
wire n_971;
wire n_2702;
wire n_3241;
wire n_946;
wire n_2906;
wire n_1303;
wire n_761;
wire n_2769;
wire n_3622;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_4095;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3897;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_4106;
wire n_795;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_1245;
wire n_838;
wire n_3215;
wire n_3969;
wire n_3336;
wire n_647;
wire n_4160;
wire n_4231;
wire n_844;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_3853;
wire n_2117;
wire n_2234;
wire n_4256;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_3553;
wire n_1561;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_3811;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_653;
wire n_2430;
wire n_3486;
wire n_1414;
wire n_3584;
wire n_4086;
wire n_752;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_3556;
wire n_2034;
wire n_576;
wire n_1028;
wire n_3836;
wire n_2106;
wire n_472;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_563;
wire n_4068;
wire n_2032;
wire n_2744;
wire n_4309;
wire n_1011;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_839;
wire n_2437;
wire n_2743;
wire n_3962;
wire n_1973;
wire n_708;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_668;
wire n_4166;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1821;
wire n_1537;
wire n_2205;
wire n_3699;
wire n_4243;
wire n_3204;
wire n_1104;
wire n_854;
wire n_1058;
wire n_3378;
wire n_4025;
wire n_2312;
wire n_498;
wire n_3404;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_3745;
wire n_3362;
wire n_4059;
wire n_1509;
wire n_4188;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_4121;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3256;
wire n_1276;
wire n_3802;
wire n_3868;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_3982;
wire n_4266;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_3796;
wire n_2999;
wire n_4115;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3697;
wire n_3643;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_3461;
wire n_3408;
wire n_1582;
wire n_492;
wire n_3680;
wire n_4265;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_2408;
wire n_4246;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2950;
wire n_2483;
wire n_1972;
wire n_719;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_3098;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_2666;
wire n_4105;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_4244;
wire n_1816;
wire n_4064;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_4049;
wire n_829;
wire n_1156;
wire n_1362;
wire n_4259;
wire n_3123;
wire n_984;
wire n_2600;
wire n_3380;
wire n_1829;
wire n_503;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_868;
wire n_3038;
wire n_570;
wire n_859;
wire n_2033;
wire n_3086;
wire n_735;
wire n_4104;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_3285;
wire n_519;
wire n_4208;
wire n_2523;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_3769;
wire n_1482;
wire n_3361;
wire n_981;
wire n_3596;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_4089;
wire n_1144;
wire n_2071;
wire n_3669;
wire n_3863;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_985;
wire n_4316;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_481;
wire n_3521;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_4061;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_4075;
wire n_3344;
wire n_2334;
wire n_3902;
wire n_4062;
wire n_3881;
wire n_3295;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_3989;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_4233;
wire n_1606;
wire n_810;
wire n_4108;
wire n_1133;
wire n_635;
wire n_1194;
wire n_3374;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_2640;
wire n_3695;
wire n_4051;
wire n_1051;
wire n_3976;
wire n_4254;
wire n_1552;
wire n_2918;
wire n_583;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_3992;
wire n_2367;
wire n_4307;
wire n_3876;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_4303;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_4293;
wire n_941;
wire n_3552;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2578;
wire n_2363;
wire n_553;
wire n_849;
wire n_2662;
wire n_3116;
wire n_3147;
wire n_3383;
wire n_3709;
wire n_753;
wire n_3925;
wire n_4091;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_4186;
wire n_467;
wire n_3187;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_2879;
wire n_861;
wire n_3717;
wire n_857;
wire n_967;
wire n_4148;
wire n_571;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_4057;
wire n_2968;
wire n_4201;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_4263;
wire n_1819;
wire n_2055;
wire n_1260;
wire n_3555;
wire n_1010;
wire n_3444;
wire n_4210;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_3955;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_3903;
wire n_730;
wire n_1311;
wire n_3945;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_4205;
wire n_2162;
wire n_3908;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_4278;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3950;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_1417;
wire n_1242;
wire n_2185;
wire n_2086;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_3833;
wire n_4281;
wire n_3815;
wire n_2774;
wire n_3896;
wire n_3039;
wire n_681;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3274;
wire n_3333;
wire n_3186;
wire n_1322;
wire n_640;
wire n_4129;
wire n_965;
wire n_1899;
wire n_1428;
wire n_4093;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_3965;
wire n_2632;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_540;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_4039;
wire n_3387;
wire n_2027;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_4197;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_629;
wire n_1621;
wire n_4275;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_4283;
wire n_900;
wire n_3504;
wire n_4194;
wire n_1449;
wire n_827;
wire n_531;
wire n_2912;
wire n_4272;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_649;
wire n_1742;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_456),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_89),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_35),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_394),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_308),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_321),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_216),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_141),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_260),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_69),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_324),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_125),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_226),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_267),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_119),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_302),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_425),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_115),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_433),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_419),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_81),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_406),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_113),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_393),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_59),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_304),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_283),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_169),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_431),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_388),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_417),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_350),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_464),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_225),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_116),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_133),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_83),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_355),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_155),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_387),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_382),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_231),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_373),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_113),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_23),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_328),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_368),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_230),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_451),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_372),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_412),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_268),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_465),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_200),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_352),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_195),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_105),
.Y(n_523)
);

BUFx10_ASAP7_75t_L g524 ( 
.A(n_13),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_386),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_43),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_88),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_385),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_230),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_103),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_340),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_20),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_212),
.Y(n_533)
);

INVx1_ASAP7_75t_SL g534 ( 
.A(n_365),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_295),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_218),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_174),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_375),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_317),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_337),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_445),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_391),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_97),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_252),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_242),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_149),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_102),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_60),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_281),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_291),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_315),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g552 ( 
.A(n_357),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_284),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_43),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_354),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_398),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_438),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_244),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_260),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_182),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_79),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_423),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_436),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_347),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_397),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_295),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_59),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_152),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_285),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_216),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_336),
.Y(n_571)
);

BUFx10_ASAP7_75t_L g572 ( 
.A(n_318),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_179),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_269),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_422),
.Y(n_575)
);

CKINVDCx14_ASAP7_75t_R g576 ( 
.A(n_26),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_461),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_310),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_23),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_301),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_66),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_173),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_228),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_25),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_44),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_253),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_70),
.Y(n_587)
);

BUFx8_ASAP7_75t_SL g588 ( 
.A(n_172),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_101),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_362),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_136),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_98),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_20),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_185),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_159),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_145),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_121),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_275),
.Y(n_598)
);

CKINVDCx16_ASAP7_75t_R g599 ( 
.A(n_261),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_156),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_127),
.Y(n_601)
);

INVx1_ASAP7_75t_SL g602 ( 
.A(n_447),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_270),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_4),
.Y(n_604)
);

CKINVDCx16_ASAP7_75t_R g605 ( 
.A(n_303),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_348),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_404),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_409),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_341),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_390),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_400),
.Y(n_611)
);

BUFx5_ASAP7_75t_L g612 ( 
.A(n_85),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_127),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_228),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_206),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_74),
.Y(n_616)
);

BUFx10_ASAP7_75t_L g617 ( 
.A(n_70),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_421),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_65),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_283),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_290),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_41),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_143),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_109),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_74),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_428),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_408),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_41),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_334),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_33),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_183),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_93),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_148),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_134),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_443),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_299),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_245),
.Y(n_637)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_411),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_466),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_239),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_157),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_30),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_289),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_459),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_343),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_166),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_77),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_426),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_136),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_255),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_279),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_252),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_202),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_366),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_117),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_55),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_294),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_235),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_441),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_237),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_454),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_279),
.Y(n_662)
);

BUFx2_ASAP7_75t_SL g663 ( 
.A(n_153),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_167),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_170),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_233),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_15),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_198),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_143),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_106),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_64),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_114),
.Y(n_672)
);

INVx1_ASAP7_75t_SL g673 ( 
.A(n_305),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_432),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_392),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_128),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_162),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_174),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_18),
.Y(n_679)
);

CKINVDCx16_ASAP7_75t_R g680 ( 
.A(n_266),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_63),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_374),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_266),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_322),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_342),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_62),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_314),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_49),
.Y(n_688)
);

CKINVDCx20_ASAP7_75t_R g689 ( 
.A(n_181),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_110),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_38),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_207),
.Y(n_692)
);

CKINVDCx14_ASAP7_75t_R g693 ( 
.A(n_178),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_281),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_414),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_167),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_68),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_405),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_12),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_182),
.Y(n_700)
);

CKINVDCx16_ASAP7_75t_R g701 ( 
.A(n_60),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_108),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_233),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_186),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_108),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_10),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_131),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_290),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_319),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_439),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_64),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_94),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_251),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_379),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_86),
.Y(n_715)
);

BUFx2_ASAP7_75t_SL g716 ( 
.A(n_53),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_6),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_178),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_220),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_395),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_44),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_371),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_10),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_103),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_194),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_238),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_30),
.Y(n_727)
);

CKINVDCx16_ASAP7_75t_R g728 ( 
.A(n_248),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_282),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_131),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_259),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_410),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_76),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_42),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_455),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_449),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_91),
.Y(n_737)
);

BUFx10_ASAP7_75t_L g738 ( 
.A(n_147),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_353),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_125),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_420),
.Y(n_741)
);

CKINVDCx16_ASAP7_75t_R g742 ( 
.A(n_293),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_112),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_80),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_65),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_282),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_284),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_416),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_267),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_235),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_138),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_46),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_286),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_165),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_227),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_185),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_82),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_294),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_229),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_446),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_148),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_659),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_612),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_612),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_612),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_612),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_588),
.Y(n_767)
);

INVxp67_ASAP7_75t_SL g768 ( 
.A(n_626),
.Y(n_768)
);

CKINVDCx14_ASAP7_75t_R g769 ( 
.A(n_576),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_612),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_467),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_612),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_471),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_477),
.Y(n_774)
);

INVxp33_ASAP7_75t_SL g775 ( 
.A(n_679),
.Y(n_775)
);

CKINVDCx20_ASAP7_75t_R g776 ( 
.A(n_495),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_612),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_485),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_612),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_612),
.Y(n_780)
);

CKINVDCx20_ASAP7_75t_R g781 ( 
.A(n_557),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_536),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_536),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_536),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_492),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_536),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_536),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_536),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_546),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_546),
.Y(n_790)
);

INVx1_ASAP7_75t_SL g791 ( 
.A(n_637),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_546),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_546),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_515),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_546),
.Y(n_795)
);

CKINVDCx20_ASAP7_75t_R g796 ( 
.A(n_565),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_637),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_546),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_496),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_569),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_569),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_498),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_569),
.Y(n_803)
);

INVxp67_ASAP7_75t_SL g804 ( 
.A(n_626),
.Y(n_804)
);

INVxp67_ASAP7_75t_SL g805 ( 
.A(n_659),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_569),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_569),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_569),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_613),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_613),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_613),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_613),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_613),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_613),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_730),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_730),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_730),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_730),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_730),
.Y(n_819)
);

INVxp33_ASAP7_75t_L g820 ( 
.A(n_758),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_730),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_615),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_615),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_646),
.Y(n_824)
);

CKINVDCx16_ASAP7_75t_R g825 ( 
.A(n_693),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_646),
.Y(n_826)
);

INVxp67_ASAP7_75t_SL g827 ( 
.A(n_515),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_606),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_683),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_683),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_705),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_705),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_749),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_749),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_553),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_553),
.Y(n_836)
);

CKINVDCx20_ASAP7_75t_R g837 ( 
.A(n_607),
.Y(n_837)
);

CKINVDCx20_ASAP7_75t_R g838 ( 
.A(n_638),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_553),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_598),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_598),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_598),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_474),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_474),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_472),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_478),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_478),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_479),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_504),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_507),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_479),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_509),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_484),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_472),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_484),
.Y(n_855)
);

CKINVDCx16_ASAP7_75t_R g856 ( 
.A(n_599),
.Y(n_856)
);

INVxp67_ASAP7_75t_SL g857 ( 
.A(n_515),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_489),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_482),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_482),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_489),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_508),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_508),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_523),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_523),
.Y(n_865)
);

INVxp67_ASAP7_75t_SL g866 ( 
.A(n_563),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_605),
.Y(n_867)
);

INVxp33_ASAP7_75t_SL g868 ( 
.A(n_758),
.Y(n_868)
);

CKINVDCx16_ASAP7_75t_R g869 ( 
.A(n_599),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_530),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_530),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_532),
.Y(n_872)
);

BUFx2_ASAP7_75t_L g873 ( 
.A(n_570),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_532),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_535),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_512),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_535),
.Y(n_877)
);

INVxp67_ASAP7_75t_L g878 ( 
.A(n_663),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_537),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_537),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_545),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_513),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_545),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_483),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_680),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_483),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_554),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_554),
.Y(n_888)
);

NOR2xp67_ASAP7_75t_L g889 ( 
.A(n_548),
.B(n_0),
.Y(n_889)
);

INVxp33_ASAP7_75t_L g890 ( 
.A(n_558),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_558),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_680),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_559),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_559),
.Y(n_894)
);

INVxp67_ASAP7_75t_SL g895 ( 
.A(n_563),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_486),
.Y(n_896)
);

INVxp67_ASAP7_75t_SL g897 ( 
.A(n_563),
.Y(n_897)
);

INVxp67_ASAP7_75t_SL g898 ( 
.A(n_629),
.Y(n_898)
);

CKINVDCx14_ASAP7_75t_R g899 ( 
.A(n_524),
.Y(n_899)
);

INVxp67_ASAP7_75t_L g900 ( 
.A(n_663),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_486),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_561),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_561),
.Y(n_903)
);

INVxp67_ASAP7_75t_SL g904 ( 
.A(n_629),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_516),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_566),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_519),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_566),
.Y(n_908)
);

INVxp33_ASAP7_75t_L g909 ( 
.A(n_579),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_579),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_784),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_784),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_782),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_782),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_788),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_788),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_783),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_800),
.Y(n_918)
);

AND2x2_ASAP7_75t_SL g919 ( 
.A(n_825),
.B(n_605),
.Y(n_919)
);

INVx6_ASAP7_75t_L g920 ( 
.A(n_762),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_783),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_800),
.Y(n_922)
);

OA21x2_ASAP7_75t_L g923 ( 
.A1(n_786),
.A2(n_497),
.B(n_490),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_827),
.B(n_570),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_786),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_794),
.B(n_556),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_801),
.Y(n_927)
);

INVxp67_ASAP7_75t_SL g928 ( 
.A(n_845),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_857),
.B(n_755),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_801),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_866),
.B(n_755),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_810),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_769),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_810),
.Y(n_934)
);

INVx5_ASAP7_75t_L g935 ( 
.A(n_794),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_787),
.Y(n_936)
);

AND2x6_ASAP7_75t_L g937 ( 
.A(n_763),
.B(n_488),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_821),
.Y(n_938)
);

INVx5_ASAP7_75t_L g939 ( 
.A(n_794),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_821),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_787),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_825),
.B(n_701),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_789),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_763),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_789),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_790),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_885),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_764),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_895),
.B(n_584),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_790),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_771),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_792),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_794),
.B(n_556),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_897),
.B(n_564),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_764),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_792),
.Y(n_956)
);

OA21x2_ASAP7_75t_L g957 ( 
.A1(n_793),
.A2(n_497),
.B(n_490),
.Y(n_957)
);

NOR2x1_ASAP7_75t_L g958 ( 
.A(n_793),
.B(n_629),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_795),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_795),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_868),
.A2(n_728),
.B1(n_742),
.B2(n_701),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_768),
.B(n_564),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_798),
.Y(n_963)
);

INVx5_ASAP7_75t_L g964 ( 
.A(n_845),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_839),
.B(n_488),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_798),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_765),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_803),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_773),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_892),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_803),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_806),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_806),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_898),
.B(n_904),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_765),
.Y(n_975)
);

BUFx12f_ASAP7_75t_L g976 ( 
.A(n_767),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_766),
.Y(n_977)
);

BUFx12f_ASAP7_75t_L g978 ( 
.A(n_774),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_807),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_766),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_770),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_SL g982 ( 
.A1(n_856),
.A2(n_550),
.B1(n_585),
.B2(n_567),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_807),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_808),
.Y(n_984)
);

BUFx8_ASAP7_75t_L g985 ( 
.A(n_797),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_808),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_809),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_839),
.B(n_842),
.Y(n_988)
);

INVx5_ASAP7_75t_L g989 ( 
.A(n_854),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_778),
.Y(n_990)
);

OAI21x1_ASAP7_75t_L g991 ( 
.A1(n_770),
.A2(n_580),
.B(n_542),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_804),
.B(n_506),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_791),
.A2(n_742),
.B1(n_728),
.B2(n_636),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_785),
.Y(n_994)
);

BUFx2_ASAP7_75t_L g995 ( 
.A(n_867),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_809),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_811),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_811),
.Y(n_998)
);

OA21x2_ASAP7_75t_L g999 ( 
.A1(n_812),
.A2(n_814),
.B(n_813),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_775),
.A2(n_664),
.B1(n_689),
.B2(n_676),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_812),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_842),
.B(n_542),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_813),
.Y(n_1003)
);

INVx5_ASAP7_75t_L g1004 ( 
.A(n_854),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_814),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_820),
.A2(n_724),
.B1(n_475),
.B2(n_668),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_815),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_815),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_772),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_816),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_816),
.Y(n_1011)
);

OAI21x1_ASAP7_75t_L g1012 ( 
.A1(n_772),
.A2(n_709),
.B(n_580),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_817),
.Y(n_1013)
);

NAND2x1p5_ASAP7_75t_L g1014 ( 
.A(n_889),
.B(n_709),
.Y(n_1014)
);

BUFx3_ASAP7_75t_L g1015 ( 
.A(n_762),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_805),
.B(n_584),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_835),
.B(n_521),
.Y(n_1017)
);

BUFx8_ASAP7_75t_L g1018 ( 
.A(n_797),
.Y(n_1018)
);

BUFx2_ASAP7_75t_L g1019 ( 
.A(n_873),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_777),
.Y(n_1020)
);

INVxp33_ASAP7_75t_SL g1021 ( 
.A(n_799),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_777),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_779),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_802),
.B(n_534),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_779),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_817),
.Y(n_1026)
);

INVx5_ASAP7_75t_L g1027 ( 
.A(n_859),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_835),
.Y(n_1028)
);

INVx2_ASAP7_75t_SL g1029 ( 
.A(n_873),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_818),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_818),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_836),
.B(n_840),
.Y(n_1032)
);

XNOR2x2_ASAP7_75t_L g1033 ( 
.A(n_843),
.B(n_586),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_819),
.Y(n_1034)
);

INVx5_ASAP7_75t_L g1035 ( 
.A(n_859),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_1019),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_928),
.Y(n_1037)
);

NAND2xp33_ASAP7_75t_SL g1038 ( 
.A(n_1029),
.B(n_668),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_911),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_1015),
.B(n_836),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_1019),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_944),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1032),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_1015),
.B(n_840),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_1015),
.B(n_1028),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1032),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_974),
.B(n_841),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_920),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_974),
.B(n_849),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_911),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_918),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_911),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_912),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_944),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_918),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_928),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_1024),
.B(n_850),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_948),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_948),
.Y(n_1059)
);

CKINVDCx6p67_ASAP7_75t_R g1060 ( 
.A(n_976),
.Y(n_1060)
);

INVx2_ASAP7_75t_SL g1061 ( 
.A(n_920),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_948),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_992),
.B(n_852),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_948),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_955),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_912),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_929),
.B(n_876),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_918),
.Y(n_1068)
);

XNOR2x2_ASAP7_75t_L g1069 ( 
.A(n_1033),
.B(n_586),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_962),
.A2(n_899),
.B1(n_869),
.B2(n_856),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_955),
.Y(n_1071)
);

OA21x2_ASAP7_75t_L g1072 ( 
.A1(n_991),
.A2(n_780),
.B(n_819),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_929),
.B(n_882),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_912),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_955),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_931),
.B(n_905),
.Y(n_1076)
);

BUFx8_ASAP7_75t_L g1077 ( 
.A(n_995),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_955),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1023),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_918),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_1028),
.B(n_841),
.Y(n_1081)
);

BUFx2_ASAP7_75t_L g1082 ( 
.A(n_970),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_SL g1083 ( 
.A1(n_982),
.A2(n_869),
.B1(n_781),
.B2(n_796),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_931),
.B(n_907),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_944),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1023),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_944),
.Y(n_1087)
);

NAND2x1_ASAP7_75t_L g1088 ( 
.A(n_999),
.B(n_923),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1023),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_949),
.B(n_860),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_918),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_949),
.B(n_860),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_920),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_918),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_991),
.A2(n_780),
.B(n_884),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1023),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_988),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_944),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_922),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_944),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_988),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_922),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1028),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_913),
.Y(n_1104)
);

NAND2xp33_ASAP7_75t_L g1105 ( 
.A(n_1014),
.B(n_499),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_913),
.Y(n_1106)
);

NOR2x1_ASAP7_75t_L g1107 ( 
.A(n_933),
.B(n_884),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1016),
.B(n_886),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_965),
.B(n_823),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_914),
.Y(n_1110)
);

CKINVDCx8_ASAP7_75t_R g1111 ( 
.A(n_995),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_922),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_914),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1016),
.B(n_886),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_917),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_917),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_921),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_938),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_921),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_965),
.B(n_823),
.Y(n_1120)
);

AND2x4_ASAP7_75t_L g1121 ( 
.A(n_965),
.B(n_829),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_925),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_924),
.B(n_896),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1014),
.B(n_1017),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_965),
.B(n_829),
.Y(n_1125)
);

INVxp67_ASAP7_75t_L g1126 ( 
.A(n_970),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_925),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_936),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_936),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_938),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_945),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_915),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_915),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_945),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_938),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_959),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_944),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_959),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_915),
.Y(n_1139)
);

INVx3_ASAP7_75t_L g1140 ( 
.A(n_915),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1014),
.B(n_896),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_960),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_960),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_966),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_966),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_967),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1014),
.B(n_901),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_998),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_998),
.Y(n_1149)
);

OA21x2_ASAP7_75t_L g1150 ( 
.A1(n_991),
.A2(n_901),
.B(n_517),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1017),
.B(n_552),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_940),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_1029),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_940),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_915),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1003),
.Y(n_1156)
);

BUFx8_ASAP7_75t_L g1157 ( 
.A(n_933),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_940),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1003),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1007),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_1029),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_924),
.B(n_602),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1007),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_941),
.Y(n_1164)
);

AND2x6_ASAP7_75t_L g1165 ( 
.A(n_1002),
.B(n_499),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1030),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_1002),
.B(n_517),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1030),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1002),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_954),
.B(n_673),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_941),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_954),
.B(n_1002),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_947),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_967),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_967),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_926),
.B(n_900),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_941),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_958),
.B(n_525),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_943),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_943),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_967),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_915),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_915),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_943),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_999),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_920),
.B(n_975),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_967),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_951),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_999),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_946),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_999),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_967),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_999),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_967),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_975),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_969),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_975),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_975),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_975),
.Y(n_1199)
);

INVxp67_ASAP7_75t_L g1200 ( 
.A(n_942),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_946),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_946),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_975),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_975),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_977),
.Y(n_1205)
);

NAND2x1_ASAP7_75t_L g1206 ( 
.A(n_923),
.B(n_525),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_956),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_977),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_956),
.Y(n_1209)
);

OR2x2_ASAP7_75t_L g1210 ( 
.A(n_947),
.B(n_878),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1012),
.A2(n_541),
.B(n_539),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_977),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_977),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_956),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_977),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_985),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_977),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_977),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_961),
.A2(n_469),
.B1(n_473),
.B2(n_468),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_920),
.B(n_528),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_980),
.Y(n_1221)
);

AND2x6_ASAP7_75t_L g1222 ( 
.A(n_926),
.B(n_539),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1021),
.B(n_990),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_919),
.B(n_572),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_980),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_980),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_980),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_953),
.B(n_822),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_980),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_980),
.B(n_531),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_927),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_980),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_981),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_981),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_981),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_927),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_963),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_981),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_981),
.B(n_540),
.Y(n_1239)
);

CKINVDCx16_ASAP7_75t_R g1240 ( 
.A(n_978),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_963),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_981),
.Y(n_1242)
);

INVx6_ASAP7_75t_L g1243 ( 
.A(n_935),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1033),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_981),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_1009),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_1033),
.Y(n_1247)
);

HB1xp67_ASAP7_75t_L g1248 ( 
.A(n_985),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1009),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1009),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1009),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1009),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_958),
.B(n_541),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1009),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1009),
.B(n_551),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1012),
.A2(n_571),
.B(n_562),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1020),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1020),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_SL g1259 ( 
.A(n_919),
.B(n_572),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_963),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1095),
.Y(n_1261)
);

INVxp33_ASAP7_75t_SL g1262 ( 
.A(n_1083),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1123),
.B(n_919),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1048),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1095),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1097),
.B(n_1020),
.Y(n_1266)
);

AND2x2_ASAP7_75t_SL g1267 ( 
.A(n_1105),
.B(n_562),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1169),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1097),
.A2(n_957),
.B1(n_923),
.B2(n_937),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1104),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1150),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1101),
.B(n_1020),
.Y(n_1272)
);

INVx1_ASAP7_75t_SL g1273 ( 
.A(n_1041),
.Y(n_1273)
);

INVx1_ASAP7_75t_SL g1274 ( 
.A(n_1082),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1104),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1106),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1057),
.B(n_994),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_1063),
.B(n_978),
.Y(n_1278)
);

INVxp67_ASAP7_75t_SL g1279 ( 
.A(n_1042),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1067),
.B(n_978),
.Y(n_1280)
);

CKINVDCx20_ASAP7_75t_R g1281 ( 
.A(n_1111),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1106),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1045),
.Y(n_1283)
);

INVx2_ASAP7_75t_SL g1284 ( 
.A(n_1153),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1110),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1110),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_SL g1287 ( 
.A(n_1223),
.B(n_976),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1123),
.B(n_923),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1101),
.B(n_1020),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1113),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1113),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1172),
.B(n_1020),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1228),
.B(n_923),
.Y(n_1293)
);

AND2x6_ASAP7_75t_L g1294 ( 
.A(n_1185),
.B(n_571),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1115),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1045),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1115),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1116),
.Y(n_1298)
);

BUFx6f_ASAP7_75t_L g1299 ( 
.A(n_1048),
.Y(n_1299)
);

AND2x6_ASAP7_75t_L g1300 ( 
.A(n_1185),
.B(n_1189),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1116),
.Y(n_1301)
);

AND2x6_ASAP7_75t_L g1302 ( 
.A(n_1189),
.B(n_575),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1049),
.B(n_776),
.Y(n_1303)
);

CKINVDCx14_ASAP7_75t_R g1304 ( 
.A(n_1060),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1117),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1172),
.B(n_1020),
.Y(n_1306)
);

BUFx4f_ASAP7_75t_L g1307 ( 
.A(n_1222),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1073),
.B(n_828),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1076),
.B(n_1084),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1117),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_1093),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1210),
.B(n_993),
.Y(n_1312)
);

CKINVDCx8_ASAP7_75t_R g1313 ( 
.A(n_1240),
.Y(n_1313)
);

XNOR2xp5_ASAP7_75t_L g1314 ( 
.A(n_1069),
.B(n_982),
.Y(n_1314)
);

INVx5_ASAP7_75t_L g1315 ( 
.A(n_1243),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1105),
.A2(n_957),
.B1(n_937),
.B2(n_993),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1119),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1228),
.B(n_957),
.Y(n_1318)
);

INVx3_ASAP7_75t_L g1319 ( 
.A(n_1150),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1119),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1148),
.Y(n_1321)
);

BUFx3_ASAP7_75t_L g1322 ( 
.A(n_1045),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1148),
.Y(n_1323)
);

INVxp33_ASAP7_75t_L g1324 ( 
.A(n_1082),
.Y(n_1324)
);

INVxp67_ASAP7_75t_SL g1325 ( 
.A(n_1042),
.Y(n_1325)
);

INVx3_ASAP7_75t_L g1326 ( 
.A(n_1150),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1058),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1150),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1103),
.Y(n_1329)
);

INVx5_ASAP7_75t_L g1330 ( 
.A(n_1243),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1103),
.Y(n_1331)
);

AOI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1176),
.A2(n_837),
.B1(n_838),
.B2(n_961),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_1188),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_SL g1334 ( 
.A(n_1162),
.B(n_985),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1200),
.B(n_1006),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1151),
.B(n_1006),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1109),
.Y(n_1337)
);

AND2x2_ASAP7_75t_SL g1338 ( 
.A(n_1244),
.B(n_575),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1109),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1109),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_SL g1341 ( 
.A(n_1170),
.B(n_985),
.Y(n_1341)
);

INVx3_ASAP7_75t_L g1342 ( 
.A(n_1072),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_1188),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1120),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1120),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1167),
.A2(n_957),
.B1(n_937),
.B2(n_577),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1124),
.B(n_1022),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1161),
.B(n_1000),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1120),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1108),
.B(n_957),
.Y(n_1350)
);

NAND2xp33_ASAP7_75t_L g1351 ( 
.A(n_1191),
.B(n_937),
.Y(n_1351)
);

INVx4_ASAP7_75t_L g1352 ( 
.A(n_1042),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1126),
.B(n_1000),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1036),
.Y(n_1354)
);

BUFx10_ASAP7_75t_L g1355 ( 
.A(n_1196),
.Y(n_1355)
);

INVx4_ASAP7_75t_L g1356 ( 
.A(n_1042),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1058),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1059),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1121),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1167),
.A2(n_937),
.B1(n_577),
.B2(n_609),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1173),
.B(n_1018),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_SL g1362 ( 
.A(n_1176),
.B(n_1018),
.Y(n_1362)
);

INVx4_ASAP7_75t_L g1363 ( 
.A(n_1042),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1040),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1121),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1043),
.A2(n_470),
.B1(n_953),
.B2(n_609),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1121),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1125),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1210),
.B(n_1018),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_1072),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1125),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_SL g1372 ( 
.A(n_1108),
.B(n_1018),
.Y(n_1372)
);

INVx1_ASAP7_75t_SL g1373 ( 
.A(n_1196),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1125),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1090),
.B(n_1092),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1069),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1167),
.A2(n_937),
.B1(n_639),
.B2(n_675),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1040),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1046),
.A2(n_578),
.B1(n_675),
.B2(n_639),
.Y(n_1379)
);

NAND3xp33_ASAP7_75t_L g1380 ( 
.A(n_1038),
.B(n_480),
.C(n_476),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1040),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1044),
.Y(n_1382)
);

INVx1_ASAP7_75t_SL g1383 ( 
.A(n_1038),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1044),
.Y(n_1384)
);

BUFx3_ASAP7_75t_L g1385 ( 
.A(n_1044),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1090),
.B(n_1022),
.Y(n_1386)
);

INVx1_ASAP7_75t_SL g1387 ( 
.A(n_1107),
.Y(n_1387)
);

INVx4_ASAP7_75t_L g1388 ( 
.A(n_1054),
.Y(n_1388)
);

INVxp67_ASAP7_75t_L g1389 ( 
.A(n_1070),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1247),
.B(n_890),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1081),
.Y(n_1391)
);

INVx4_ASAP7_75t_L g1392 ( 
.A(n_1054),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1039),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1059),
.Y(n_1394)
);

AND2x6_ASAP7_75t_L g1395 ( 
.A(n_1191),
.B(n_1193),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1114),
.B(n_909),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1062),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1062),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1039),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_SL g1400 ( 
.A(n_1114),
.B(n_1092),
.Y(n_1400)
);

AOI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1047),
.A2(n_538),
.B1(n_590),
.B2(n_555),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1047),
.B(n_1037),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1064),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1219),
.B(n_716),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1050),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1064),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1050),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1081),
.B(n_1037),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1224),
.B(n_716),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_SL g1410 ( 
.A(n_1056),
.B(n_608),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1259),
.B(n_976),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1122),
.B(n_481),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1193),
.B(n_1022),
.Y(n_1413)
);

INVx4_ASAP7_75t_L g1414 ( 
.A(n_1054),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1065),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1065),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1071),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1081),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1141),
.B(n_1022),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1052),
.Y(n_1420)
);

INVxp67_ASAP7_75t_SL g1421 ( 
.A(n_1054),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1052),
.Y(n_1422)
);

OAI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1147),
.A2(n_695),
.B1(n_714),
.B2(n_578),
.Y(n_1423)
);

INVx2_ASAP7_75t_SL g1424 ( 
.A(n_1178),
.Y(n_1424)
);

INVx3_ASAP7_75t_L g1425 ( 
.A(n_1072),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1127),
.B(n_1022),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1072),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1128),
.B(n_1022),
.Y(n_1428)
);

BUFx10_ASAP7_75t_L g1429 ( 
.A(n_1178),
.Y(n_1429)
);

INVx4_ASAP7_75t_L g1430 ( 
.A(n_1054),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1129),
.B(n_1022),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1131),
.B(n_1025),
.Y(n_1432)
);

INVx5_ASAP7_75t_L g1433 ( 
.A(n_1243),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1053),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1071),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1053),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1075),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1066),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1066),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1074),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1074),
.Y(n_1441)
);

INVx4_ASAP7_75t_L g1442 ( 
.A(n_1085),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1134),
.B(n_1025),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1099),
.Y(n_1444)
);

INVx1_ASAP7_75t_SL g1445 ( 
.A(n_1060),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1093),
.B(n_695),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1165),
.A2(n_937),
.B1(n_735),
.B2(n_736),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1136),
.B(n_487),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1075),
.Y(n_1449)
);

INVxp67_ASAP7_75t_SL g1450 ( 
.A(n_1085),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1099),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1102),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1102),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1077),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1112),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1216),
.B(n_843),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1165),
.A2(n_937),
.B1(n_735),
.B2(n_736),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1112),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1178),
.B(n_844),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_SL g1460 ( 
.A(n_1253),
.B(n_610),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1157),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1078),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1138),
.B(n_1025),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_1157),
.Y(n_1464)
);

INVx2_ASAP7_75t_SL g1465 ( 
.A(n_1253),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1118),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_L g1467 ( 
.A(n_1142),
.B(n_491),
.Y(n_1467)
);

BUFx10_ASAP7_75t_L g1468 ( 
.A(n_1253),
.Y(n_1468)
);

NAND2xp33_ASAP7_75t_L g1469 ( 
.A(n_1165),
.B(n_937),
.Y(n_1469)
);

INVx4_ASAP7_75t_L g1470 ( 
.A(n_1085),
.Y(n_1470)
);

INVx4_ASAP7_75t_L g1471 ( 
.A(n_1085),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1078),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1079),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1079),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1143),
.B(n_611),
.Y(n_1475)
);

INVxp33_ASAP7_75t_SL g1476 ( 
.A(n_1248),
.Y(n_1476)
);

INVx3_ASAP7_75t_L g1477 ( 
.A(n_1088),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1118),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1144),
.B(n_618),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1086),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1145),
.B(n_844),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1086),
.Y(n_1482)
);

NAND2x1_ASAP7_75t_L g1483 ( 
.A(n_1132),
.B(n_1025),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1149),
.B(n_1025),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1156),
.B(n_1025),
.Y(n_1485)
);

BUFx6f_ASAP7_75t_L g1486 ( 
.A(n_1088),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1216),
.B(n_846),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1077),
.Y(n_1488)
);

INVxp67_ASAP7_75t_SL g1489 ( 
.A(n_1085),
.Y(n_1489)
);

INVx4_ASAP7_75t_L g1490 ( 
.A(n_1087),
.Y(n_1490)
);

INVx4_ASAP7_75t_L g1491 ( 
.A(n_1087),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1159),
.B(n_493),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1160),
.B(n_846),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1163),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1166),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1168),
.Y(n_1496)
);

OR2x6_ASAP7_75t_L g1497 ( 
.A(n_1206),
.B(n_714),
.Y(n_1497)
);

INVxp33_ASAP7_75t_L g1498 ( 
.A(n_1111),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1089),
.B(n_1025),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_L g1500 ( 
.A(n_1087),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1130),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1089),
.B(n_935),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1157),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1096),
.B(n_935),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1096),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_SL g1506 ( 
.A(n_1424),
.B(n_1186),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1375),
.B(n_1222),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1359),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1408),
.B(n_1222),
.Y(n_1509)
);

NOR2xp67_ASAP7_75t_L g1510 ( 
.A(n_1333),
.B(n_1220),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1408),
.B(n_1222),
.Y(n_1511)
);

NAND3xp33_ASAP7_75t_L g1512 ( 
.A(n_1336),
.B(n_1348),
.C(n_1335),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1359),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_SL g1514 ( 
.A(n_1424),
.B(n_1194),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1465),
.A2(n_1206),
.B1(n_1061),
.B2(n_1230),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1396),
.B(n_524),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1376),
.A2(n_1222),
.B1(n_1165),
.B2(n_591),
.Y(n_1517)
);

OAI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1465),
.A2(n_741),
.B1(n_739),
.B2(n_1239),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1270),
.Y(n_1519)
);

BUFx2_ASAP7_75t_L g1520 ( 
.A(n_1273),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1274),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1376),
.A2(n_1222),
.B1(n_1165),
.B2(n_591),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1277),
.B(n_1255),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1408),
.B(n_1459),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1459),
.B(n_1194),
.Y(n_1525)
);

NOR3xp33_ASAP7_75t_L g1526 ( 
.A(n_1303),
.B(n_741),
.C(n_739),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1309),
.B(n_1195),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1365),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1353),
.B(n_1390),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_SL g1530 ( 
.A(n_1284),
.B(n_1429),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1275),
.B(n_1195),
.Y(n_1531)
);

INVxp67_ASAP7_75t_SL g1532 ( 
.A(n_1486),
.Y(n_1532)
);

NAND3xp33_ASAP7_75t_L g1533 ( 
.A(n_1314),
.B(n_1077),
.C(n_500),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1275),
.B(n_1197),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_SL g1535 ( 
.A(n_1284),
.B(n_1061),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1365),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1282),
.B(n_1197),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_R g1538 ( 
.A(n_1333),
.B(n_1165),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1270),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_SL g1540 ( 
.A(n_1429),
.B(n_1468),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1367),
.Y(n_1541)
);

NOR3xp33_ASAP7_75t_L g1542 ( 
.A(n_1308),
.B(n_501),
.C(n_494),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1367),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1276),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1276),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1286),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1282),
.B(n_1198),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1285),
.B(n_1198),
.Y(n_1548)
);

BUFx6f_ASAP7_75t_L g1549 ( 
.A(n_1283),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_L g1550 ( 
.A(n_1390),
.B(n_1199),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_SL g1551 ( 
.A(n_1429),
.B(n_1199),
.Y(n_1551)
);

A2O1A1Ixp33_ASAP7_75t_L g1552 ( 
.A1(n_1263),
.A2(n_1211),
.B(n_1256),
.C(n_1012),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1285),
.B(n_1204),
.Y(n_1553)
);

O2A1O1Ixp33_ASAP7_75t_L g1554 ( 
.A1(n_1400),
.A2(n_1171),
.B(n_1177),
.C(n_1164),
.Y(n_1554)
);

NOR2x1p5_ASAP7_75t_L g1555 ( 
.A(n_1461),
.B(n_502),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1396),
.B(n_524),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1337),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1286),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1291),
.B(n_1204),
.Y(n_1559)
);

INVxp67_ASAP7_75t_SL g1560 ( 
.A(n_1486),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1263),
.B(n_1205),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1291),
.B(n_1205),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1312),
.B(n_1208),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1298),
.B(n_1208),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1290),
.Y(n_1565)
);

INVx3_ASAP7_75t_L g1566 ( 
.A(n_1283),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1338),
.A2(n_593),
.B1(n_600),
.B2(n_595),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1298),
.B(n_1235),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1301),
.B(n_1235),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1338),
.A2(n_593),
.B1(n_600),
.B2(n_595),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1290),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1312),
.B(n_1238),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1339),
.Y(n_1573)
);

NOR2x1p5_ASAP7_75t_L g1574 ( 
.A(n_1461),
.B(n_503),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1354),
.B(n_847),
.Y(n_1575)
);

O2A1O1Ixp5_ASAP7_75t_L g1576 ( 
.A1(n_1301),
.A2(n_1242),
.B(n_1245),
.C(n_1238),
.Y(n_1576)
);

BUFx5_ASAP7_75t_L g1577 ( 
.A(n_1300),
.Y(n_1577)
);

INVx3_ASAP7_75t_L g1578 ( 
.A(n_1296),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1320),
.B(n_1242),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1320),
.B(n_1245),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1321),
.B(n_1249),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1267),
.A2(n_1293),
.B1(n_1318),
.B2(n_1288),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1321),
.B(n_1249),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1323),
.B(n_1250),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1340),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1389),
.B(n_1250),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1344),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1323),
.B(n_1251),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1402),
.B(n_1251),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1347),
.A2(n_1098),
.B(n_1087),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1345),
.Y(n_1591)
);

INVx2_ASAP7_75t_SL g1592 ( 
.A(n_1456),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1387),
.B(n_1254),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1295),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1468),
.B(n_1254),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1383),
.B(n_1258),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1295),
.B(n_1258),
.Y(n_1597)
);

XOR2x2_ASAP7_75t_L g1598 ( 
.A(n_1314),
.B(n_1),
.Y(n_1598)
);

NAND2xp33_ASAP7_75t_L g1599 ( 
.A(n_1300),
.B(n_1087),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1404),
.B(n_1174),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1324),
.B(n_524),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1297),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1456),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1404),
.B(n_1175),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_SL g1605 ( 
.A(n_1468),
.B(n_935),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1349),
.Y(n_1606)
);

INVx4_ASAP7_75t_L g1607 ( 
.A(n_1296),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1409),
.B(n_1203),
.Y(n_1608)
);

NOR2xp67_ASAP7_75t_L g1609 ( 
.A(n_1343),
.B(n_847),
.Y(n_1609)
);

AO22x2_ASAP7_75t_L g1610 ( 
.A1(n_1409),
.A2(n_616),
.B1(n_620),
.B2(n_604),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_SL g1611 ( 
.A(n_1486),
.B(n_1098),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1368),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1371),
.Y(n_1613)
);

BUFx3_ASAP7_75t_L g1614 ( 
.A(n_1355),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1487),
.B(n_1212),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1267),
.A2(n_1217),
.B1(n_1218),
.B2(n_1215),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1297),
.B(n_1227),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_SL g1618 ( 
.A(n_1343),
.B(n_572),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1374),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1487),
.B(n_1332),
.Y(n_1620)
);

AOI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1391),
.A2(n_1225),
.B1(n_1226),
.B2(n_1221),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1305),
.B(n_1233),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1418),
.B(n_1364),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1327),
.Y(n_1624)
);

AOI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1378),
.A2(n_1232),
.B1(n_1257),
.B2(n_1229),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_SL g1626 ( 
.A(n_1418),
.B(n_1364),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1486),
.B(n_1098),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1305),
.B(n_1051),
.Y(n_1628)
);

INVxp67_ASAP7_75t_L g1629 ( 
.A(n_1412),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1310),
.B(n_1051),
.Y(n_1630)
);

O2A1O1Ixp33_ASAP7_75t_L g1631 ( 
.A1(n_1366),
.A2(n_1171),
.B(n_1177),
.C(n_1164),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1327),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1373),
.B(n_617),
.Y(n_1633)
);

NAND2xp33_ASAP7_75t_L g1634 ( 
.A(n_1300),
.B(n_1098),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1486),
.B(n_1098),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1357),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1357),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1310),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1385),
.B(n_935),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_SL g1640 ( 
.A(n_1385),
.B(n_935),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1317),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_SL g1642 ( 
.A(n_1322),
.B(n_935),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1317),
.B(n_1051),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1268),
.B(n_1055),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1358),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1494),
.B(n_1495),
.Y(n_1646)
);

NOR2xp67_ASAP7_75t_L g1647 ( 
.A(n_1411),
.B(n_848),
.Y(n_1647)
);

INVx8_ASAP7_75t_L g1648 ( 
.A(n_1300),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1358),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1300),
.B(n_1055),
.Y(n_1650)
);

NOR2xp67_ASAP7_75t_L g1651 ( 
.A(n_1369),
.B(n_848),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1498),
.B(n_1496),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1293),
.A2(n_604),
.B1(n_620),
.B2(n_616),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1394),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1394),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_SL g1656 ( 
.A(n_1322),
.B(n_939),
.Y(n_1656)
);

AOI22xp33_ASAP7_75t_L g1657 ( 
.A1(n_1318),
.A2(n_647),
.B1(n_650),
.B2(n_632),
.Y(n_1657)
);

INVxp67_ASAP7_75t_L g1658 ( 
.A(n_1448),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1397),
.Y(n_1659)
);

BUFx3_ASAP7_75t_L g1660 ( 
.A(n_1355),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_SL g1661 ( 
.A(n_1292),
.B(n_1100),
.Y(n_1661)
);

NAND2xp33_ASAP7_75t_L g1662 ( 
.A(n_1300),
.B(n_1100),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1397),
.Y(n_1663)
);

NOR3xp33_ASAP7_75t_L g1664 ( 
.A(n_1362),
.B(n_510),
.C(n_505),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_SL g1665 ( 
.A(n_1306),
.B(n_1100),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1398),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1398),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1395),
.B(n_1055),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1395),
.B(n_1068),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1381),
.A2(n_1080),
.B1(n_1091),
.B2(n_1068),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1403),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1395),
.B(n_1068),
.Y(n_1672)
);

OAI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1346),
.A2(n_1091),
.B1(n_1094),
.B2(n_1080),
.Y(n_1673)
);

OR2x6_ASAP7_75t_L g1674 ( 
.A(n_1503),
.B(n_1211),
.Y(n_1674)
);

AOI22x1_ASAP7_75t_L g1675 ( 
.A1(n_1288),
.A2(n_1236),
.B1(n_1231),
.B2(n_1133),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1403),
.Y(n_1676)
);

INVx8_ASAP7_75t_L g1677 ( 
.A(n_1395),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1355),
.B(n_617),
.Y(n_1678)
);

INVx2_ASAP7_75t_SL g1679 ( 
.A(n_1481),
.Y(n_1679)
);

OAI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1382),
.A2(n_647),
.B1(n_650),
.B2(n_632),
.Y(n_1680)
);

O2A1O1Ixp5_ASAP7_75t_L g1681 ( 
.A1(n_1266),
.A2(n_1091),
.B(n_1094),
.C(n_1080),
.Y(n_1681)
);

OAI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1413),
.A2(n_1256),
.B(n_1133),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1481),
.B(n_617),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_SL g1684 ( 
.A(n_1287),
.B(n_939),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1395),
.B(n_1094),
.Y(n_1685)
);

INVxp67_ASAP7_75t_L g1686 ( 
.A(n_1467),
.Y(n_1686)
);

BUFx6f_ASAP7_75t_L g1687 ( 
.A(n_1500),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1386),
.A2(n_1137),
.B(n_1100),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1406),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1406),
.Y(n_1690)
);

BUFx3_ASAP7_75t_L g1691 ( 
.A(n_1281),
.Y(n_1691)
);

BUFx6f_ASAP7_75t_L g1692 ( 
.A(n_1500),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1415),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1350),
.A2(n_665),
.B1(n_667),
.B2(n_662),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1395),
.B(n_1231),
.Y(n_1695)
);

NOR3xp33_ASAP7_75t_L g1696 ( 
.A(n_1334),
.B(n_514),
.C(n_511),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1415),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1280),
.B(n_851),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1493),
.B(n_617),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1416),
.Y(n_1700)
);

INVxp67_ASAP7_75t_L g1701 ( 
.A(n_1492),
.Y(n_1701)
);

OAI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1384),
.A2(n_665),
.B1(n_667),
.B2(n_662),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1329),
.B(n_1132),
.Y(n_1703)
);

BUFx5_ASAP7_75t_L g1704 ( 
.A(n_1294),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1331),
.B(n_1272),
.Y(n_1705)
);

INVxp67_ASAP7_75t_L g1706 ( 
.A(n_1380),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1289),
.B(n_1132),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1350),
.B(n_1133),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1416),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1477),
.B(n_1417),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1477),
.B(n_1139),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_SL g1712 ( 
.A(n_1361),
.B(n_939),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1477),
.B(n_1139),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1417),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1435),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1401),
.B(n_939),
.Y(n_1716)
);

NOR2xp33_ASAP7_75t_L g1717 ( 
.A(n_1278),
.B(n_1100),
.Y(n_1717)
);

NOR2xp67_ASAP7_75t_L g1718 ( 
.A(n_1341),
.B(n_1464),
.Y(n_1718)
);

BUFx10_ASAP7_75t_L g1719 ( 
.A(n_1464),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_1281),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1435),
.Y(n_1721)
);

INVx2_ASAP7_75t_SL g1722 ( 
.A(n_1493),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1437),
.Y(n_1723)
);

NAND2xp33_ASAP7_75t_L g1724 ( 
.A(n_1294),
.B(n_1302),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1437),
.B(n_1231),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1449),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_SL g1727 ( 
.A(n_1460),
.B(n_939),
.Y(n_1727)
);

OAI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1269),
.A2(n_1146),
.B1(n_1181),
.B2(n_1137),
.Y(n_1728)
);

INVx2_ASAP7_75t_SL g1729 ( 
.A(n_1446),
.Y(n_1729)
);

INVxp67_ASAP7_75t_L g1730 ( 
.A(n_1379),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_SL g1731 ( 
.A(n_1307),
.B(n_1137),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1449),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1462),
.B(n_1236),
.Y(n_1733)
);

INVx2_ASAP7_75t_SL g1734 ( 
.A(n_1446),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1462),
.B(n_1472),
.Y(n_1735)
);

BUFx3_ASAP7_75t_L g1736 ( 
.A(n_1503),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1472),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1473),
.B(n_1236),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1473),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1445),
.B(n_738),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_L g1741 ( 
.A(n_1410),
.B(n_1137),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1294),
.A2(n_669),
.B1(n_672),
.B2(n_670),
.Y(n_1742)
);

AOI221xp5_ASAP7_75t_L g1743 ( 
.A1(n_1262),
.A2(n_672),
.B1(n_678),
.B2(n_670),
.C(n_669),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1474),
.B(n_1139),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1474),
.B(n_1140),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1480),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1480),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_L g1748 ( 
.A(n_1372),
.B(n_1137),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1482),
.B(n_1140),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1523),
.B(n_1294),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1645),
.Y(n_1751)
);

BUFx12f_ASAP7_75t_L g1752 ( 
.A(n_1719),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1645),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1649),
.Y(n_1754)
);

BUFx3_ASAP7_75t_L g1755 ( 
.A(n_1520),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1649),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1654),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1654),
.Y(n_1758)
);

AOI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1512),
.A2(n_1529),
.B1(n_1620),
.B2(n_1523),
.Y(n_1759)
);

AND2x4_ASAP7_75t_L g1760 ( 
.A(n_1679),
.B(n_1446),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1563),
.B(n_1294),
.Y(n_1761)
);

AOI21xp5_ASAP7_75t_L g1762 ( 
.A1(n_1532),
.A2(n_1356),
.B(n_1352),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1666),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1529),
.B(n_1262),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1567),
.A2(n_1316),
.B1(n_1302),
.B2(n_1294),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_1720),
.Y(n_1766)
);

AOI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1620),
.A2(n_1629),
.B1(n_1686),
.B2(n_1658),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1666),
.Y(n_1768)
);

INVxp67_ASAP7_75t_L g1769 ( 
.A(n_1521),
.Y(n_1769)
);

BUFx4f_ASAP7_75t_L g1770 ( 
.A(n_1549),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1676),
.Y(n_1771)
);

NAND2xp33_ASAP7_75t_L g1772 ( 
.A(n_1577),
.B(n_1302),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1676),
.Y(n_1773)
);

AO22x1_ASAP7_75t_L g1774 ( 
.A1(n_1526),
.A2(n_1476),
.B1(n_1488),
.B2(n_1454),
.Y(n_1774)
);

NAND2xp33_ASAP7_75t_L g1775 ( 
.A(n_1577),
.B(n_1302),
.Y(n_1775)
);

INVx3_ASAP7_75t_L g1776 ( 
.A(n_1687),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_R g1777 ( 
.A(n_1614),
.B(n_1304),
.Y(n_1777)
);

BUFx6f_ASAP7_75t_L g1778 ( 
.A(n_1687),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_SL g1779 ( 
.A(n_1577),
.B(n_1307),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1693),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1693),
.Y(n_1781)
);

OAI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1722),
.A2(n_1497),
.B1(n_1307),
.B2(n_1482),
.Y(n_1782)
);

INVx3_ASAP7_75t_L g1783 ( 
.A(n_1687),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1697),
.Y(n_1784)
);

INVx5_ASAP7_75t_L g1785 ( 
.A(n_1648),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1563),
.B(n_1302),
.Y(n_1786)
);

CKINVDCx5p33_ASAP7_75t_R g1787 ( 
.A(n_1691),
.Y(n_1787)
);

INVx3_ASAP7_75t_L g1788 ( 
.A(n_1687),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_1691),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1697),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1709),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1709),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1714),
.Y(n_1793)
);

BUFx3_ASAP7_75t_L g1794 ( 
.A(n_1736),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1603),
.B(n_1454),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_SL g1796 ( 
.A(n_1577),
.B(n_1505),
.Y(n_1796)
);

BUFx3_ASAP7_75t_L g1797 ( 
.A(n_1736),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_SL g1798 ( 
.A(n_1577),
.B(n_1500),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1714),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1721),
.Y(n_1800)
);

OR2x6_ASAP7_75t_L g1801 ( 
.A(n_1648),
.B(n_1488),
.Y(n_1801)
);

BUFx3_ASAP7_75t_L g1802 ( 
.A(n_1614),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1721),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1519),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1624),
.Y(n_1805)
);

OR2x2_ASAP7_75t_SL g1806 ( 
.A(n_1533),
.B(n_1313),
.Y(n_1806)
);

INVx3_ASAP7_75t_L g1807 ( 
.A(n_1692),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1519),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1632),
.Y(n_1809)
);

AO22x1_ASAP7_75t_L g1810 ( 
.A1(n_1696),
.A2(n_1476),
.B1(n_1302),
.B2(n_520),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1567),
.A2(n_1423),
.B1(n_1497),
.B2(n_678),
.Y(n_1811)
);

AND2x6_ASAP7_75t_L g1812 ( 
.A(n_1509),
.B(n_1328),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1539),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1572),
.B(n_1342),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1636),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1572),
.B(n_1342),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1550),
.B(n_1342),
.Y(n_1817)
);

INVxp67_ASAP7_75t_L g1818 ( 
.A(n_1652),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1550),
.B(n_1370),
.Y(n_1819)
);

INVx3_ASAP7_75t_L g1820 ( 
.A(n_1692),
.Y(n_1820)
);

NOR3xp33_ASAP7_75t_SL g1821 ( 
.A(n_1743),
.B(n_522),
.C(n_518),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1701),
.B(n_1370),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_SL g1823 ( 
.A1(n_1618),
.A2(n_572),
.B1(n_738),
.B2(n_527),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1539),
.Y(n_1824)
);

INVx3_ASAP7_75t_L g1825 ( 
.A(n_1692),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_SL g1826 ( 
.A(n_1577),
.B(n_1500),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1637),
.Y(n_1827)
);

NAND2xp33_ASAP7_75t_SL g1828 ( 
.A(n_1538),
.B(n_1328),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_SL g1829 ( 
.A(n_1524),
.B(n_1500),
.Y(n_1829)
);

BUFx3_ASAP7_75t_L g1830 ( 
.A(n_1660),
.Y(n_1830)
);

AOI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1542),
.A2(n_1475),
.B1(n_1479),
.B2(n_1351),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1655),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1646),
.B(n_1370),
.Y(n_1833)
);

OAI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1582),
.A2(n_1560),
.B1(n_1561),
.B2(n_1730),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1646),
.B(n_1425),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1544),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1615),
.B(n_1425),
.Y(n_1837)
);

OAI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1582),
.A2(n_1351),
.B(n_1419),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1615),
.B(n_1425),
.Y(n_1839)
);

AOI22xp5_ASAP7_75t_SL g1840 ( 
.A1(n_1598),
.A2(n_529),
.B1(n_543),
.B2(n_533),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1596),
.B(n_1427),
.Y(n_1841)
);

NAND3xp33_ASAP7_75t_SL g1842 ( 
.A(n_1570),
.B(n_1313),
.C(n_544),
.Y(n_1842)
);

AOI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1706),
.A2(n_1497),
.B1(n_1469),
.B2(n_1428),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_SL g1844 ( 
.A(n_1517),
.B(n_1426),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1516),
.B(n_738),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1596),
.B(n_1427),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1586),
.B(n_1561),
.Y(n_1847)
);

AOI21xp5_ASAP7_75t_L g1848 ( 
.A1(n_1599),
.A2(n_1356),
.B(n_1352),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1659),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1586),
.B(n_1427),
.Y(n_1850)
);

AND2x4_ASAP7_75t_L g1851 ( 
.A(n_1607),
.B(n_1264),
.Y(n_1851)
);

OAI21xp33_ASAP7_75t_L g1852 ( 
.A1(n_1570),
.A2(n_547),
.B(n_526),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1653),
.A2(n_1497),
.B1(n_690),
.B2(n_697),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_1660),
.Y(n_1854)
);

INVxp67_ASAP7_75t_L g1855 ( 
.A(n_1575),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1600),
.B(n_1271),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1544),
.Y(n_1857)
);

BUFx3_ASAP7_75t_L g1858 ( 
.A(n_1549),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1600),
.B(n_1604),
.Y(n_1859)
);

BUFx3_ASAP7_75t_L g1860 ( 
.A(n_1549),
.Y(n_1860)
);

BUFx3_ASAP7_75t_L g1861 ( 
.A(n_1549),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1592),
.B(n_1431),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1663),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1604),
.B(n_1271),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1667),
.Y(n_1865)
);

CKINVDCx5p33_ASAP7_75t_R g1866 ( 
.A(n_1719),
.Y(n_1866)
);

INVxp67_ASAP7_75t_L g1867 ( 
.A(n_1633),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1671),
.Y(n_1868)
);

BUFx6f_ASAP7_75t_L g1869 ( 
.A(n_1692),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1545),
.Y(n_1870)
);

NOR2xp33_ASAP7_75t_L g1871 ( 
.A(n_1593),
.B(n_1432),
.Y(n_1871)
);

INVxp67_ASAP7_75t_L g1872 ( 
.A(n_1601),
.Y(n_1872)
);

AOI22xp33_ASAP7_75t_L g1873 ( 
.A1(n_1653),
.A2(n_1657),
.B1(n_1694),
.B2(n_1742),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1593),
.B(n_1443),
.Y(n_1874)
);

INVx3_ASAP7_75t_L g1875 ( 
.A(n_1648),
.Y(n_1875)
);

NOR2x1_ASAP7_75t_L g1876 ( 
.A(n_1510),
.B(n_1490),
.Y(n_1876)
);

AOI22xp5_ASAP7_75t_L g1877 ( 
.A1(n_1647),
.A2(n_1469),
.B1(n_1485),
.B2(n_1484),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1545),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_SL g1879 ( 
.A(n_1517),
.B(n_1463),
.Y(n_1879)
);

OR2x2_ASAP7_75t_SL g1880 ( 
.A(n_1698),
.B(n_690),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1689),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1546),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_SL g1883 ( 
.A(n_1522),
.B(n_1299),
.Y(n_1883)
);

AOI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1651),
.A2(n_1664),
.B1(n_1734),
.B2(n_1729),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_1538),
.Y(n_1885)
);

BUFx2_ASAP7_75t_L g1886 ( 
.A(n_1740),
.Y(n_1886)
);

AOI22xp33_ASAP7_75t_L g1887 ( 
.A1(n_1657),
.A2(n_697),
.B1(n_702),
.B2(n_686),
.Y(n_1887)
);

AOI21xp5_ASAP7_75t_L g1888 ( 
.A1(n_1634),
.A2(n_1356),
.B(n_1352),
.Y(n_1888)
);

AND2x6_ASAP7_75t_L g1889 ( 
.A(n_1511),
.B(n_1271),
.Y(n_1889)
);

NOR2x1p5_ASAP7_75t_L g1890 ( 
.A(n_1678),
.B(n_549),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1546),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1522),
.B(n_1507),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1662),
.A2(n_1388),
.B(n_1363),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1556),
.B(n_1326),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1690),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1558),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1608),
.B(n_1705),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1608),
.B(n_1319),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1683),
.B(n_738),
.Y(n_1899)
);

OAI22xp5_ASAP7_75t_L g1900 ( 
.A1(n_1710),
.A2(n_1325),
.B1(n_1421),
.B2(n_1279),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1700),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1715),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1558),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1694),
.A2(n_702),
.B1(n_711),
.B2(n_686),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1723),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1699),
.B(n_1319),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1726),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1732),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1557),
.B(n_1319),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1573),
.B(n_1326),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1565),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_SL g1912 ( 
.A(n_1704),
.B(n_1264),
.Y(n_1912)
);

INVx2_ASAP7_75t_SL g1913 ( 
.A(n_1555),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_SL g1914 ( 
.A(n_1704),
.B(n_1264),
.Y(n_1914)
);

AOI22xp33_ASAP7_75t_L g1915 ( 
.A1(n_1742),
.A2(n_727),
.B1(n_731),
.B2(n_711),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1585),
.B(n_1326),
.Y(n_1916)
);

AND2x4_ASAP7_75t_SL g1917 ( 
.A(n_1607),
.B(n_1264),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1565),
.Y(n_1918)
);

INVx3_ASAP7_75t_L g1919 ( 
.A(n_1677),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1587),
.B(n_1393),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1737),
.Y(n_1921)
);

BUFx2_ASAP7_75t_L g1922 ( 
.A(n_1674),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1739),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_SL g1924 ( 
.A(n_1704),
.B(n_1299),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1746),
.Y(n_1925)
);

CKINVDCx5p33_ASAP7_75t_R g1926 ( 
.A(n_1574),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1591),
.B(n_1393),
.Y(n_1927)
);

CKINVDCx5p33_ASAP7_75t_R g1928 ( 
.A(n_1674),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1747),
.Y(n_1929)
);

INVx2_ASAP7_75t_SL g1930 ( 
.A(n_1610),
.Y(n_1930)
);

INVx5_ASAP7_75t_L g1931 ( 
.A(n_1677),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1571),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1530),
.B(n_1264),
.Y(n_1933)
);

AOI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1623),
.A2(n_1311),
.B1(n_1299),
.B2(n_635),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1571),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1594),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1606),
.B(n_1399),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1612),
.B(n_1399),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1613),
.B(n_1405),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1594),
.Y(n_1940)
);

NOR2xp33_ASAP7_75t_L g1941 ( 
.A(n_1619),
.B(n_1499),
.Y(n_1941)
);

NOR3xp33_ASAP7_75t_SL g1942 ( 
.A(n_1680),
.B(n_568),
.C(n_560),
.Y(n_1942)
);

INVx4_ASAP7_75t_L g1943 ( 
.A(n_1677),
.Y(n_1943)
);

NOR2x2_ASAP7_75t_L g1944 ( 
.A(n_1674),
.B(n_1602),
.Y(n_1944)
);

NAND2x1p5_ASAP7_75t_L g1945 ( 
.A(n_1566),
.B(n_1363),
.Y(n_1945)
);

AOI22xp5_ASAP7_75t_L g1946 ( 
.A1(n_1626),
.A2(n_1540),
.B1(n_1717),
.B2(n_1748),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1602),
.Y(n_1947)
);

INVx3_ASAP7_75t_L g1948 ( 
.A(n_1566),
.Y(n_1948)
);

BUFx3_ASAP7_75t_L g1949 ( 
.A(n_1578),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1638),
.Y(n_1950)
);

AOI22xp5_ASAP7_75t_L g1951 ( 
.A1(n_1717),
.A2(n_1311),
.B1(n_1299),
.B2(n_644),
.Y(n_1951)
);

INVx2_ASAP7_75t_SL g1952 ( 
.A(n_1610),
.Y(n_1952)
);

BUFx6f_ASAP7_75t_L g1953 ( 
.A(n_1578),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1638),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1641),
.Y(n_1955)
);

NOR2xp67_ASAP7_75t_L g1956 ( 
.A(n_1609),
.B(n_1405),
.Y(n_1956)
);

INVx2_ASAP7_75t_SL g1957 ( 
.A(n_1610),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1641),
.Y(n_1958)
);

NAND2xp33_ASAP7_75t_SL g1959 ( 
.A(n_1873),
.B(n_1735),
.Y(n_1959)
);

NAND2xp33_ASAP7_75t_SL g1960 ( 
.A(n_1873),
.B(n_1765),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_SL g1961 ( 
.A(n_1759),
.B(n_1718),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_SL g1962 ( 
.A(n_1767),
.B(n_1764),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_SL g1963 ( 
.A(n_1764),
.B(n_1513),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1886),
.B(n_1508),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1859),
.B(n_1525),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_SL g1966 ( 
.A(n_1755),
.B(n_1528),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_SL g1967 ( 
.A(n_1755),
.B(n_1541),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_SL g1968 ( 
.A(n_1867),
.B(n_1543),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1899),
.B(n_1535),
.Y(n_1969)
);

NAND2xp33_ASAP7_75t_SL g1970 ( 
.A(n_1765),
.B(n_1611),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_SL g1971 ( 
.A(n_1818),
.B(n_1536),
.Y(n_1971)
);

AND2x4_ASAP7_75t_L g1972 ( 
.A(n_1943),
.B(n_1785),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_SL g1973 ( 
.A(n_1766),
.B(n_1748),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_SL g1974 ( 
.A(n_1855),
.B(n_1551),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_SL g1975 ( 
.A(n_1787),
.B(n_1551),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_SL g1976 ( 
.A(n_1789),
.B(n_1595),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_SL g1977 ( 
.A(n_1872),
.B(n_1595),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_SL g1978 ( 
.A(n_1769),
.B(n_1518),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_SL g1979 ( 
.A(n_1760),
.B(n_1702),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_SL g1980 ( 
.A(n_1760),
.B(n_1704),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_SL g1981 ( 
.A(n_1795),
.B(n_1704),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_SL g1982 ( 
.A(n_1821),
.B(n_1704),
.Y(n_1982)
);

NAND2xp33_ASAP7_75t_SL g1983 ( 
.A(n_1847),
.B(n_1611),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_SL g1984 ( 
.A(n_1823),
.B(n_1741),
.Y(n_1984)
);

NAND2xp33_ASAP7_75t_SL g1985 ( 
.A(n_1943),
.B(n_1627),
.Y(n_1985)
);

AND2x4_ASAP7_75t_L g1986 ( 
.A(n_1785),
.B(n_1514),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_SL g1987 ( 
.A(n_1897),
.B(n_1741),
.Y(n_1987)
);

NAND2xp33_ASAP7_75t_SL g1988 ( 
.A(n_1777),
.B(n_1885),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_SL g1989 ( 
.A(n_1770),
.B(n_1527),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_SL g1990 ( 
.A(n_1770),
.B(n_1650),
.Y(n_1990)
);

NAND2xp33_ASAP7_75t_SL g1991 ( 
.A(n_1777),
.B(n_1684),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1871),
.B(n_1708),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_SL g1993 ( 
.A(n_1942),
.B(n_1834),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1854),
.B(n_1668),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_SL g1995 ( 
.A(n_1884),
.B(n_1669),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1871),
.B(n_1589),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_SL g1997 ( 
.A(n_1794),
.B(n_1672),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_SL g1998 ( 
.A(n_1794),
.B(n_1685),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_SL g1999 ( 
.A(n_1797),
.B(n_1695),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1874),
.B(n_1531),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_SL g2001 ( 
.A(n_1797),
.B(n_1712),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1874),
.B(n_1534),
.Y(n_2002)
);

NAND2xp33_ASAP7_75t_SL g2003 ( 
.A(n_1890),
.B(n_1731),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_SL g2004 ( 
.A(n_1845),
.B(n_1621),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1894),
.B(n_1537),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_SL g2006 ( 
.A(n_1750),
.B(n_1625),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_SL g2007 ( 
.A(n_1946),
.B(n_1514),
.Y(n_2007)
);

AND2x4_ASAP7_75t_L g2008 ( 
.A(n_1785),
.B(n_1639),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_SL g2009 ( 
.A(n_1862),
.B(n_1547),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_SL g2010 ( 
.A(n_1956),
.B(n_1548),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1894),
.B(n_1553),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_SL g2012 ( 
.A(n_1831),
.B(n_1559),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_SL g2013 ( 
.A(n_1802),
.B(n_1562),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_SL g2014 ( 
.A(n_1802),
.B(n_1564),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1941),
.B(n_1568),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_SL g2016 ( 
.A(n_1830),
.B(n_1569),
.Y(n_2016)
);

NAND2xp33_ASAP7_75t_SL g2017 ( 
.A(n_1866),
.B(n_1731),
.Y(n_2017)
);

NAND2xp33_ASAP7_75t_SL g2018 ( 
.A(n_1913),
.B(n_1627),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1840),
.B(n_851),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_SL g2020 ( 
.A(n_1830),
.B(n_1579),
.Y(n_2020)
);

NAND2xp33_ASAP7_75t_SL g2021 ( 
.A(n_1883),
.B(n_1635),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_SL g2022 ( 
.A(n_1953),
.B(n_1580),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_SL g2023 ( 
.A(n_1953),
.B(n_1761),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1941),
.B(n_1581),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_SL g2025 ( 
.A(n_1953),
.B(n_1583),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1906),
.B(n_1584),
.Y(n_2026)
);

NAND2xp33_ASAP7_75t_SL g2027 ( 
.A(n_1883),
.B(n_1635),
.Y(n_2027)
);

NAND2xp33_ASAP7_75t_SL g2028 ( 
.A(n_1786),
.B(n_1728),
.Y(n_2028)
);

NAND2xp33_ASAP7_75t_SL g2029 ( 
.A(n_1853),
.B(n_1616),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_SL g2030 ( 
.A(n_1953),
.B(n_1588),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_SL g2031 ( 
.A(n_1805),
.B(n_1299),
.Y(n_2031)
);

NAND2xp33_ASAP7_75t_SL g2032 ( 
.A(n_1853),
.B(n_1363),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1809),
.B(n_1597),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_SL g2034 ( 
.A(n_1815),
.B(n_1311),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_SL g2035 ( 
.A(n_1827),
.B(n_1311),
.Y(n_2035)
);

NAND2xp33_ASAP7_75t_SL g2036 ( 
.A(n_1875),
.B(n_1388),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_SL g2037 ( 
.A(n_1832),
.B(n_1311),
.Y(n_2037)
);

NAND2xp33_ASAP7_75t_SL g2038 ( 
.A(n_1875),
.B(n_1388),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1849),
.B(n_1707),
.Y(n_2039)
);

NAND2xp33_ASAP7_75t_SL g2040 ( 
.A(n_1919),
.B(n_1392),
.Y(n_2040)
);

NAND2xp33_ASAP7_75t_SL g2041 ( 
.A(n_1919),
.B(n_1392),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_SL g2042 ( 
.A(n_1863),
.B(n_1644),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_SL g2043 ( 
.A(n_1865),
.B(n_1703),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_SL g2044 ( 
.A(n_1868),
.B(n_1515),
.Y(n_2044)
);

NAND2xp33_ASAP7_75t_SL g2045 ( 
.A(n_1778),
.B(n_1392),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_SL g2046 ( 
.A(n_1881),
.B(n_1670),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_SL g2047 ( 
.A(n_1895),
.B(n_1617),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_1901),
.B(n_1622),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1902),
.B(n_1905),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_SL g2050 ( 
.A(n_1907),
.B(n_1725),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1908),
.B(n_1661),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_SL g2052 ( 
.A(n_1921),
.B(n_1733),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1923),
.B(n_1661),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_SL g2054 ( 
.A(n_1925),
.B(n_1929),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_SL g2055 ( 
.A(n_1949),
.B(n_1738),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_SL g2056 ( 
.A(n_1949),
.B(n_1744),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_SL g2057 ( 
.A(n_1851),
.B(n_1745),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_SL g2058 ( 
.A(n_1851),
.B(n_1749),
.Y(n_2058)
);

NAND2xp33_ASAP7_75t_SL g2059 ( 
.A(n_1778),
.B(n_1414),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_SL g2060 ( 
.A(n_1948),
.B(n_1628),
.Y(n_2060)
);

NAND2xp33_ASAP7_75t_SL g2061 ( 
.A(n_1778),
.B(n_1414),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_SL g2062 ( 
.A(n_1948),
.B(n_1858),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_SL g2063 ( 
.A(n_1858),
.B(n_1860),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_1930),
.B(n_853),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_SL g2065 ( 
.A(n_1860),
.B(n_1643),
.Y(n_2065)
);

NAND2xp33_ASAP7_75t_SL g2066 ( 
.A(n_1778),
.B(n_1414),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_SL g2067 ( 
.A(n_1861),
.B(n_1630),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_SL g2068 ( 
.A(n_1861),
.B(n_1727),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_SL g2069 ( 
.A(n_1852),
.B(n_1711),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_SL g2070 ( 
.A(n_1933),
.B(n_1713),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_SL g2071 ( 
.A(n_1933),
.B(n_1430),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_SL g2072 ( 
.A(n_1785),
.B(n_1931),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1822),
.B(n_1952),
.Y(n_2073)
);

NAND2xp33_ASAP7_75t_SL g2074 ( 
.A(n_1869),
.B(n_1430),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_SL g2075 ( 
.A(n_1931),
.B(n_1430),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1957),
.B(n_1665),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_SL g2077 ( 
.A(n_1931),
.B(n_1442),
.Y(n_2077)
);

NAND2xp33_ASAP7_75t_SL g2078 ( 
.A(n_1869),
.B(n_1442),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1833),
.B(n_1665),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1835),
.B(n_1506),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1887),
.B(n_1506),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_SL g2082 ( 
.A(n_1931),
.B(n_1442),
.Y(n_2082)
);

AND2x4_ASAP7_75t_L g2083 ( 
.A(n_1801),
.B(n_1922),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_SL g2084 ( 
.A(n_1782),
.B(n_1470),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_SL g2085 ( 
.A(n_1782),
.B(n_1470),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_SL g2086 ( 
.A(n_1843),
.B(n_1470),
.Y(n_2086)
);

OR2x2_ASAP7_75t_L g2087 ( 
.A(n_1880),
.B(n_1640),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_SL g2088 ( 
.A(n_1751),
.B(n_1471),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_SL g2089 ( 
.A(n_1753),
.B(n_1754),
.Y(n_2089)
);

NAND2xp33_ASAP7_75t_SL g2090 ( 
.A(n_1928),
.B(n_1605),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_1801),
.B(n_853),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1887),
.B(n_1407),
.Y(n_2092)
);

NAND2xp33_ASAP7_75t_SL g2093 ( 
.A(n_1926),
.B(n_1642),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_SL g2094 ( 
.A(n_1756),
.B(n_1471),
.Y(n_2094)
);

NAND2xp33_ASAP7_75t_SL g2095 ( 
.A(n_1869),
.B(n_1656),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_SL g2096 ( 
.A(n_1757),
.B(n_1471),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_SL g2097 ( 
.A(n_1758),
.B(n_1490),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_SL g2098 ( 
.A(n_1768),
.B(n_1490),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_SL g2099 ( 
.A(n_1771),
.B(n_1491),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_SL g2100 ( 
.A(n_1773),
.B(n_1491),
.Y(n_2100)
);

NAND2xp33_ASAP7_75t_SL g2101 ( 
.A(n_1869),
.B(n_1491),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_SL g2102 ( 
.A(n_1784),
.B(n_1554),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_SL g2103 ( 
.A(n_1790),
.B(n_1673),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_SL g2104 ( 
.A(n_1792),
.B(n_1688),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_SL g2105 ( 
.A(n_1793),
.B(n_1631),
.Y(n_2105)
);

NAND2xp33_ASAP7_75t_SL g2106 ( 
.A(n_1904),
.B(n_1716),
.Y(n_2106)
);

NAND2xp33_ASAP7_75t_SL g2107 ( 
.A(n_1904),
.B(n_1261),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_1841),
.B(n_1407),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1846),
.B(n_1420),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_SL g2110 ( 
.A(n_1763),
.B(n_1420),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_SL g2111 ( 
.A(n_1763),
.B(n_1780),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_SL g2112 ( 
.A(n_1780),
.B(n_1781),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_SL g2113 ( 
.A(n_1781),
.B(n_1422),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_SL g2114 ( 
.A(n_1791),
.B(n_1422),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_SL g2115 ( 
.A(n_1791),
.B(n_1434),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_SL g2116 ( 
.A(n_1799),
.B(n_1800),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_SL g2117 ( 
.A(n_1799),
.B(n_1434),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_SL g2118 ( 
.A(n_1800),
.B(n_1436),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_SL g2119 ( 
.A(n_1803),
.B(n_1436),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_SL g2120 ( 
.A(n_1803),
.B(n_1438),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_SL g2121 ( 
.A(n_1838),
.B(n_1438),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_SL g2122 ( 
.A(n_1811),
.B(n_1439),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_SL g2123 ( 
.A(n_1811),
.B(n_1439),
.Y(n_2123)
);

NAND2xp33_ASAP7_75t_SL g2124 ( 
.A(n_1779),
.B(n_1261),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_SL g2125 ( 
.A(n_1752),
.B(n_1440),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_SL g2126 ( 
.A(n_1752),
.B(n_1440),
.Y(n_2126)
);

NOR2xp33_ASAP7_75t_L g2127 ( 
.A(n_1842),
.B(n_1441),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_SL g2128 ( 
.A(n_1876),
.B(n_1441),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_1856),
.B(n_1444),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_SL g2130 ( 
.A(n_1951),
.B(n_1444),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1864),
.B(n_1451),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1814),
.B(n_1451),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_SL g2133 ( 
.A(n_1920),
.B(n_1452),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_SL g2134 ( 
.A(n_1927),
.B(n_1452),
.Y(n_2134)
);

NAND2xp33_ASAP7_75t_SL g2135 ( 
.A(n_1779),
.B(n_1265),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_1801),
.B(n_855),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_SL g2137 ( 
.A(n_1937),
.B(n_1453),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_SL g2138 ( 
.A(n_1938),
.B(n_1453),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_1816),
.B(n_1455),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_SL g2140 ( 
.A(n_1939),
.B(n_1455),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_SL g2141 ( 
.A(n_1934),
.B(n_1458),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_SL g2142 ( 
.A(n_1917),
.B(n_1458),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_1915),
.B(n_855),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_SL g2144 ( 
.A(n_1917),
.B(n_1466),
.Y(n_2144)
);

NAND2xp33_ASAP7_75t_SL g2145 ( 
.A(n_1850),
.B(n_1724),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_SL g2146 ( 
.A(n_1804),
.B(n_1466),
.Y(n_2146)
);

NAND2xp33_ASAP7_75t_SL g2147 ( 
.A(n_1837),
.B(n_1265),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1817),
.B(n_1478),
.Y(n_2148)
);

AND2x4_ASAP7_75t_L g2149 ( 
.A(n_1776),
.B(n_1450),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_SL g2150 ( 
.A(n_1804),
.B(n_1478),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_SL g2151 ( 
.A(n_1958),
.B(n_1501),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_SL g2152 ( 
.A(n_1958),
.B(n_1808),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_SL g2153 ( 
.A(n_1808),
.B(n_1501),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_SL g2154 ( 
.A(n_1955),
.B(n_1682),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_SL g2155 ( 
.A(n_1955),
.B(n_1590),
.Y(n_2155)
);

NAND2xp33_ASAP7_75t_SL g2156 ( 
.A(n_1839),
.B(n_1483),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_SL g2157 ( 
.A(n_1954),
.B(n_1576),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_SL g2158 ( 
.A(n_1954),
.B(n_627),
.Y(n_2158)
);

NAND2xp33_ASAP7_75t_SL g2159 ( 
.A(n_1898),
.B(n_1483),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_1819),
.B(n_1489),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1813),
.B(n_1360),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_SL g2162 ( 
.A(n_1813),
.B(n_645),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_1915),
.B(n_858),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_SL g2164 ( 
.A(n_1824),
.B(n_648),
.Y(n_2164)
);

NAND2xp33_ASAP7_75t_SL g2165 ( 
.A(n_1798),
.B(n_1447),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_SL g2166 ( 
.A(n_1824),
.B(n_654),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_SL g2167 ( 
.A(n_1836),
.B(n_661),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_1950),
.B(n_858),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_SL g2169 ( 
.A(n_1836),
.B(n_674),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_1857),
.B(n_1377),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_SL g2171 ( 
.A(n_1857),
.B(n_682),
.Y(n_2171)
);

NAND2xp33_ASAP7_75t_SL g2172 ( 
.A(n_1798),
.B(n_1457),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_SL g2173 ( 
.A(n_1870),
.B(n_684),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_1870),
.B(n_1552),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_SL g2175 ( 
.A(n_1878),
.B(n_1882),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_SL g2176 ( 
.A(n_1878),
.B(n_685),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_SL g2177 ( 
.A(n_1882),
.B(n_687),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_1891),
.B(n_1675),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_SL g2179 ( 
.A(n_1891),
.B(n_698),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_1896),
.B(n_1502),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_SL g2181 ( 
.A(n_1896),
.B(n_710),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_SL g2182 ( 
.A(n_1903),
.B(n_720),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_SL g2183 ( 
.A(n_1903),
.B(n_722),
.Y(n_2183)
);

NAND2xp33_ASAP7_75t_SL g2184 ( 
.A(n_1826),
.B(n_1892),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_SL g2185 ( 
.A(n_1911),
.B(n_732),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_SL g2186 ( 
.A(n_1911),
.B(n_748),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_SL g2187 ( 
.A(n_1918),
.B(n_760),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_SL g2188 ( 
.A(n_1918),
.B(n_573),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_SL g2189 ( 
.A(n_1935),
.B(n_574),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_SL g2190 ( 
.A(n_1935),
.B(n_581),
.Y(n_2190)
);

CKINVDCx20_ASAP7_75t_R g2191 ( 
.A(n_1988),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1962),
.B(n_1774),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_SL g2193 ( 
.A(n_2000),
.B(n_1892),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_2152),
.Y(n_2194)
);

AND2x2_ASAP7_75t_L g2195 ( 
.A(n_2019),
.B(n_1810),
.Y(n_2195)
);

HB1xp67_ASAP7_75t_L g2196 ( 
.A(n_1964),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2049),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_1965),
.B(n_1936),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_1996),
.B(n_1936),
.Y(n_2199)
);

AOI22xp5_ASAP7_75t_L g2200 ( 
.A1(n_2003),
.A2(n_1829),
.B1(n_1775),
.B2(n_1772),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_2175),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_2111),
.Y(n_2202)
);

INVxp33_ASAP7_75t_SL g2203 ( 
.A(n_1969),
.Y(n_2203)
);

AND3x1_ASAP7_75t_SL g2204 ( 
.A(n_1993),
.B(n_731),
.C(n_727),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2002),
.B(n_1963),
.Y(n_2205)
);

AND2x4_ASAP7_75t_L g2206 ( 
.A(n_2083),
.B(n_1776),
.Y(n_2206)
);

INVxp67_ASAP7_75t_L g2207 ( 
.A(n_2091),
.Y(n_2207)
);

AOI22xp33_ASAP7_75t_L g2208 ( 
.A1(n_1960),
.A2(n_753),
.B1(n_759),
.B2(n_750),
.Y(n_2208)
);

AND2x4_ASAP7_75t_L g2209 ( 
.A(n_2083),
.B(n_1783),
.Y(n_2209)
);

OR2x6_ASAP7_75t_L g2210 ( 
.A(n_2083),
.B(n_1829),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2009),
.B(n_1932),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2015),
.B(n_1940),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_2024),
.B(n_1987),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_1961),
.B(n_1947),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2136),
.B(n_861),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2064),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_2168),
.B(n_861),
.Y(n_2217)
);

INVxp67_ASAP7_75t_L g2218 ( 
.A(n_1973),
.Y(n_2218)
);

OAI21xp5_ASAP7_75t_L g2219 ( 
.A1(n_2012),
.A2(n_1877),
.B(n_1844),
.Y(n_2219)
);

AND3x1_ASAP7_75t_SL g2220 ( 
.A(n_1960),
.B(n_753),
.C(n_750),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_2112),
.Y(n_2221)
);

INVxp67_ASAP7_75t_L g2222 ( 
.A(n_1975),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_2116),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_1992),
.B(n_1909),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_2087),
.B(n_862),
.Y(n_2225)
);

INVxp67_ASAP7_75t_L g2226 ( 
.A(n_1976),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2054),
.Y(n_2227)
);

AOI22xp33_ASAP7_75t_L g2228 ( 
.A1(n_2029),
.A2(n_761),
.B1(n_759),
.B2(n_1844),
.Y(n_2228)
);

AND2x2_ASAP7_75t_SL g2229 ( 
.A(n_2143),
.B(n_1944),
.Y(n_2229)
);

AND3x1_ASAP7_75t_SL g2230 ( 
.A(n_1984),
.B(n_761),
.C(n_862),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2073),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_2174),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2089),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2051),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2039),
.B(n_1910),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2033),
.B(n_1916),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_1978),
.B(n_1783),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2163),
.B(n_1971),
.Y(n_2238)
);

BUFx12f_ASAP7_75t_L g2239 ( 
.A(n_2008),
.Y(n_2239)
);

NOR2xp33_ASAP7_75t_R g2240 ( 
.A(n_2017),
.B(n_1828),
.Y(n_2240)
);

AND2x4_ASAP7_75t_L g2241 ( 
.A(n_1972),
.B(n_1788),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_SL g2242 ( 
.A(n_1959),
.B(n_1900),
.Y(n_2242)
);

BUFx6f_ASAP7_75t_L g2243 ( 
.A(n_1972),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_SL g2244 ( 
.A(n_1959),
.B(n_1828),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2053),
.Y(n_2245)
);

AND2x2_ASAP7_75t_L g2246 ( 
.A(n_1974),
.B(n_863),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_2178),
.Y(n_2247)
);

NAND2x1p5_ASAP7_75t_L g2248 ( 
.A(n_1972),
.B(n_1826),
.Y(n_2248)
);

BUFx6f_ASAP7_75t_L g2249 ( 
.A(n_2072),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_1966),
.B(n_863),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2076),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_2004),
.B(n_1788),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_SL g2253 ( 
.A(n_2005),
.B(n_1848),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_1967),
.B(n_864),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_1977),
.B(n_1807),
.Y(n_2255)
);

NAND2xp33_ASAP7_75t_L g2256 ( 
.A(n_2032),
.B(n_1812),
.Y(n_2256)
);

AOI22xp5_ASAP7_75t_L g2257 ( 
.A1(n_2093),
.A2(n_2090),
.B1(n_2029),
.B2(n_2018),
.Y(n_2257)
);

AND3x1_ASAP7_75t_SL g2258 ( 
.A(n_1991),
.B(n_865),
.C(n_864),
.Y(n_2258)
);

AOI22xp33_ASAP7_75t_L g2259 ( 
.A1(n_2106),
.A2(n_1879),
.B1(n_583),
.B2(n_587),
.Y(n_2259)
);

CKINVDCx5p33_ASAP7_75t_R g2260 ( 
.A(n_1994),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2047),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_2146),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2048),
.Y(n_2263)
);

INVx1_ASAP7_75t_SL g2264 ( 
.A(n_2063),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2080),
.B(n_1807),
.Y(n_2265)
);

BUFx6f_ASAP7_75t_L g2266 ( 
.A(n_2008),
.Y(n_2266)
);

AOI22xp5_ASAP7_75t_L g2267 ( 
.A1(n_1979),
.A2(n_1879),
.B1(n_1796),
.B2(n_1812),
.Y(n_2267)
);

AND2x2_ASAP7_75t_L g2268 ( 
.A(n_1968),
.B(n_865),
.Y(n_2268)
);

OR2x2_ASAP7_75t_L g2269 ( 
.A(n_2188),
.B(n_1806),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_2150),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2110),
.Y(n_2271)
);

INVx5_ASAP7_75t_L g2272 ( 
.A(n_1986),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_2189),
.B(n_870),
.Y(n_2273)
);

AOI21xp5_ASAP7_75t_L g2274 ( 
.A1(n_2032),
.A2(n_1893),
.B(n_1888),
.Y(n_2274)
);

AOI22xp33_ASAP7_75t_L g2275 ( 
.A1(n_1970),
.A2(n_589),
.B1(n_592),
.B2(n_582),
.Y(n_2275)
);

INVx3_ASAP7_75t_L g2276 ( 
.A(n_2149),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2113),
.Y(n_2277)
);

INVx1_ASAP7_75t_SL g2278 ( 
.A(n_2062),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_2011),
.B(n_1820),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2114),
.Y(n_2280)
);

INVx5_ASAP7_75t_L g2281 ( 
.A(n_1986),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_2151),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2013),
.B(n_1820),
.Y(n_2283)
);

BUFx6f_ASAP7_75t_L g2284 ( 
.A(n_2008),
.Y(n_2284)
);

HB1xp67_ASAP7_75t_L g2285 ( 
.A(n_2014),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2153),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_SL g2287 ( 
.A(n_2127),
.B(n_1796),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2115),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_2016),
.B(n_1825),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_2020),
.B(n_1825),
.Y(n_2290)
);

OAI22xp5_ASAP7_75t_SL g2291 ( 
.A1(n_2081),
.A2(n_596),
.B1(n_597),
.B2(n_594),
.Y(n_2291)
);

CKINVDCx16_ASAP7_75t_R g2292 ( 
.A(n_2149),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_SL g2293 ( 
.A(n_2007),
.B(n_1945),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_SL g2294 ( 
.A(n_1983),
.B(n_1995),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2117),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2026),
.B(n_1812),
.Y(n_2296)
);

INVx4_ASAP7_75t_L g2297 ( 
.A(n_2149),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2118),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_1989),
.B(n_2079),
.Y(n_2299)
);

AND2x2_ASAP7_75t_L g2300 ( 
.A(n_2190),
.B(n_870),
.Y(n_2300)
);

INVx3_ASAP7_75t_L g2301 ( 
.A(n_1986),
.Y(n_2301)
);

NOR2xp33_ASAP7_75t_L g2302 ( 
.A(n_2006),
.B(n_1912),
.Y(n_2302)
);

AND2x4_ASAP7_75t_L g2303 ( 
.A(n_1980),
.B(n_1912),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2050),
.B(n_1812),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_2119),
.Y(n_2305)
);

AND2x4_ASAP7_75t_L g2306 ( 
.A(n_1990),
.B(n_2057),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2120),
.Y(n_2307)
);

BUFx6f_ASAP7_75t_L g2308 ( 
.A(n_1997),
.Y(n_2308)
);

AND2x2_ASAP7_75t_L g2309 ( 
.A(n_2125),
.B(n_871),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2180),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_2126),
.B(n_871),
.Y(n_2311)
);

AND2x2_ASAP7_75t_L g2312 ( 
.A(n_2001),
.B(n_1998),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_1999),
.B(n_872),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2052),
.B(n_1812),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2043),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2042),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2105),
.Y(n_2317)
);

NOR2xp33_ASAP7_75t_L g2318 ( 
.A(n_2070),
.B(n_1914),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2133),
.Y(n_2319)
);

NOR2xp33_ASAP7_75t_R g2320 ( 
.A(n_1970),
.B(n_1889),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2160),
.B(n_601),
.Y(n_2321)
);

INVx1_ASAP7_75t_SL g2322 ( 
.A(n_1981),
.Y(n_2322)
);

OAI22xp5_ASAP7_75t_SL g2323 ( 
.A1(n_2092),
.A2(n_614),
.B1(n_619),
.B2(n_603),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2023),
.B(n_621),
.Y(n_2324)
);

OAI21xp5_ASAP7_75t_L g2325 ( 
.A1(n_2010),
.A2(n_1681),
.B(n_1762),
.Y(n_2325)
);

INVx5_ASAP7_75t_L g2326 ( 
.A(n_2045),
.Y(n_2326)
);

BUFx2_ASAP7_75t_L g2327 ( 
.A(n_2095),
.Y(n_2327)
);

BUFx8_ASAP7_75t_L g2328 ( 
.A(n_1985),
.Y(n_2328)
);

INVx1_ASAP7_75t_SL g2329 ( 
.A(n_2055),
.Y(n_2329)
);

INVx1_ASAP7_75t_SL g2330 ( 
.A(n_2056),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_2157),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_2154),
.Y(n_2332)
);

HB1xp67_ASAP7_75t_L g2333 ( 
.A(n_2022),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2155),
.Y(n_2334)
);

NOR2xp33_ASAP7_75t_R g2335 ( 
.A(n_1983),
.B(n_1889),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_2058),
.B(n_622),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2158),
.B(n_623),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2187),
.B(n_624),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2162),
.B(n_872),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2134),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2102),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2186),
.B(n_625),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_2164),
.B(n_874),
.Y(n_2343)
);

OAI21xp5_ASAP7_75t_L g2344 ( 
.A1(n_2069),
.A2(n_1924),
.B(n_1914),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_2137),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_SL g2346 ( 
.A(n_2184),
.B(n_1945),
.Y(n_2346)
);

NOR2xp33_ASAP7_75t_L g2347 ( 
.A(n_2046),
.B(n_1924),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_2138),
.Y(n_2348)
);

OAI22xp5_ASAP7_75t_L g2349 ( 
.A1(n_2084),
.A2(n_630),
.B1(n_631),
.B2(n_628),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_2140),
.Y(n_2350)
);

AND2x4_ASAP7_75t_L g2351 ( 
.A(n_2071),
.B(n_1889),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2025),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2104),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2166),
.B(n_633),
.Y(n_2354)
);

CKINVDCx20_ASAP7_75t_R g2355 ( 
.A(n_2167),
.Y(n_2355)
);

OAI22xp5_ASAP7_75t_SL g2356 ( 
.A1(n_2132),
.A2(n_640),
.B1(n_641),
.B2(n_634),
.Y(n_2356)
);

CKINVDCx5p33_ASAP7_75t_R g2357 ( 
.A(n_2169),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2171),
.B(n_2173),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_2103),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2030),
.Y(n_2360)
);

AOI22xp33_ASAP7_75t_L g2361 ( 
.A1(n_2184),
.A2(n_2028),
.B1(n_2021),
.B2(n_2027),
.Y(n_2361)
);

AOI22xp33_ASAP7_75t_L g2362 ( 
.A1(n_2028),
.A2(n_643),
.B1(n_649),
.B2(n_642),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_2176),
.B(n_651),
.Y(n_2363)
);

AOI22xp33_ASAP7_75t_L g2364 ( 
.A1(n_2021),
.A2(n_653),
.B1(n_655),
.B2(n_652),
.Y(n_2364)
);

AND3x1_ASAP7_75t_SL g2365 ( 
.A(n_2027),
.B(n_875),
.C(n_874),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2031),
.Y(n_2366)
);

NOR2xp33_ASAP7_75t_R g2367 ( 
.A(n_1985),
.B(n_1889),
.Y(n_2367)
);

NAND2x1p5_ASAP7_75t_L g2368 ( 
.A(n_2075),
.B(n_1146),
.Y(n_2368)
);

CKINVDCx5p33_ASAP7_75t_R g2369 ( 
.A(n_2177),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2108),
.Y(n_2370)
);

OAI21xp5_ASAP7_75t_L g2371 ( 
.A1(n_2044),
.A2(n_1889),
.B(n_1504),
.Y(n_2371)
);

AND2x4_ASAP7_75t_L g2372 ( 
.A(n_2068),
.B(n_300),
.Y(n_2372)
);

HB1xp67_ASAP7_75t_L g2373 ( 
.A(n_2065),
.Y(n_2373)
);

BUFx6f_ASAP7_75t_L g2374 ( 
.A(n_2077),
.Y(n_2374)
);

AOI22xp5_ASAP7_75t_L g2375 ( 
.A1(n_1982),
.A2(n_657),
.B1(n_658),
.B2(n_656),
.Y(n_2375)
);

INVx2_ASAP7_75t_L g2376 ( 
.A(n_2109),
.Y(n_2376)
);

AND2x2_ASAP7_75t_L g2377 ( 
.A(n_2179),
.B(n_875),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2185),
.B(n_877),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2129),
.Y(n_2379)
);

CKINVDCx20_ASAP7_75t_R g2380 ( 
.A(n_2181),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_SL g2381 ( 
.A(n_2086),
.B(n_877),
.Y(n_2381)
);

AO22x1_ASAP7_75t_L g2382 ( 
.A1(n_2161),
.A2(n_666),
.B1(n_671),
.B2(n_660),
.Y(n_2382)
);

AND2x2_ASAP7_75t_L g2383 ( 
.A(n_2182),
.B(n_879),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2183),
.B(n_677),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2034),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2035),
.Y(n_2386)
);

AND2x2_ASAP7_75t_L g2387 ( 
.A(n_2067),
.B(n_879),
.Y(n_2387)
);

AND2x2_ASAP7_75t_L g2388 ( 
.A(n_2170),
.B(n_880),
.Y(n_2388)
);

AOI22xp33_ASAP7_75t_L g2389 ( 
.A1(n_2165),
.A2(n_688),
.B1(n_691),
.B2(n_681),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2037),
.Y(n_2390)
);

OAI22xp5_ASAP7_75t_L g2391 ( 
.A1(n_2085),
.A2(n_694),
.B1(n_696),
.B2(n_692),
.Y(n_2391)
);

AND2x2_ASAP7_75t_L g2392 ( 
.A(n_2060),
.B(n_880),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_2122),
.B(n_881),
.Y(n_2393)
);

AND2x2_ASAP7_75t_L g2394 ( 
.A(n_2123),
.B(n_881),
.Y(n_2394)
);

CKINVDCx5p33_ASAP7_75t_R g2395 ( 
.A(n_2045),
.Y(n_2395)
);

NOR2xp67_ASAP7_75t_L g2396 ( 
.A(n_2088),
.B(n_306),
.Y(n_2396)
);

INVx3_ASAP7_75t_L g2397 ( 
.A(n_2139),
.Y(n_2397)
);

BUFx6f_ASAP7_75t_L g2398 ( 
.A(n_2082),
.Y(n_2398)
);

CKINVDCx5p33_ASAP7_75t_R g2399 ( 
.A(n_2059),
.Y(n_2399)
);

CKINVDCx16_ASAP7_75t_R g2400 ( 
.A(n_2059),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_L g2401 ( 
.A(n_2148),
.B(n_699),
.Y(n_2401)
);

CKINVDCx5p33_ASAP7_75t_R g2402 ( 
.A(n_2061),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2131),
.B(n_700),
.Y(n_2403)
);

AOI22xp33_ASAP7_75t_L g2404 ( 
.A1(n_2165),
.A2(n_704),
.B1(n_706),
.B2(n_703),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_2121),
.B(n_707),
.Y(n_2405)
);

NOR2xp33_ASAP7_75t_L g2406 ( 
.A(n_2130),
.B(n_708),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2128),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2141),
.B(n_712),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_2142),
.B(n_713),
.Y(n_2409)
);

INVx1_ASAP7_75t_SL g2410 ( 
.A(n_2144),
.Y(n_2410)
);

AND2x2_ASAP7_75t_L g2411 ( 
.A(n_2094),
.B(n_883),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2096),
.B(n_715),
.Y(n_2412)
);

HB1xp67_ASAP7_75t_L g2413 ( 
.A(n_2097),
.Y(n_2413)
);

AOI22xp33_ASAP7_75t_L g2414 ( 
.A1(n_2172),
.A2(n_718),
.B1(n_719),
.B2(n_717),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_SL g2415 ( 
.A(n_2145),
.B(n_883),
.Y(n_2415)
);

BUFx3_ASAP7_75t_L g2416 ( 
.A(n_2061),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2098),
.B(n_721),
.Y(n_2417)
);

AND2x2_ASAP7_75t_L g2418 ( 
.A(n_2099),
.B(n_887),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_2100),
.Y(n_2419)
);

AOI22xp5_ASAP7_75t_L g2420 ( 
.A1(n_2172),
.A2(n_725),
.B1(n_726),
.B2(n_723),
.Y(n_2420)
);

AOI22xp33_ASAP7_75t_L g2421 ( 
.A1(n_2107),
.A2(n_733),
.B1(n_734),
.B2(n_729),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2066),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2066),
.Y(n_2423)
);

AOI22xp5_ASAP7_75t_L g2424 ( 
.A1(n_2145),
.A2(n_740),
.B1(n_743),
.B2(n_737),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2074),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2156),
.B(n_744),
.Y(n_2426)
);

NOR2x1_ASAP7_75t_L g2427 ( 
.A(n_2074),
.B(n_887),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2078),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_2156),
.B(n_745),
.Y(n_2429)
);

CKINVDCx5p33_ASAP7_75t_R g2430 ( 
.A(n_2078),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2159),
.B(n_746),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2101),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2159),
.B(n_747),
.Y(n_2433)
);

NOR2xp67_ASAP7_75t_L g2434 ( 
.A(n_2036),
.B(n_307),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_2147),
.B(n_751),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2147),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2124),
.B(n_752),
.Y(n_2437)
);

AND2x6_ASAP7_75t_L g2438 ( 
.A(n_2036),
.B(n_1146),
.Y(n_2438)
);

CKINVDCx12_ASAP7_75t_R g2439 ( 
.A(n_2038),
.Y(n_2439)
);

OR2x2_ASAP7_75t_L g2440 ( 
.A(n_2135),
.B(n_888),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2038),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2040),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2040),
.B(n_754),
.Y(n_2443)
);

AND2x2_ASAP7_75t_L g2444 ( 
.A(n_2041),
.B(n_888),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2041),
.B(n_756),
.Y(n_2445)
);

BUFx2_ASAP7_75t_L g2446 ( 
.A(n_2083),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2049),
.Y(n_2447)
);

BUFx3_ASAP7_75t_L g2448 ( 
.A(n_2083),
.Y(n_2448)
);

AND2x2_ASAP7_75t_L g2449 ( 
.A(n_1962),
.B(n_891),
.Y(n_2449)
);

AND2x2_ASAP7_75t_L g2450 ( 
.A(n_1962),
.B(n_891),
.Y(n_2450)
);

INVx2_ASAP7_75t_L g2451 ( 
.A(n_2152),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2049),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_1962),
.B(n_757),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_1962),
.B(n_893),
.Y(n_2454)
);

AOI22xp33_ASAP7_75t_L g2455 ( 
.A1(n_1960),
.A2(n_894),
.B1(n_902),
.B2(n_893),
.Y(n_2455)
);

INVx3_ASAP7_75t_L g2456 ( 
.A(n_1972),
.Y(n_2456)
);

INVxp67_ASAP7_75t_L g2457 ( 
.A(n_1964),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_1962),
.B(n_894),
.Y(n_2458)
);

BUFx8_ASAP7_75t_L g2459 ( 
.A(n_2243),
.Y(n_2459)
);

BUFx12f_ASAP7_75t_L g2460 ( 
.A(n_2357),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2231),
.Y(n_2461)
);

AO21x2_ASAP7_75t_L g2462 ( 
.A1(n_2274),
.A2(n_903),
.B(n_902),
.Y(n_2462)
);

OAI21x1_ASAP7_75t_L g2463 ( 
.A1(n_2325),
.A2(n_1180),
.B(n_1179),
.Y(n_2463)
);

HB1xp67_ASAP7_75t_L g2464 ( 
.A(n_2196),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2251),
.Y(n_2465)
);

BUFx3_ASAP7_75t_L g2466 ( 
.A(n_2448),
.Y(n_2466)
);

AO21x1_ASAP7_75t_L g2467 ( 
.A1(n_2242),
.A2(n_906),
.B(n_903),
.Y(n_2467)
);

INVx5_ASAP7_75t_SL g2468 ( 
.A(n_2210),
.Y(n_2468)
);

INVx1_ASAP7_75t_SL g2469 ( 
.A(n_2203),
.Y(n_2469)
);

AOI22xp5_ASAP7_75t_L g2470 ( 
.A1(n_2195),
.A2(n_2355),
.B1(n_2380),
.B2(n_2369),
.Y(n_2470)
);

OA21x2_ASAP7_75t_L g2471 ( 
.A1(n_2294),
.A2(n_908),
.B(n_906),
.Y(n_2471)
);

HB1xp67_ASAP7_75t_L g2472 ( 
.A(n_2285),
.Y(n_2472)
);

OAI21x1_ASAP7_75t_L g2473 ( 
.A1(n_2436),
.A2(n_2371),
.B(n_2253),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2332),
.Y(n_2474)
);

INVx2_ASAP7_75t_SL g2475 ( 
.A(n_2272),
.Y(n_2475)
);

INVx4_ASAP7_75t_L g2476 ( 
.A(n_2326),
.Y(n_2476)
);

BUFx12f_ASAP7_75t_SL g2477 ( 
.A(n_2243),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2261),
.Y(n_2478)
);

HB1xp67_ASAP7_75t_L g2479 ( 
.A(n_2373),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2263),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2332),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_2205),
.B(n_908),
.Y(n_2482)
);

OAI21x1_ASAP7_75t_L g2483 ( 
.A1(n_2436),
.A2(n_1180),
.B(n_1179),
.Y(n_2483)
);

BUFx4_ASAP7_75t_SL g2484 ( 
.A(n_2191),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_L g2485 ( 
.A(n_2213),
.B(n_910),
.Y(n_2485)
);

BUFx2_ASAP7_75t_R g2486 ( 
.A(n_2399),
.Y(n_2486)
);

BUFx6f_ASAP7_75t_L g2487 ( 
.A(n_2266),
.Y(n_2487)
);

INVx5_ASAP7_75t_L g2488 ( 
.A(n_2438),
.Y(n_2488)
);

INVx4_ASAP7_75t_L g2489 ( 
.A(n_2326),
.Y(n_2489)
);

BUFx3_ASAP7_75t_L g2490 ( 
.A(n_2448),
.Y(n_2490)
);

AOI22xp33_ASAP7_75t_L g2491 ( 
.A1(n_2389),
.A2(n_910),
.B1(n_824),
.B2(n_826),
.Y(n_2491)
);

BUFx6f_ASAP7_75t_L g2492 ( 
.A(n_2266),
.Y(n_2492)
);

OAI21x1_ASAP7_75t_L g2493 ( 
.A1(n_2253),
.A2(n_1190),
.B(n_1184),
.Y(n_2493)
);

NAND2x1p5_ASAP7_75t_L g2494 ( 
.A(n_2326),
.B(n_1184),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2197),
.B(n_822),
.Y(n_2495)
);

NAND2x1p5_ASAP7_75t_L g2496 ( 
.A(n_2326),
.B(n_1190),
.Y(n_2496)
);

BUFx3_ASAP7_75t_L g2497 ( 
.A(n_2446),
.Y(n_2497)
);

INVx4_ASAP7_75t_L g2498 ( 
.A(n_2243),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_2331),
.Y(n_2499)
);

BUFx6f_ASAP7_75t_L g2500 ( 
.A(n_2266),
.Y(n_2500)
);

BUFx6f_ASAP7_75t_L g2501 ( 
.A(n_2266),
.Y(n_2501)
);

INVx1_ASAP7_75t_SL g2502 ( 
.A(n_2203),
.Y(n_2502)
);

OAI21x1_ASAP7_75t_L g2503 ( 
.A1(n_2344),
.A2(n_1202),
.B(n_1201),
.Y(n_2503)
);

BUFx6f_ASAP7_75t_L g2504 ( 
.A(n_2284),
.Y(n_2504)
);

INVx2_ASAP7_75t_SL g2505 ( 
.A(n_2272),
.Y(n_2505)
);

INVxp67_ASAP7_75t_L g2506 ( 
.A(n_2225),
.Y(n_2506)
);

OAI21x1_ASAP7_75t_L g2507 ( 
.A1(n_2346),
.A2(n_1202),
.B(n_1201),
.Y(n_2507)
);

OAI21xp5_ASAP7_75t_L g2508 ( 
.A1(n_2259),
.A2(n_826),
.B(n_824),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2447),
.Y(n_2509)
);

BUFx2_ASAP7_75t_L g2510 ( 
.A(n_2210),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2452),
.Y(n_2511)
);

AO21x2_ASAP7_75t_L g2512 ( 
.A1(n_2294),
.A2(n_831),
.B(n_830),
.Y(n_2512)
);

OAI21xp5_ASAP7_75t_L g2513 ( 
.A1(n_2259),
.A2(n_831),
.B(n_830),
.Y(n_2513)
);

INVx3_ASAP7_75t_L g2514 ( 
.A(n_2303),
.Y(n_2514)
);

INVx3_ASAP7_75t_SL g2515 ( 
.A(n_2369),
.Y(n_2515)
);

OAI21x1_ASAP7_75t_L g2516 ( 
.A1(n_2346),
.A2(n_1209),
.B(n_1207),
.Y(n_2516)
);

AND2x2_ASAP7_75t_L g2517 ( 
.A(n_2301),
.B(n_832),
.Y(n_2517)
);

BUFx8_ASAP7_75t_L g2518 ( 
.A(n_2243),
.Y(n_2518)
);

OR2x2_ASAP7_75t_L g2519 ( 
.A(n_2296),
.B(n_832),
.Y(n_2519)
);

AO21x2_ASAP7_75t_L g2520 ( 
.A1(n_2242),
.A2(n_834),
.B(n_833),
.Y(n_2520)
);

BUFx3_ASAP7_75t_L g2521 ( 
.A(n_2239),
.Y(n_2521)
);

OAI21x1_ASAP7_75t_L g2522 ( 
.A1(n_2353),
.A2(n_2219),
.B(n_2334),
.Y(n_2522)
);

OAI21x1_ASAP7_75t_SL g2523 ( 
.A1(n_2257),
.A2(n_834),
.B(n_833),
.Y(n_2523)
);

AOI22x1_ASAP7_75t_L g2524 ( 
.A1(n_2317),
.A2(n_1209),
.B1(n_1214),
.B2(n_1207),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2227),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2331),
.Y(n_2526)
);

INVx1_ASAP7_75t_SL g2527 ( 
.A(n_2260),
.Y(n_2527)
);

OAI21x1_ASAP7_75t_L g2528 ( 
.A1(n_2353),
.A2(n_1237),
.B(n_1214),
.Y(n_2528)
);

AO21x1_ASAP7_75t_L g2529 ( 
.A1(n_2244),
.A2(n_1241),
.B(n_1237),
.Y(n_2529)
);

OAI21x1_ASAP7_75t_L g2530 ( 
.A1(n_2334),
.A2(n_1260),
.B(n_1241),
.Y(n_2530)
);

BUFx6f_ASAP7_75t_L g2531 ( 
.A(n_2284),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2315),
.Y(n_2532)
);

BUFx12f_ASAP7_75t_L g2533 ( 
.A(n_2269),
.Y(n_2533)
);

INVx3_ASAP7_75t_L g2534 ( 
.A(n_2303),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2247),
.Y(n_2535)
);

OAI21x1_ASAP7_75t_L g2536 ( 
.A1(n_2361),
.A2(n_1260),
.B(n_1155),
.Y(n_2536)
);

OAI21x1_ASAP7_75t_L g2537 ( 
.A1(n_2361),
.A2(n_1155),
.B(n_1140),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2247),
.Y(n_2538)
);

HB1xp67_ASAP7_75t_L g2539 ( 
.A(n_2333),
.Y(n_2539)
);

BUFx6f_ASAP7_75t_L g2540 ( 
.A(n_2284),
.Y(n_2540)
);

INVxp67_ASAP7_75t_SL g2541 ( 
.A(n_2397),
.Y(n_2541)
);

OAI21xp5_ASAP7_75t_L g2542 ( 
.A1(n_2406),
.A2(n_1135),
.B(n_1130),
.Y(n_2542)
);

BUFx12f_ASAP7_75t_L g2543 ( 
.A(n_2215),
.Y(n_2543)
);

AO21x1_ASAP7_75t_L g2544 ( 
.A1(n_2244),
.A2(n_0),
.B(n_1),
.Y(n_2544)
);

INVx1_ASAP7_75t_SL g2545 ( 
.A(n_2264),
.Y(n_2545)
);

INVx5_ASAP7_75t_L g2546 ( 
.A(n_2438),
.Y(n_2546)
);

BUFx6f_ASAP7_75t_L g2547 ( 
.A(n_2284),
.Y(n_2547)
);

OAI21x1_ASAP7_75t_L g2548 ( 
.A1(n_2441),
.A2(n_1182),
.B(n_1155),
.Y(n_2548)
);

INVx3_ASAP7_75t_L g2549 ( 
.A(n_2303),
.Y(n_2549)
);

AOI21xp5_ASAP7_75t_L g2550 ( 
.A1(n_2256),
.A2(n_1330),
.B(n_1315),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2316),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2341),
.Y(n_2552)
);

AND2x2_ASAP7_75t_L g2553 ( 
.A(n_2301),
.B(n_2),
.Y(n_2553)
);

BUFx8_ASAP7_75t_SL g2554 ( 
.A(n_2191),
.Y(n_2554)
);

OAI21x1_ASAP7_75t_L g2555 ( 
.A1(n_2442),
.A2(n_1183),
.B(n_1182),
.Y(n_2555)
);

OR2x6_ASAP7_75t_L g2556 ( 
.A(n_2210),
.B(n_1135),
.Y(n_2556)
);

AO21x2_ASAP7_75t_L g2557 ( 
.A1(n_2335),
.A2(n_1154),
.B(n_1152),
.Y(n_2557)
);

NOR2xp67_ASAP7_75t_L g2558 ( 
.A(n_2218),
.B(n_309),
.Y(n_2558)
);

AOI22xp33_ASAP7_75t_L g2559 ( 
.A1(n_2389),
.A2(n_952),
.B1(n_996),
.B2(n_950),
.Y(n_2559)
);

BUFx12f_ASAP7_75t_L g2560 ( 
.A(n_2372),
.Y(n_2560)
);

BUFx2_ASAP7_75t_L g2561 ( 
.A(n_2306),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_L g2562 ( 
.A(n_2234),
.B(n_2),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2232),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2216),
.Y(n_2564)
);

BUFx6f_ASAP7_75t_L g2565 ( 
.A(n_2272),
.Y(n_2565)
);

HB1xp67_ASAP7_75t_L g2566 ( 
.A(n_2329),
.Y(n_2566)
);

BUFx3_ASAP7_75t_L g2567 ( 
.A(n_2239),
.Y(n_2567)
);

INVx4_ASAP7_75t_L g2568 ( 
.A(n_2416),
.Y(n_2568)
);

OAI21xp5_ASAP7_75t_L g2569 ( 
.A1(n_2406),
.A2(n_1154),
.B(n_1152),
.Y(n_2569)
);

OAI21xp5_ASAP7_75t_L g2570 ( 
.A1(n_2404),
.A2(n_1158),
.B(n_1182),
.Y(n_2570)
);

INVx8_ASAP7_75t_L g2571 ( 
.A(n_2241),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2245),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2341),
.Y(n_2573)
);

INVx2_ASAP7_75t_L g2574 ( 
.A(n_2232),
.Y(n_2574)
);

AND2x2_ASAP7_75t_L g2575 ( 
.A(n_2397),
.B(n_3),
.Y(n_2575)
);

NOR2xp33_ASAP7_75t_L g2576 ( 
.A(n_2192),
.B(n_311),
.Y(n_2576)
);

NOR2xp33_ASAP7_75t_L g2577 ( 
.A(n_2222),
.B(n_312),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2233),
.Y(n_2578)
);

BUFx2_ASAP7_75t_R g2579 ( 
.A(n_2399),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2194),
.Y(n_2580)
);

HB1xp67_ASAP7_75t_L g2581 ( 
.A(n_2330),
.Y(n_2581)
);

AO21x2_ASAP7_75t_L g2582 ( 
.A1(n_2335),
.A2(n_1158),
.B(n_971),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_2194),
.Y(n_2583)
);

OAI21xp5_ASAP7_75t_L g2584 ( 
.A1(n_2404),
.A2(n_1183),
.B(n_971),
.Y(n_2584)
);

OAI21xp5_ASAP7_75t_L g2585 ( 
.A1(n_2414),
.A2(n_1183),
.B(n_971),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2299),
.B(n_3),
.Y(n_2586)
);

INVx4_ASAP7_75t_L g2587 ( 
.A(n_2416),
.Y(n_2587)
);

OAI21xp5_ASAP7_75t_L g2588 ( 
.A1(n_2414),
.A2(n_972),
.B(n_968),
.Y(n_2588)
);

AO21x2_ASAP7_75t_L g2589 ( 
.A1(n_2287),
.A2(n_972),
.B(n_968),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2359),
.Y(n_2590)
);

AND2x4_ASAP7_75t_L g2591 ( 
.A(n_2272),
.B(n_313),
.Y(n_2591)
);

BUFx4f_ASAP7_75t_L g2592 ( 
.A(n_2438),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2449),
.B(n_4),
.Y(n_2593)
);

AOI22xp33_ASAP7_75t_L g2594 ( 
.A1(n_2229),
.A2(n_952),
.B1(n_996),
.B2(n_950),
.Y(n_2594)
);

AND2x4_ASAP7_75t_L g2595 ( 
.A(n_2281),
.B(n_316),
.Y(n_2595)
);

AO21x2_ASAP7_75t_L g2596 ( 
.A1(n_2287),
.A2(n_972),
.B(n_968),
.Y(n_2596)
);

INVxp67_ASAP7_75t_SL g2597 ( 
.A(n_2265),
.Y(n_2597)
);

INVx2_ASAP7_75t_L g2598 ( 
.A(n_2201),
.Y(n_2598)
);

OAI21x1_ASAP7_75t_L g2599 ( 
.A1(n_2200),
.A2(n_979),
.B(n_973),
.Y(n_2599)
);

BUFx2_ASAP7_75t_SL g2600 ( 
.A(n_2438),
.Y(n_2600)
);

BUFx3_ASAP7_75t_L g2601 ( 
.A(n_2206),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2201),
.Y(n_2602)
);

OAI21xp5_ASAP7_75t_L g2603 ( 
.A1(n_2453),
.A2(n_979),
.B(n_973),
.Y(n_2603)
);

CKINVDCx5p33_ASAP7_75t_R g2604 ( 
.A(n_2355),
.Y(n_2604)
);

INVx4_ASAP7_75t_L g2605 ( 
.A(n_2395),
.Y(n_2605)
);

INVx4_ASAP7_75t_L g2606 ( 
.A(n_2402),
.Y(n_2606)
);

OAI21x1_ASAP7_75t_L g2607 ( 
.A1(n_2304),
.A2(n_979),
.B(n_973),
.Y(n_2607)
);

AND2x4_ASAP7_75t_L g2608 ( 
.A(n_2281),
.B(n_320),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2450),
.B(n_5),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2202),
.Y(n_2610)
);

NAND2x1p5_ASAP7_75t_L g2611 ( 
.A(n_2293),
.B(n_1146),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2238),
.B(n_5),
.Y(n_2612)
);

INVx1_ASAP7_75t_SL g2613 ( 
.A(n_2206),
.Y(n_2613)
);

INVx8_ASAP7_75t_L g2614 ( 
.A(n_2241),
.Y(n_2614)
);

AND2x2_ASAP7_75t_L g2615 ( 
.A(n_2302),
.B(n_6),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_2310),
.B(n_7),
.Y(n_2616)
);

INVx3_ASAP7_75t_L g2617 ( 
.A(n_2351),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2352),
.Y(n_2618)
);

OAI21x1_ASAP7_75t_L g2619 ( 
.A1(n_2314),
.A2(n_984),
.B(n_983),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2360),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_2310),
.B(n_7),
.Y(n_2621)
);

AO21x2_ASAP7_75t_L g2622 ( 
.A1(n_2320),
.A2(n_2256),
.B(n_2293),
.Y(n_2622)
);

AO21x2_ASAP7_75t_L g2623 ( 
.A1(n_2320),
.A2(n_984),
.B(n_983),
.Y(n_2623)
);

AO21x2_ASAP7_75t_L g2624 ( 
.A1(n_2367),
.A2(n_984),
.B(n_983),
.Y(n_2624)
);

AND2x2_ASAP7_75t_L g2625 ( 
.A(n_2302),
.B(n_2370),
.Y(n_2625)
);

BUFx2_ASAP7_75t_R g2626 ( 
.A(n_2430),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2202),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2211),
.Y(n_2628)
);

OAI21x1_ASAP7_75t_L g2629 ( 
.A1(n_2415),
.A2(n_987),
.B(n_986),
.Y(n_2629)
);

BUFx10_ASAP7_75t_L g2630 ( 
.A(n_2372),
.Y(n_2630)
);

INVx3_ASAP7_75t_L g2631 ( 
.A(n_2351),
.Y(n_2631)
);

OAI21x1_ASAP7_75t_L g2632 ( 
.A1(n_2415),
.A2(n_2359),
.B(n_2422),
.Y(n_2632)
);

BUFx8_ASAP7_75t_L g2633 ( 
.A(n_2327),
.Y(n_2633)
);

AO21x2_ASAP7_75t_L g2634 ( 
.A1(n_2367),
.A2(n_987),
.B(n_986),
.Y(n_2634)
);

AOI22x1_ASAP7_75t_L g2635 ( 
.A1(n_2372),
.A2(n_987),
.B1(n_1001),
.B2(n_986),
.Y(n_2635)
);

OA21x2_ASAP7_75t_L g2636 ( 
.A1(n_2193),
.A2(n_2267),
.B(n_2347),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2221),
.Y(n_2637)
);

BUFx4_ASAP7_75t_SL g2638 ( 
.A(n_2380),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_L g2639 ( 
.A(n_2212),
.B(n_8),
.Y(n_2639)
);

INVx2_ASAP7_75t_L g2640 ( 
.A(n_2221),
.Y(n_2640)
);

BUFx2_ASAP7_75t_SL g2641 ( 
.A(n_2438),
.Y(n_2641)
);

BUFx2_ASAP7_75t_R g2642 ( 
.A(n_2456),
.Y(n_2642)
);

BUFx3_ASAP7_75t_L g2643 ( 
.A(n_2206),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2223),
.Y(n_2644)
);

CKINVDCx20_ASAP7_75t_R g2645 ( 
.A(n_2292),
.Y(n_2645)
);

OAI21x1_ASAP7_75t_L g2646 ( 
.A1(n_2423),
.A2(n_1008),
.B(n_1001),
.Y(n_2646)
);

OAI21x1_ASAP7_75t_SL g2647 ( 
.A1(n_2214),
.A2(n_1008),
.B(n_1001),
.Y(n_2647)
);

BUFx4_ASAP7_75t_SL g2648 ( 
.A(n_2432),
.Y(n_2648)
);

BUFx8_ASAP7_75t_SL g2649 ( 
.A(n_2209),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2223),
.Y(n_2650)
);

BUFx2_ASAP7_75t_R g2651 ( 
.A(n_2456),
.Y(n_2651)
);

OAI21x1_ASAP7_75t_L g2652 ( 
.A1(n_2425),
.A2(n_1010),
.B(n_1008),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2388),
.B(n_8),
.Y(n_2653)
);

BUFx2_ASAP7_75t_R g2654 ( 
.A(n_2193),
.Y(n_2654)
);

INVx2_ASAP7_75t_L g2655 ( 
.A(n_2451),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2451),
.Y(n_2656)
);

OAI21x1_ASAP7_75t_SL g2657 ( 
.A1(n_2252),
.A2(n_1011),
.B(n_1010),
.Y(n_2657)
);

INVx6_ASAP7_75t_L g2658 ( 
.A(n_2281),
.Y(n_2658)
);

AO21x2_ASAP7_75t_L g2659 ( 
.A1(n_2240),
.A2(n_2429),
.B(n_2426),
.Y(n_2659)
);

INVx3_ASAP7_75t_L g2660 ( 
.A(n_2351),
.Y(n_2660)
);

BUFx6f_ASAP7_75t_L g2661 ( 
.A(n_2281),
.Y(n_2661)
);

OAI21x1_ASAP7_75t_L g2662 ( 
.A1(n_2428),
.A2(n_1011),
.B(n_1010),
.Y(n_2662)
);

OAI21x1_ASAP7_75t_L g2663 ( 
.A1(n_2248),
.A2(n_1013),
.B(n_1011),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2370),
.Y(n_2664)
);

NOR2xp67_ASAP7_75t_L g2665 ( 
.A(n_2457),
.B(n_323),
.Y(n_2665)
);

INVx3_ASAP7_75t_L g2666 ( 
.A(n_2248),
.Y(n_2666)
);

CKINVDCx14_ASAP7_75t_R g2667 ( 
.A(n_2209),
.Y(n_2667)
);

BUFx12f_ASAP7_75t_L g2668 ( 
.A(n_2209),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_L g2669 ( 
.A(n_2226),
.B(n_2279),
.Y(n_2669)
);

NOR2x1_ASAP7_75t_SL g2670 ( 
.A(n_2440),
.B(n_1146),
.Y(n_2670)
);

NOR2xp33_ASAP7_75t_L g2671 ( 
.A(n_2207),
.B(n_325),
.Y(n_2671)
);

OR2x6_ASAP7_75t_L g2672 ( 
.A(n_2306),
.B(n_1013),
.Y(n_2672)
);

OAI21x1_ASAP7_75t_L g2673 ( 
.A1(n_2345),
.A2(n_1026),
.B(n_1013),
.Y(n_2673)
);

INVx5_ASAP7_75t_L g2674 ( 
.A(n_2400),
.Y(n_2674)
);

OAI21x1_ASAP7_75t_L g2675 ( 
.A1(n_2345),
.A2(n_1031),
.B(n_1026),
.Y(n_2675)
);

HB1xp67_ASAP7_75t_L g2676 ( 
.A(n_2308),
.Y(n_2676)
);

BUFx10_ASAP7_75t_L g2677 ( 
.A(n_2241),
.Y(n_2677)
);

OAI21x1_ASAP7_75t_L g2678 ( 
.A1(n_2348),
.A2(n_1031),
.B(n_1026),
.Y(n_2678)
);

INVx1_ASAP7_75t_SL g2679 ( 
.A(n_2229),
.Y(n_2679)
);

AOI21xp5_ASAP7_75t_L g2680 ( 
.A1(n_2236),
.A2(n_1330),
.B(n_1315),
.Y(n_2680)
);

OAI21x1_ASAP7_75t_L g2681 ( 
.A1(n_2348),
.A2(n_1034),
.B(n_1031),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2366),
.Y(n_2682)
);

BUFx6f_ASAP7_75t_L g2683 ( 
.A(n_2306),
.Y(n_2683)
);

AOI22x1_ASAP7_75t_L g2684 ( 
.A1(n_2444),
.A2(n_1034),
.B1(n_1187),
.B2(n_1181),
.Y(n_2684)
);

BUFx4_ASAP7_75t_SL g2685 ( 
.A(n_2385),
.Y(n_2685)
);

INVx2_ASAP7_75t_L g2686 ( 
.A(n_2376),
.Y(n_2686)
);

OAI21x1_ASAP7_75t_L g2687 ( 
.A1(n_2350),
.A2(n_1034),
.B(n_916),
.Y(n_2687)
);

AOI22x1_ASAP7_75t_L g2688 ( 
.A1(n_2410),
.A2(n_1187),
.B1(n_1192),
.B2(n_1181),
.Y(n_2688)
);

OR3x4_ASAP7_75t_SL g2689 ( 
.A(n_2204),
.B(n_9),
.C(n_11),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2376),
.Y(n_2690)
);

OAI21x1_ASAP7_75t_L g2691 ( 
.A1(n_2350),
.A2(n_916),
.B(n_1181),
.Y(n_2691)
);

BUFx3_ASAP7_75t_L g2692 ( 
.A(n_2249),
.Y(n_2692)
);

AND2x2_ASAP7_75t_SL g2693 ( 
.A(n_2228),
.B(n_9),
.Y(n_2693)
);

INVxp67_ASAP7_75t_SL g2694 ( 
.A(n_2379),
.Y(n_2694)
);

BUFx3_ASAP7_75t_L g2695 ( 
.A(n_2249),
.Y(n_2695)
);

BUFx2_ASAP7_75t_L g2696 ( 
.A(n_2308),
.Y(n_2696)
);

BUFx5_ASAP7_75t_L g2697 ( 
.A(n_2319),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2386),
.Y(n_2698)
);

BUFx2_ASAP7_75t_SL g2699 ( 
.A(n_2249),
.Y(n_2699)
);

AO21x2_ASAP7_75t_L g2700 ( 
.A1(n_2240),
.A2(n_327),
.B(n_326),
.Y(n_2700)
);

OAI21xp5_ASAP7_75t_L g2701 ( 
.A1(n_2362),
.A2(n_916),
.B(n_939),
.Y(n_2701)
);

BUFx3_ASAP7_75t_L g2702 ( 
.A(n_2249),
.Y(n_2702)
);

INVx2_ASAP7_75t_SL g2703 ( 
.A(n_2308),
.Y(n_2703)
);

OAI21x1_ASAP7_75t_SL g2704 ( 
.A1(n_2237),
.A2(n_330),
.B(n_329),
.Y(n_2704)
);

AO21x2_ASAP7_75t_L g2705 ( 
.A1(n_2431),
.A2(n_332),
.B(n_331),
.Y(n_2705)
);

INVx4_ASAP7_75t_L g2706 ( 
.A(n_2374),
.Y(n_2706)
);

NOR2xp33_ASAP7_75t_L g2707 ( 
.A(n_2321),
.B(n_333),
.Y(n_2707)
);

AOI21x1_ASAP7_75t_L g2708 ( 
.A1(n_2381),
.A2(n_1187),
.B(n_1181),
.Y(n_2708)
);

BUFx3_ASAP7_75t_L g2709 ( 
.A(n_2308),
.Y(n_2709)
);

OA21x2_ASAP7_75t_L g2710 ( 
.A1(n_2347),
.A2(n_930),
.B(n_927),
.Y(n_2710)
);

AO21x2_ASAP7_75t_L g2711 ( 
.A1(n_2433),
.A2(n_2381),
.B(n_2435),
.Y(n_2711)
);

BUFx3_ASAP7_75t_L g2712 ( 
.A(n_2276),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2454),
.B(n_11),
.Y(n_2713)
);

AND2x4_ASAP7_75t_L g2714 ( 
.A(n_2276),
.B(n_335),
.Y(n_2714)
);

INVx4_ASAP7_75t_L g2715 ( 
.A(n_2374),
.Y(n_2715)
);

NOR2xp33_ASAP7_75t_L g2716 ( 
.A(n_2401),
.B(n_338),
.Y(n_2716)
);

BUFx2_ASAP7_75t_L g2717 ( 
.A(n_2312),
.Y(n_2717)
);

BUFx3_ASAP7_75t_L g2718 ( 
.A(n_2297),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2390),
.Y(n_2719)
);

AND2x4_ASAP7_75t_L g2720 ( 
.A(n_2297),
.B(n_339),
.Y(n_2720)
);

AOI21x1_ASAP7_75t_L g2721 ( 
.A1(n_2434),
.A2(n_1192),
.B(n_1187),
.Y(n_2721)
);

AOI22xp33_ASAP7_75t_L g2722 ( 
.A1(n_2693),
.A2(n_2275),
.B1(n_2364),
.B2(n_2362),
.Y(n_2722)
);

INVx2_ASAP7_75t_L g2723 ( 
.A(n_2509),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2525),
.Y(n_2724)
);

INVx4_ASAP7_75t_L g2725 ( 
.A(n_2543),
.Y(n_2725)
);

CKINVDCx20_ASAP7_75t_R g2726 ( 
.A(n_2554),
.Y(n_2726)
);

CKINVDCx11_ASAP7_75t_R g2727 ( 
.A(n_2515),
.Y(n_2727)
);

INVx6_ASAP7_75t_L g2728 ( 
.A(n_2633),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2578),
.Y(n_2729)
);

OAI22xp33_ASAP7_75t_L g2730 ( 
.A1(n_2679),
.A2(n_2420),
.B1(n_2458),
.B2(n_2358),
.Y(n_2730)
);

INVx6_ASAP7_75t_L g2731 ( 
.A(n_2633),
.Y(n_2731)
);

INVx6_ASAP7_75t_L g2732 ( 
.A(n_2633),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2682),
.Y(n_2733)
);

AOI21xp5_ASAP7_75t_L g2734 ( 
.A1(n_2550),
.A2(n_2228),
.B(n_2235),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_2597),
.B(n_2379),
.Y(n_2735)
);

BUFx4f_ASAP7_75t_SL g2736 ( 
.A(n_2645),
.Y(n_2736)
);

INVx1_ASAP7_75t_SL g2737 ( 
.A(n_2696),
.Y(n_2737)
);

BUFx8_ASAP7_75t_L g2738 ( 
.A(n_2460),
.Y(n_2738)
);

AOI22xp33_ASAP7_75t_SL g2739 ( 
.A1(n_2693),
.A2(n_2328),
.B1(n_2445),
.B2(n_2443),
.Y(n_2739)
);

NAND2x1p5_ASAP7_75t_L g2740 ( 
.A(n_2488),
.B(n_2322),
.Y(n_2740)
);

INVx4_ASAP7_75t_L g2741 ( 
.A(n_2543),
.Y(n_2741)
);

AOI22xp33_ASAP7_75t_L g2742 ( 
.A1(n_2560),
.A2(n_2275),
.B1(n_2364),
.B2(n_2208),
.Y(n_2742)
);

INVx6_ASAP7_75t_L g2743 ( 
.A(n_2605),
.Y(n_2743)
);

OAI22xp5_ASAP7_75t_L g2744 ( 
.A1(n_2506),
.A2(n_2208),
.B1(n_2421),
.B2(n_2455),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2625),
.B(n_2318),
.Y(n_2745)
);

BUFx8_ASAP7_75t_L g2746 ( 
.A(n_2460),
.Y(n_2746)
);

AOI22xp33_ASAP7_75t_L g2747 ( 
.A1(n_2560),
.A2(n_2291),
.B1(n_2421),
.B2(n_2328),
.Y(n_2747)
);

INVxp67_ASAP7_75t_SL g2748 ( 
.A(n_2694),
.Y(n_2748)
);

BUFx8_ASAP7_75t_L g2749 ( 
.A(n_2615),
.Y(n_2749)
);

INVx3_ASAP7_75t_L g2750 ( 
.A(n_2709),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2698),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2625),
.B(n_2318),
.Y(n_2752)
);

BUFx6f_ASAP7_75t_L g2753 ( 
.A(n_2709),
.Y(n_2753)
);

BUFx3_ASAP7_75t_L g2754 ( 
.A(n_2649),
.Y(n_2754)
);

AOI22xp33_ASAP7_75t_SL g2755 ( 
.A1(n_2700),
.A2(n_2328),
.B1(n_2437),
.B2(n_2391),
.Y(n_2755)
);

OAI22xp33_ASAP7_75t_L g2756 ( 
.A1(n_2515),
.A2(n_2424),
.B1(n_2408),
.B2(n_2278),
.Y(n_2756)
);

BUFx3_ASAP7_75t_L g2757 ( 
.A(n_2649),
.Y(n_2757)
);

HB1xp67_ASAP7_75t_L g2758 ( 
.A(n_2472),
.Y(n_2758)
);

OAI21xp5_ASAP7_75t_SL g2759 ( 
.A1(n_2470),
.A2(n_2455),
.B(n_2349),
.Y(n_2759)
);

BUFx2_ASAP7_75t_L g2760 ( 
.A(n_2696),
.Y(n_2760)
);

INVx2_ASAP7_75t_L g2761 ( 
.A(n_2511),
.Y(n_2761)
);

BUFx2_ASAP7_75t_L g2762 ( 
.A(n_2676),
.Y(n_2762)
);

BUFx4f_ASAP7_75t_SL g2763 ( 
.A(n_2645),
.Y(n_2763)
);

AOI22xp33_ASAP7_75t_L g2764 ( 
.A1(n_2533),
.A2(n_2323),
.B1(n_2273),
.B2(n_2300),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2719),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2478),
.Y(n_2766)
);

AOI22xp33_ASAP7_75t_L g2767 ( 
.A1(n_2533),
.A2(n_2339),
.B1(n_2377),
.B2(n_2343),
.Y(n_2767)
);

HB1xp67_ASAP7_75t_L g2768 ( 
.A(n_2479),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2480),
.Y(n_2769)
);

AOI22xp33_ASAP7_75t_L g2770 ( 
.A1(n_2659),
.A2(n_2378),
.B1(n_2383),
.B2(n_2246),
.Y(n_2770)
);

BUFx6f_ASAP7_75t_L g2771 ( 
.A(n_2487),
.Y(n_2771)
);

AOI22xp5_ASAP7_75t_L g2772 ( 
.A1(n_2659),
.A2(n_2204),
.B1(n_2230),
.B2(n_2258),
.Y(n_2772)
);

AOI22xp33_ASAP7_75t_L g2773 ( 
.A1(n_2659),
.A2(n_2576),
.B1(n_2707),
.B2(n_2716),
.Y(n_2773)
);

INVx6_ASAP7_75t_L g2774 ( 
.A(n_2605),
.Y(n_2774)
);

CKINVDCx5p33_ASAP7_75t_R g2775 ( 
.A(n_2554),
.Y(n_2775)
);

BUFx2_ASAP7_75t_L g2776 ( 
.A(n_2717),
.Y(n_2776)
);

AOI21xp33_ASAP7_75t_L g2777 ( 
.A1(n_2711),
.A2(n_2405),
.B(n_2340),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2532),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2551),
.Y(n_2779)
);

OAI21xp5_ASAP7_75t_L g2780 ( 
.A1(n_2701),
.A2(n_2427),
.B(n_2396),
.Y(n_2780)
);

AOI22xp33_ASAP7_75t_L g2781 ( 
.A1(n_2683),
.A2(n_2217),
.B1(n_2394),
.B2(n_2393),
.Y(n_2781)
);

AOI22xp33_ASAP7_75t_L g2782 ( 
.A1(n_2683),
.A2(n_2313),
.B1(n_2387),
.B2(n_2392),
.Y(n_2782)
);

AOI22xp33_ASAP7_75t_L g2783 ( 
.A1(n_2683),
.A2(n_2356),
.B1(n_2418),
.B2(n_2411),
.Y(n_2783)
);

CKINVDCx20_ASAP7_75t_R g2784 ( 
.A(n_2667),
.Y(n_2784)
);

OAI22xp5_ASAP7_75t_L g2785 ( 
.A1(n_2592),
.A2(n_2654),
.B1(n_2593),
.B2(n_2609),
.Y(n_2785)
);

CKINVDCx20_ASAP7_75t_R g2786 ( 
.A(n_2667),
.Y(n_2786)
);

OAI22xp5_ASAP7_75t_L g2787 ( 
.A1(n_2592),
.A2(n_2224),
.B1(n_2198),
.B2(n_2199),
.Y(n_2787)
);

BUFx12f_ASAP7_75t_L g2788 ( 
.A(n_2604),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2461),
.Y(n_2789)
);

BUFx12f_ASAP7_75t_L g2790 ( 
.A(n_2604),
.Y(n_2790)
);

CKINVDCx16_ASAP7_75t_R g2791 ( 
.A(n_2668),
.Y(n_2791)
);

AOI22xp33_ASAP7_75t_SL g2792 ( 
.A1(n_2700),
.A2(n_2398),
.B1(n_2374),
.B2(n_2230),
.Y(n_2792)
);

BUFx4f_ASAP7_75t_L g2793 ( 
.A(n_2689),
.Y(n_2793)
);

OAI21xp5_ASAP7_75t_L g2794 ( 
.A1(n_2632),
.A2(n_2324),
.B(n_2336),
.Y(n_2794)
);

BUFx6f_ASAP7_75t_L g2795 ( 
.A(n_2487),
.Y(n_2795)
);

AOI22xp33_ASAP7_75t_L g2796 ( 
.A1(n_2683),
.A2(n_2398),
.B1(n_2374),
.B2(n_2338),
.Y(n_2796)
);

AOI22xp33_ASAP7_75t_SL g2797 ( 
.A1(n_2700),
.A2(n_2398),
.B1(n_2220),
.B2(n_2413),
.Y(n_2797)
);

AND2x4_ASAP7_75t_L g2798 ( 
.A(n_2561),
.B(n_2398),
.Y(n_2798)
);

CKINVDCx5p33_ASAP7_75t_R g2799 ( 
.A(n_2484),
.Y(n_2799)
);

OAI21xp5_ASAP7_75t_SL g2800 ( 
.A1(n_2615),
.A2(n_2375),
.B(n_2342),
.Y(n_2800)
);

BUFx4f_ASAP7_75t_L g2801 ( 
.A(n_2689),
.Y(n_2801)
);

AOI22xp33_ASAP7_75t_L g2802 ( 
.A1(n_2683),
.A2(n_2354),
.B1(n_2363),
.B2(n_2337),
.Y(n_2802)
);

CKINVDCx20_ASAP7_75t_R g2803 ( 
.A(n_2527),
.Y(n_2803)
);

AOI22xp33_ASAP7_75t_L g2804 ( 
.A1(n_2711),
.A2(n_2510),
.B1(n_2544),
.B2(n_2630),
.Y(n_2804)
);

BUFx4f_ASAP7_75t_L g2805 ( 
.A(n_2591),
.Y(n_2805)
);

AOI22xp33_ASAP7_75t_L g2806 ( 
.A1(n_2711),
.A2(n_2384),
.B1(n_2250),
.B2(n_2254),
.Y(n_2806)
);

BUFx12f_ASAP7_75t_L g2807 ( 
.A(n_2605),
.Y(n_2807)
);

OAI22xp5_ASAP7_75t_L g2808 ( 
.A1(n_2592),
.A2(n_2403),
.B1(n_2255),
.B2(n_2268),
.Y(n_2808)
);

BUFx2_ASAP7_75t_L g2809 ( 
.A(n_2717),
.Y(n_2809)
);

AOI22xp33_ASAP7_75t_L g2810 ( 
.A1(n_2510),
.A2(n_2311),
.B1(n_2309),
.B2(n_2412),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2552),
.Y(n_2811)
);

AOI22xp33_ASAP7_75t_SL g2812 ( 
.A1(n_2674),
.A2(n_2220),
.B1(n_2365),
.B2(n_2407),
.Y(n_2812)
);

INVx6_ASAP7_75t_L g2813 ( 
.A(n_2606),
.Y(n_2813)
);

BUFx2_ASAP7_75t_L g2814 ( 
.A(n_2692),
.Y(n_2814)
);

OAI22xp33_ASAP7_75t_L g2815 ( 
.A1(n_2674),
.A2(n_2417),
.B1(n_2409),
.B2(n_2289),
.Y(n_2815)
);

CKINVDCx5p33_ASAP7_75t_R g2816 ( 
.A(n_2638),
.Y(n_2816)
);

AOI22xp33_ASAP7_75t_L g2817 ( 
.A1(n_2544),
.A2(n_2419),
.B1(n_2277),
.B2(n_2280),
.Y(n_2817)
);

OAI22xp5_ASAP7_75t_L g2818 ( 
.A1(n_2713),
.A2(n_2674),
.B1(n_2639),
.B2(n_2586),
.Y(n_2818)
);

AOI22xp33_ASAP7_75t_L g2819 ( 
.A1(n_2630),
.A2(n_2419),
.B1(n_2288),
.B2(n_2295),
.Y(n_2819)
);

INVx2_ASAP7_75t_L g2820 ( 
.A(n_2465),
.Y(n_2820)
);

BUFx3_ASAP7_75t_L g2821 ( 
.A(n_2521),
.Y(n_2821)
);

OAI22xp5_ASAP7_75t_L g2822 ( 
.A1(n_2674),
.A2(n_2298),
.B1(n_2307),
.B2(n_2271),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_2572),
.Y(n_2823)
);

BUFx6f_ASAP7_75t_SL g2824 ( 
.A(n_2521),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2618),
.Y(n_2825)
);

INVx6_ASAP7_75t_L g2826 ( 
.A(n_2606),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2552),
.Y(n_2827)
);

CKINVDCx20_ASAP7_75t_R g2828 ( 
.A(n_2601),
.Y(n_2828)
);

AND2x2_ASAP7_75t_L g2829 ( 
.A(n_2561),
.B(n_2514),
.Y(n_2829)
);

AOI22xp5_ASAP7_75t_L g2830 ( 
.A1(n_2577),
.A2(n_2258),
.B1(n_2382),
.B2(n_2365),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2620),
.Y(n_2831)
);

AOI22xp33_ASAP7_75t_L g2832 ( 
.A1(n_2630),
.A2(n_2270),
.B1(n_2282),
.B2(n_2262),
.Y(n_2832)
);

OAI22xp5_ASAP7_75t_L g2833 ( 
.A1(n_2674),
.A2(n_2290),
.B1(n_2283),
.B2(n_2270),
.Y(n_2833)
);

AOI22xp33_ASAP7_75t_SL g2834 ( 
.A1(n_2704),
.A2(n_2368),
.B1(n_2282),
.B2(n_2286),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2590),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2590),
.Y(n_2836)
);

AOI22xp33_ASAP7_75t_L g2837 ( 
.A1(n_2672),
.A2(n_2286),
.B1(n_2305),
.B2(n_2262),
.Y(n_2837)
);

AOI22xp33_ASAP7_75t_SL g2838 ( 
.A1(n_2704),
.A2(n_2368),
.B1(n_2305),
.B2(n_2439),
.Y(n_2838)
);

INVx2_ASAP7_75t_L g2839 ( 
.A(n_2564),
.Y(n_2839)
);

OAI21xp5_ASAP7_75t_SL g2840 ( 
.A1(n_2491),
.A2(n_2653),
.B(n_2594),
.Y(n_2840)
);

INVx1_ASAP7_75t_SL g2841 ( 
.A(n_2539),
.Y(n_2841)
);

CKINVDCx11_ASAP7_75t_R g2842 ( 
.A(n_2469),
.Y(n_2842)
);

AOI22xp33_ASAP7_75t_L g2843 ( 
.A1(n_2672),
.A2(n_952),
.B1(n_996),
.B2(n_950),
.Y(n_2843)
);

OAI22xp33_ASAP7_75t_L g2844 ( 
.A1(n_2502),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_2844)
);

INVx6_ASAP7_75t_L g2845 ( 
.A(n_2606),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2541),
.B(n_14),
.Y(n_2846)
);

INVx2_ASAP7_75t_L g2847 ( 
.A(n_2474),
.Y(n_2847)
);

AOI22xp33_ASAP7_75t_L g2848 ( 
.A1(n_2672),
.A2(n_952),
.B1(n_996),
.B2(n_950),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2474),
.Y(n_2849)
);

AOI22xp33_ASAP7_75t_L g2850 ( 
.A1(n_2672),
.A2(n_952),
.B1(n_996),
.B2(n_950),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2481),
.Y(n_2851)
);

OAI22xp5_ASAP7_75t_L g2852 ( 
.A1(n_2669),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_2852)
);

CKINVDCx6p67_ASAP7_75t_R g2853 ( 
.A(n_2567),
.Y(n_2853)
);

AOI22xp33_ASAP7_75t_L g2854 ( 
.A1(n_2617),
.A2(n_952),
.B1(n_996),
.B2(n_950),
.Y(n_2854)
);

BUFx3_ASAP7_75t_L g2855 ( 
.A(n_2567),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2664),
.B(n_16),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2481),
.Y(n_2857)
);

INVx6_ASAP7_75t_L g2858 ( 
.A(n_2459),
.Y(n_2858)
);

CKINVDCx6p67_ASAP7_75t_R g2859 ( 
.A(n_2545),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2664),
.B(n_17),
.Y(n_2860)
);

INVx6_ASAP7_75t_L g2861 ( 
.A(n_2459),
.Y(n_2861)
);

OAI22xp33_ASAP7_75t_L g2862 ( 
.A1(n_2568),
.A2(n_21),
.B1(n_18),
.B2(n_19),
.Y(n_2862)
);

CKINVDCx11_ASAP7_75t_R g2863 ( 
.A(n_2668),
.Y(n_2863)
);

INVx1_ASAP7_75t_SL g2864 ( 
.A(n_2464),
.Y(n_2864)
);

BUFx3_ASAP7_75t_L g2865 ( 
.A(n_2692),
.Y(n_2865)
);

INVx4_ASAP7_75t_L g2866 ( 
.A(n_2568),
.Y(n_2866)
);

AOI22xp33_ASAP7_75t_L g2867 ( 
.A1(n_2617),
.A2(n_2660),
.B1(n_2631),
.B2(n_2534),
.Y(n_2867)
);

INVx6_ASAP7_75t_L g2868 ( 
.A(n_2459),
.Y(n_2868)
);

OAI22xp5_ASAP7_75t_L g2869 ( 
.A1(n_2562),
.A2(n_22),
.B1(n_19),
.B2(n_21),
.Y(n_2869)
);

CKINVDCx11_ASAP7_75t_R g2870 ( 
.A(n_2677),
.Y(n_2870)
);

INVx5_ASAP7_75t_L g2871 ( 
.A(n_2488),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2580),
.Y(n_2872)
);

AND2x2_ASAP7_75t_L g2873 ( 
.A(n_2514),
.B(n_22),
.Y(n_2873)
);

OAI22xp5_ASAP7_75t_L g2874 ( 
.A1(n_2612),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_2874)
);

CKINVDCx11_ASAP7_75t_R g2875 ( 
.A(n_2677),
.Y(n_2875)
);

INVx1_ASAP7_75t_SL g2876 ( 
.A(n_2566),
.Y(n_2876)
);

OAI22x1_ASAP7_75t_SL g2877 ( 
.A1(n_2648),
.A2(n_28),
.B1(n_24),
.B2(n_27),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2580),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_2686),
.Y(n_2879)
);

BUFx6f_ASAP7_75t_L g2880 ( 
.A(n_2487),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2686),
.Y(n_2881)
);

AND2x2_ASAP7_75t_L g2882 ( 
.A(n_2514),
.B(n_27),
.Y(n_2882)
);

AOI22xp33_ASAP7_75t_L g2883 ( 
.A1(n_2617),
.A2(n_1005),
.B1(n_997),
.B2(n_927),
.Y(n_2883)
);

NAND2x1p5_ASAP7_75t_L g2884 ( 
.A(n_2488),
.B(n_927),
.Y(n_2884)
);

BUFx2_ASAP7_75t_L g2885 ( 
.A(n_2695),
.Y(n_2885)
);

OAI22xp5_ASAP7_75t_L g2886 ( 
.A1(n_2488),
.A2(n_31),
.B1(n_28),
.B2(n_29),
.Y(n_2886)
);

BUFx4_ASAP7_75t_SL g2887 ( 
.A(n_2695),
.Y(n_2887)
);

BUFx12f_ASAP7_75t_L g2888 ( 
.A(n_2591),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2583),
.Y(n_2889)
);

OAI22xp33_ASAP7_75t_L g2890 ( 
.A1(n_2568),
.A2(n_32),
.B1(n_29),
.B2(n_31),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2583),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_L g2892 ( 
.A(n_2690),
.B(n_32),
.Y(n_2892)
);

AOI22xp33_ASAP7_75t_L g2893 ( 
.A1(n_2631),
.A2(n_1005),
.B1(n_997),
.B2(n_927),
.Y(n_2893)
);

BUFx2_ASAP7_75t_L g2894 ( 
.A(n_2702),
.Y(n_2894)
);

NAND2x1p5_ASAP7_75t_L g2895 ( 
.A(n_2488),
.B(n_927),
.Y(n_2895)
);

BUFx3_ASAP7_75t_L g2896 ( 
.A(n_2702),
.Y(n_2896)
);

BUFx12f_ASAP7_75t_L g2897 ( 
.A(n_2591),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2690),
.B(n_33),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2598),
.Y(n_2899)
);

OAI22xp5_ASAP7_75t_L g2900 ( 
.A1(n_2546),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_2900)
);

OAI22xp33_ASAP7_75t_L g2901 ( 
.A1(n_2587),
.A2(n_37),
.B1(n_34),
.B2(n_36),
.Y(n_2901)
);

OAI21xp5_ASAP7_75t_L g2902 ( 
.A1(n_2632),
.A2(n_916),
.B(n_939),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_L g2903 ( 
.A(n_2628),
.B(n_37),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2598),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2602),
.Y(n_2905)
);

BUFx2_ASAP7_75t_L g2906 ( 
.A(n_2466),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2602),
.Y(n_2907)
);

AOI22xp33_ASAP7_75t_L g2908 ( 
.A1(n_2631),
.A2(n_1005),
.B1(n_997),
.B2(n_932),
.Y(n_2908)
);

INVx4_ASAP7_75t_L g2909 ( 
.A(n_2587),
.Y(n_2909)
);

NAND2x1p5_ASAP7_75t_L g2910 ( 
.A(n_2546),
.B(n_930),
.Y(n_2910)
);

BUFx3_ASAP7_75t_L g2911 ( 
.A(n_2581),
.Y(n_2911)
);

AOI22xp33_ASAP7_75t_L g2912 ( 
.A1(n_2660),
.A2(n_1005),
.B1(n_997),
.B2(n_932),
.Y(n_2912)
);

INVx3_ASAP7_75t_L g2913 ( 
.A(n_2587),
.Y(n_2913)
);

INVx1_ASAP7_75t_SL g2914 ( 
.A(n_2497),
.Y(n_2914)
);

BUFx8_ASAP7_75t_L g2915 ( 
.A(n_2575),
.Y(n_2915)
);

INVx5_ASAP7_75t_L g2916 ( 
.A(n_2546),
.Y(n_2916)
);

BUFx6f_ASAP7_75t_L g2917 ( 
.A(n_2487),
.Y(n_2917)
);

AOI22xp33_ASAP7_75t_SL g2918 ( 
.A1(n_2636),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_2918)
);

BUFx3_ASAP7_75t_L g2919 ( 
.A(n_2497),
.Y(n_2919)
);

OAI21xp5_ASAP7_75t_SL g2920 ( 
.A1(n_2508),
.A2(n_39),
.B(n_40),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2610),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2610),
.Y(n_2922)
);

INVx2_ASAP7_75t_L g2923 ( 
.A(n_2627),
.Y(n_2923)
);

BUFx2_ASAP7_75t_SL g2924 ( 
.A(n_2703),
.Y(n_2924)
);

AOI22xp33_ASAP7_75t_L g2925 ( 
.A1(n_2660),
.A2(n_1005),
.B1(n_997),
.B2(n_932),
.Y(n_2925)
);

OAI22xp5_ASAP7_75t_L g2926 ( 
.A1(n_2546),
.A2(n_46),
.B1(n_42),
.B2(n_45),
.Y(n_2926)
);

OAI21xp5_ASAP7_75t_SL g2927 ( 
.A1(n_2513),
.A2(n_45),
.B(n_47),
.Y(n_2927)
);

CKINVDCx20_ASAP7_75t_R g2928 ( 
.A(n_2601),
.Y(n_2928)
);

CKINVDCx11_ASAP7_75t_R g2929 ( 
.A(n_2677),
.Y(n_2929)
);

OAI22xp5_ASAP7_75t_L g2930 ( 
.A1(n_2546),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2627),
.Y(n_2931)
);

AOI22xp33_ASAP7_75t_L g2932 ( 
.A1(n_2534),
.A2(n_1005),
.B1(n_997),
.B2(n_932),
.Y(n_2932)
);

BUFx3_ASAP7_75t_L g2933 ( 
.A(n_2466),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2640),
.Y(n_2934)
);

AOI22xp5_ASAP7_75t_L g2935 ( 
.A1(n_2558),
.A2(n_932),
.B1(n_934),
.B2(n_930),
.Y(n_2935)
);

CKINVDCx6p67_ASAP7_75t_R g2936 ( 
.A(n_2490),
.Y(n_2936)
);

AOI22xp33_ASAP7_75t_L g2937 ( 
.A1(n_2534),
.A2(n_932),
.B1(n_934),
.B2(n_930),
.Y(n_2937)
);

CKINVDCx10_ASAP7_75t_R g2938 ( 
.A(n_2685),
.Y(n_2938)
);

INVx6_ASAP7_75t_L g2939 ( 
.A(n_2518),
.Y(n_2939)
);

INVx2_ASAP7_75t_L g2940 ( 
.A(n_2640),
.Y(n_2940)
);

BUFx3_ASAP7_75t_L g2941 ( 
.A(n_2490),
.Y(n_2941)
);

INVx4_ASAP7_75t_L g2942 ( 
.A(n_2595),
.Y(n_2942)
);

INVx6_ASAP7_75t_L g2943 ( 
.A(n_2518),
.Y(n_2943)
);

CKINVDCx11_ASAP7_75t_R g2944 ( 
.A(n_2487),
.Y(n_2944)
);

INVx3_ASAP7_75t_SL g2945 ( 
.A(n_2703),
.Y(n_2945)
);

BUFx12f_ASAP7_75t_L g2946 ( 
.A(n_2595),
.Y(n_2946)
);

BUFx6f_ASAP7_75t_L g2947 ( 
.A(n_2492),
.Y(n_2947)
);

INVx2_ASAP7_75t_L g2948 ( 
.A(n_2839),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_L g2949 ( 
.A(n_2748),
.B(n_2636),
.Y(n_2949)
);

AOI222xp33_ASAP7_75t_SL g2950 ( 
.A1(n_2877),
.A2(n_51),
.B1(n_53),
.B2(n_48),
.C1(n_50),
.C2(n_52),
.Y(n_2950)
);

A2O1A1Ixp33_ASAP7_75t_L g2951 ( 
.A1(n_2793),
.A2(n_2665),
.B(n_2671),
.C(n_2595),
.Y(n_2951)
);

A2O1A1Ixp33_ASAP7_75t_L g2952 ( 
.A1(n_2793),
.A2(n_2801),
.B(n_2927),
.C(n_2920),
.Y(n_2952)
);

AOI22xp5_ASAP7_75t_L g2953 ( 
.A1(n_2722),
.A2(n_2622),
.B1(n_2636),
.B2(n_2720),
.Y(n_2953)
);

AOI21xp5_ASAP7_75t_L g2954 ( 
.A1(n_2734),
.A2(n_2680),
.B(n_2489),
.Y(n_2954)
);

A2O1A1Ixp33_ASAP7_75t_L g2955 ( 
.A1(n_2801),
.A2(n_2608),
.B(n_2720),
.C(n_2641),
.Y(n_2955)
);

AOI221xp5_ASAP7_75t_L g2956 ( 
.A1(n_2852),
.A2(n_2621),
.B1(n_2616),
.B2(n_2485),
.C(n_2482),
.Y(n_2956)
);

BUFx2_ASAP7_75t_L g2957 ( 
.A(n_2906),
.Y(n_2957)
);

INVx2_ASAP7_75t_L g2958 ( 
.A(n_2825),
.Y(n_2958)
);

OAI22xp5_ASAP7_75t_L g2959 ( 
.A1(n_2920),
.A2(n_2651),
.B1(n_2642),
.B2(n_2486),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2724),
.Y(n_2960)
);

OAI21xp5_ASAP7_75t_L g2961 ( 
.A1(n_2927),
.A2(n_2473),
.B(n_2522),
.Y(n_2961)
);

INVx2_ASAP7_75t_L g2962 ( 
.A(n_2723),
.Y(n_2962)
);

OA21x2_ASAP7_75t_L g2963 ( 
.A1(n_2777),
.A2(n_2473),
.B(n_2607),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2729),
.Y(n_2964)
);

BUFx3_ASAP7_75t_L g2965 ( 
.A(n_2799),
.Y(n_2965)
);

OAI221xp5_ASAP7_75t_L g2966 ( 
.A1(n_2773),
.A2(n_2519),
.B1(n_2495),
.B2(n_2613),
.C(n_2706),
.Y(n_2966)
);

AOI22xp33_ASAP7_75t_L g2967 ( 
.A1(n_2739),
.A2(n_2622),
.B1(n_2523),
.B2(n_2549),
.Y(n_2967)
);

AOI21xp5_ASAP7_75t_L g2968 ( 
.A1(n_2734),
.A2(n_2489),
.B(n_2476),
.Y(n_2968)
);

AOI21xp5_ASAP7_75t_L g2969 ( 
.A1(n_2780),
.A2(n_2489),
.B(n_2476),
.Y(n_2969)
);

AOI221xp5_ASAP7_75t_L g2970 ( 
.A1(n_2852),
.A2(n_2575),
.B1(n_2553),
.B2(n_2523),
.C(n_2573),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_L g2971 ( 
.A(n_2733),
.B(n_2751),
.Y(n_2971)
);

AND2x2_ASAP7_75t_L g2972 ( 
.A(n_2776),
.B(n_2809),
.Y(n_2972)
);

AOI21xp5_ASAP7_75t_L g2973 ( 
.A1(n_2780),
.A2(n_2476),
.B(n_2622),
.Y(n_2973)
);

AOI21xp5_ASAP7_75t_L g2974 ( 
.A1(n_2805),
.A2(n_2467),
.B(n_2705),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2765),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2766),
.Y(n_2976)
);

OR2x6_ASAP7_75t_L g2977 ( 
.A(n_2740),
.B(n_2600),
.Y(n_2977)
);

INVx2_ASAP7_75t_L g2978 ( 
.A(n_2761),
.Y(n_2978)
);

INVx2_ASAP7_75t_L g2979 ( 
.A(n_2789),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2769),
.B(n_2697),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2778),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2820),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2779),
.Y(n_2983)
);

BUFx3_ASAP7_75t_L g2984 ( 
.A(n_2736),
.Y(n_2984)
);

AND2x4_ASAP7_75t_SL g2985 ( 
.A(n_2859),
.B(n_2492),
.Y(n_2985)
);

NOR4xp25_ASAP7_75t_L g2986 ( 
.A(n_2869),
.B(n_2553),
.C(n_2519),
.D(n_2637),
.Y(n_2986)
);

OAI21x1_ASAP7_75t_L g2987 ( 
.A1(n_2902),
.A2(n_2619),
.B(n_2607),
.Y(n_2987)
);

OAI22xp5_ASAP7_75t_L g2988 ( 
.A1(n_2742),
.A2(n_2579),
.B1(n_2641),
.B2(n_2600),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2831),
.Y(n_2989)
);

OAI21xp5_ASAP7_75t_L g2990 ( 
.A1(n_2759),
.A2(n_2522),
.B(n_2635),
.Y(n_2990)
);

INVx2_ASAP7_75t_L g2991 ( 
.A(n_2823),
.Y(n_2991)
);

AOI21xp5_ASAP7_75t_L g2992 ( 
.A1(n_2805),
.A2(n_2467),
.B(n_2705),
.Y(n_2992)
);

OAI21xp5_ASAP7_75t_L g2993 ( 
.A1(n_2759),
.A2(n_2635),
.B(n_2611),
.Y(n_2993)
);

OAI221xp5_ASAP7_75t_L g2994 ( 
.A1(n_2800),
.A2(n_2715),
.B1(n_2706),
.B2(n_2666),
.C(n_2643),
.Y(n_2994)
);

OAI22xp5_ASAP7_75t_L g2995 ( 
.A1(n_2918),
.A2(n_2468),
.B1(n_2626),
.B2(n_2556),
.Y(n_2995)
);

AND2x2_ASAP7_75t_L g2996 ( 
.A(n_2829),
.B(n_2549),
.Y(n_2996)
);

HB1xp67_ASAP7_75t_L g2997 ( 
.A(n_2758),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2811),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2841),
.B(n_2697),
.Y(n_2999)
);

OAI221xp5_ASAP7_75t_SL g3000 ( 
.A1(n_2800),
.A2(n_2559),
.B1(n_2556),
.B2(n_2549),
.C(n_2650),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2827),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2762),
.Y(n_3002)
);

NAND2x1_ASAP7_75t_L g3003 ( 
.A(n_2866),
.B(n_2658),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2760),
.Y(n_3004)
);

AND2x4_ASAP7_75t_L g3005 ( 
.A(n_2737),
.B(n_2666),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_L g3006 ( 
.A(n_2841),
.B(n_2697),
.Y(n_3006)
);

INVx2_ASAP7_75t_L g3007 ( 
.A(n_2847),
.Y(n_3007)
);

AO21x2_ASAP7_75t_L g3008 ( 
.A1(n_2777),
.A2(n_2647),
.B(n_2657),
.Y(n_3008)
);

INVx3_ASAP7_75t_L g3009 ( 
.A(n_2933),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2864),
.B(n_2697),
.Y(n_3010)
);

AOI21xp5_ASAP7_75t_L g3011 ( 
.A1(n_2787),
.A2(n_2705),
.B(n_2608),
.Y(n_3011)
);

OA21x2_ASAP7_75t_L g3012 ( 
.A1(n_2804),
.A2(n_2619),
.B(n_2555),
.Y(n_3012)
);

OR2x6_ASAP7_75t_L g3013 ( 
.A(n_2740),
.B(n_2833),
.Y(n_3013)
);

OAI22xp5_ASAP7_75t_L g3014 ( 
.A1(n_2744),
.A2(n_2468),
.B1(n_2556),
.B2(n_2471),
.Y(n_3014)
);

OAI21xp5_ASAP7_75t_L g3015 ( 
.A1(n_2755),
.A2(n_2611),
.B(n_2608),
.Y(n_3015)
);

INVx6_ASAP7_75t_L g3016 ( 
.A(n_2738),
.Y(n_3016)
);

AO22x1_ASAP7_75t_L g3017 ( 
.A1(n_2738),
.A2(n_2518),
.B1(n_2715),
.B2(n_2706),
.Y(n_3017)
);

CKINVDCx5p33_ASAP7_75t_R g3018 ( 
.A(n_2938),
.Y(n_3018)
);

AND2x2_ASAP7_75t_L g3019 ( 
.A(n_2768),
.B(n_2864),
.Y(n_3019)
);

INVx3_ASAP7_75t_L g3020 ( 
.A(n_2941),
.Y(n_3020)
);

NOR2xp33_ASAP7_75t_L g3021 ( 
.A(n_2763),
.B(n_2643),
.Y(n_3021)
);

BUFx3_ASAP7_75t_L g3022 ( 
.A(n_2816),
.Y(n_3022)
);

AND2x4_ASAP7_75t_L g3023 ( 
.A(n_2737),
.B(n_2666),
.Y(n_3023)
);

AOI21xp5_ASAP7_75t_L g3024 ( 
.A1(n_2787),
.A2(n_2462),
.B(n_2494),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2835),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_SL g3026 ( 
.A(n_2808),
.B(n_2718),
.Y(n_3026)
);

AO21x2_ASAP7_75t_L g3027 ( 
.A1(n_2902),
.A2(n_2647),
.B(n_2657),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2836),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2849),
.Y(n_3029)
);

AOI21xp5_ASAP7_75t_L g3030 ( 
.A1(n_2730),
.A2(n_2462),
.B(n_2494),
.Y(n_3030)
);

A2O1A1Ixp33_ASAP7_75t_L g3031 ( 
.A1(n_2830),
.A2(n_2720),
.B(n_2714),
.C(n_2718),
.Y(n_3031)
);

OA21x2_ASAP7_75t_L g3032 ( 
.A1(n_2794),
.A2(n_2555),
.B(n_2548),
.Y(n_3032)
);

OAI21x1_ASAP7_75t_SL g3033 ( 
.A1(n_2772),
.A2(n_2670),
.B(n_2715),
.Y(n_3033)
);

AO21x2_ASAP7_75t_L g3034 ( 
.A1(n_2794),
.A2(n_2462),
.B(n_2670),
.Y(n_3034)
);

AOI22xp33_ASAP7_75t_L g3035 ( 
.A1(n_2818),
.A2(n_2808),
.B1(n_2744),
.B2(n_2785),
.Y(n_3035)
);

A2O1A1Ixp33_ASAP7_75t_L g3036 ( 
.A1(n_2840),
.A2(n_2714),
.B(n_2505),
.C(n_2475),
.Y(n_3036)
);

OA21x2_ASAP7_75t_L g3037 ( 
.A1(n_2817),
.A2(n_2548),
.B(n_2599),
.Y(n_3037)
);

OAI211xp5_ASAP7_75t_L g3038 ( 
.A1(n_2869),
.A2(n_2656),
.B(n_2655),
.C(n_2644),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2851),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2857),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_2735),
.B(n_2697),
.Y(n_3041)
);

OAI21x1_ASAP7_75t_L g3042 ( 
.A1(n_2833),
.A2(n_2708),
.B(n_2652),
.Y(n_3042)
);

AO21x2_ASAP7_75t_L g3043 ( 
.A1(n_2815),
.A2(n_2529),
.B(n_2708),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_SL g3044 ( 
.A(n_2818),
.B(n_2697),
.Y(n_3044)
);

OAI21x1_ASAP7_75t_SL g3045 ( 
.A1(n_2886),
.A2(n_2655),
.B(n_2644),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2872),
.Y(n_3046)
);

OAI22xp5_ASAP7_75t_L g3047 ( 
.A1(n_2747),
.A2(n_2468),
.B1(n_2556),
.B2(n_2471),
.Y(n_3047)
);

A2O1A1Ixp33_ASAP7_75t_L g3048 ( 
.A1(n_2840),
.A2(n_2797),
.B(n_2792),
.C(n_2785),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2735),
.B(n_2745),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_SL g3050 ( 
.A(n_2791),
.B(n_2697),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_2745),
.B(n_2535),
.Y(n_3051)
);

OAI21x1_ASAP7_75t_L g3052 ( 
.A1(n_2822),
.A2(n_2652),
.B(n_2646),
.Y(n_3052)
);

OA21x2_ASAP7_75t_L g3053 ( 
.A1(n_2770),
.A2(n_2806),
.B(n_2867),
.Y(n_3053)
);

INVx4_ASAP7_75t_L g3054 ( 
.A(n_2728),
.Y(n_3054)
);

AOI21xp5_ASAP7_75t_L g3055 ( 
.A1(n_2871),
.A2(n_2496),
.B(n_2494),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_2752),
.B(n_2535),
.Y(n_3056)
);

OAI22xp5_ASAP7_75t_SL g3057 ( 
.A1(n_2726),
.A2(n_2658),
.B1(n_2699),
.B2(n_2661),
.Y(n_3057)
);

INVx2_ASAP7_75t_L g3058 ( 
.A(n_2922),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2878),
.Y(n_3059)
);

OAI22xp5_ASAP7_75t_L g3060 ( 
.A1(n_2886),
.A2(n_2468),
.B1(n_2471),
.B2(n_2699),
.Y(n_3060)
);

INVx1_ASAP7_75t_SL g3061 ( 
.A(n_2876),
.Y(n_3061)
);

OR2x2_ASAP7_75t_L g3062 ( 
.A(n_2752),
.B(n_2499),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_L g3063 ( 
.A(n_2889),
.B(n_2538),
.Y(n_3063)
);

AO31x2_ASAP7_75t_L g3064 ( 
.A1(n_2822),
.A2(n_2529),
.A3(n_2526),
.B(n_2499),
.Y(n_3064)
);

OAI21x1_ASAP7_75t_SL g3065 ( 
.A1(n_2900),
.A2(n_2538),
.B(n_2526),
.Y(n_3065)
);

INVx2_ASAP7_75t_L g3066 ( 
.A(n_2923),
.Y(n_3066)
);

INVx2_ASAP7_75t_L g3067 ( 
.A(n_2940),
.Y(n_3067)
);

AO21x2_ASAP7_75t_L g3068 ( 
.A1(n_2846),
.A2(n_2596),
.B(n_2589),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_L g3069 ( 
.A(n_2891),
.B(n_2563),
.Y(n_3069)
);

A2O1A1Ixp33_ASAP7_75t_L g3070 ( 
.A1(n_2764),
.A2(n_2714),
.B(n_2475),
.C(n_2505),
.Y(n_3070)
);

INVx3_ASAP7_75t_L g3071 ( 
.A(n_2743),
.Y(n_3071)
);

OAI22xp33_ASAP7_75t_L g3072 ( 
.A1(n_2900),
.A2(n_2658),
.B1(n_2661),
.B2(n_2565),
.Y(n_3072)
);

HB1xp67_ASAP7_75t_L g3073 ( 
.A(n_2876),
.Y(n_3073)
);

OAI22xp33_ASAP7_75t_L g3074 ( 
.A1(n_2926),
.A2(n_2658),
.B1(n_2661),
.B2(n_2565),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_L g3075 ( 
.A(n_2899),
.B(n_2563),
.Y(n_3075)
);

AOI22xp33_ASAP7_75t_L g3076 ( 
.A1(n_2756),
.A2(n_2571),
.B1(n_2614),
.B2(n_2517),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2904),
.Y(n_3077)
);

NAND2x1p5_ASAP7_75t_L g3078 ( 
.A(n_2871),
.B(n_2565),
.Y(n_3078)
);

AOI21xp5_ASAP7_75t_L g3079 ( 
.A1(n_2871),
.A2(n_2496),
.B(n_2520),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2905),
.Y(n_3080)
);

AOI21xp5_ASAP7_75t_SL g3081 ( 
.A1(n_2926),
.A2(n_2661),
.B(n_2565),
.Y(n_3081)
);

AND2x4_ASAP7_75t_L g3082 ( 
.A(n_2798),
.B(n_2492),
.Y(n_3082)
);

CKINVDCx20_ASAP7_75t_R g3083 ( 
.A(n_2803),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_L g3084 ( 
.A(n_2907),
.B(n_2921),
.Y(n_3084)
);

INVx2_ASAP7_75t_L g3085 ( 
.A(n_2931),
.Y(n_3085)
);

OR2x2_ASAP7_75t_L g3086 ( 
.A(n_2911),
.B(n_2934),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2879),
.Y(n_3087)
);

AND2x2_ASAP7_75t_L g3088 ( 
.A(n_2919),
.B(n_2492),
.Y(n_3088)
);

OAI21x1_ASAP7_75t_L g3089 ( 
.A1(n_2884),
.A2(n_2662),
.B(n_2646),
.Y(n_3089)
);

AO21x2_ASAP7_75t_L g3090 ( 
.A1(n_2846),
.A2(n_2596),
.B(n_2589),
.Y(n_3090)
);

OAI221xp5_ASAP7_75t_L g3091 ( 
.A1(n_2802),
.A2(n_2712),
.B1(n_2611),
.B2(n_2603),
.C(n_2517),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_L g3092 ( 
.A(n_2881),
.B(n_2574),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_2914),
.B(n_2574),
.Y(n_3093)
);

AOI21xp5_ASAP7_75t_L g3094 ( 
.A1(n_2871),
.A2(n_2496),
.B(n_2520),
.Y(n_3094)
);

BUFx3_ASAP7_75t_L g3095 ( 
.A(n_2788),
.Y(n_3095)
);

AOI21xp5_ASAP7_75t_L g3096 ( 
.A1(n_2916),
.A2(n_2520),
.B(n_2565),
.Y(n_3096)
);

AOI21xp5_ASAP7_75t_L g3097 ( 
.A1(n_2916),
.A2(n_2661),
.B(n_2688),
.Y(n_3097)
);

OAI21xp5_ASAP7_75t_L g3098 ( 
.A1(n_2930),
.A2(n_2569),
.B(n_2542),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2856),
.Y(n_3099)
);

AOI21xp5_ASAP7_75t_L g3100 ( 
.A1(n_2916),
.A2(n_2688),
.B(n_2512),
.Y(n_3100)
);

BUFx2_ASAP7_75t_L g3101 ( 
.A(n_2814),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2856),
.Y(n_3102)
);

AOI21xp5_ASAP7_75t_L g3103 ( 
.A1(n_2916),
.A2(n_2512),
.B(n_2684),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2914),
.B(n_2589),
.Y(n_3104)
);

INVx2_ASAP7_75t_L g3105 ( 
.A(n_2885),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_2903),
.B(n_2596),
.Y(n_3106)
);

CKINVDCx20_ASAP7_75t_R g3107 ( 
.A(n_2727),
.Y(n_3107)
);

OAI221xp5_ASAP7_75t_L g3108 ( 
.A1(n_2767),
.A2(n_2712),
.B1(n_2498),
.B2(n_2500),
.C(n_2501),
.Y(n_3108)
);

INVx2_ASAP7_75t_L g3109 ( 
.A(n_2894),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_2903),
.B(n_2512),
.Y(n_3110)
);

NOR2xp33_ASAP7_75t_L g3111 ( 
.A(n_2842),
.B(n_2571),
.Y(n_3111)
);

AOI21xp5_ASAP7_75t_L g3112 ( 
.A1(n_2935),
.A2(n_2684),
.B(n_2557),
.Y(n_3112)
);

AOI221xp5_ASAP7_75t_L g3113 ( 
.A1(n_2844),
.A2(n_2500),
.B1(n_2504),
.B2(n_2501),
.C(n_2492),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_2860),
.B(n_2710),
.Y(n_3114)
);

NOR2xp67_ASAP7_75t_L g3115 ( 
.A(n_2725),
.B(n_2498),
.Y(n_3115)
);

AND2x2_ASAP7_75t_L g3116 ( 
.A(n_2798),
.B(n_2500),
.Y(n_3116)
);

AOI21xp5_ASAP7_75t_L g3117 ( 
.A1(n_2884),
.A2(n_2910),
.B(n_2895),
.Y(n_3117)
);

NAND2x1_ASAP7_75t_L g3118 ( 
.A(n_2866),
.B(n_2500),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2860),
.Y(n_3119)
);

OAI21x1_ASAP7_75t_L g3120 ( 
.A1(n_2895),
.A2(n_2662),
.B(n_2599),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2892),
.Y(n_3121)
);

CKINVDCx5p33_ASAP7_75t_R g3122 ( 
.A(n_2775),
.Y(n_3122)
);

CKINVDCx8_ASAP7_75t_R g3123 ( 
.A(n_2753),
.Y(n_3123)
);

BUFx3_ASAP7_75t_L g3124 ( 
.A(n_2790),
.Y(n_3124)
);

OAI21x1_ASAP7_75t_L g3125 ( 
.A1(n_2910),
.A2(n_2463),
.B(n_2691),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2892),
.Y(n_3126)
);

OAI21x1_ASAP7_75t_L g3127 ( 
.A1(n_2819),
.A2(n_2463),
.B(n_2691),
.Y(n_3127)
);

INVx4_ASAP7_75t_L g3128 ( 
.A(n_2728),
.Y(n_3128)
);

AO21x2_ASAP7_75t_L g3129 ( 
.A1(n_2898),
.A2(n_2623),
.B(n_2624),
.Y(n_3129)
);

INVx1_ASAP7_75t_SL g3130 ( 
.A(n_2945),
.Y(n_3130)
);

A2O1A1Ixp33_ASAP7_75t_L g3131 ( 
.A1(n_2874),
.A2(n_2571),
.B(n_2614),
.C(n_2588),
.Y(n_3131)
);

AOI22xp33_ASAP7_75t_L g3132 ( 
.A1(n_2930),
.A2(n_2614),
.B1(n_2571),
.B2(n_2501),
.Y(n_3132)
);

INVx2_ASAP7_75t_L g3133 ( 
.A(n_2750),
.Y(n_3133)
);

HB1xp67_ASAP7_75t_L g3134 ( 
.A(n_2750),
.Y(n_3134)
);

NOR2xp33_ASAP7_75t_L g3135 ( 
.A(n_2807),
.B(n_2614),
.Y(n_3135)
);

AO21x2_ASAP7_75t_L g3136 ( 
.A1(n_2898),
.A2(n_2623),
.B(n_2624),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2913),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2913),
.Y(n_3138)
);

OAI22xp33_ASAP7_75t_L g3139 ( 
.A1(n_2874),
.A2(n_2501),
.B1(n_2504),
.B2(n_2500),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2924),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_L g3141 ( 
.A(n_2832),
.B(n_2771),
.Y(n_3141)
);

O2A1O1Ixp33_ASAP7_75t_L g3142 ( 
.A1(n_2862),
.A2(n_2623),
.B(n_2634),
.C(n_2624),
.Y(n_3142)
);

OR2x2_ASAP7_75t_L g3143 ( 
.A(n_2865),
.B(n_2501),
.Y(n_3143)
);

AOI21xp5_ASAP7_75t_L g3144 ( 
.A1(n_2838),
.A2(n_2557),
.B(n_2634),
.Y(n_3144)
);

AND2x2_ASAP7_75t_L g3145 ( 
.A(n_2896),
.B(n_2504),
.Y(n_3145)
);

INVx1_ASAP7_75t_L g3146 ( 
.A(n_2873),
.Y(n_3146)
);

AOI21x1_ASAP7_75t_L g3147 ( 
.A1(n_2882),
.A2(n_2721),
.B(n_2710),
.Y(n_3147)
);

CKINVDCx6p67_ASAP7_75t_R g3148 ( 
.A(n_2824),
.Y(n_3148)
);

OAI211xp5_ASAP7_75t_L g3149 ( 
.A1(n_3035),
.A2(n_2783),
.B(n_2812),
.C(n_2810),
.Y(n_3149)
);

AOI22xp33_ASAP7_75t_L g3150 ( 
.A1(n_2959),
.A2(n_2749),
.B1(n_2915),
.B2(n_2901),
.Y(n_3150)
);

AOI22xp33_ASAP7_75t_L g3151 ( 
.A1(n_2959),
.A2(n_2956),
.B1(n_3098),
.B2(n_2995),
.Y(n_3151)
);

AND2x2_ASAP7_75t_L g3152 ( 
.A(n_2972),
.B(n_2725),
.Y(n_3152)
);

AOI22xp33_ASAP7_75t_L g3153 ( 
.A1(n_3098),
.A2(n_2890),
.B1(n_2749),
.B2(n_2915),
.Y(n_3153)
);

INVx4_ASAP7_75t_L g3154 ( 
.A(n_3016),
.Y(n_3154)
);

OAI221xp5_ASAP7_75t_L g3155 ( 
.A1(n_2952),
.A2(n_2796),
.B1(n_2782),
.B2(n_2781),
.C(n_2834),
.Y(n_3155)
);

OAI211xp5_ASAP7_75t_L g3156 ( 
.A1(n_3048),
.A2(n_2837),
.B(n_2875),
.C(n_2870),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2960),
.Y(n_3157)
);

NAND2xp5_ASAP7_75t_L g3158 ( 
.A(n_3049),
.B(n_3073),
.Y(n_3158)
);

INVx2_ASAP7_75t_L g3159 ( 
.A(n_3101),
.Y(n_3159)
);

OAI211xp5_ASAP7_75t_L g3160 ( 
.A1(n_3044),
.A2(n_2929),
.B(n_2863),
.C(n_2741),
.Y(n_3160)
);

AO222x2_ASAP7_75t_L g3161 ( 
.A1(n_2950),
.A2(n_52),
.B1(n_55),
.B2(n_50),
.C1(n_51),
.C2(n_54),
.Y(n_3161)
);

AND2x4_ASAP7_75t_L g3162 ( 
.A(n_3140),
.B(n_2821),
.Y(n_3162)
);

NOR2xp33_ASAP7_75t_SL g3163 ( 
.A(n_3107),
.B(n_2746),
.Y(n_3163)
);

OAI22xp5_ASAP7_75t_L g3164 ( 
.A1(n_3131),
.A2(n_2732),
.B1(n_2731),
.B2(n_2784),
.Y(n_3164)
);

AOI21xp5_ASAP7_75t_L g3165 ( 
.A1(n_3011),
.A2(n_2942),
.B(n_2741),
.Y(n_3165)
);

OAI22xp5_ASAP7_75t_L g3166 ( 
.A1(n_3031),
.A2(n_2732),
.B1(n_2731),
.B2(n_2786),
.Y(n_3166)
);

BUFx12f_ASAP7_75t_L g3167 ( 
.A(n_3018),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2964),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2975),
.Y(n_3169)
);

OAI221xp5_ASAP7_75t_SL g3170 ( 
.A1(n_2950),
.A2(n_2757),
.B1(n_2754),
.B2(n_2853),
.C(n_2848),
.Y(n_3170)
);

AOI33xp33_ASAP7_75t_L g3171 ( 
.A1(n_2986),
.A2(n_2850),
.A3(n_2843),
.B1(n_57),
.B2(n_61),
.B3(n_54),
.Y(n_3171)
);

OR2x6_ASAP7_75t_L g3172 ( 
.A(n_2973),
.B(n_2909),
.Y(n_3172)
);

OR2x2_ASAP7_75t_L g3173 ( 
.A(n_3049),
.B(n_2936),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_SL g3174 ( 
.A(n_3054),
.B(n_2753),
.Y(n_3174)
);

AND2x2_ASAP7_75t_L g3175 ( 
.A(n_2957),
.B(n_2855),
.Y(n_3175)
);

INVx2_ASAP7_75t_L g3176 ( 
.A(n_3133),
.Y(n_3176)
);

AOI22xp5_ASAP7_75t_L g3177 ( 
.A1(n_2995),
.A2(n_2828),
.B1(n_2928),
.B2(n_2824),
.Y(n_3177)
);

AOI221xp5_ASAP7_75t_L g3178 ( 
.A1(n_3139),
.A2(n_2753),
.B1(n_2909),
.B2(n_2795),
.C(n_2880),
.Y(n_3178)
);

AOI22xp33_ASAP7_75t_L g3179 ( 
.A1(n_2988),
.A2(n_2897),
.B1(n_2946),
.B2(n_2888),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2976),
.Y(n_3180)
);

AO21x2_ASAP7_75t_L g3181 ( 
.A1(n_2949),
.A2(n_2557),
.B(n_2634),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_L g3182 ( 
.A(n_3061),
.B(n_2743),
.Y(n_3182)
);

AOI22xp33_ASAP7_75t_L g3183 ( 
.A1(n_2988),
.A2(n_2942),
.B1(n_2774),
.B2(n_2826),
.Y(n_3183)
);

INVx3_ASAP7_75t_L g3184 ( 
.A(n_3071),
.Y(n_3184)
);

BUFx3_ASAP7_75t_L g3185 ( 
.A(n_2984),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_3061),
.B(n_2774),
.Y(n_3186)
);

OAI22xp33_ASAP7_75t_L g3187 ( 
.A1(n_2953),
.A2(n_2826),
.B1(n_2845),
.B2(n_2813),
.Y(n_3187)
);

AOI221xp5_ASAP7_75t_L g3188 ( 
.A1(n_3099),
.A2(n_2880),
.B1(n_2917),
.B2(n_2795),
.C(n_2771),
.Y(n_3188)
);

AOI22xp33_ASAP7_75t_L g3189 ( 
.A1(n_2966),
.A2(n_2813),
.B1(n_2845),
.B2(n_2746),
.Y(n_3189)
);

AND2x4_ASAP7_75t_SL g3190 ( 
.A(n_3083),
.B(n_2504),
.Y(n_3190)
);

OAI221xp5_ASAP7_75t_L g3191 ( 
.A1(n_3070),
.A2(n_2861),
.B1(n_2939),
.B2(n_2868),
.C(n_2858),
.Y(n_3191)
);

NAND3xp33_ASAP7_75t_L g3192 ( 
.A(n_2961),
.B(n_3026),
.C(n_3110),
.Y(n_3192)
);

AOI22xp33_ASAP7_75t_SL g3193 ( 
.A1(n_3053),
.A2(n_2861),
.B1(n_2868),
.B2(n_2858),
.Y(n_3193)
);

AOI22xp33_ASAP7_75t_L g3194 ( 
.A1(n_3053),
.A2(n_2943),
.B1(n_2939),
.B2(n_2531),
.Y(n_3194)
);

AOI22xp33_ASAP7_75t_L g3195 ( 
.A1(n_2994),
.A2(n_2943),
.B1(n_2531),
.B2(n_2540),
.Y(n_3195)
);

AOI221xp5_ASAP7_75t_SL g3196 ( 
.A1(n_3036),
.A2(n_2880),
.B1(n_2917),
.B2(n_2795),
.C(n_2771),
.Y(n_3196)
);

OAI221xp5_ASAP7_75t_L g3197 ( 
.A1(n_3076),
.A2(n_2498),
.B1(n_2947),
.B2(n_2917),
.C(n_2531),
.Y(n_3197)
);

AOI22xp33_ASAP7_75t_L g3198 ( 
.A1(n_3091),
.A2(n_2504),
.B1(n_2540),
.B2(n_2531),
.Y(n_3198)
);

AOI22xp33_ASAP7_75t_L g3199 ( 
.A1(n_3047),
.A2(n_2531),
.B1(n_2547),
.B2(n_2540),
.Y(n_3199)
);

A2O1A1Ixp33_ASAP7_75t_L g3200 ( 
.A1(n_3000),
.A2(n_2887),
.B(n_2547),
.C(n_2540),
.Y(n_3200)
);

AOI22xp33_ASAP7_75t_L g3201 ( 
.A1(n_3047),
.A2(n_3015),
.B1(n_2970),
.B2(n_3108),
.Y(n_3201)
);

AOI22xp33_ASAP7_75t_SL g3202 ( 
.A1(n_3038),
.A2(n_2547),
.B1(n_2540),
.B2(n_2582),
.Y(n_3202)
);

AND2x2_ASAP7_75t_L g3203 ( 
.A(n_2996),
.B(n_2944),
.Y(n_3203)
);

OAI211xp5_ASAP7_75t_L g3204 ( 
.A1(n_3113),
.A2(n_3081),
.B(n_2961),
.C(n_2993),
.Y(n_3204)
);

OAI22xp5_ASAP7_75t_L g3205 ( 
.A1(n_3132),
.A2(n_2951),
.B1(n_2955),
.B2(n_2967),
.Y(n_3205)
);

OAI22xp5_ASAP7_75t_L g3206 ( 
.A1(n_3015),
.A2(n_2547),
.B1(n_2854),
.B2(n_2947),
.Y(n_3206)
);

OAI221xp5_ASAP7_75t_L g3207 ( 
.A1(n_3102),
.A2(n_2947),
.B1(n_2547),
.B2(n_2932),
.C(n_2893),
.Y(n_3207)
);

AOI22xp33_ASAP7_75t_L g3208 ( 
.A1(n_2993),
.A2(n_2477),
.B1(n_2582),
.B2(n_2584),
.Y(n_3208)
);

AOI222xp33_ASAP7_75t_L g3209 ( 
.A1(n_3014),
.A2(n_2585),
.B1(n_57),
.B2(n_58),
.C1(n_61),
.C2(n_62),
.Y(n_3209)
);

OR2x2_ASAP7_75t_L g3210 ( 
.A(n_2997),
.B(n_2710),
.Y(n_3210)
);

A2O1A1Ixp33_ASAP7_75t_L g3211 ( 
.A1(n_2969),
.A2(n_2537),
.B(n_2570),
.C(n_2477),
.Y(n_3211)
);

AOI22xp33_ASAP7_75t_L g3212 ( 
.A1(n_3014),
.A2(n_2582),
.B1(n_2908),
.B2(n_2883),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_2981),
.Y(n_3213)
);

AOI22xp33_ASAP7_75t_SL g3214 ( 
.A1(n_3060),
.A2(n_2537),
.B1(n_2524),
.B2(n_2536),
.Y(n_3214)
);

HB1xp67_ASAP7_75t_L g3215 ( 
.A(n_2949),
.Y(n_3215)
);

OAI21xp33_ASAP7_75t_L g3216 ( 
.A1(n_3110),
.A2(n_2925),
.B(n_2912),
.Y(n_3216)
);

AOI22xp33_ASAP7_75t_L g3217 ( 
.A1(n_3030),
.A2(n_2937),
.B1(n_2524),
.B2(n_2503),
.Y(n_3217)
);

INVx1_ASAP7_75t_L g3218 ( 
.A(n_2983),
.Y(n_3218)
);

OAI22xp33_ASAP7_75t_L g3219 ( 
.A1(n_3148),
.A2(n_2721),
.B1(n_63),
.B2(n_56),
.Y(n_3219)
);

OAI22xp5_ASAP7_75t_L g3220 ( 
.A1(n_3057),
.A2(n_2536),
.B1(n_2663),
.B2(n_66),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_L g3221 ( 
.A(n_3019),
.B(n_2687),
.Y(n_3221)
);

HB1xp67_ASAP7_75t_L g3222 ( 
.A(n_3041),
.Y(n_3222)
);

AOI22xp33_ASAP7_75t_L g3223 ( 
.A1(n_3119),
.A2(n_2503),
.B1(n_2687),
.B2(n_2675),
.Y(n_3223)
);

AOI22xp33_ASAP7_75t_SL g3224 ( 
.A1(n_3060),
.A2(n_67),
.B1(n_56),
.B2(n_58),
.Y(n_3224)
);

INVx2_ASAP7_75t_SL g3225 ( 
.A(n_3016),
.Y(n_3225)
);

AOI22xp33_ASAP7_75t_L g3226 ( 
.A1(n_3121),
.A2(n_2663),
.B1(n_2629),
.B2(n_2493),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_L g3227 ( 
.A(n_3126),
.B(n_2493),
.Y(n_3227)
);

AOI22xp33_ASAP7_75t_L g3228 ( 
.A1(n_3013),
.A2(n_2629),
.B1(n_2507),
.B2(n_2516),
.Y(n_3228)
);

OAI22xp5_ASAP7_75t_SL g3229 ( 
.A1(n_3054),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_3051),
.B(n_2673),
.Y(n_3230)
);

AOI21xp5_ASAP7_75t_L g3231 ( 
.A1(n_2968),
.A2(n_2516),
.B(n_2507),
.Y(n_3231)
);

OA21x2_ASAP7_75t_L g3232 ( 
.A1(n_2980),
.A2(n_2675),
.B(n_2673),
.Y(n_3232)
);

AOI22xp33_ASAP7_75t_L g3233 ( 
.A1(n_2990),
.A2(n_2681),
.B1(n_2678),
.B2(n_2528),
.Y(n_3233)
);

AOI22xp33_ASAP7_75t_SL g3234 ( 
.A1(n_2990),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_3234)
);

OAI22xp5_ASAP7_75t_L g3235 ( 
.A1(n_3130),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_3235)
);

AOI22xp33_ASAP7_75t_L g3236 ( 
.A1(n_3072),
.A2(n_2681),
.B1(n_2678),
.B2(n_2528),
.Y(n_3236)
);

OAI22xp5_ASAP7_75t_L g3237 ( 
.A1(n_3130),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_3237)
);

OAI221xp5_ASAP7_75t_L g3238 ( 
.A1(n_3013),
.A2(n_79),
.B1(n_75),
.B2(n_78),
.C(n_80),
.Y(n_3238)
);

OAI22xp33_ASAP7_75t_L g3239 ( 
.A1(n_3128),
.A2(n_82),
.B1(n_78),
.B2(n_81),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_2989),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_2998),
.Y(n_3241)
);

AOI22xp33_ASAP7_75t_L g3242 ( 
.A1(n_3013),
.A2(n_2530),
.B1(n_2483),
.B2(n_932),
.Y(n_3242)
);

AO21x2_ASAP7_75t_L g3243 ( 
.A1(n_2954),
.A2(n_3033),
.B(n_2992),
.Y(n_3243)
);

CKINVDCx5p33_ASAP7_75t_R g3244 ( 
.A(n_3122),
.Y(n_3244)
);

AND2x4_ASAP7_75t_L g3245 ( 
.A(n_3005),
.B(n_2483),
.Y(n_3245)
);

OAI21x1_ASAP7_75t_L g3246 ( 
.A1(n_3096),
.A2(n_2530),
.B(n_83),
.Y(n_3246)
);

AOI22xp33_ASAP7_75t_SL g3247 ( 
.A1(n_3045),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_3247)
);

AND2x4_ASAP7_75t_L g3248 ( 
.A(n_3005),
.B(n_3023),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_3105),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_3001),
.Y(n_3250)
);

BUFx2_ASAP7_75t_L g3251 ( 
.A(n_3071),
.Y(n_3251)
);

OR2x2_ASAP7_75t_L g3252 ( 
.A(n_3041),
.B(n_84),
.Y(n_3252)
);

OR2x2_ASAP7_75t_L g3253 ( 
.A(n_3002),
.B(n_3004),
.Y(n_3253)
);

OAI22xp5_ASAP7_75t_L g3254 ( 
.A1(n_3074),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_3254)
);

INVxp33_ASAP7_75t_L g3255 ( 
.A(n_3111),
.Y(n_3255)
);

BUFx3_ASAP7_75t_L g3256 ( 
.A(n_2965),
.Y(n_3256)
);

OAI21xp33_ASAP7_75t_L g3257 ( 
.A1(n_3106),
.A2(n_87),
.B(n_90),
.Y(n_3257)
);

OAI211xp5_ASAP7_75t_L g3258 ( 
.A1(n_3142),
.A2(n_92),
.B(n_90),
.C(n_91),
.Y(n_3258)
);

AOI22xp33_ASAP7_75t_L g3259 ( 
.A1(n_3146),
.A2(n_934),
.B1(n_930),
.B2(n_1187),
.Y(n_3259)
);

AND2x2_ASAP7_75t_L g3260 ( 
.A(n_3109),
.B(n_92),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_L g3261 ( 
.A(n_3051),
.B(n_93),
.Y(n_3261)
);

OAI221xp5_ASAP7_75t_L g3262 ( 
.A1(n_3141),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.C(n_97),
.Y(n_3262)
);

OAI221xp5_ASAP7_75t_L g3263 ( 
.A1(n_3141),
.A2(n_95),
.B1(n_96),
.B2(n_98),
.C(n_99),
.Y(n_3263)
);

OA21x2_ASAP7_75t_L g3264 ( 
.A1(n_2980),
.A2(n_99),
.B(n_100),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_3025),
.Y(n_3265)
);

INVx2_ASAP7_75t_L g3266 ( 
.A(n_3085),
.Y(n_3266)
);

OAI22xp5_ASAP7_75t_L g3267 ( 
.A1(n_3128),
.A2(n_102),
.B1(n_100),
.B2(n_101),
.Y(n_3267)
);

AOI21xp5_ASAP7_75t_L g3268 ( 
.A1(n_2974),
.A2(n_934),
.B(n_930),
.Y(n_3268)
);

CKINVDCx5p33_ASAP7_75t_R g3269 ( 
.A(n_3022),
.Y(n_3269)
);

INVx3_ASAP7_75t_L g3270 ( 
.A(n_3009),
.Y(n_3270)
);

AND2x2_ASAP7_75t_L g3271 ( 
.A(n_3134),
.B(n_3116),
.Y(n_3271)
);

AND2x2_ASAP7_75t_SL g3272 ( 
.A(n_2985),
.B(n_104),
.Y(n_3272)
);

OAI22xp5_ASAP7_75t_SL g3273 ( 
.A1(n_3095),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_3273)
);

AOI22xp33_ASAP7_75t_L g3274 ( 
.A1(n_3024),
.A2(n_110),
.B1(n_107),
.B2(n_109),
.Y(n_3274)
);

AOI21x1_ASAP7_75t_L g3275 ( 
.A1(n_3017),
.A2(n_107),
.B(n_111),
.Y(n_3275)
);

HB1xp67_ASAP7_75t_L g3276 ( 
.A(n_3028),
.Y(n_3276)
);

INVx1_ASAP7_75t_SL g3277 ( 
.A(n_3009),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_2971),
.Y(n_3278)
);

BUFx3_ASAP7_75t_L g3279 ( 
.A(n_3124),
.Y(n_3279)
);

AO21x2_ASAP7_75t_L g3280 ( 
.A1(n_3114),
.A2(n_111),
.B(n_112),
.Y(n_3280)
);

BUFx6f_ASAP7_75t_L g3281 ( 
.A(n_3003),
.Y(n_3281)
);

AOI22xp33_ASAP7_75t_L g3282 ( 
.A1(n_3065),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_3282)
);

AND2x2_ASAP7_75t_L g3283 ( 
.A(n_3020),
.B(n_3088),
.Y(n_3283)
);

OAI22xp5_ASAP7_75t_L g3284 ( 
.A1(n_3123),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_3284)
);

AOI22xp33_ASAP7_75t_L g3285 ( 
.A1(n_3144),
.A2(n_121),
.B1(n_118),
.B2(n_120),
.Y(n_3285)
);

NAND3xp33_ASAP7_75t_L g3286 ( 
.A(n_3106),
.B(n_934),
.C(n_930),
.Y(n_3286)
);

BUFx2_ASAP7_75t_L g3287 ( 
.A(n_3023),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_2971),
.Y(n_3288)
);

AOI221xp5_ASAP7_75t_L g3289 ( 
.A1(n_2999),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.C(n_124),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_3056),
.B(n_122),
.Y(n_3290)
);

NAND2x1_ASAP7_75t_L g3291 ( 
.A(n_2977),
.B(n_3020),
.Y(n_3291)
);

INVx11_ASAP7_75t_L g3292 ( 
.A(n_3021),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_3029),
.Y(n_3293)
);

OAI22xp5_ASAP7_75t_L g3294 ( 
.A1(n_2977),
.A2(n_126),
.B1(n_123),
.B2(n_124),
.Y(n_3294)
);

OAI21xp33_ASAP7_75t_SL g3295 ( 
.A1(n_3050),
.A2(n_126),
.B(n_128),
.Y(n_3295)
);

OA21x2_ASAP7_75t_L g3296 ( 
.A1(n_3114),
.A2(n_129),
.B(n_130),
.Y(n_3296)
);

OAI22xp5_ASAP7_75t_L g3297 ( 
.A1(n_2977),
.A2(n_132),
.B1(n_129),
.B2(n_130),
.Y(n_3297)
);

CKINVDCx5p33_ASAP7_75t_R g3298 ( 
.A(n_3145),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_3056),
.B(n_132),
.Y(n_3299)
);

A2O1A1Ixp33_ASAP7_75t_L g3300 ( 
.A1(n_3115),
.A2(n_135),
.B(n_133),
.C(n_134),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_3039),
.Y(n_3301)
);

AOI22xp5_ASAP7_75t_L g3302 ( 
.A1(n_3135),
.A2(n_3027),
.B1(n_3082),
.B2(n_3008),
.Y(n_3302)
);

AOI221xp5_ASAP7_75t_L g3303 ( 
.A1(n_2999),
.A2(n_135),
.B1(n_137),
.B2(n_138),
.C(n_139),
.Y(n_3303)
);

AOI22xp33_ASAP7_75t_L g3304 ( 
.A1(n_3027),
.A2(n_934),
.B1(n_1213),
.B2(n_1192),
.Y(n_3304)
);

BUFx12f_ASAP7_75t_L g3305 ( 
.A(n_3086),
.Y(n_3305)
);

OAI22xp5_ASAP7_75t_L g3306 ( 
.A1(n_3117),
.A2(n_140),
.B1(n_137),
.B2(n_139),
.Y(n_3306)
);

INVx2_ASAP7_75t_L g3307 ( 
.A(n_2948),
.Y(n_3307)
);

NOR2x1_ASAP7_75t_SL g3308 ( 
.A(n_3006),
.B(n_140),
.Y(n_3308)
);

AOI22xp33_ASAP7_75t_L g3309 ( 
.A1(n_3082),
.A2(n_934),
.B1(n_1213),
.B2(n_1192),
.Y(n_3309)
);

OAI221xp5_ASAP7_75t_L g3310 ( 
.A1(n_3006),
.A2(n_141),
.B1(n_142),
.B2(n_144),
.C(n_145),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_3276),
.Y(n_3311)
);

AND2x2_ASAP7_75t_L g3312 ( 
.A(n_3215),
.B(n_3034),
.Y(n_3312)
);

BUFx2_ASAP7_75t_L g3313 ( 
.A(n_3172),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_3276),
.Y(n_3314)
);

AND2x2_ASAP7_75t_L g3315 ( 
.A(n_3215),
.B(n_3222),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_3241),
.Y(n_3316)
);

AND2x2_ASAP7_75t_L g3317 ( 
.A(n_3287),
.B(n_3137),
.Y(n_3317)
);

INVx2_ASAP7_75t_L g3318 ( 
.A(n_3296),
.Y(n_3318)
);

AOI22xp33_ASAP7_75t_L g3319 ( 
.A1(n_3151),
.A2(n_3008),
.B1(n_3034),
.B2(n_3129),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_3250),
.Y(n_3320)
);

INVx4_ASAP7_75t_R g3321 ( 
.A(n_3225),
.Y(n_3321)
);

AND2x2_ASAP7_75t_L g3322 ( 
.A(n_3222),
.B(n_3138),
.Y(n_3322)
);

OR2x2_ASAP7_75t_L g3323 ( 
.A(n_3192),
.B(n_3062),
.Y(n_3323)
);

AND2x2_ASAP7_75t_L g3324 ( 
.A(n_3172),
.B(n_2958),
.Y(n_3324)
);

INVx1_ASAP7_75t_SL g3325 ( 
.A(n_3251),
.Y(n_3325)
);

BUFx2_ASAP7_75t_L g3326 ( 
.A(n_3172),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_3265),
.Y(n_3327)
);

AND2x2_ASAP7_75t_L g3328 ( 
.A(n_3243),
.B(n_3271),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_3293),
.Y(n_3329)
);

INVx2_ASAP7_75t_L g3330 ( 
.A(n_3296),
.Y(n_3330)
);

AND2x4_ASAP7_75t_L g3331 ( 
.A(n_3243),
.B(n_3010),
.Y(n_3331)
);

INVx2_ASAP7_75t_L g3332 ( 
.A(n_3264),
.Y(n_3332)
);

AND2x4_ASAP7_75t_L g3333 ( 
.A(n_3291),
.B(n_3010),
.Y(n_3333)
);

INVx2_ASAP7_75t_L g3334 ( 
.A(n_3264),
.Y(n_3334)
);

HB1xp67_ASAP7_75t_L g3335 ( 
.A(n_3280),
.Y(n_3335)
);

INVx4_ASAP7_75t_L g3336 ( 
.A(n_3154),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3301),
.Y(n_3337)
);

INVx2_ASAP7_75t_L g3338 ( 
.A(n_3280),
.Y(n_3338)
);

AND2x4_ASAP7_75t_L g3339 ( 
.A(n_3281),
.B(n_3007),
.Y(n_3339)
);

HB1xp67_ASAP7_75t_L g3340 ( 
.A(n_3210),
.Y(n_3340)
);

HB1xp67_ASAP7_75t_L g3341 ( 
.A(n_3278),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_3157),
.Y(n_3342)
);

AND2x2_ASAP7_75t_L g3343 ( 
.A(n_3193),
.B(n_2962),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3168),
.Y(n_3344)
);

INVx2_ASAP7_75t_L g3345 ( 
.A(n_3288),
.Y(n_3345)
);

INVx2_ASAP7_75t_L g3346 ( 
.A(n_3169),
.Y(n_3346)
);

AND2x2_ASAP7_75t_L g3347 ( 
.A(n_3193),
.B(n_2978),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_L g3348 ( 
.A(n_3158),
.B(n_2979),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_3180),
.Y(n_3349)
);

AO21x2_ASAP7_75t_L g3350 ( 
.A1(n_3268),
.A2(n_3100),
.B(n_3103),
.Y(n_3350)
);

INVx2_ASAP7_75t_L g3351 ( 
.A(n_3213),
.Y(n_3351)
);

AND2x2_ASAP7_75t_L g3352 ( 
.A(n_3159),
.B(n_3248),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_3218),
.Y(n_3353)
);

BUFx3_ASAP7_75t_L g3354 ( 
.A(n_3167),
.Y(n_3354)
);

HB1xp67_ASAP7_75t_L g3355 ( 
.A(n_3240),
.Y(n_3355)
);

AND2x2_ASAP7_75t_L g3356 ( 
.A(n_3248),
.B(n_2982),
.Y(n_3356)
);

OAI21xp33_ASAP7_75t_L g3357 ( 
.A1(n_3151),
.A2(n_3093),
.B(n_3104),
.Y(n_3357)
);

AND2x2_ASAP7_75t_L g3358 ( 
.A(n_3249),
.B(n_2991),
.Y(n_3358)
);

AND2x4_ASAP7_75t_L g3359 ( 
.A(n_3281),
.B(n_3058),
.Y(n_3359)
);

OR2x2_ASAP7_75t_L g3360 ( 
.A(n_3252),
.B(n_3307),
.Y(n_3360)
);

AND2x2_ASAP7_75t_L g3361 ( 
.A(n_3184),
.B(n_3143),
.Y(n_3361)
);

INVx2_ASAP7_75t_L g3362 ( 
.A(n_3266),
.Y(n_3362)
);

AND2x2_ASAP7_75t_L g3363 ( 
.A(n_3184),
.B(n_3066),
.Y(n_3363)
);

AND2x2_ASAP7_75t_L g3364 ( 
.A(n_3283),
.B(n_3067),
.Y(n_3364)
);

AND2x2_ASAP7_75t_L g3365 ( 
.A(n_3152),
.B(n_3270),
.Y(n_3365)
);

AND2x2_ASAP7_75t_L g3366 ( 
.A(n_3270),
.B(n_3087),
.Y(n_3366)
);

INVx1_ASAP7_75t_SL g3367 ( 
.A(n_3277),
.Y(n_3367)
);

INVx2_ASAP7_75t_L g3368 ( 
.A(n_3181),
.Y(n_3368)
);

INVx11_ASAP7_75t_L g3369 ( 
.A(n_3305),
.Y(n_3369)
);

HB1xp67_ASAP7_75t_L g3370 ( 
.A(n_3230),
.Y(n_3370)
);

AND2x2_ASAP7_75t_L g3371 ( 
.A(n_3175),
.B(n_3040),
.Y(n_3371)
);

BUFx3_ASAP7_75t_L g3372 ( 
.A(n_3154),
.Y(n_3372)
);

AND2x2_ASAP7_75t_L g3373 ( 
.A(n_3194),
.B(n_2963),
.Y(n_3373)
);

AND2x2_ASAP7_75t_L g3374 ( 
.A(n_3176),
.B(n_2963),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_L g3375 ( 
.A(n_3261),
.B(n_3046),
.Y(n_3375)
);

AOI22xp33_ASAP7_75t_L g3376 ( 
.A1(n_3209),
.A2(n_3129),
.B1(n_3136),
.B2(n_3037),
.Y(n_3376)
);

AND2x2_ASAP7_75t_L g3377 ( 
.A(n_3173),
.B(n_3059),
.Y(n_3377)
);

NOR2xp33_ASAP7_75t_SL g3378 ( 
.A(n_3170),
.B(n_3191),
.Y(n_3378)
);

INVx2_ASAP7_75t_L g3379 ( 
.A(n_3181),
.Y(n_3379)
);

INVx2_ASAP7_75t_L g3380 ( 
.A(n_3308),
.Y(n_3380)
);

AND2x2_ASAP7_75t_L g3381 ( 
.A(n_3302),
.B(n_3077),
.Y(n_3381)
);

AND2x2_ASAP7_75t_L g3382 ( 
.A(n_3199),
.B(n_3080),
.Y(n_3382)
);

INVx2_ASAP7_75t_SL g3383 ( 
.A(n_3281),
.Y(n_3383)
);

AND2x2_ASAP7_75t_L g3384 ( 
.A(n_3253),
.B(n_3064),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3227),
.Y(n_3385)
);

INVx2_ASAP7_75t_L g3386 ( 
.A(n_3221),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3290),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_3299),
.Y(n_3388)
);

BUFx2_ASAP7_75t_L g3389 ( 
.A(n_3281),
.Y(n_3389)
);

INVx1_ASAP7_75t_L g3390 ( 
.A(n_3245),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_3245),
.Y(n_3391)
);

BUFx4f_ASAP7_75t_SL g3392 ( 
.A(n_3185),
.Y(n_3392)
);

HB1xp67_ASAP7_75t_L g3393 ( 
.A(n_3246),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3182),
.Y(n_3394)
);

BUFx3_ASAP7_75t_L g3395 ( 
.A(n_3279),
.Y(n_3395)
);

OR2x2_ASAP7_75t_L g3396 ( 
.A(n_3186),
.B(n_3093),
.Y(n_3396)
);

HB1xp67_ASAP7_75t_L g3397 ( 
.A(n_3260),
.Y(n_3397)
);

INVx2_ASAP7_75t_L g3398 ( 
.A(n_3232),
.Y(n_3398)
);

INVx3_ASAP7_75t_L g3399 ( 
.A(n_3162),
.Y(n_3399)
);

INVx3_ASAP7_75t_L g3400 ( 
.A(n_3162),
.Y(n_3400)
);

AND2x2_ASAP7_75t_L g3401 ( 
.A(n_3201),
.B(n_3064),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_3174),
.Y(n_3402)
);

INVx2_ASAP7_75t_L g3403 ( 
.A(n_3232),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_L g3404 ( 
.A(n_3204),
.B(n_3084),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_3202),
.Y(n_3405)
);

AND2x2_ASAP7_75t_L g3406 ( 
.A(n_3202),
.B(n_3064),
.Y(n_3406)
);

AOI22xp33_ASAP7_75t_L g3407 ( 
.A1(n_3285),
.A2(n_3262),
.B1(n_3263),
.B2(n_3205),
.Y(n_3407)
);

AND2x2_ASAP7_75t_L g3408 ( 
.A(n_3196),
.B(n_3012),
.Y(n_3408)
);

AND2x4_ASAP7_75t_L g3409 ( 
.A(n_3165),
.B(n_3104),
.Y(n_3409)
);

INVx2_ASAP7_75t_SL g3410 ( 
.A(n_3292),
.Y(n_3410)
);

INVx2_ASAP7_75t_L g3411 ( 
.A(n_3275),
.Y(n_3411)
);

AND2x2_ASAP7_75t_L g3412 ( 
.A(n_3203),
.B(n_3078),
.Y(n_3412)
);

INVx2_ASAP7_75t_L g3413 ( 
.A(n_3286),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_3188),
.Y(n_3414)
);

INVx2_ASAP7_75t_L g3415 ( 
.A(n_3272),
.Y(n_3415)
);

INVxp67_ASAP7_75t_L g3416 ( 
.A(n_3238),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_3187),
.Y(n_3417)
);

AND2x4_ASAP7_75t_L g3418 ( 
.A(n_3190),
.B(n_3118),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_3187),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_3216),
.B(n_3084),
.Y(n_3420)
);

AND2x2_ASAP7_75t_L g3421 ( 
.A(n_3195),
.B(n_3012),
.Y(n_3421)
);

AND2x2_ASAP7_75t_L g3422 ( 
.A(n_3298),
.B(n_3032),
.Y(n_3422)
);

AND2x2_ASAP7_75t_SL g3423 ( 
.A(n_3171),
.B(n_3037),
.Y(n_3423)
);

INVx2_ASAP7_75t_L g3424 ( 
.A(n_3272),
.Y(n_3424)
);

AND2x2_ASAP7_75t_L g3425 ( 
.A(n_3255),
.B(n_3032),
.Y(n_3425)
);

BUFx3_ASAP7_75t_L g3426 ( 
.A(n_3256),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3206),
.Y(n_3427)
);

AND2x2_ASAP7_75t_L g3428 ( 
.A(n_3178),
.B(n_3043),
.Y(n_3428)
);

AND2x2_ASAP7_75t_L g3429 ( 
.A(n_3198),
.B(n_3043),
.Y(n_3429)
);

AND2x2_ASAP7_75t_L g3430 ( 
.A(n_3211),
.B(n_3136),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_3197),
.Y(n_3431)
);

AND2x2_ASAP7_75t_L g3432 ( 
.A(n_3200),
.B(n_3068),
.Y(n_3432)
);

INVx3_ASAP7_75t_L g3433 ( 
.A(n_3269),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_3160),
.Y(n_3434)
);

INVx2_ASAP7_75t_L g3435 ( 
.A(n_3310),
.Y(n_3435)
);

AND2x2_ASAP7_75t_L g3436 ( 
.A(n_3177),
.B(n_3068),
.Y(n_3436)
);

AND2x2_ASAP7_75t_L g3437 ( 
.A(n_3214),
.B(n_3090),
.Y(n_3437)
);

CKINVDCx20_ASAP7_75t_R g3438 ( 
.A(n_3244),
.Y(n_3438)
);

BUFx6f_ASAP7_75t_L g3439 ( 
.A(n_3234),
.Y(n_3439)
);

INVxp67_ASAP7_75t_L g3440 ( 
.A(n_3306),
.Y(n_3440)
);

AND2x2_ASAP7_75t_L g3441 ( 
.A(n_3214),
.B(n_3090),
.Y(n_3441)
);

INVx2_ASAP7_75t_L g3442 ( 
.A(n_3294),
.Y(n_3442)
);

INVx3_ASAP7_75t_L g3443 ( 
.A(n_3372),
.Y(n_3443)
);

OAI31xp33_ASAP7_75t_L g3444 ( 
.A1(n_3378),
.A2(n_3156),
.A3(n_3407),
.B(n_3435),
.Y(n_3444)
);

INVx1_ASAP7_75t_L g3445 ( 
.A(n_3355),
.Y(n_3445)
);

HB1xp67_ASAP7_75t_L g3446 ( 
.A(n_3318),
.Y(n_3446)
);

A2O1A1Ixp33_ASAP7_75t_L g3447 ( 
.A1(n_3439),
.A2(n_3170),
.B(n_3161),
.C(n_3258),
.Y(n_3447)
);

INVx3_ASAP7_75t_L g3448 ( 
.A(n_3372),
.Y(n_3448)
);

A2O1A1Ixp33_ASAP7_75t_L g3449 ( 
.A1(n_3439),
.A2(n_3257),
.B(n_3150),
.C(n_3149),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_3355),
.Y(n_3450)
);

A2O1A1Ixp33_ASAP7_75t_L g3451 ( 
.A1(n_3439),
.A2(n_3300),
.B(n_3285),
.C(n_3153),
.Y(n_3451)
);

NOR2xp33_ASAP7_75t_L g3452 ( 
.A(n_3416),
.B(n_3163),
.Y(n_3452)
);

OR2x2_ASAP7_75t_L g3453 ( 
.A(n_3323),
.B(n_3063),
.Y(n_3453)
);

AND2x4_ASAP7_75t_L g3454 ( 
.A(n_3399),
.B(n_3183),
.Y(n_3454)
);

INVxp67_ASAP7_75t_SL g3455 ( 
.A(n_3335),
.Y(n_3455)
);

INVx2_ASAP7_75t_L g3456 ( 
.A(n_3374),
.Y(n_3456)
);

AND2x2_ASAP7_75t_L g3457 ( 
.A(n_3352),
.B(n_3189),
.Y(n_3457)
);

AND2x2_ASAP7_75t_L g3458 ( 
.A(n_3352),
.B(n_3164),
.Y(n_3458)
);

AND2x2_ASAP7_75t_L g3459 ( 
.A(n_3352),
.B(n_3179),
.Y(n_3459)
);

NAND4xp25_ASAP7_75t_L g3460 ( 
.A(n_3378),
.B(n_3234),
.C(n_3303),
.D(n_3289),
.Y(n_3460)
);

A2O1A1Ixp33_ASAP7_75t_L g3461 ( 
.A1(n_3439),
.A2(n_3153),
.B(n_3166),
.C(n_3274),
.Y(n_3461)
);

AOI22xp33_ASAP7_75t_L g3462 ( 
.A1(n_3439),
.A2(n_3274),
.B1(n_3224),
.B2(n_3229),
.Y(n_3462)
);

BUFx6f_ASAP7_75t_L g3463 ( 
.A(n_3354),
.Y(n_3463)
);

OAI21xp5_ASAP7_75t_L g3464 ( 
.A1(n_3416),
.A2(n_3224),
.B(n_3247),
.Y(n_3464)
);

OA21x2_ASAP7_75t_L g3465 ( 
.A1(n_3405),
.A2(n_3231),
.B(n_3282),
.Y(n_3465)
);

BUFx2_ASAP7_75t_L g3466 ( 
.A(n_3372),
.Y(n_3466)
);

O2A1O1Ixp5_ASAP7_75t_L g3467 ( 
.A1(n_3435),
.A2(n_3239),
.B(n_3219),
.C(n_3254),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3316),
.Y(n_3468)
);

AOI21xp5_ASAP7_75t_L g3469 ( 
.A1(n_3423),
.A2(n_3219),
.B(n_3239),
.Y(n_3469)
);

NAND3xp33_ASAP7_75t_L g3470 ( 
.A(n_3439),
.B(n_3247),
.C(n_3282),
.Y(n_3470)
);

BUFx3_ASAP7_75t_L g3471 ( 
.A(n_3354),
.Y(n_3471)
);

AOI22xp33_ASAP7_75t_L g3472 ( 
.A1(n_3439),
.A2(n_3273),
.B1(n_3284),
.B2(n_3155),
.Y(n_3472)
);

INVx2_ASAP7_75t_SL g3473 ( 
.A(n_3369),
.Y(n_3473)
);

OAI221xp5_ASAP7_75t_L g3474 ( 
.A1(n_3435),
.A2(n_3295),
.B1(n_3235),
.B2(n_3237),
.C(n_3297),
.Y(n_3474)
);

AND2x4_ASAP7_75t_L g3475 ( 
.A(n_3399),
.B(n_3063),
.Y(n_3475)
);

OAI22xp5_ASAP7_75t_SL g3476 ( 
.A1(n_3434),
.A2(n_3267),
.B1(n_3208),
.B2(n_3207),
.Y(n_3476)
);

BUFx3_ASAP7_75t_L g3477 ( 
.A(n_3354),
.Y(n_3477)
);

OAI21xp5_ASAP7_75t_L g3478 ( 
.A1(n_3401),
.A2(n_3208),
.B(n_3212),
.Y(n_3478)
);

HB1xp67_ASAP7_75t_L g3479 ( 
.A(n_3318),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_L g3480 ( 
.A(n_3404),
.B(n_3212),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3316),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3320),
.Y(n_3482)
);

INVx2_ASAP7_75t_SL g3483 ( 
.A(n_3369),
.Y(n_3483)
);

INVx2_ASAP7_75t_L g3484 ( 
.A(n_3339),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_L g3485 ( 
.A(n_3404),
.B(n_3069),
.Y(n_3485)
);

AOI21xp5_ASAP7_75t_L g3486 ( 
.A1(n_3423),
.A2(n_3097),
.B(n_3220),
.Y(n_3486)
);

AO21x2_ASAP7_75t_L g3487 ( 
.A1(n_3335),
.A2(n_3094),
.B(n_3079),
.Y(n_3487)
);

BUFx3_ASAP7_75t_L g3488 ( 
.A(n_3395),
.Y(n_3488)
);

INVx2_ASAP7_75t_L g3489 ( 
.A(n_3374),
.Y(n_3489)
);

A2O1A1Ixp33_ASAP7_75t_L g3490 ( 
.A1(n_3423),
.A2(n_3217),
.B(n_3112),
.C(n_3055),
.Y(n_3490)
);

OA21x2_ASAP7_75t_L g3491 ( 
.A1(n_3405),
.A2(n_3042),
.B(n_3052),
.Y(n_3491)
);

AOI221xp5_ASAP7_75t_L g3492 ( 
.A1(n_3401),
.A2(n_3217),
.B1(n_3304),
.B2(n_3069),
.C(n_3075),
.Y(n_3492)
);

HB1xp67_ASAP7_75t_L g3493 ( 
.A(n_3318),
.Y(n_3493)
);

HB1xp67_ASAP7_75t_L g3494 ( 
.A(n_3330),
.Y(n_3494)
);

AO21x2_ASAP7_75t_L g3495 ( 
.A1(n_3338),
.A2(n_3075),
.B(n_3092),
.Y(n_3495)
);

AND2x6_ASAP7_75t_L g3496 ( 
.A(n_3380),
.B(n_3078),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3320),
.Y(n_3497)
);

INVx2_ASAP7_75t_L g3498 ( 
.A(n_3374),
.Y(n_3498)
);

INVx3_ASAP7_75t_L g3499 ( 
.A(n_3336),
.Y(n_3499)
);

AND2x2_ASAP7_75t_L g3500 ( 
.A(n_3399),
.B(n_3092),
.Y(n_3500)
);

AOI21xp33_ASAP7_75t_L g3501 ( 
.A1(n_3401),
.A2(n_3236),
.B(n_3259),
.Y(n_3501)
);

OAI22xp5_ASAP7_75t_L g3502 ( 
.A1(n_3376),
.A2(n_3242),
.B1(n_3236),
.B2(n_3228),
.Y(n_3502)
);

OA21x2_ASAP7_75t_L g3503 ( 
.A1(n_3398),
.A2(n_3127),
.B(n_3233),
.Y(n_3503)
);

INVx2_ASAP7_75t_SL g3504 ( 
.A(n_3321),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_3327),
.Y(n_3505)
);

INVx2_ASAP7_75t_L g3506 ( 
.A(n_3346),
.Y(n_3506)
);

INVx2_ASAP7_75t_L g3507 ( 
.A(n_3346),
.Y(n_3507)
);

HB1xp67_ASAP7_75t_L g3508 ( 
.A(n_3330),
.Y(n_3508)
);

AOI211xp5_ASAP7_75t_L g3509 ( 
.A1(n_3430),
.A2(n_2987),
.B(n_146),
.C(n_142),
.Y(n_3509)
);

AND2x2_ASAP7_75t_L g3510 ( 
.A(n_3399),
.B(n_3233),
.Y(n_3510)
);

OAI221xp5_ASAP7_75t_L g3511 ( 
.A1(n_3319),
.A2(n_3309),
.B1(n_3226),
.B2(n_3223),
.C(n_3147),
.Y(n_3511)
);

BUFx3_ASAP7_75t_L g3512 ( 
.A(n_3395),
.Y(n_3512)
);

INVx4_ASAP7_75t_R g3513 ( 
.A(n_3410),
.Y(n_3513)
);

NAND4xp25_ASAP7_75t_L g3514 ( 
.A(n_3440),
.B(n_3223),
.C(n_147),
.D(n_144),
.Y(n_3514)
);

OAI21xp5_ASAP7_75t_L g3515 ( 
.A1(n_3430),
.A2(n_3120),
.B(n_3125),
.Y(n_3515)
);

HB1xp67_ASAP7_75t_L g3516 ( 
.A(n_3330),
.Y(n_3516)
);

AND2x4_ASAP7_75t_L g3517 ( 
.A(n_3400),
.B(n_3089),
.Y(n_3517)
);

INVx2_ASAP7_75t_L g3518 ( 
.A(n_3346),
.Y(n_3518)
);

BUFx3_ASAP7_75t_L g3519 ( 
.A(n_3395),
.Y(n_3519)
);

INVx2_ASAP7_75t_L g3520 ( 
.A(n_3351),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_3420),
.B(n_146),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3327),
.Y(n_3522)
);

INVx2_ASAP7_75t_L g3523 ( 
.A(n_3351),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3329),
.Y(n_3524)
);

NOR2xp33_ASAP7_75t_L g3525 ( 
.A(n_3440),
.B(n_149),
.Y(n_3525)
);

INVx2_ASAP7_75t_L g3526 ( 
.A(n_3351),
.Y(n_3526)
);

NAND3xp33_ASAP7_75t_L g3527 ( 
.A(n_3430),
.B(n_150),
.C(n_151),
.Y(n_3527)
);

INVx3_ASAP7_75t_L g3528 ( 
.A(n_3336),
.Y(n_3528)
);

AOI21xp5_ASAP7_75t_L g3529 ( 
.A1(n_3420),
.A2(n_150),
.B(n_151),
.Y(n_3529)
);

AOI221xp5_ASAP7_75t_L g3530 ( 
.A1(n_3428),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.C(n_155),
.Y(n_3530)
);

OAI21xp5_ASAP7_75t_L g3531 ( 
.A1(n_3428),
.A2(n_154),
.B(n_156),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3329),
.Y(n_3532)
);

AOI222xp33_ASAP7_75t_L g3533 ( 
.A1(n_3442),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.C1(n_160),
.C2(n_161),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3337),
.Y(n_3534)
);

BUFx2_ASAP7_75t_L g3535 ( 
.A(n_3336),
.Y(n_3535)
);

OAI21x1_ASAP7_75t_L g3536 ( 
.A1(n_3400),
.A2(n_158),
.B(n_160),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3337),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_3342),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3387),
.B(n_161),
.Y(n_3539)
);

HB1xp67_ASAP7_75t_L g3540 ( 
.A(n_3332),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3342),
.Y(n_3541)
);

OA21x2_ASAP7_75t_L g3542 ( 
.A1(n_3398),
.A2(n_162),
.B(n_163),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_3344),
.Y(n_3543)
);

OAI21x1_ASAP7_75t_L g3544 ( 
.A1(n_3400),
.A2(n_163),
.B(n_164),
.Y(n_3544)
);

AOI21xp5_ASAP7_75t_L g3545 ( 
.A1(n_3411),
.A2(n_164),
.B(n_165),
.Y(n_3545)
);

INVx2_ASAP7_75t_L g3546 ( 
.A(n_3315),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3344),
.Y(n_3547)
);

AOI211xp5_ASAP7_75t_L g3548 ( 
.A1(n_3436),
.A2(n_166),
.B(n_168),
.C(n_169),
.Y(n_3548)
);

AOI22xp33_ASAP7_75t_L g3549 ( 
.A1(n_3442),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_3549)
);

AND2x2_ASAP7_75t_L g3550 ( 
.A(n_3400),
.B(n_171),
.Y(n_3550)
);

AOI21xp5_ASAP7_75t_L g3551 ( 
.A1(n_3411),
.A2(n_172),
.B(n_173),
.Y(n_3551)
);

INVx2_ASAP7_75t_SL g3552 ( 
.A(n_3321),
.Y(n_3552)
);

INVx4_ASAP7_75t_L g3553 ( 
.A(n_3433),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_3387),
.B(n_175),
.Y(n_3554)
);

OAI211xp5_ASAP7_75t_L g3555 ( 
.A1(n_3428),
.A2(n_175),
.B(n_176),
.C(n_177),
.Y(n_3555)
);

INVx1_ASAP7_75t_L g3556 ( 
.A(n_3349),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3349),
.Y(n_3557)
);

AOI22xp33_ASAP7_75t_L g3558 ( 
.A1(n_3442),
.A2(n_176),
.B1(n_177),
.B2(n_179),
.Y(n_3558)
);

AND2x2_ASAP7_75t_L g3559 ( 
.A(n_3365),
.B(n_180),
.Y(n_3559)
);

INVx2_ASAP7_75t_L g3560 ( 
.A(n_3315),
.Y(n_3560)
);

INVx2_ASAP7_75t_SL g3561 ( 
.A(n_3426),
.Y(n_3561)
);

AOI22xp5_ASAP7_75t_L g3562 ( 
.A1(n_3434),
.A2(n_180),
.B1(n_181),
.B2(n_183),
.Y(n_3562)
);

AOI22xp5_ASAP7_75t_L g3563 ( 
.A1(n_3427),
.A2(n_3431),
.B1(n_3414),
.B2(n_3419),
.Y(n_3563)
);

INVx2_ASAP7_75t_L g3564 ( 
.A(n_3339),
.Y(n_3564)
);

AND2x2_ASAP7_75t_L g3565 ( 
.A(n_3365),
.B(n_184),
.Y(n_3565)
);

OAI21xp5_ASAP7_75t_L g3566 ( 
.A1(n_3411),
.A2(n_184),
.B(n_186),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3353),
.Y(n_3567)
);

AND2x4_ASAP7_75t_L g3568 ( 
.A(n_3383),
.B(n_187),
.Y(n_3568)
);

NOR2xp33_ASAP7_75t_L g3569 ( 
.A(n_3463),
.B(n_3433),
.Y(n_3569)
);

AND2x2_ASAP7_75t_L g3570 ( 
.A(n_3553),
.B(n_3328),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3446),
.Y(n_3571)
);

AND2x2_ASAP7_75t_L g3572 ( 
.A(n_3553),
.B(n_3328),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3469),
.B(n_3380),
.Y(n_3573)
);

INVx4_ASAP7_75t_L g3574 ( 
.A(n_3463),
.Y(n_3574)
);

INVxp67_ASAP7_75t_L g3575 ( 
.A(n_3466),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3446),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_3563),
.B(n_3380),
.Y(n_3577)
);

OAI22xp5_ASAP7_75t_L g3578 ( 
.A1(n_3447),
.A2(n_3415),
.B1(n_3424),
.B2(n_3431),
.Y(n_3578)
);

INVx2_ASAP7_75t_L g3579 ( 
.A(n_3479),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3480),
.B(n_3388),
.Y(n_3580)
);

HB1xp67_ASAP7_75t_L g3581 ( 
.A(n_3479),
.Y(n_3581)
);

INVx2_ASAP7_75t_L g3582 ( 
.A(n_3493),
.Y(n_3582)
);

OAI33xp33_ASAP7_75t_L g3583 ( 
.A1(n_3470),
.A2(n_3332),
.A3(n_3334),
.B1(n_3338),
.B2(n_3388),
.B3(n_3419),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3493),
.Y(n_3584)
);

OAI21xp33_ASAP7_75t_L g3585 ( 
.A1(n_3447),
.A2(n_3436),
.B(n_3417),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3494),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3494),
.Y(n_3587)
);

NOR2xp33_ASAP7_75t_R g3588 ( 
.A(n_3463),
.B(n_3410),
.Y(n_3588)
);

INVx2_ASAP7_75t_L g3589 ( 
.A(n_3508),
.Y(n_3589)
);

INVx2_ASAP7_75t_L g3590 ( 
.A(n_3508),
.Y(n_3590)
);

HB1xp67_ASAP7_75t_L g3591 ( 
.A(n_3516),
.Y(n_3591)
);

AND2x2_ASAP7_75t_L g3592 ( 
.A(n_3504),
.B(n_3328),
.Y(n_3592)
);

AND2x4_ASAP7_75t_L g3593 ( 
.A(n_3552),
.B(n_3336),
.Y(n_3593)
);

AO21x2_ASAP7_75t_L g3594 ( 
.A1(n_3455),
.A2(n_3338),
.B(n_3334),
.Y(n_3594)
);

AND2x2_ASAP7_75t_L g3595 ( 
.A(n_3484),
.B(n_3313),
.Y(n_3595)
);

NOR2x1_ASAP7_75t_SL g3596 ( 
.A(n_3487),
.B(n_3343),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_3516),
.Y(n_3597)
);

AND2x2_ASAP7_75t_L g3598 ( 
.A(n_3564),
.B(n_3313),
.Y(n_3598)
);

AND2x2_ASAP7_75t_L g3599 ( 
.A(n_3443),
.B(n_3448),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_3540),
.Y(n_3600)
);

AND2x2_ASAP7_75t_L g3601 ( 
.A(n_3443),
.B(n_3448),
.Y(n_3601)
);

INVx2_ASAP7_75t_L g3602 ( 
.A(n_3540),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_3468),
.Y(n_3603)
);

HB1xp67_ASAP7_75t_L g3604 ( 
.A(n_3542),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_L g3605 ( 
.A(n_3550),
.B(n_3414),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3481),
.Y(n_3606)
);

AO21x2_ASAP7_75t_L g3607 ( 
.A1(n_3455),
.A2(n_3334),
.B(n_3332),
.Y(n_3607)
);

AND2x2_ASAP7_75t_L g3608 ( 
.A(n_3459),
.B(n_3326),
.Y(n_3608)
);

AND2x2_ASAP7_75t_L g3609 ( 
.A(n_3458),
.B(n_3326),
.Y(n_3609)
);

OAI21xp33_ASAP7_75t_L g3610 ( 
.A1(n_3460),
.A2(n_3436),
.B(n_3417),
.Y(n_3610)
);

HB1xp67_ASAP7_75t_L g3611 ( 
.A(n_3542),
.Y(n_3611)
);

BUFx3_ASAP7_75t_L g3612 ( 
.A(n_3471),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_3482),
.Y(n_3613)
);

AND2x4_ASAP7_75t_L g3614 ( 
.A(n_3499),
.B(n_3383),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3497),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3505),
.Y(n_3616)
);

HB1xp67_ASAP7_75t_L g3617 ( 
.A(n_3542),
.Y(n_3617)
);

AND2x2_ASAP7_75t_L g3618 ( 
.A(n_3457),
.B(n_3431),
.Y(n_3618)
);

INVx2_ASAP7_75t_L g3619 ( 
.A(n_3488),
.Y(n_3619)
);

INVx3_ASAP7_75t_L g3620 ( 
.A(n_3463),
.Y(n_3620)
);

NAND3xp33_ASAP7_75t_L g3621 ( 
.A(n_3509),
.B(n_3393),
.C(n_3437),
.Y(n_3621)
);

AND2x4_ASAP7_75t_L g3622 ( 
.A(n_3499),
.B(n_3383),
.Y(n_3622)
);

INVx2_ASAP7_75t_L g3623 ( 
.A(n_3488),
.Y(n_3623)
);

AND2x2_ASAP7_75t_L g3624 ( 
.A(n_3454),
.B(n_3510),
.Y(n_3624)
);

NOR2xp33_ASAP7_75t_L g3625 ( 
.A(n_3471),
.B(n_3433),
.Y(n_3625)
);

BUFx3_ASAP7_75t_L g3626 ( 
.A(n_3477),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3522),
.Y(n_3627)
);

HB1xp67_ASAP7_75t_L g3628 ( 
.A(n_3512),
.Y(n_3628)
);

INVx2_ASAP7_75t_L g3629 ( 
.A(n_3512),
.Y(n_3629)
);

INVx1_ASAP7_75t_L g3630 ( 
.A(n_3524),
.Y(n_3630)
);

NAND3xp33_ASAP7_75t_L g3631 ( 
.A(n_3444),
.B(n_3393),
.C(n_3437),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3532),
.Y(n_3632)
);

INVx3_ASAP7_75t_L g3633 ( 
.A(n_3519),
.Y(n_3633)
);

AO21x2_ASAP7_75t_L g3634 ( 
.A1(n_3527),
.A2(n_3406),
.B(n_3314),
.Y(n_3634)
);

INVx2_ASAP7_75t_L g3635 ( 
.A(n_3519),
.Y(n_3635)
);

INVxp67_ASAP7_75t_L g3636 ( 
.A(n_3452),
.Y(n_3636)
);

AND2x2_ASAP7_75t_L g3637 ( 
.A(n_3454),
.B(n_3389),
.Y(n_3637)
);

AND2x2_ASAP7_75t_L g3638 ( 
.A(n_3500),
.B(n_3389),
.Y(n_3638)
);

CKINVDCx16_ASAP7_75t_R g3639 ( 
.A(n_3477),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3534),
.Y(n_3640)
);

AND2x2_ASAP7_75t_L g3641 ( 
.A(n_3535),
.B(n_3390),
.Y(n_3641)
);

INVx1_ASAP7_75t_L g3642 ( 
.A(n_3537),
.Y(n_3642)
);

AND2x2_ASAP7_75t_L g3643 ( 
.A(n_3561),
.B(n_3390),
.Y(n_3643)
);

OR2x2_ASAP7_75t_L g3644 ( 
.A(n_3485),
.B(n_3323),
.Y(n_3644)
);

AOI22xp33_ASAP7_75t_L g3645 ( 
.A1(n_3472),
.A2(n_3429),
.B1(n_3441),
.B2(n_3437),
.Y(n_3645)
);

NAND2xp5_ASAP7_75t_L g3646 ( 
.A(n_3449),
.B(n_3427),
.Y(n_3646)
);

OR2x2_ASAP7_75t_L g3647 ( 
.A(n_3453),
.B(n_3360),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3538),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_3541),
.Y(n_3649)
);

OAI31xp33_ASAP7_75t_L g3650 ( 
.A1(n_3461),
.A2(n_3449),
.A3(n_3451),
.B(n_3490),
.Y(n_3650)
);

AND2x2_ASAP7_75t_L g3651 ( 
.A(n_3546),
.B(n_3391),
.Y(n_3651)
);

INVxp67_ASAP7_75t_SL g3652 ( 
.A(n_3452),
.Y(n_3652)
);

OAI22xp5_ASAP7_75t_L g3653 ( 
.A1(n_3462),
.A2(n_3415),
.B1(n_3424),
.B2(n_3325),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_L g3654 ( 
.A(n_3486),
.B(n_3397),
.Y(n_3654)
);

INVx3_ASAP7_75t_L g3655 ( 
.A(n_3528),
.Y(n_3655)
);

AND2x2_ASAP7_75t_L g3656 ( 
.A(n_3546),
.B(n_3560),
.Y(n_3656)
);

OR2x2_ASAP7_75t_L g3657 ( 
.A(n_3465),
.B(n_3360),
.Y(n_3657)
);

INVx1_ASAP7_75t_L g3658 ( 
.A(n_3543),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_3547),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3548),
.B(n_3397),
.Y(n_3660)
);

INVx1_ASAP7_75t_L g3661 ( 
.A(n_3556),
.Y(n_3661)
);

NOR2xp33_ASAP7_75t_L g3662 ( 
.A(n_3473),
.B(n_3433),
.Y(n_3662)
);

AOI22xp33_ASAP7_75t_L g3663 ( 
.A1(n_3472),
.A2(n_3429),
.B1(n_3441),
.B2(n_3406),
.Y(n_3663)
);

INVx5_ASAP7_75t_L g3664 ( 
.A(n_3528),
.Y(n_3664)
);

INVx5_ASAP7_75t_L g3665 ( 
.A(n_3496),
.Y(n_3665)
);

HB1xp67_ASAP7_75t_L g3666 ( 
.A(n_3445),
.Y(n_3666)
);

NAND2xp5_ASAP7_75t_L g3667 ( 
.A(n_3478),
.B(n_3415),
.Y(n_3667)
);

A2O1A1Ixp33_ASAP7_75t_SL g3668 ( 
.A1(n_3531),
.A2(n_3441),
.B(n_3413),
.C(n_3406),
.Y(n_3668)
);

AOI221xp5_ASAP7_75t_L g3669 ( 
.A1(n_3464),
.A2(n_3429),
.B1(n_3357),
.B2(n_3432),
.C(n_3331),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_L g3670 ( 
.A(n_3521),
.B(n_3559),
.Y(n_3670)
);

AOI31xp33_ASAP7_75t_L g3671 ( 
.A1(n_3462),
.A2(n_3410),
.A3(n_3424),
.B(n_3325),
.Y(n_3671)
);

AND2x2_ASAP7_75t_L g3672 ( 
.A(n_3560),
.B(n_3391),
.Y(n_3672)
);

INVx2_ASAP7_75t_L g3673 ( 
.A(n_3456),
.Y(n_3673)
);

INVx4_ASAP7_75t_L g3674 ( 
.A(n_3568),
.Y(n_3674)
);

OR2x2_ASAP7_75t_L g3675 ( 
.A(n_3465),
.B(n_3394),
.Y(n_3675)
);

NAND3xp33_ASAP7_75t_L g3676 ( 
.A(n_3490),
.B(n_3432),
.C(n_3413),
.Y(n_3676)
);

INVx2_ASAP7_75t_L g3677 ( 
.A(n_3456),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3557),
.Y(n_3678)
);

INVx3_ASAP7_75t_L g3679 ( 
.A(n_3496),
.Y(n_3679)
);

BUFx2_ASAP7_75t_L g3680 ( 
.A(n_3568),
.Y(n_3680)
);

INVx2_ASAP7_75t_L g3681 ( 
.A(n_3489),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_3567),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3450),
.Y(n_3683)
);

AND2x2_ASAP7_75t_L g3684 ( 
.A(n_3624),
.B(n_3475),
.Y(n_3684)
);

OR2x2_ASAP7_75t_L g3685 ( 
.A(n_3644),
.B(n_3489),
.Y(n_3685)
);

HB1xp67_ASAP7_75t_L g3686 ( 
.A(n_3680),
.Y(n_3686)
);

AND2x4_ASAP7_75t_L g3687 ( 
.A(n_3612),
.B(n_3483),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_L g3688 ( 
.A(n_3618),
.B(n_3525),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_3581),
.Y(n_3689)
);

NAND2xp5_ASAP7_75t_L g3690 ( 
.A(n_3652),
.B(n_3525),
.Y(n_3690)
);

AND2x2_ASAP7_75t_L g3691 ( 
.A(n_3624),
.B(n_3475),
.Y(n_3691)
);

BUFx2_ASAP7_75t_L g3692 ( 
.A(n_3588),
.Y(n_3692)
);

OAI21xp33_ASAP7_75t_L g3693 ( 
.A1(n_3585),
.A2(n_3461),
.B(n_3451),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3591),
.Y(n_3694)
);

AND2x2_ASAP7_75t_L g3695 ( 
.A(n_3639),
.B(n_3381),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3579),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3579),
.Y(n_3697)
);

INVx2_ASAP7_75t_L g3698 ( 
.A(n_3607),
.Y(n_3698)
);

NAND2xp33_ASAP7_75t_R g3699 ( 
.A(n_3588),
.B(n_3633),
.Y(n_3699)
);

NAND4xp25_ASAP7_75t_L g3700 ( 
.A(n_3650),
.B(n_3467),
.C(n_3530),
.D(n_3514),
.Y(n_3700)
);

INVx4_ASAP7_75t_L g3701 ( 
.A(n_3574),
.Y(n_3701)
);

INVx1_ASAP7_75t_L g3702 ( 
.A(n_3582),
.Y(n_3702)
);

INVx2_ASAP7_75t_L g3703 ( 
.A(n_3607),
.Y(n_3703)
);

HB1xp67_ASAP7_75t_L g3704 ( 
.A(n_3628),
.Y(n_3704)
);

AND2x2_ASAP7_75t_L g3705 ( 
.A(n_3608),
.B(n_3381),
.Y(n_3705)
);

NAND3x1_ASAP7_75t_L g3706 ( 
.A(n_3646),
.B(n_3529),
.C(n_3467),
.Y(n_3706)
);

NAND2xp5_ASAP7_75t_L g3707 ( 
.A(n_3578),
.B(n_3539),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_3671),
.B(n_3554),
.Y(n_3708)
);

AND2x2_ASAP7_75t_L g3709 ( 
.A(n_3608),
.B(n_3381),
.Y(n_3709)
);

OR2x2_ASAP7_75t_L g3710 ( 
.A(n_3657),
.B(n_3498),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3582),
.Y(n_3711)
);

AND2x2_ASAP7_75t_L g3712 ( 
.A(n_3609),
.B(n_3425),
.Y(n_3712)
);

INVx2_ASAP7_75t_L g3713 ( 
.A(n_3594),
.Y(n_3713)
);

NOR2xp67_ASAP7_75t_L g3714 ( 
.A(n_3674),
.B(n_3343),
.Y(n_3714)
);

AND2x2_ASAP7_75t_L g3715 ( 
.A(n_3609),
.B(n_3425),
.Y(n_3715)
);

AND2x2_ASAP7_75t_L g3716 ( 
.A(n_3637),
.B(n_3599),
.Y(n_3716)
);

AND2x2_ASAP7_75t_L g3717 ( 
.A(n_3599),
.B(n_3425),
.Y(n_3717)
);

NAND2xp33_ASAP7_75t_R g3718 ( 
.A(n_3633),
.B(n_3465),
.Y(n_3718)
);

AND2x2_ASAP7_75t_L g3719 ( 
.A(n_3601),
.B(n_3515),
.Y(n_3719)
);

INVx2_ASAP7_75t_L g3720 ( 
.A(n_3594),
.Y(n_3720)
);

AND2x2_ASAP7_75t_L g3721 ( 
.A(n_3601),
.B(n_3331),
.Y(n_3721)
);

AND2x4_ASAP7_75t_L g3722 ( 
.A(n_3612),
.B(n_3506),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_3589),
.Y(n_3723)
);

INVxp67_ASAP7_75t_L g3724 ( 
.A(n_3626),
.Y(n_3724)
);

NAND2xp5_ASAP7_75t_L g3725 ( 
.A(n_3636),
.B(n_3575),
.Y(n_3725)
);

NAND2xp5_ASAP7_75t_L g3726 ( 
.A(n_3674),
.B(n_3565),
.Y(n_3726)
);

AND2x2_ASAP7_75t_L g3727 ( 
.A(n_3626),
.B(n_3593),
.Y(n_3727)
);

AND2x2_ASAP7_75t_L g3728 ( 
.A(n_3593),
.B(n_3331),
.Y(n_3728)
);

AND2x2_ASAP7_75t_L g3729 ( 
.A(n_3593),
.B(n_3331),
.Y(n_3729)
);

HB1xp67_ASAP7_75t_L g3730 ( 
.A(n_3589),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_L g3731 ( 
.A(n_3674),
.B(n_3545),
.Y(n_3731)
);

AND2x2_ASAP7_75t_L g3732 ( 
.A(n_3592),
.B(n_3343),
.Y(n_3732)
);

AND2x4_ASAP7_75t_L g3733 ( 
.A(n_3620),
.B(n_3506),
.Y(n_3733)
);

AND2x4_ASAP7_75t_L g3734 ( 
.A(n_3620),
.B(n_3507),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_3590),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3590),
.Y(n_3736)
);

AND2x2_ASAP7_75t_L g3737 ( 
.A(n_3592),
.B(n_3347),
.Y(n_3737)
);

AND2x2_ASAP7_75t_L g3738 ( 
.A(n_3633),
.B(n_3347),
.Y(n_3738)
);

NAND2xp5_ASAP7_75t_L g3739 ( 
.A(n_3653),
.B(n_3551),
.Y(n_3739)
);

INVx4_ASAP7_75t_L g3740 ( 
.A(n_3574),
.Y(n_3740)
);

INVx2_ASAP7_75t_L g3741 ( 
.A(n_3620),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3602),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3602),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3571),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3576),
.Y(n_3745)
);

HB1xp67_ASAP7_75t_L g3746 ( 
.A(n_3604),
.Y(n_3746)
);

AND2x2_ASAP7_75t_L g3747 ( 
.A(n_3638),
.B(n_3347),
.Y(n_3747)
);

INVx2_ASAP7_75t_L g3748 ( 
.A(n_3574),
.Y(n_3748)
);

INVx2_ASAP7_75t_L g3749 ( 
.A(n_3664),
.Y(n_3749)
);

AND2x2_ASAP7_75t_L g3750 ( 
.A(n_3638),
.B(n_3409),
.Y(n_3750)
);

AND2x2_ASAP7_75t_L g3751 ( 
.A(n_3619),
.B(n_3409),
.Y(n_3751)
);

BUFx2_ASAP7_75t_L g3752 ( 
.A(n_3634),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3584),
.Y(n_3753)
);

INVx2_ASAP7_75t_L g3754 ( 
.A(n_3664),
.Y(n_3754)
);

OR2x2_ASAP7_75t_L g3755 ( 
.A(n_3647),
.B(n_3498),
.Y(n_3755)
);

AND2x2_ASAP7_75t_L g3756 ( 
.A(n_3619),
.B(n_3409),
.Y(n_3756)
);

AND2x2_ASAP7_75t_L g3757 ( 
.A(n_3623),
.B(n_3409),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_L g3758 ( 
.A(n_3573),
.B(n_3562),
.Y(n_3758)
);

AOI22xp33_ASAP7_75t_L g3759 ( 
.A1(n_3621),
.A2(n_3476),
.B1(n_3502),
.B2(n_3501),
.Y(n_3759)
);

INVx2_ASAP7_75t_L g3760 ( 
.A(n_3664),
.Y(n_3760)
);

AND2x2_ASAP7_75t_L g3761 ( 
.A(n_3623),
.B(n_3517),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3586),
.Y(n_3762)
);

OR2x2_ASAP7_75t_L g3763 ( 
.A(n_3675),
.B(n_3507),
.Y(n_3763)
);

INVx2_ASAP7_75t_L g3764 ( 
.A(n_3664),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_3587),
.Y(n_3765)
);

NAND5xp2_ASAP7_75t_L g3766 ( 
.A(n_3645),
.B(n_3533),
.C(n_3474),
.D(n_3555),
.E(n_3566),
.Y(n_3766)
);

HB1xp67_ASAP7_75t_L g3767 ( 
.A(n_3611),
.Y(n_3767)
);

AND2x2_ASAP7_75t_L g3768 ( 
.A(n_3629),
.B(n_3517),
.Y(n_3768)
);

AND2x2_ASAP7_75t_SL g3769 ( 
.A(n_3663),
.B(n_3549),
.Y(n_3769)
);

OR2x2_ASAP7_75t_L g3770 ( 
.A(n_3634),
.B(n_3518),
.Y(n_3770)
);

AND2x2_ASAP7_75t_L g3771 ( 
.A(n_3629),
.B(n_3432),
.Y(n_3771)
);

INVx2_ASAP7_75t_L g3772 ( 
.A(n_3664),
.Y(n_3772)
);

OR2x2_ASAP7_75t_L g3773 ( 
.A(n_3580),
.B(n_3518),
.Y(n_3773)
);

NOR4xp25_ASAP7_75t_SL g3774 ( 
.A(n_3669),
.B(n_3610),
.C(n_3600),
.D(n_3597),
.Y(n_3774)
);

INVx2_ASAP7_75t_L g3775 ( 
.A(n_3655),
.Y(n_3775)
);

OR2x2_ASAP7_75t_L g3776 ( 
.A(n_3666),
.B(n_3520),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3686),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3730),
.Y(n_3778)
);

AND2x2_ASAP7_75t_L g3779 ( 
.A(n_3716),
.B(n_3625),
.Y(n_3779)
);

OR2x2_ASAP7_75t_L g3780 ( 
.A(n_3688),
.B(n_3667),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3704),
.Y(n_3781)
);

XNOR2x2_ASAP7_75t_L g3782 ( 
.A(n_3700),
.B(n_3631),
.Y(n_3782)
);

INVx2_ASAP7_75t_L g3783 ( 
.A(n_3716),
.Y(n_3783)
);

INVxp67_ASAP7_75t_L g3784 ( 
.A(n_3699),
.Y(n_3784)
);

NOR2x1_ASAP7_75t_L g3785 ( 
.A(n_3752),
.B(n_3676),
.Y(n_3785)
);

NOR2x1_ASAP7_75t_L g3786 ( 
.A(n_3752),
.B(n_3569),
.Y(n_3786)
);

INVx1_ASAP7_75t_SL g3787 ( 
.A(n_3692),
.Y(n_3787)
);

NOR3xp33_ASAP7_75t_L g3788 ( 
.A(n_3693),
.B(n_3583),
.C(n_3569),
.Y(n_3788)
);

INVx2_ASAP7_75t_L g3789 ( 
.A(n_3687),
.Y(n_3789)
);

INVx2_ASAP7_75t_SL g3790 ( 
.A(n_3727),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_3746),
.Y(n_3791)
);

INVx3_ASAP7_75t_SL g3792 ( 
.A(n_3687),
.Y(n_3792)
);

AOI22xp5_ASAP7_75t_L g3793 ( 
.A1(n_3706),
.A2(n_3660),
.B1(n_3663),
.B2(n_3645),
.Y(n_3793)
);

XNOR2xp5_ASAP7_75t_L g3794 ( 
.A(n_3706),
.B(n_3605),
.Y(n_3794)
);

INVx1_ASAP7_75t_SL g3795 ( 
.A(n_3692),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_L g3796 ( 
.A(n_3769),
.B(n_3635),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_3767),
.Y(n_3797)
);

NAND2xp5_ASAP7_75t_L g3798 ( 
.A(n_3769),
.B(n_3635),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_L g3799 ( 
.A(n_3759),
.B(n_3668),
.Y(n_3799)
);

NAND4xp75_ASAP7_75t_L g3800 ( 
.A(n_3714),
.B(n_3654),
.C(n_3570),
.D(n_3572),
.Y(n_3800)
);

INVx1_ASAP7_75t_L g3801 ( 
.A(n_3689),
.Y(n_3801)
);

AND2x2_ASAP7_75t_L g3802 ( 
.A(n_3687),
.B(n_3684),
.Y(n_3802)
);

INVx2_ASAP7_75t_L g3803 ( 
.A(n_3701),
.Y(n_3803)
);

OAI22xp5_ASAP7_75t_SL g3804 ( 
.A1(n_3758),
.A2(n_3392),
.B1(n_3558),
.B2(n_3549),
.Y(n_3804)
);

AND2x2_ASAP7_75t_L g3805 ( 
.A(n_3684),
.B(n_3625),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_3689),
.Y(n_3806)
);

NAND2xp5_ASAP7_75t_L g3807 ( 
.A(n_3694),
.B(n_3668),
.Y(n_3807)
);

INVx1_ASAP7_75t_L g3808 ( 
.A(n_3694),
.Y(n_3808)
);

AND2x2_ASAP7_75t_L g3809 ( 
.A(n_3691),
.B(n_3662),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_L g3810 ( 
.A(n_3724),
.B(n_3577),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_L g3811 ( 
.A(n_3727),
.B(n_3670),
.Y(n_3811)
);

NAND4xp75_ASAP7_75t_L g3812 ( 
.A(n_3774),
.B(n_3738),
.C(n_3739),
.D(n_3708),
.Y(n_3812)
);

INVx1_ASAP7_75t_SL g3813 ( 
.A(n_3738),
.Y(n_3813)
);

NAND4xp75_ASAP7_75t_SL g3814 ( 
.A(n_3695),
.B(n_3747),
.C(n_3719),
.D(n_3570),
.Y(n_3814)
);

AND2x2_ASAP7_75t_L g3815 ( 
.A(n_3691),
.B(n_3662),
.Y(n_3815)
);

INVx1_ASAP7_75t_L g3816 ( 
.A(n_3696),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3696),
.Y(n_3817)
);

INVx1_ASAP7_75t_L g3818 ( 
.A(n_3697),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3697),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_3690),
.B(n_3641),
.Y(n_3820)
);

AND2x2_ASAP7_75t_L g3821 ( 
.A(n_3695),
.B(n_3643),
.Y(n_3821)
);

AND2x2_ASAP7_75t_L g3822 ( 
.A(n_3747),
.B(n_3643),
.Y(n_3822)
);

OAI21xp33_ASAP7_75t_L g3823 ( 
.A1(n_3766),
.A2(n_3558),
.B(n_3617),
.Y(n_3823)
);

INVx1_ASAP7_75t_L g3824 ( 
.A(n_3702),
.Y(n_3824)
);

INVx2_ASAP7_75t_L g3825 ( 
.A(n_3701),
.Y(n_3825)
);

INVx2_ASAP7_75t_L g3826 ( 
.A(n_3701),
.Y(n_3826)
);

NAND4xp75_ASAP7_75t_SL g3827 ( 
.A(n_3719),
.B(n_3572),
.C(n_3598),
.D(n_3595),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3702),
.Y(n_3828)
);

INVx2_ASAP7_75t_L g3829 ( 
.A(n_3740),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_L g3830 ( 
.A(n_3748),
.B(n_3641),
.Y(n_3830)
);

INVxp67_ASAP7_75t_L g3831 ( 
.A(n_3718),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_L g3832 ( 
.A(n_3748),
.B(n_3683),
.Y(n_3832)
);

INVx1_ASAP7_75t_SL g3833 ( 
.A(n_3722),
.Y(n_3833)
);

BUFx3_ASAP7_75t_L g3834 ( 
.A(n_3726),
.Y(n_3834)
);

CKINVDCx14_ASAP7_75t_R g3835 ( 
.A(n_3725),
.Y(n_3835)
);

INVxp67_ASAP7_75t_SL g3836 ( 
.A(n_3749),
.Y(n_3836)
);

NOR3xp33_ASAP7_75t_SL g3837 ( 
.A(n_3707),
.B(n_3606),
.C(n_3603),
.Y(n_3837)
);

INVx2_ASAP7_75t_L g3838 ( 
.A(n_3740),
.Y(n_3838)
);

XOR2x2_ASAP7_75t_L g3839 ( 
.A(n_3731),
.B(n_3596),
.Y(n_3839)
);

XOR2x2_ASAP7_75t_L g3840 ( 
.A(n_3732),
.B(n_3426),
.Y(n_3840)
);

INVx3_ASAP7_75t_L g3841 ( 
.A(n_3740),
.Y(n_3841)
);

NAND4xp75_ASAP7_75t_L g3842 ( 
.A(n_3698),
.B(n_3595),
.C(n_3598),
.D(n_3656),
.Y(n_3842)
);

NAND4xp75_ASAP7_75t_L g3843 ( 
.A(n_3698),
.B(n_3656),
.C(n_3677),
.D(n_3673),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3711),
.Y(n_3844)
);

INVx2_ASAP7_75t_L g3845 ( 
.A(n_3775),
.Y(n_3845)
);

NOR4xp25_ASAP7_75t_L g3846 ( 
.A(n_3703),
.B(n_3613),
.C(n_3616),
.D(n_3615),
.Y(n_3846)
);

NAND4xp75_ASAP7_75t_SL g3847 ( 
.A(n_3732),
.B(n_3491),
.C(n_3503),
.D(n_3408),
.Y(n_3847)
);

INVx2_ASAP7_75t_L g3848 ( 
.A(n_3775),
.Y(n_3848)
);

BUFx6f_ASAP7_75t_L g3849 ( 
.A(n_3749),
.Y(n_3849)
);

INVx4_ASAP7_75t_L g3850 ( 
.A(n_3754),
.Y(n_3850)
);

OAI22xp5_ASAP7_75t_L g3851 ( 
.A1(n_3703),
.A2(n_3413),
.B1(n_3408),
.B2(n_3492),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_3711),
.Y(n_3852)
);

HB1xp67_ASAP7_75t_L g3853 ( 
.A(n_3754),
.Y(n_3853)
);

INVx2_ASAP7_75t_L g3854 ( 
.A(n_3760),
.Y(n_3854)
);

NAND4xp25_ASAP7_75t_L g3855 ( 
.A(n_3744),
.B(n_3655),
.C(n_3682),
.D(n_3630),
.Y(n_3855)
);

AND2x4_ASAP7_75t_L g3856 ( 
.A(n_3741),
.B(n_3614),
.Y(n_3856)
);

INVx1_ASAP7_75t_L g3857 ( 
.A(n_3723),
.Y(n_3857)
);

BUFx3_ASAP7_75t_L g3858 ( 
.A(n_3722),
.Y(n_3858)
);

NOR2xp33_ASAP7_75t_L g3859 ( 
.A(n_3685),
.B(n_3426),
.Y(n_3859)
);

NAND4xp75_ASAP7_75t_SL g3860 ( 
.A(n_3737),
.B(n_3491),
.C(n_3503),
.D(n_3408),
.Y(n_3860)
);

AND2x4_ASAP7_75t_L g3861 ( 
.A(n_3741),
.B(n_3614),
.Y(n_3861)
);

NAND2xp5_ASAP7_75t_L g3862 ( 
.A(n_3723),
.B(n_3627),
.Y(n_3862)
);

NAND4xp75_ASAP7_75t_L g3863 ( 
.A(n_3713),
.B(n_3677),
.C(n_3681),
.D(n_3673),
.Y(n_3863)
);

NAND3xp33_ASAP7_75t_L g3864 ( 
.A(n_3713),
.B(n_3720),
.C(n_3744),
.Y(n_3864)
);

XOR2x2_ASAP7_75t_L g3865 ( 
.A(n_3737),
.B(n_3513),
.Y(n_3865)
);

OR2x2_ASAP7_75t_L g3866 ( 
.A(n_3685),
.B(n_3632),
.Y(n_3866)
);

NOR2xp33_ASAP7_75t_L g3867 ( 
.A(n_3745),
.B(n_3438),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3735),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_L g3869 ( 
.A(n_3735),
.B(n_3640),
.Y(n_3869)
);

INVx1_ASAP7_75t_L g3870 ( 
.A(n_3785),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_3864),
.Y(n_3871)
);

INVx2_ASAP7_75t_L g3872 ( 
.A(n_3858),
.Y(n_3872)
);

INVx2_ASAP7_75t_SL g3873 ( 
.A(n_3802),
.Y(n_3873)
);

NAND2xp5_ASAP7_75t_L g3874 ( 
.A(n_3787),
.B(n_3795),
.Y(n_3874)
);

INVx1_ASAP7_75t_L g3875 ( 
.A(n_3864),
.Y(n_3875)
);

INVx2_ASAP7_75t_L g3876 ( 
.A(n_3792),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3853),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3813),
.Y(n_3878)
);

OR2x2_ASAP7_75t_L g3879 ( 
.A(n_3796),
.B(n_3755),
.Y(n_3879)
);

OR2x2_ASAP7_75t_L g3880 ( 
.A(n_3798),
.B(n_3787),
.Y(n_3880)
);

OR2x6_ASAP7_75t_L g3881 ( 
.A(n_3784),
.B(n_3760),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_3836),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_3795),
.B(n_3790),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_3813),
.Y(n_3884)
);

AOI21xp5_ASAP7_75t_L g3885 ( 
.A1(n_3794),
.A2(n_3823),
.B(n_3799),
.Y(n_3885)
);

NAND2xp5_ASAP7_75t_L g3886 ( 
.A(n_3789),
.B(n_3722),
.Y(n_3886)
);

INVx1_ASAP7_75t_SL g3887 ( 
.A(n_3821),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3777),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3833),
.Y(n_3889)
);

AND2x2_ASAP7_75t_L g3890 ( 
.A(n_3779),
.B(n_3705),
.Y(n_3890)
);

INVx2_ASAP7_75t_L g3891 ( 
.A(n_3856),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_3833),
.Y(n_3892)
);

OR2x2_ASAP7_75t_L g3893 ( 
.A(n_3783),
.B(n_3755),
.Y(n_3893)
);

AND2x2_ASAP7_75t_L g3894 ( 
.A(n_3805),
.B(n_3705),
.Y(n_3894)
);

NAND2x1p5_ASAP7_75t_L g3895 ( 
.A(n_3841),
.B(n_3536),
.Y(n_3895)
);

AND2x4_ASAP7_75t_L g3896 ( 
.A(n_3809),
.B(n_3764),
.Y(n_3896)
);

AND2x4_ASAP7_75t_L g3897 ( 
.A(n_3815),
.B(n_3764),
.Y(n_3897)
);

AND2x2_ASAP7_75t_L g3898 ( 
.A(n_3822),
.B(n_3709),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_3781),
.Y(n_3899)
);

AND2x4_ASAP7_75t_L g3900 ( 
.A(n_3856),
.B(n_3772),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_3778),
.Y(n_3901)
);

OR2x2_ASAP7_75t_L g3902 ( 
.A(n_3820),
.B(n_3811),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_L g3903 ( 
.A(n_3835),
.B(n_3709),
.Y(n_3903)
);

INVxp67_ASAP7_75t_L g3904 ( 
.A(n_3867),
.Y(n_3904)
);

NAND2xp5_ASAP7_75t_L g3905 ( 
.A(n_3793),
.B(n_3745),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_3793),
.B(n_3753),
.Y(n_3906)
);

INVxp67_ASAP7_75t_L g3907 ( 
.A(n_3800),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3849),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_L g3909 ( 
.A(n_3831),
.B(n_3753),
.Y(n_3909)
);

NAND2xp5_ASAP7_75t_L g3910 ( 
.A(n_3788),
.B(n_3762),
.Y(n_3910)
);

AND2x4_ASAP7_75t_L g3911 ( 
.A(n_3861),
.B(n_3772),
.Y(n_3911)
);

INVx1_ASAP7_75t_L g3912 ( 
.A(n_3791),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3849),
.Y(n_3913)
);

NAND2xp5_ASAP7_75t_L g3914 ( 
.A(n_3823),
.B(n_3762),
.Y(n_3914)
);

NAND2x1_ASAP7_75t_L g3915 ( 
.A(n_3861),
.B(n_3655),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3849),
.Y(n_3916)
);

OR2x2_ASAP7_75t_L g3917 ( 
.A(n_3810),
.B(n_3710),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3854),
.Y(n_3918)
);

AND2x2_ASAP7_75t_L g3919 ( 
.A(n_3834),
.B(n_3761),
.Y(n_3919)
);

NAND2xp5_ASAP7_75t_L g3920 ( 
.A(n_3859),
.B(n_3765),
.Y(n_3920)
);

NAND2xp5_ASAP7_75t_L g3921 ( 
.A(n_3797),
.B(n_3765),
.Y(n_3921)
);

INVx2_ASAP7_75t_L g3922 ( 
.A(n_3840),
.Y(n_3922)
);

NAND3xp33_ASAP7_75t_L g3923 ( 
.A(n_3837),
.B(n_3720),
.C(n_3736),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3845),
.Y(n_3924)
);

AND2x2_ASAP7_75t_L g3925 ( 
.A(n_3865),
.B(n_3761),
.Y(n_3925)
);

NOR2xp33_ASAP7_75t_SL g3926 ( 
.A(n_3842),
.B(n_3665),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3848),
.Y(n_3927)
);

INVx2_ASAP7_75t_SL g3928 ( 
.A(n_3841),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3801),
.Y(n_3929)
);

INVx2_ASAP7_75t_L g3930 ( 
.A(n_3850),
.Y(n_3930)
);

AND2x2_ASAP7_75t_L g3931 ( 
.A(n_3830),
.B(n_3768),
.Y(n_3931)
);

NOR2xp33_ASAP7_75t_L g3932 ( 
.A(n_3799),
.B(n_3773),
.Y(n_3932)
);

OAI21xp33_ASAP7_75t_L g3933 ( 
.A1(n_3807),
.A2(n_3756),
.B(n_3751),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_3850),
.B(n_3751),
.Y(n_3934)
);

INVx2_ASAP7_75t_L g3935 ( 
.A(n_3803),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3806),
.Y(n_3936)
);

NAND2x1p5_ASAP7_75t_L g3937 ( 
.A(n_3786),
.B(n_3544),
.Y(n_3937)
);

INVx3_ASAP7_75t_L g3938 ( 
.A(n_3825),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_L g3939 ( 
.A(n_3826),
.B(n_3756),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3808),
.Y(n_3940)
);

NOR2x1p5_ASAP7_75t_SL g3941 ( 
.A(n_3812),
.B(n_3770),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3816),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3817),
.Y(n_3943)
);

INVx2_ASAP7_75t_SL g3944 ( 
.A(n_3866),
.Y(n_3944)
);

BUFx3_ASAP7_75t_L g3945 ( 
.A(n_3829),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3818),
.Y(n_3946)
);

AOI22xp5_ASAP7_75t_L g3947 ( 
.A1(n_3804),
.A2(n_3851),
.B1(n_3843),
.B2(n_3807),
.Y(n_3947)
);

OR2x2_ASAP7_75t_L g3948 ( 
.A(n_3780),
.B(n_3832),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_3838),
.B(n_3757),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3819),
.Y(n_3950)
);

INVxp33_ASAP7_75t_L g3951 ( 
.A(n_3839),
.Y(n_3951)
);

INVx1_ASAP7_75t_SL g3952 ( 
.A(n_3814),
.Y(n_3952)
);

AND2x2_ASAP7_75t_L g3953 ( 
.A(n_3824),
.B(n_3768),
.Y(n_3953)
);

INVxp67_ASAP7_75t_L g3954 ( 
.A(n_3863),
.Y(n_3954)
);

OR2x2_ASAP7_75t_L g3955 ( 
.A(n_3855),
.B(n_3782),
.Y(n_3955)
);

AND2x2_ASAP7_75t_L g3956 ( 
.A(n_3828),
.B(n_3757),
.Y(n_3956)
);

AND2x2_ASAP7_75t_L g3957 ( 
.A(n_3844),
.B(n_3750),
.Y(n_3957)
);

OR2x2_ASAP7_75t_L g3958 ( 
.A(n_3855),
.B(n_3710),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_L g3959 ( 
.A(n_3894),
.B(n_3804),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3877),
.Y(n_3960)
);

AOI22xp5_ASAP7_75t_L g3961 ( 
.A1(n_3907),
.A2(n_3851),
.B1(n_3771),
.B2(n_3728),
.Y(n_3961)
);

INVx1_ASAP7_75t_L g3962 ( 
.A(n_3877),
.Y(n_3962)
);

OAI21xp5_ASAP7_75t_L g3963 ( 
.A1(n_3885),
.A2(n_3846),
.B(n_3770),
.Y(n_3963)
);

INVx1_ASAP7_75t_SL g3964 ( 
.A(n_3880),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3874),
.Y(n_3965)
);

INVxp67_ASAP7_75t_L g3966 ( 
.A(n_3926),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_3878),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_3878),
.Y(n_3968)
);

OAI21xp5_ASAP7_75t_L g3969 ( 
.A1(n_3947),
.A2(n_3910),
.B(n_3955),
.Y(n_3969)
);

OAI21xp33_ASAP7_75t_L g3970 ( 
.A1(n_3941),
.A2(n_3951),
.B(n_3903),
.Y(n_3970)
);

NOR2x1_ASAP7_75t_R g3971 ( 
.A(n_3945),
.B(n_3862),
.Y(n_3971)
);

INVxp67_ASAP7_75t_SL g3972 ( 
.A(n_3915),
.Y(n_3972)
);

AOI21xp5_ASAP7_75t_L g3973 ( 
.A1(n_3905),
.A2(n_3846),
.B(n_3862),
.Y(n_3973)
);

OAI211xp5_ASAP7_75t_SL g3974 ( 
.A1(n_3954),
.A2(n_3869),
.B(n_3857),
.C(n_3868),
.Y(n_3974)
);

OAI21xp33_ASAP7_75t_L g3975 ( 
.A1(n_3952),
.A2(n_3771),
.B(n_3750),
.Y(n_3975)
);

OAI21xp5_ASAP7_75t_L g3976 ( 
.A1(n_3906),
.A2(n_3869),
.B(n_3742),
.Y(n_3976)
);

AOI22xp5_ASAP7_75t_L g3977 ( 
.A1(n_3871),
.A2(n_3875),
.B1(n_3870),
.B2(n_3873),
.Y(n_3977)
);

HB1xp67_ASAP7_75t_L g3978 ( 
.A(n_3881),
.Y(n_3978)
);

INVx1_ASAP7_75t_L g3979 ( 
.A(n_3889),
.Y(n_3979)
);

AOI22xp5_ASAP7_75t_L g3980 ( 
.A1(n_3871),
.A2(n_3728),
.B1(n_3729),
.B2(n_3721),
.Y(n_3980)
);

INVxp67_ASAP7_75t_SL g3981 ( 
.A(n_3870),
.Y(n_3981)
);

OAI21xp5_ASAP7_75t_L g3982 ( 
.A1(n_3914),
.A2(n_3742),
.B(n_3736),
.Y(n_3982)
);

XOR2x2_ASAP7_75t_L g3983 ( 
.A(n_3925),
.B(n_3827),
.Y(n_3983)
);

AOI22xp33_ASAP7_75t_L g3984 ( 
.A1(n_3875),
.A2(n_3712),
.B1(n_3715),
.B2(n_3665),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3892),
.Y(n_3985)
);

INVx1_ASAP7_75t_L g3986 ( 
.A(n_3883),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3882),
.Y(n_3987)
);

INVx1_ASAP7_75t_SL g3988 ( 
.A(n_3919),
.Y(n_3988)
);

AND2x2_ASAP7_75t_L g3989 ( 
.A(n_3890),
.B(n_3712),
.Y(n_3989)
);

INVx2_ASAP7_75t_L g3990 ( 
.A(n_3900),
.Y(n_3990)
);

INVxp67_ASAP7_75t_L g3991 ( 
.A(n_3881),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3893),
.Y(n_3992)
);

INVx1_ASAP7_75t_L g3993 ( 
.A(n_3884),
.Y(n_3993)
);

INVx2_ASAP7_75t_SL g3994 ( 
.A(n_3900),
.Y(n_3994)
);

OAI211xp5_ASAP7_75t_SL g3995 ( 
.A1(n_3904),
.A2(n_3852),
.B(n_3743),
.C(n_3763),
.Y(n_3995)
);

INVx1_ASAP7_75t_L g3996 ( 
.A(n_3944),
.Y(n_3996)
);

AOI22xp5_ASAP7_75t_L g3997 ( 
.A1(n_3887),
.A2(n_3729),
.B1(n_3721),
.B2(n_3715),
.Y(n_3997)
);

INVx1_ASAP7_75t_L g3998 ( 
.A(n_3891),
.Y(n_3998)
);

INVx1_ASAP7_75t_L g3999 ( 
.A(n_3911),
.Y(n_3999)
);

XNOR2x1_ASAP7_75t_L g4000 ( 
.A(n_3876),
.B(n_3847),
.Y(n_4000)
);

NAND3xp33_ASAP7_75t_L g4001 ( 
.A(n_3923),
.B(n_3743),
.C(n_3763),
.Y(n_4001)
);

OAI21xp5_ASAP7_75t_L g4002 ( 
.A1(n_3937),
.A2(n_3776),
.B(n_3622),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_3911),
.Y(n_4003)
);

OAI22xp5_ASAP7_75t_L g4004 ( 
.A1(n_3922),
.A2(n_3665),
.B1(n_3776),
.B2(n_3679),
.Y(n_4004)
);

NAND3xp33_ASAP7_75t_L g4005 ( 
.A(n_3932),
.B(n_3773),
.C(n_3665),
.Y(n_4005)
);

AOI22xp5_ASAP7_75t_L g4006 ( 
.A1(n_3898),
.A2(n_3622),
.B1(n_3614),
.B2(n_3717),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3953),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_3957),
.Y(n_4008)
);

INVx1_ASAP7_75t_SL g4009 ( 
.A(n_3879),
.Y(n_4009)
);

INVx1_ASAP7_75t_L g4010 ( 
.A(n_3956),
.Y(n_4010)
);

AOI21xp5_ASAP7_75t_L g4011 ( 
.A1(n_3958),
.A2(n_3622),
.B(n_3733),
.Y(n_4011)
);

INVxp67_ASAP7_75t_L g4012 ( 
.A(n_3934),
.Y(n_4012)
);

AND2x2_ASAP7_75t_L g4013 ( 
.A(n_3931),
.B(n_3717),
.Y(n_4013)
);

AOI21xp33_ASAP7_75t_SL g4014 ( 
.A1(n_3917),
.A2(n_3679),
.B(n_3733),
.Y(n_4014)
);

OAI211xp5_ASAP7_75t_L g4015 ( 
.A1(n_3933),
.A2(n_3665),
.B(n_3679),
.C(n_3860),
.Y(n_4015)
);

OAI21xp5_ASAP7_75t_L g4016 ( 
.A1(n_3909),
.A2(n_3734),
.B(n_3733),
.Y(n_4016)
);

INVx1_ASAP7_75t_L g4017 ( 
.A(n_3918),
.Y(n_4017)
);

AOI221xp5_ASAP7_75t_L g4018 ( 
.A1(n_3899),
.A2(n_3888),
.B1(n_3912),
.B2(n_3901),
.C(n_3921),
.Y(n_4018)
);

O2A1O1Ixp33_ASAP7_75t_L g4019 ( 
.A1(n_3912),
.A2(n_3642),
.B(n_3649),
.C(n_3648),
.Y(n_4019)
);

NAND3xp33_ASAP7_75t_L g4020 ( 
.A(n_3901),
.B(n_3734),
.C(n_3659),
.Y(n_4020)
);

AOI21xp33_ASAP7_75t_SL g4021 ( 
.A1(n_3948),
.A2(n_3734),
.B(n_3661),
.Y(n_4021)
);

INVx1_ASAP7_75t_L g4022 ( 
.A(n_3908),
.Y(n_4022)
);

O2A1O1Ixp33_ASAP7_75t_SL g4023 ( 
.A1(n_3886),
.A2(n_3367),
.B(n_3678),
.C(n_3658),
.Y(n_4023)
);

OAI21xp33_ASAP7_75t_L g4024 ( 
.A1(n_3872),
.A2(n_3681),
.B(n_3672),
.Y(n_4024)
);

OAI22xp33_ASAP7_75t_L g4025 ( 
.A1(n_3895),
.A2(n_3367),
.B1(n_3402),
.B2(n_3511),
.Y(n_4025)
);

BUFx2_ASAP7_75t_SL g4026 ( 
.A(n_3930),
.Y(n_4026)
);

AOI22xp5_ASAP7_75t_L g4027 ( 
.A1(n_3896),
.A2(n_3897),
.B1(n_3928),
.B2(n_3939),
.Y(n_4027)
);

INVx1_ASAP7_75t_L g4028 ( 
.A(n_3913),
.Y(n_4028)
);

AOI21xp33_ASAP7_75t_L g4029 ( 
.A1(n_3902),
.A2(n_3487),
.B(n_3491),
.Y(n_4029)
);

INVx1_ASAP7_75t_L g4030 ( 
.A(n_3916),
.Y(n_4030)
);

NOR2xp33_ASAP7_75t_L g4031 ( 
.A(n_3949),
.B(n_3920),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_3896),
.B(n_3651),
.Y(n_4032)
);

OAI221xp5_ASAP7_75t_SL g4033 ( 
.A1(n_3935),
.A2(n_3357),
.B1(n_3373),
.B2(n_3421),
.C(n_3402),
.Y(n_4033)
);

OAI21xp5_ASAP7_75t_L g4034 ( 
.A1(n_3897),
.A2(n_3927),
.B(n_3924),
.Y(n_4034)
);

XNOR2xp5_ASAP7_75t_L g4035 ( 
.A(n_3938),
.B(n_3412),
.Y(n_4035)
);

NAND3xp33_ASAP7_75t_SL g4036 ( 
.A(n_3929),
.B(n_3373),
.C(n_3421),
.Y(n_4036)
);

INVx1_ASAP7_75t_L g4037 ( 
.A(n_3946),
.Y(n_4037)
);

XOR2x2_ASAP7_75t_L g4038 ( 
.A(n_3936),
.B(n_3412),
.Y(n_4038)
);

XOR2x2_ASAP7_75t_L g4039 ( 
.A(n_3940),
.B(n_3373),
.Y(n_4039)
);

OAI22xp33_ASAP7_75t_L g4040 ( 
.A1(n_3938),
.A2(n_3421),
.B1(n_3314),
.B2(n_3311),
.Y(n_4040)
);

AOI22xp33_ASAP7_75t_SL g4041 ( 
.A1(n_3942),
.A2(n_3943),
.B1(n_3950),
.B2(n_3946),
.Y(n_4041)
);

INVxp67_ASAP7_75t_L g4042 ( 
.A(n_3971),
.Y(n_4042)
);

AOI21xp5_ASAP7_75t_L g4043 ( 
.A1(n_3973),
.A2(n_3950),
.B(n_3375),
.Y(n_4043)
);

NAND2xp5_ASAP7_75t_SL g4044 ( 
.A(n_4035),
.B(n_3651),
.Y(n_4044)
);

OAI211xp5_ASAP7_75t_SL g4045 ( 
.A1(n_3969),
.A2(n_3375),
.B(n_3394),
.C(n_3379),
.Y(n_4045)
);

AOI22xp5_ASAP7_75t_L g4046 ( 
.A1(n_3970),
.A2(n_3496),
.B1(n_3672),
.B2(n_3503),
.Y(n_4046)
);

OAI322xp33_ASAP7_75t_L g4047 ( 
.A1(n_3977),
.A2(n_3368),
.A3(n_3379),
.B1(n_3311),
.B2(n_3398),
.C1(n_3403),
.C2(n_3526),
.Y(n_4047)
);

NOR2xp33_ASAP7_75t_L g4048 ( 
.A(n_3991),
.B(n_3496),
.Y(n_4048)
);

OAI32xp33_ASAP7_75t_L g4049 ( 
.A1(n_3963),
.A2(n_3368),
.A3(n_3379),
.B1(n_3403),
.B2(n_3312),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_3999),
.Y(n_4050)
);

AOI221xp5_ASAP7_75t_L g4051 ( 
.A1(n_4001),
.A2(n_3368),
.B1(n_3403),
.B2(n_3312),
.C(n_3526),
.Y(n_4051)
);

OAI21xp33_ASAP7_75t_SL g4052 ( 
.A1(n_3972),
.A2(n_3523),
.B(n_3520),
.Y(n_4052)
);

NAND2xp5_ASAP7_75t_L g4053 ( 
.A(n_3994),
.B(n_3496),
.Y(n_4053)
);

NAND2xp5_ASAP7_75t_L g4054 ( 
.A(n_3978),
.B(n_3315),
.Y(n_4054)
);

BUFx2_ASAP7_75t_L g4055 ( 
.A(n_4002),
.Y(n_4055)
);

NAND3x2_ASAP7_75t_L g4056 ( 
.A(n_3989),
.B(n_3333),
.C(n_3422),
.Y(n_4056)
);

INVx1_ASAP7_75t_L g4057 ( 
.A(n_4003),
.Y(n_4057)
);

INVx2_ASAP7_75t_L g4058 ( 
.A(n_3990),
.Y(n_4058)
);

OAI22xp33_ASAP7_75t_L g4059 ( 
.A1(n_3964),
.A2(n_3523),
.B1(n_3340),
.B2(n_3341),
.Y(n_4059)
);

NOR2xp33_ASAP7_75t_L g4060 ( 
.A(n_3988),
.B(n_3386),
.Y(n_4060)
);

INVx1_ASAP7_75t_L g4061 ( 
.A(n_4032),
.Y(n_4061)
);

AOI22xp5_ASAP7_75t_L g4062 ( 
.A1(n_3975),
.A2(n_3422),
.B1(n_3333),
.B2(n_3350),
.Y(n_4062)
);

INVx1_ASAP7_75t_L g4063 ( 
.A(n_3981),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_3988),
.Y(n_4064)
);

NOR2xp67_ASAP7_75t_L g4065 ( 
.A(n_4027),
.B(n_3341),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_L g4066 ( 
.A(n_4011),
.B(n_3370),
.Y(n_4066)
);

AOI21xp33_ASAP7_75t_SL g4067 ( 
.A1(n_4000),
.A2(n_187),
.B(n_188),
.Y(n_4067)
);

NAND3xp33_ASAP7_75t_L g4068 ( 
.A(n_4018),
.B(n_3312),
.C(n_188),
.Y(n_4068)
);

INVx1_ASAP7_75t_SL g4069 ( 
.A(n_4026),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_4020),
.Y(n_4070)
);

INVx1_ASAP7_75t_L g4071 ( 
.A(n_4020),
.Y(n_4071)
);

INVx1_ASAP7_75t_L g4072 ( 
.A(n_4008),
.Y(n_4072)
);

INVx1_ASAP7_75t_L g4073 ( 
.A(n_3996),
.Y(n_4073)
);

NAND2xp5_ASAP7_75t_L g4074 ( 
.A(n_4013),
.B(n_3370),
.Y(n_4074)
);

INVx1_ASAP7_75t_L g4075 ( 
.A(n_3967),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_3968),
.Y(n_4076)
);

AND2x2_ASAP7_75t_L g4077 ( 
.A(n_4009),
.B(n_3361),
.Y(n_4077)
);

NAND3xp33_ASAP7_75t_L g4078 ( 
.A(n_4001),
.B(n_4041),
.C(n_3976),
.Y(n_4078)
);

INVx1_ASAP7_75t_L g4079 ( 
.A(n_4007),
.Y(n_4079)
);

OAI22xp5_ASAP7_75t_L g4080 ( 
.A1(n_3997),
.A2(n_3422),
.B1(n_3333),
.B2(n_3386),
.Y(n_4080)
);

AND2x2_ASAP7_75t_L g4081 ( 
.A(n_4010),
.B(n_3361),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_3980),
.B(n_3386),
.Y(n_4082)
);

INVx2_ASAP7_75t_SL g4083 ( 
.A(n_4038),
.Y(n_4083)
);

INVx1_ASAP7_75t_L g4084 ( 
.A(n_3979),
.Y(n_4084)
);

INVx1_ASAP7_75t_L g4085 ( 
.A(n_3985),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_L g4086 ( 
.A(n_3961),
.B(n_3385),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_3992),
.Y(n_4087)
);

INVx1_ASAP7_75t_L g4088 ( 
.A(n_3998),
.Y(n_4088)
);

O2A1O1Ixp33_ASAP7_75t_SL g4089 ( 
.A1(n_4015),
.A2(n_3340),
.B(n_3353),
.C(n_3345),
.Y(n_4089)
);

INVx1_ASAP7_75t_L g4090 ( 
.A(n_3960),
.Y(n_4090)
);

NAND2xp5_ASAP7_75t_L g4091 ( 
.A(n_3965),
.B(n_3385),
.Y(n_4091)
);

AOI21xp5_ASAP7_75t_L g4092 ( 
.A1(n_4023),
.A2(n_3495),
.B(n_3348),
.Y(n_4092)
);

INVx1_ASAP7_75t_L g4093 ( 
.A(n_3962),
.Y(n_4093)
);

OR2x2_ASAP7_75t_L g4094 ( 
.A(n_3986),
.B(n_3396),
.Y(n_4094)
);

AND2x2_ASAP7_75t_L g4095 ( 
.A(n_3966),
.B(n_3377),
.Y(n_4095)
);

AND2x4_ASAP7_75t_L g4096 ( 
.A(n_4034),
.B(n_3333),
.Y(n_4096)
);

AND2x2_ASAP7_75t_L g4097 ( 
.A(n_4012),
.B(n_3993),
.Y(n_4097)
);

OAI21xp33_ASAP7_75t_L g4098 ( 
.A1(n_3983),
.A2(n_3324),
.B(n_3382),
.Y(n_4098)
);

OAI21xp5_ASAP7_75t_L g4099 ( 
.A1(n_4005),
.A2(n_3324),
.B(n_3382),
.Y(n_4099)
);

INVx1_ASAP7_75t_L g4100 ( 
.A(n_4037),
.Y(n_4100)
);

OAI21xp5_ASAP7_75t_L g4101 ( 
.A1(n_4005),
.A2(n_3324),
.B(n_3382),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_3987),
.Y(n_4102)
);

AOI222xp33_ASAP7_75t_L g4103 ( 
.A1(n_4036),
.A2(n_3384),
.B1(n_3377),
.B2(n_3322),
.C1(n_3359),
.C2(n_3339),
.Y(n_4103)
);

AOI22xp5_ASAP7_75t_L g4104 ( 
.A1(n_4031),
.A2(n_3350),
.B1(n_3418),
.B2(n_3339),
.Y(n_4104)
);

AOI21xp5_ASAP7_75t_L g4105 ( 
.A1(n_4025),
.A2(n_3495),
.B(n_3348),
.Y(n_4105)
);

AO22x1_ASAP7_75t_L g4106 ( 
.A1(n_4016),
.A2(n_3982),
.B1(n_3959),
.B2(n_4022),
.Y(n_4106)
);

INVx1_ASAP7_75t_SL g4107 ( 
.A(n_4069),
.Y(n_4107)
);

AOI221xp5_ASAP7_75t_L g4108 ( 
.A1(n_4078),
.A2(n_3974),
.B1(n_4021),
.B2(n_4014),
.C(n_4004),
.Y(n_4108)
);

OA21x2_ASAP7_75t_L g4109 ( 
.A1(n_4078),
.A2(n_4030),
.B(n_4028),
.Y(n_4109)
);

NAND2xp5_ASAP7_75t_L g4110 ( 
.A(n_4069),
.B(n_4024),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_L g4111 ( 
.A(n_4106),
.B(n_4017),
.Y(n_4111)
);

OAI21xp33_ASAP7_75t_L g4112 ( 
.A1(n_4098),
.A2(n_4006),
.B(n_3984),
.Y(n_4112)
);

AOI22xp5_ASAP7_75t_L g4113 ( 
.A1(n_4042),
.A2(n_4039),
.B1(n_3995),
.B2(n_4040),
.Y(n_4113)
);

OAI21xp33_ASAP7_75t_L g4114 ( 
.A1(n_4083),
.A2(n_4033),
.B(n_4019),
.Y(n_4114)
);

AOI22xp5_ASAP7_75t_L g4115 ( 
.A1(n_4048),
.A2(n_4029),
.B1(n_3418),
.B2(n_3350),
.Y(n_4115)
);

AOI22xp5_ASAP7_75t_SL g4116 ( 
.A1(n_4070),
.A2(n_3418),
.B1(n_3359),
.B2(n_3384),
.Y(n_4116)
);

INVx1_ASAP7_75t_L g4117 ( 
.A(n_4077),
.Y(n_4117)
);

INVx2_ASAP7_75t_SL g4118 ( 
.A(n_4096),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_4064),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_L g4120 ( 
.A(n_4071),
.B(n_3384),
.Y(n_4120)
);

OAI22xp5_ASAP7_75t_L g4121 ( 
.A1(n_4068),
.A2(n_3396),
.B1(n_3359),
.B2(n_3345),
.Y(n_4121)
);

AOI22xp33_ASAP7_75t_L g4122 ( 
.A1(n_4055),
.A2(n_3350),
.B1(n_3418),
.B2(n_3359),
.Y(n_4122)
);

NAND4xp25_ASAP7_75t_L g4123 ( 
.A(n_4065),
.B(n_3377),
.C(n_3356),
.D(n_3317),
.Y(n_4123)
);

AOI21xp33_ASAP7_75t_SL g4124 ( 
.A1(n_4068),
.A2(n_189),
.B(n_190),
.Y(n_4124)
);

INVxp67_ASAP7_75t_L g4125 ( 
.A(n_4054),
.Y(n_4125)
);

AND2x2_ASAP7_75t_L g4126 ( 
.A(n_4081),
.B(n_3371),
.Y(n_4126)
);

AOI22xp33_ASAP7_75t_L g4127 ( 
.A1(n_4073),
.A2(n_3345),
.B1(n_3362),
.B2(n_3356),
.Y(n_4127)
);

O2A1O1Ixp33_ASAP7_75t_L g4128 ( 
.A1(n_4067),
.A2(n_3362),
.B(n_190),
.C(n_191),
.Y(n_4128)
);

AOI22xp5_ASAP7_75t_L g4129 ( 
.A1(n_4044),
.A2(n_3317),
.B1(n_3322),
.B2(n_3362),
.Y(n_4129)
);

AOI211xp5_ASAP7_75t_L g4130 ( 
.A1(n_4049),
.A2(n_3322),
.B(n_3356),
.C(n_192),
.Y(n_4130)
);

AOI221xp5_ASAP7_75t_L g4131 ( 
.A1(n_4043),
.A2(n_3366),
.B1(n_3363),
.B2(n_3371),
.C(n_3358),
.Y(n_4131)
);

INVx1_ASAP7_75t_SL g4132 ( 
.A(n_4096),
.Y(n_4132)
);

NOR3xp33_ASAP7_75t_L g4133 ( 
.A(n_4087),
.B(n_3366),
.C(n_3363),
.Y(n_4133)
);

XOR2x2_ASAP7_75t_L g4134 ( 
.A(n_4095),
.B(n_189),
.Y(n_4134)
);

OAI22xp5_ASAP7_75t_SL g4135 ( 
.A1(n_4063),
.A2(n_4058),
.B1(n_4057),
.B2(n_4050),
.Y(n_4135)
);

AO221x1_ASAP7_75t_L g4136 ( 
.A1(n_4059),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.C(n_194),
.Y(n_4136)
);

AOI22xp5_ASAP7_75t_L g4137 ( 
.A1(n_4056),
.A2(n_3358),
.B1(n_3364),
.B2(n_196),
.Y(n_4137)
);

INVx2_ASAP7_75t_L g4138 ( 
.A(n_4097),
.Y(n_4138)
);

INVx3_ASAP7_75t_L g4139 ( 
.A(n_4072),
.Y(n_4139)
);

NAND2xp5_ASAP7_75t_L g4140 ( 
.A(n_4079),
.B(n_3358),
.Y(n_4140)
);

INVxp67_ASAP7_75t_L g4141 ( 
.A(n_4053),
.Y(n_4141)
);

INVxp67_ASAP7_75t_SL g4142 ( 
.A(n_4066),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_4094),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_4075),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_4076),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_4088),
.Y(n_4146)
);

NAND2xp5_ASAP7_75t_L g4147 ( 
.A(n_4084),
.B(n_3364),
.Y(n_4147)
);

INVxp67_ASAP7_75t_L g4148 ( 
.A(n_4060),
.Y(n_4148)
);

INVxp67_ASAP7_75t_L g4149 ( 
.A(n_4085),
.Y(n_4149)
);

NOR2xp33_ASAP7_75t_L g4150 ( 
.A(n_4061),
.B(n_193),
.Y(n_4150)
);

INVx1_ASAP7_75t_L g4151 ( 
.A(n_4090),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_L g4152 ( 
.A(n_4102),
.B(n_195),
.Y(n_4152)
);

AOI22xp5_ASAP7_75t_L g4153 ( 
.A1(n_4080),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_4093),
.Y(n_4154)
);

AOI22xp33_ASAP7_75t_SL g4155 ( 
.A1(n_4099),
.A2(n_197),
.B1(n_199),
.B2(n_200),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_L g4156 ( 
.A(n_4100),
.B(n_199),
.Y(n_4156)
);

NAND2xp5_ASAP7_75t_L g4157 ( 
.A(n_4086),
.B(n_201),
.Y(n_4157)
);

AOI21xp33_ASAP7_75t_L g4158 ( 
.A1(n_4052),
.A2(n_201),
.B(n_202),
.Y(n_4158)
);

OAI21xp5_ASAP7_75t_L g4159 ( 
.A1(n_4105),
.A2(n_203),
.B(n_204),
.Y(n_4159)
);

AOI221xp5_ASAP7_75t_L g4160 ( 
.A1(n_4045),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.C(n_206),
.Y(n_4160)
);

AOI211xp5_ASAP7_75t_L g4161 ( 
.A1(n_4089),
.A2(n_205),
.B(n_207),
.C(n_208),
.Y(n_4161)
);

INVx2_ASAP7_75t_L g4162 ( 
.A(n_4074),
.Y(n_4162)
);

OAI22xp5_ASAP7_75t_L g4163 ( 
.A1(n_4046),
.A2(n_4062),
.B1(n_4082),
.B2(n_4101),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_4091),
.Y(n_4164)
);

OAI211xp5_ASAP7_75t_SL g4165 ( 
.A1(n_4103),
.A2(n_208),
.B(n_209),
.C(n_210),
.Y(n_4165)
);

BUFx6f_ASAP7_75t_L g4166 ( 
.A(n_4047),
.Y(n_4166)
);

NOR3x1_ASAP7_75t_L g4167 ( 
.A(n_4136),
.B(n_4110),
.C(n_4118),
.Y(n_4167)
);

NOR2xp33_ASAP7_75t_L g4168 ( 
.A(n_4107),
.B(n_4047),
.Y(n_4168)
);

INVx1_ASAP7_75t_L g4169 ( 
.A(n_4135),
.Y(n_4169)
);

NOR2xp33_ASAP7_75t_L g4170 ( 
.A(n_4132),
.B(n_4092),
.Y(n_4170)
);

NAND3xp33_ASAP7_75t_SL g4171 ( 
.A(n_4108),
.B(n_4051),
.C(n_4104),
.Y(n_4171)
);

AOI21xp5_ASAP7_75t_L g4172 ( 
.A1(n_4111),
.A2(n_209),
.B(n_210),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_4117),
.Y(n_4173)
);

AND3x1_ASAP7_75t_L g4174 ( 
.A(n_4114),
.B(n_211),
.C(n_212),
.Y(n_4174)
);

NOR3xp33_ASAP7_75t_L g4175 ( 
.A(n_4112),
.B(n_211),
.C(n_213),
.Y(n_4175)
);

NAND2xp5_ASAP7_75t_L g4176 ( 
.A(n_4155),
.B(n_213),
.Y(n_4176)
);

AOI21xp5_ASAP7_75t_L g4177 ( 
.A1(n_4142),
.A2(n_214),
.B(n_215),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_4134),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_L g4179 ( 
.A(n_4139),
.B(n_214),
.Y(n_4179)
);

NOR2x1_ASAP7_75t_L g4180 ( 
.A(n_4139),
.B(n_215),
.Y(n_4180)
);

NAND2xp5_ASAP7_75t_L g4181 ( 
.A(n_4124),
.B(n_217),
.Y(n_4181)
);

NAND2xp5_ASAP7_75t_L g4182 ( 
.A(n_4109),
.B(n_217),
.Y(n_4182)
);

AOI221xp5_ASAP7_75t_L g4183 ( 
.A1(n_4166),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.C(n_221),
.Y(n_4183)
);

INVx1_ASAP7_75t_SL g4184 ( 
.A(n_4109),
.Y(n_4184)
);

AOI221xp5_ASAP7_75t_SL g4185 ( 
.A1(n_4163),
.A2(n_219),
.B1(n_221),
.B2(n_222),
.C(n_223),
.Y(n_4185)
);

AOI221xp5_ASAP7_75t_L g4186 ( 
.A1(n_4166),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.C(n_225),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_4119),
.Y(n_4187)
);

NAND3x1_ASAP7_75t_L g4188 ( 
.A(n_4113),
.B(n_224),
.C(n_226),
.Y(n_4188)
);

NOR2x1_ASAP7_75t_L g4189 ( 
.A(n_4143),
.B(n_227),
.Y(n_4189)
);

NOR2x1_ASAP7_75t_L g4190 ( 
.A(n_4138),
.B(n_229),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_4156),
.Y(n_4191)
);

NAND2xp5_ASAP7_75t_L g4192 ( 
.A(n_4161),
.B(n_231),
.Y(n_4192)
);

NOR2xp33_ASAP7_75t_L g4193 ( 
.A(n_4148),
.B(n_232),
.Y(n_4193)
);

AOI211xp5_ASAP7_75t_L g4194 ( 
.A1(n_4165),
.A2(n_232),
.B(n_234),
.C(n_236),
.Y(n_4194)
);

INVxp33_ASAP7_75t_SL g4195 ( 
.A(n_4150),
.Y(n_4195)
);

AO22x1_ASAP7_75t_L g4196 ( 
.A1(n_4166),
.A2(n_4159),
.B1(n_4146),
.B2(n_4162),
.Y(n_4196)
);

AOI21xp5_ASAP7_75t_L g4197 ( 
.A1(n_4128),
.A2(n_234),
.B(n_236),
.Y(n_4197)
);

NOR2xp33_ASAP7_75t_L g4198 ( 
.A(n_4125),
.B(n_237),
.Y(n_4198)
);

INVx2_ASAP7_75t_L g4199 ( 
.A(n_4126),
.Y(n_4199)
);

NAND3xp33_ASAP7_75t_L g4200 ( 
.A(n_4160),
.B(n_238),
.C(n_239),
.Y(n_4200)
);

NAND2xp5_ASAP7_75t_L g4201 ( 
.A(n_4130),
.B(n_240),
.Y(n_4201)
);

NAND2xp5_ASAP7_75t_SL g4202 ( 
.A(n_4116),
.B(n_240),
.Y(n_4202)
);

AOI221xp5_ASAP7_75t_L g4203 ( 
.A1(n_4158),
.A2(n_4120),
.B1(n_4149),
.B2(n_4141),
.C(n_4154),
.Y(n_4203)
);

NOR2xp33_ASAP7_75t_L g4204 ( 
.A(n_4147),
.B(n_241),
.Y(n_4204)
);

OA21x2_ASAP7_75t_SL g4205 ( 
.A1(n_4157),
.A2(n_241),
.B(n_242),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_4152),
.Y(n_4206)
);

NAND3xp33_ASAP7_75t_L g4207 ( 
.A(n_4153),
.B(n_243),
.C(n_244),
.Y(n_4207)
);

BUFx4f_ASAP7_75t_SL g4208 ( 
.A(n_4144),
.Y(n_4208)
);

NAND2xp5_ASAP7_75t_L g4209 ( 
.A(n_4137),
.B(n_243),
.Y(n_4209)
);

AOI21xp5_ASAP7_75t_L g4210 ( 
.A1(n_4140),
.A2(n_245),
.B(n_246),
.Y(n_4210)
);

OA22x2_ASAP7_75t_SL g4211 ( 
.A1(n_4145),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.Y(n_4211)
);

AND2x2_ASAP7_75t_L g4212 ( 
.A(n_4133),
.B(n_247),
.Y(n_4212)
);

XOR2x2_ASAP7_75t_L g4213 ( 
.A(n_4151),
.B(n_249),
.Y(n_4213)
);

AOI221xp5_ASAP7_75t_L g4214 ( 
.A1(n_4164),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.C(n_253),
.Y(n_4214)
);

AOI221x1_ASAP7_75t_L g4215 ( 
.A1(n_4121),
.A2(n_250),
.B1(n_254),
.B2(n_255),
.C(n_256),
.Y(n_4215)
);

NAND2xp5_ASAP7_75t_SL g4216 ( 
.A(n_4122),
.B(n_254),
.Y(n_4216)
);

AOI22xp5_ASAP7_75t_L g4217 ( 
.A1(n_4175),
.A2(n_4123),
.B1(n_4115),
.B2(n_4129),
.Y(n_4217)
);

NAND3xp33_ASAP7_75t_L g4218 ( 
.A(n_4183),
.B(n_4127),
.C(n_4131),
.Y(n_4218)
);

OAI21xp33_ASAP7_75t_L g4219 ( 
.A1(n_4168),
.A2(n_256),
.B(n_257),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_L g4220 ( 
.A(n_4196),
.B(n_257),
.Y(n_4220)
);

NAND3xp33_ASAP7_75t_L g4221 ( 
.A(n_4186),
.B(n_4215),
.C(n_4170),
.Y(n_4221)
);

O2A1O1Ixp5_ASAP7_75t_L g4222 ( 
.A1(n_4182),
.A2(n_258),
.B(n_259),
.C(n_261),
.Y(n_4222)
);

OAI211xp5_ASAP7_75t_SL g4223 ( 
.A1(n_4203),
.A2(n_258),
.B(n_262),
.C(n_263),
.Y(n_4223)
);

INVx1_ASAP7_75t_SL g4224 ( 
.A(n_4208),
.Y(n_4224)
);

AOI221xp5_ASAP7_75t_L g4225 ( 
.A1(n_4184),
.A2(n_262),
.B1(n_263),
.B2(n_264),
.C(n_265),
.Y(n_4225)
);

AOI221xp5_ASAP7_75t_L g4226 ( 
.A1(n_4184),
.A2(n_4169),
.B1(n_4171),
.B2(n_4174),
.C(n_4185),
.Y(n_4226)
);

AOI221xp5_ASAP7_75t_L g4227 ( 
.A1(n_4172),
.A2(n_264),
.B1(n_265),
.B2(n_268),
.C(n_269),
.Y(n_4227)
);

AOI21xp5_ASAP7_75t_L g4228 ( 
.A1(n_4202),
.A2(n_4197),
.B(n_4216),
.Y(n_4228)
);

AOI221xp5_ASAP7_75t_L g4229 ( 
.A1(n_4173),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.C(n_273),
.Y(n_4229)
);

NAND3xp33_ASAP7_75t_SL g4230 ( 
.A(n_4194),
.B(n_271),
.C(n_272),
.Y(n_4230)
);

OAI211xp5_ASAP7_75t_L g4231 ( 
.A1(n_4189),
.A2(n_273),
.B(n_274),
.C(n_275),
.Y(n_4231)
);

AOI22xp5_ASAP7_75t_L g4232 ( 
.A1(n_4188),
.A2(n_274),
.B1(n_276),
.B2(n_277),
.Y(n_4232)
);

NAND4xp25_ASAP7_75t_L g4233 ( 
.A(n_4167),
.B(n_276),
.C(n_277),
.D(n_278),
.Y(n_4233)
);

OAI221xp5_ASAP7_75t_L g4234 ( 
.A1(n_4201),
.A2(n_278),
.B1(n_280),
.B2(n_285),
.C(n_286),
.Y(n_4234)
);

AOI22xp5_ASAP7_75t_L g4235 ( 
.A1(n_4199),
.A2(n_280),
.B1(n_287),
.B2(n_288),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_4180),
.Y(n_4236)
);

AOI211x1_ASAP7_75t_L g4237 ( 
.A1(n_4200),
.A2(n_287),
.B(n_288),
.C(n_289),
.Y(n_4237)
);

OAI22xp5_ASAP7_75t_L g4238 ( 
.A1(n_4178),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_4238)
);

NOR2xp33_ASAP7_75t_L g4239 ( 
.A(n_4195),
.B(n_292),
.Y(n_4239)
);

OAI21xp5_ASAP7_75t_L g4240 ( 
.A1(n_4190),
.A2(n_296),
.B(n_297),
.Y(n_4240)
);

OAI21xp5_ASAP7_75t_L g4241 ( 
.A1(n_4177),
.A2(n_4210),
.B(n_4179),
.Y(n_4241)
);

AOI211xp5_ASAP7_75t_L g4242 ( 
.A1(n_4193),
.A2(n_296),
.B(n_297),
.C(n_298),
.Y(n_4242)
);

O2A1O1Ixp5_ASAP7_75t_L g4243 ( 
.A1(n_4187),
.A2(n_298),
.B(n_299),
.C(n_344),
.Y(n_4243)
);

INVx2_ASAP7_75t_L g4244 ( 
.A(n_4211),
.Y(n_4244)
);

INVx2_ASAP7_75t_SL g4245 ( 
.A(n_4213),
.Y(n_4245)
);

NAND2xp5_ASAP7_75t_L g4246 ( 
.A(n_4212),
.B(n_345),
.Y(n_4246)
);

NAND3xp33_ASAP7_75t_L g4247 ( 
.A(n_4198),
.B(n_1035),
.C(n_1027),
.Y(n_4247)
);

NOR2xp33_ASAP7_75t_R g4248 ( 
.A(n_4192),
.B(n_346),
.Y(n_4248)
);

AOI21xp33_ASAP7_75t_SL g4249 ( 
.A1(n_4179),
.A2(n_349),
.B(n_351),
.Y(n_4249)
);

AOI211xp5_ASAP7_75t_L g4250 ( 
.A1(n_4209),
.A2(n_356),
.B(n_358),
.C(n_359),
.Y(n_4250)
);

AOI211xp5_ASAP7_75t_L g4251 ( 
.A1(n_4204),
.A2(n_360),
.B(n_361),
.C(n_363),
.Y(n_4251)
);

A2O1A1Ixp33_ASAP7_75t_L g4252 ( 
.A1(n_4214),
.A2(n_364),
.B(n_367),
.C(n_369),
.Y(n_4252)
);

AOI21xp5_ASAP7_75t_L g4253 ( 
.A1(n_4181),
.A2(n_370),
.B(n_376),
.Y(n_4253)
);

INVx2_ASAP7_75t_L g4254 ( 
.A(n_4244),
.Y(n_4254)
);

INVx1_ASAP7_75t_SL g4255 ( 
.A(n_4236),
.Y(n_4255)
);

INVx1_ASAP7_75t_L g4256 ( 
.A(n_4220),
.Y(n_4256)
);

INVx1_ASAP7_75t_L g4257 ( 
.A(n_4232),
.Y(n_4257)
);

INVx1_ASAP7_75t_L g4258 ( 
.A(n_4222),
.Y(n_4258)
);

INVx2_ASAP7_75t_SL g4259 ( 
.A(n_4224),
.Y(n_4259)
);

OAI22xp5_ASAP7_75t_L g4260 ( 
.A1(n_4217),
.A2(n_4207),
.B1(n_4176),
.B2(n_4191),
.Y(n_4260)
);

NAND4xp75_ASAP7_75t_L g4261 ( 
.A(n_4226),
.B(n_4206),
.C(n_4205),
.D(n_380),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_4238),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_4231),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_4239),
.Y(n_4264)
);

AO22x1_ASAP7_75t_L g4265 ( 
.A1(n_4240),
.A2(n_377),
.B1(n_378),
.B2(n_381),
.Y(n_4265)
);

INVxp33_ASAP7_75t_SL g4266 ( 
.A(n_4248),
.Y(n_4266)
);

OAI22xp5_ASAP7_75t_L g4267 ( 
.A1(n_4221),
.A2(n_383),
.B1(n_384),
.B2(n_389),
.Y(n_4267)
);

O2A1O1Ixp33_ASAP7_75t_SL g4268 ( 
.A1(n_4245),
.A2(n_396),
.B(n_399),
.C(n_401),
.Y(n_4268)
);

AOI22xp5_ASAP7_75t_L g4269 ( 
.A1(n_4233),
.A2(n_402),
.B1(n_403),
.B2(n_407),
.Y(n_4269)
);

INVx1_ASAP7_75t_L g4270 ( 
.A(n_4246),
.Y(n_4270)
);

A2O1A1Ixp33_ASAP7_75t_L g4271 ( 
.A1(n_4243),
.A2(n_4225),
.B(n_4219),
.C(n_4228),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_4237),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_4241),
.Y(n_4273)
);

AOI22xp5_ASAP7_75t_L g4274 ( 
.A1(n_4230),
.A2(n_413),
.B1(n_415),
.B2(n_418),
.Y(n_4274)
);

INVxp67_ASAP7_75t_L g4275 ( 
.A(n_4234),
.Y(n_4275)
);

OAI22xp5_ASAP7_75t_L g4276 ( 
.A1(n_4218),
.A2(n_424),
.B1(n_427),
.B2(n_429),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_4241),
.Y(n_4277)
);

AOI221xp5_ASAP7_75t_L g4278 ( 
.A1(n_4255),
.A2(n_4223),
.B1(n_4227),
.B2(n_4247),
.C(n_4249),
.Y(n_4278)
);

OAI221xp5_ASAP7_75t_L g4279 ( 
.A1(n_4255),
.A2(n_4252),
.B1(n_4242),
.B2(n_4253),
.C(n_4229),
.Y(n_4279)
);

NAND2xp33_ASAP7_75t_R g4280 ( 
.A(n_4266),
.B(n_4250),
.Y(n_4280)
);

NAND2xp5_ASAP7_75t_L g4281 ( 
.A(n_4259),
.B(n_4235),
.Y(n_4281)
);

BUFx2_ASAP7_75t_L g4282 ( 
.A(n_4258),
.Y(n_4282)
);

AOI211xp5_ASAP7_75t_SL g4283 ( 
.A1(n_4260),
.A2(n_4251),
.B(n_434),
.C(n_435),
.Y(n_4283)
);

AOI222xp33_ASAP7_75t_L g4284 ( 
.A1(n_4273),
.A2(n_430),
.B1(n_437),
.B2(n_440),
.C1(n_442),
.C2(n_444),
.Y(n_4284)
);

NOR2xp33_ASAP7_75t_R g4285 ( 
.A(n_4263),
.B(n_448),
.Y(n_4285)
);

AOI222xp33_ASAP7_75t_L g4286 ( 
.A1(n_4277),
.A2(n_450),
.B1(n_452),
.B2(n_453),
.C1(n_457),
.C2(n_458),
.Y(n_4286)
);

AOI211x1_ASAP7_75t_SL g4287 ( 
.A1(n_4271),
.A2(n_460),
.B(n_462),
.C(n_463),
.Y(n_4287)
);

AOI31xp33_ASAP7_75t_L g4288 ( 
.A1(n_4262),
.A2(n_964),
.A3(n_989),
.B(n_1004),
.Y(n_4288)
);

NAND2xp5_ASAP7_75t_SL g4289 ( 
.A(n_4254),
.B(n_964),
.Y(n_4289)
);

AOI21xp33_ASAP7_75t_SL g4290 ( 
.A1(n_4272),
.A2(n_964),
.B(n_989),
.Y(n_4290)
);

AOI221xp5_ASAP7_75t_L g4291 ( 
.A1(n_4257),
.A2(n_1234),
.B1(n_1252),
.B2(n_1246),
.C(n_1213),
.Y(n_4291)
);

AOI22xp5_ASAP7_75t_L g4292 ( 
.A1(n_4261),
.A2(n_964),
.B1(n_989),
.B2(n_1004),
.Y(n_4292)
);

NAND2xp5_ASAP7_75t_SL g4293 ( 
.A(n_4274),
.B(n_964),
.Y(n_4293)
);

NAND2x1_ASAP7_75t_L g4294 ( 
.A(n_4282),
.B(n_4264),
.Y(n_4294)
);

INVx2_ASAP7_75t_SL g4295 ( 
.A(n_4285),
.Y(n_4295)
);

OAI22xp5_ASAP7_75t_L g4296 ( 
.A1(n_4279),
.A2(n_4269),
.B1(n_4275),
.B2(n_4256),
.Y(n_4296)
);

AOI221xp5_ASAP7_75t_L g4297 ( 
.A1(n_4278),
.A2(n_4276),
.B1(n_4267),
.B2(n_4268),
.C(n_4270),
.Y(n_4297)
);

AOI221xp5_ASAP7_75t_L g4298 ( 
.A1(n_4281),
.A2(n_4265),
.B1(n_1234),
.B2(n_1246),
.C(n_1252),
.Y(n_4298)
);

OAI211xp5_ASAP7_75t_SL g4299 ( 
.A1(n_4292),
.A2(n_964),
.B(n_989),
.C(n_1004),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_4287),
.Y(n_4300)
);

HB1xp67_ASAP7_75t_L g4301 ( 
.A(n_4280),
.Y(n_4301)
);

INVx1_ASAP7_75t_SL g4302 ( 
.A(n_4293),
.Y(n_4302)
);

AO221x1_ASAP7_75t_L g4303 ( 
.A1(n_4290),
.A2(n_1234),
.B1(n_1252),
.B2(n_1246),
.C(n_1213),
.Y(n_4303)
);

NAND4xp25_ASAP7_75t_L g4304 ( 
.A(n_4283),
.B(n_964),
.C(n_989),
.D(n_1004),
.Y(n_4304)
);

NOR2x1_ASAP7_75t_L g4305 ( 
.A(n_4294),
.B(n_4288),
.Y(n_4305)
);

AOI21xp5_ASAP7_75t_L g4306 ( 
.A1(n_4296),
.A2(n_4289),
.B(n_4291),
.Y(n_4306)
);

AND3x4_ASAP7_75t_L g4307 ( 
.A(n_4301),
.B(n_4286),
.C(n_4284),
.Y(n_4307)
);

AOI222xp33_ASAP7_75t_L g4308 ( 
.A1(n_4297),
.A2(n_989),
.B1(n_1004),
.B2(n_1027),
.C1(n_1035),
.C2(n_1192),
.Y(n_4308)
);

INVxp67_ASAP7_75t_SL g4309 ( 
.A(n_4300),
.Y(n_4309)
);

AOI21xp5_ASAP7_75t_L g4310 ( 
.A1(n_4295),
.A2(n_989),
.B(n_1004),
.Y(n_4310)
);

AND2x2_ASAP7_75t_L g4311 ( 
.A(n_4302),
.B(n_1004),
.Y(n_4311)
);

XNOR2x1_ASAP7_75t_L g4312 ( 
.A(n_4307),
.B(n_4304),
.Y(n_4312)
);

OAI22xp5_ASAP7_75t_L g4313 ( 
.A1(n_4309),
.A2(n_4298),
.B1(n_4303),
.B2(n_4299),
.Y(n_4313)
);

AND2x2_ASAP7_75t_L g4314 ( 
.A(n_4305),
.B(n_1027),
.Y(n_4314)
);

HB1xp67_ASAP7_75t_L g4315 ( 
.A(n_4311),
.Y(n_4315)
);

OR2x2_ASAP7_75t_L g4316 ( 
.A(n_4306),
.B(n_4310),
.Y(n_4316)
);

AOI22xp5_ASAP7_75t_L g4317 ( 
.A1(n_4312),
.A2(n_4308),
.B1(n_1035),
.B2(n_1027),
.Y(n_4317)
);

AND2x4_ASAP7_75t_L g4318 ( 
.A(n_4315),
.B(n_1252),
.Y(n_4318)
);

NOR2xp67_ASAP7_75t_L g4319 ( 
.A(n_4317),
.B(n_4313),
.Y(n_4319)
);

OR4x1_ASAP7_75t_L g4320 ( 
.A(n_4318),
.B(n_4316),
.C(n_4314),
.D(n_1027),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_4320),
.Y(n_4321)
);

NAND2xp5_ASAP7_75t_L g4322 ( 
.A(n_4321),
.B(n_4319),
.Y(n_4322)
);

NAND4xp25_ASAP7_75t_SL g4323 ( 
.A(n_4322),
.B(n_1027),
.C(n_1035),
.D(n_1213),
.Y(n_4323)
);

AOI22xp33_ASAP7_75t_L g4324 ( 
.A1(n_4323),
.A2(n_1252),
.B1(n_1246),
.B2(n_1234),
.Y(n_4324)
);

INVx1_ASAP7_75t_L g4325 ( 
.A(n_4324),
.Y(n_4325)
);

NAND2xp5_ASAP7_75t_SL g4326 ( 
.A(n_4325),
.B(n_1027),
.Y(n_4326)
);

OAI21xp5_ASAP7_75t_SL g4327 ( 
.A1(n_4326),
.A2(n_1234),
.B(n_1246),
.Y(n_4327)
);

HB1xp67_ASAP7_75t_L g4328 ( 
.A(n_4327),
.Y(n_4328)
);

OR2x6_ASAP7_75t_L g4329 ( 
.A(n_4328),
.B(n_1035),
.Y(n_4329)
);

AOI21xp5_ASAP7_75t_L g4330 ( 
.A1(n_4329),
.A2(n_1035),
.B(n_1315),
.Y(n_4330)
);

AOI211xp5_ASAP7_75t_L g4331 ( 
.A1(n_4330),
.A2(n_1035),
.B(n_1433),
.C(n_1330),
.Y(n_4331)
);


endmodule