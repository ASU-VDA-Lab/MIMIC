module fake_jpeg_2719_n_204 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_204);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_7),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_28),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_9),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_6),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_14),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_2),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_45),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_19),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_21),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_14),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_1),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_77),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_1),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_2),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_78),
.B(n_60),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_3),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_60),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_86),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_56),
.C(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_88),
.B(n_98),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_72),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_93),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_55),
.B1(n_56),
.B2(n_70),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_63),
.B1(n_59),
.B2(n_64),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_58),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_55),
.B1(n_72),
.B2(n_66),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_82),
.B1(n_64),
.B2(n_71),
.Y(n_103)
);

CKINVDCx6p67_ASAP7_75t_R g97 ( 
.A(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_66),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_63),
.B1(n_76),
.B2(n_82),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_107),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_97),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_105),
.B(n_57),
.Y(n_133)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_110),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_136)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_97),
.A2(n_71),
.B1(n_59),
.B2(n_62),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_111),
.A2(n_114),
.B(n_95),
.Y(n_123)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_113),
.Y(n_141)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_67),
.B(n_69),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_73),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_118),
.Y(n_140)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_96),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_68),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_65),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_126),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_52),
.B(n_91),
.C(n_57),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_125),
.B(n_128),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_96),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_114),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_4),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_130),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_4),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_5),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_132),
.B(n_135),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_133),
.Y(n_153)
);

NAND2xp33_ASAP7_75t_SL g134 ( 
.A(n_117),
.B(n_27),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_SL g148 ( 
.A1(n_134),
.A2(n_32),
.B(n_49),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_103),
.B(n_5),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_103),
.B(n_10),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_138),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_10),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_111),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_11),
.Y(n_146)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_141),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_147),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_152),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_31),
.C(n_48),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_158),
.C(n_119),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_131),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_151),
.A2(n_155),
.B1(n_160),
.B2(n_162),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_12),
.Y(n_152)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_164),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_35),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_131),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_123),
.B(n_36),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_119),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_131),
.A2(n_17),
.B1(n_18),
.B2(n_20),
.Y(n_162)
);

NAND2x1p5_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_22),
.Y(n_163)
);

A2O1A1O1Ixp25_ASAP7_75t_L g166 ( 
.A1(n_163),
.A2(n_134),
.B(n_136),
.C(n_34),
.D(n_37),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_120),
.B(n_24),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_168),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_120),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_25),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_171),
.B(n_177),
.Y(n_181)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_174),
.C(n_158),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_L g175 ( 
.A1(n_159),
.A2(n_30),
.B1(n_38),
.B2(n_39),
.Y(n_175)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_157),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_44),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_178),
.B(n_50),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_159),
.A2(n_46),
.B(n_47),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_166),
.B(n_175),
.Y(n_182)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_144),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_179),
.B(n_163),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_184),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_165),
.Y(n_191)
);

INVxp33_ASAP7_75t_SL g190 ( 
.A(n_185),
.Y(n_190)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_190),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_192),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_187),
.A2(n_170),
.B1(n_143),
.B2(n_161),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_193),
.A2(n_169),
.B1(n_188),
.B2(n_184),
.Y(n_197)
);

AO221x1_ASAP7_75t_L g195 ( 
.A1(n_190),
.A2(n_181),
.B1(n_176),
.B2(n_170),
.C(n_148),
.Y(n_195)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_195),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_194),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_198),
.A2(n_196),
.B(n_197),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_199),
.C(n_173),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_201),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_202),
.A2(n_189),
.B1(n_167),
.B2(n_174),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_203),
.B(n_149),
.Y(n_204)
);


endmodule