module fake_jpeg_1937_n_261 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_261);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_261;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_2),
.B(n_1),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_25),
.B(n_14),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_50),
.Y(n_79)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_52),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_25),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_21),
.B(n_7),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_53),
.B(n_54),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_21),
.B(n_13),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_55),
.B(n_57),
.Y(n_97)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_SL g93 ( 
.A(n_56),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_22),
.B(n_6),
.C(n_10),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_58),
.B(n_61),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_64),
.Y(n_91)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_62),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_73),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_18),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_18),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_67),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_15),
.B(n_6),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_66),
.B(n_40),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_15),
.B(n_28),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_69),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_17),
.B(n_5),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_17),
.B(n_5),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_71),
.Y(n_111)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_72),
.A2(n_26),
.B1(n_36),
.B2(n_29),
.Y(n_74)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_22),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_78),
.B(n_84),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_39),
.B1(n_36),
.B2(n_29),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_81),
.A2(n_83),
.B1(n_87),
.B2(n_89),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_58),
.A2(n_39),
.B1(n_20),
.B2(n_27),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_38),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_53),
.A2(n_36),
.B1(n_29),
.B2(n_38),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_85),
.A2(n_88),
.B1(n_103),
.B2(n_107),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_73),
.A2(n_33),
.B1(n_28),
.B2(n_27),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_86),
.A2(n_110),
.B1(n_55),
.B2(n_81),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_56),
.A2(n_72),
.B1(n_62),
.B2(n_64),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_66),
.A2(n_37),
.B1(n_23),
.B2(n_33),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_41),
.A2(n_20),
.B1(n_19),
.B2(n_23),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_59),
.A2(n_37),
.B(n_19),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_SL g116 ( 
.A1(n_95),
.A2(n_98),
.B(n_100),
.C(n_112),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_63),
.A2(n_16),
.B1(n_31),
.B2(n_0),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_42),
.A2(n_16),
.B1(n_1),
.B2(n_31),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_99),
.A2(n_104),
.B1(n_109),
.B2(n_106),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_46),
.A2(n_16),
.B1(n_4),
.B2(n_8),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_47),
.A2(n_16),
.B1(n_9),
.B2(n_10),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_60),
.A2(n_16),
.B1(n_9),
.B2(n_12),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_3),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_115),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_49),
.A2(n_3),
.B1(n_12),
.B2(n_51),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_68),
.A2(n_71),
.B1(n_61),
.B2(n_44),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_113),
.B(n_43),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_55),
.B(n_44),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_91),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_117),
.B(n_124),
.Y(n_162)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_118),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_45),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_120),
.B(n_122),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_55),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_143),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_44),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_50),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_125),
.B(n_126),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_79),
.B(n_50),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_50),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_127),
.Y(n_156)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_131),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_132),
.A2(n_115),
.B1(n_90),
.B2(n_76),
.Y(n_180)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_77),
.Y(n_135)
);

BUFx24_ASAP7_75t_SL g157 ( 
.A(n_135),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_140),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_121),
.B1(n_100),
.B2(n_147),
.Y(n_170)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_82),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_141),
.Y(n_168)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_82),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

AOI21xp33_ASAP7_75t_L g158 ( 
.A1(n_144),
.A2(n_150),
.B(n_152),
.Y(n_158)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_76),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_146),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_104),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_78),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_149),
.Y(n_174)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_106),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_96),
.B(n_88),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_90),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_108),
.B(n_111),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_148),
.A2(n_97),
.B1(n_80),
.B2(n_75),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_154),
.A2(n_159),
.B1(n_161),
.B2(n_170),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_116),
.A2(n_80),
.B1(n_75),
.B2(n_85),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_123),
.A2(n_104),
.B(n_95),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_160),
.A2(n_164),
.B(n_153),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_116),
.A2(n_99),
.B1(n_105),
.B2(n_98),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_SL g166 ( 
.A1(n_116),
.A2(n_98),
.B(n_93),
.C(n_112),
.Y(n_166)
);

A2O1A1O1Ixp25_ASAP7_75t_L g199 ( 
.A1(n_166),
.A2(n_161),
.B(n_164),
.C(n_172),
.D(n_179),
.Y(n_199)
);

AO21x2_ASAP7_75t_L g172 ( 
.A1(n_139),
.A2(n_110),
.B(n_98),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_172),
.A2(n_177),
.B1(n_131),
.B2(n_140),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_119),
.A2(n_116),
.B1(n_136),
.B2(n_142),
.Y(n_177)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_179),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_180),
.Y(n_187)
);

NOR3xp33_ASAP7_75t_SL g182 ( 
.A(n_165),
.B(n_136),
.C(n_128),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_182),
.B(n_186),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_145),
.C(n_133),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_190),
.C(n_192),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_184),
.A2(n_185),
.B1(n_180),
.B2(n_175),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_177),
.A2(n_149),
.B1(n_141),
.B2(n_130),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_129),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_151),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_188),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_162),
.B(n_143),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_189),
.B(n_191),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_137),
.C(n_114),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_118),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_114),
.C(n_176),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_114),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_193),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_194),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_195),
.B(n_198),
.Y(n_213)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_199),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_159),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_155),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_200),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_155),
.B(n_178),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_201),
.A2(n_172),
.B1(n_178),
.B2(n_175),
.Y(n_210)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_184),
.A2(n_166),
.B1(n_172),
.B2(n_158),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_207),
.A2(n_188),
.B(n_201),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_210),
.B(n_183),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_189),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_214),
.B(n_216),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_198),
.A2(n_172),
.B1(n_166),
.B2(n_173),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_215),
.A2(n_217),
.B1(n_181),
.B2(n_196),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_186),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_187),
.A2(n_167),
.B1(n_173),
.B2(n_169),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_214),
.A2(n_181),
.B1(n_199),
.B2(n_182),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_218),
.A2(n_229),
.B(n_219),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_212),
.A2(n_185),
.B1(n_203),
.B2(n_216),
.Y(n_221)
);

NAND4xp25_ASAP7_75t_SL g230 ( 
.A(n_221),
.B(n_206),
.C(n_217),
.D(n_208),
.Y(n_230)
);

AOI21xp33_ASAP7_75t_L g222 ( 
.A1(n_212),
.A2(n_195),
.B(n_193),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_227),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_203),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_215),
.A2(n_197),
.B1(n_191),
.B2(n_192),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_202),
.B(n_190),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_226),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_197),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_188),
.C(n_200),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_209),
.Y(n_232)
);

NOR3xp33_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_231),
.C(n_237),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_236),
.C(n_227),
.Y(n_245)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_233),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_224),
.Y(n_239)
);

AOI322xp5_ASAP7_75t_L g236 ( 
.A1(n_229),
.A2(n_203),
.A3(n_205),
.B1(n_202),
.B2(n_213),
.C1(n_211),
.C2(n_207),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_225),
.A2(n_204),
.B(n_155),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_235),
.Y(n_247)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_233),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_243),
.Y(n_246)
);

NOR2xp67_ASAP7_75t_SL g243 ( 
.A(n_231),
.B(n_228),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_237),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_245),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_247),
.A2(n_249),
.B(n_250),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_240),
.A2(n_238),
.B1(n_218),
.B2(n_220),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_232),
.C(n_226),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_246),
.A2(n_241),
.B(n_234),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_253),
.Y(n_257)
);

AO21x1_ASAP7_75t_L g253 ( 
.A1(n_248),
.A2(n_241),
.B(n_220),
.Y(n_253)
);

OAI221xp5_ASAP7_75t_L g254 ( 
.A1(n_250),
.A2(n_230),
.B1(n_204),
.B2(n_171),
.C(n_167),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_254),
.B(n_194),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_249),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_256),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_257),
.A2(n_247),
.B(n_163),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_258),
.B(n_168),
.C(n_171),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_259),
.Y(n_261)
);


endmodule