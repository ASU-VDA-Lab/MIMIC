module fake_jpeg_2658_n_517 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_517);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_517;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_5),
.B(n_17),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_56),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_35),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_57),
.B(n_65),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_1),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_58),
.B(n_93),
.Y(n_171)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_59),
.Y(n_133)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_61),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_62),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g151 ( 
.A(n_63),
.Y(n_151)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_64),
.Y(n_140)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_67),
.Y(n_157)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_30),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_70),
.B(n_71),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_27),
.B(n_1),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_72),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_73),
.Y(n_173)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_74),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_37),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_75),
.B(n_79),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_77),
.Y(n_159)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_78),
.Y(n_182)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_80),
.Y(n_174)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_81),
.Y(n_186)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_82),
.B(n_87),
.Y(n_156)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_24),
.Y(n_84)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx11_ASAP7_75t_L g169 ( 
.A(n_86),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_27),
.Y(n_87)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

BUFx24_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_89),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_90),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_91),
.Y(n_166)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_92),
.Y(n_158)
);

NAND2xp33_ASAP7_75t_SL g93 ( 
.A(n_18),
.B(n_36),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_94),
.Y(n_172)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_34),
.Y(n_96)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_96),
.Y(n_175)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_97),
.B(n_120),
.Y(n_161)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_18),
.Y(n_98)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_99),
.Y(n_192)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_23),
.Y(n_100)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_100),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_24),
.Y(n_101)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_101),
.Y(n_187)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_25),
.B(n_1),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_2),
.Y(n_141)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g185 ( 
.A(n_104),
.Y(n_185)
);

BUFx12_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_105),
.Y(n_131)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_21),
.Y(n_107)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_29),
.Y(n_108)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_109),
.Y(n_160)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_21),
.Y(n_110)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_110),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_21),
.Y(n_111)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_43),
.Y(n_113)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_113),
.Y(n_168)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_43),
.Y(n_114)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_29),
.Y(n_115)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_115),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_31),
.Y(n_116)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_116),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_45),
.Y(n_117)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_117),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_45),
.Y(n_118)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_118),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_119),
.Y(n_197)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_39),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_58),
.A2(n_111),
.B1(n_118),
.B2(n_117),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_121),
.A2(n_126),
.B1(n_144),
.B2(n_91),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_28),
.B1(n_54),
.B2(n_53),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_76),
.B(n_55),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_134),
.B(n_162),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_113),
.A2(n_28),
.B1(n_54),
.B2(n_53),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_139),
.A2(n_179),
.B1(n_194),
.B2(n_198),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_141),
.B(n_150),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_101),
.A2(n_55),
.B1(n_42),
.B2(n_39),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g241 ( 
.A1(n_142),
.A2(n_143),
.B1(n_146),
.B2(n_154),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_63),
.A2(n_42),
.B1(n_44),
.B2(n_50),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_72),
.A2(n_52),
.B1(n_20),
.B2(n_50),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_63),
.A2(n_52),
.B1(n_20),
.B2(n_48),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_84),
.B(n_48),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_99),
.B(n_44),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_99),
.B(n_33),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_176),
.B(n_178),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_56),
.B(n_26),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_102),
.A2(n_33),
.B1(n_26),
.B2(n_31),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_73),
.B(n_2),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_189),
.B(n_190),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_78),
.B(n_2),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_119),
.B(n_46),
.C(n_31),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_12),
.C(n_13),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_61),
.A2(n_46),
.B1(n_51),
.B2(n_7),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_SL g195 ( 
.A(n_89),
.Y(n_195)
);

INVx11_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_62),
.B(n_4),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_199),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_109),
.A2(n_46),
.B1(n_51),
.B2(n_7),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_67),
.B(n_4),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_77),
.Y(n_200)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_200),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_202),
.B(n_207),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_195),
.A2(n_88),
.B1(n_107),
.B2(n_114),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_203),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_151),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_205),
.B(n_210),
.Y(n_295)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_137),
.Y(n_206)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_206),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_154),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_171),
.A2(n_94),
.B1(n_90),
.B2(n_105),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_208),
.A2(n_214),
.B1(n_232),
.B2(n_234),
.Y(n_315)
);

A2O1A1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_171),
.A2(n_51),
.B(n_5),
.C(n_8),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_142),
.A2(n_168),
.B1(n_164),
.B2(n_167),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_213),
.A2(n_228),
.B1(n_262),
.B2(n_263),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_139),
.A2(n_51),
.B1(n_5),
.B2(n_9),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_155),
.Y(n_215)
);

INVx6_ASAP7_75t_L g288 ( 
.A(n_215),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_148),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_216),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_153),
.A2(n_4),
.B1(n_9),
.B2(n_10),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_217),
.A2(n_220),
.B1(n_258),
.B2(n_261),
.Y(n_283)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_129),
.Y(n_218)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_218),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_123),
.B(n_9),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_219),
.B(n_267),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_183),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_220)
);

XNOR2x1_ASAP7_75t_L g314 ( 
.A(n_221),
.B(n_228),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_155),
.Y(n_222)
);

INVx6_ASAP7_75t_L g308 ( 
.A(n_222),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_161),
.B(n_16),
.C(n_14),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_223),
.B(n_158),
.C(n_147),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_156),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_224),
.B(n_236),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_184),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_226),
.Y(n_312)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_138),
.Y(n_227)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_227),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_188),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_160),
.Y(n_229)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_229),
.Y(n_291)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_181),
.Y(n_230)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_230),
.Y(n_292)
);

AOI32xp33_ASAP7_75t_L g231 ( 
.A1(n_122),
.A2(n_14),
.A3(n_15),
.B1(n_16),
.B2(n_175),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_231),
.B(n_237),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_194),
.A2(n_163),
.B1(n_145),
.B2(n_136),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_146),
.A2(n_143),
.B1(n_191),
.B2(n_125),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_173),
.Y(n_235)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_235),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_131),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_127),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_175),
.Y(n_238)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_238),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_192),
.Y(n_239)
);

BUFx2_ASAP7_75t_SL g280 ( 
.A(n_239),
.Y(n_280)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_124),
.Y(n_240)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_240),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_241),
.Y(n_287)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_128),
.Y(n_242)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_242),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_181),
.Y(n_243)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_243),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_130),
.B(n_132),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_244),
.Y(n_304)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_133),
.Y(n_246)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_246),
.Y(n_294)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_182),
.Y(n_247)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_247),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_131),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_248),
.B(n_250),
.Y(n_286)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_133),
.Y(n_249)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_249),
.Y(n_307)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_140),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_157),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_251),
.B(n_253),
.Y(n_284)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_140),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_135),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_254),
.B(n_255),
.Y(n_310)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_157),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_151),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_256),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_159),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_257),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_170),
.A2(n_174),
.B1(n_186),
.B2(n_149),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_L g259 ( 
.A1(n_159),
.A2(n_172),
.B1(n_166),
.B2(n_165),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_259),
.A2(n_169),
.B1(n_185),
.B2(n_267),
.Y(n_274)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_165),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_260),
.Y(n_316)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_152),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_177),
.A2(n_197),
.B1(n_201),
.B2(n_149),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_192),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_166),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_265),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_201),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_187),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_266),
.B(n_268),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_180),
.B(n_172),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_180),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_209),
.A2(n_185),
.B(n_187),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_269),
.B(n_314),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_270),
.B(n_247),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_209),
.A2(n_169),
.B1(n_147),
.B2(n_158),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_272),
.A2(n_318),
.B1(n_212),
.B2(n_266),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_274),
.A2(n_284),
.B1(n_310),
.B2(n_293),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_204),
.A2(n_185),
.B1(n_252),
.B2(n_245),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_281),
.A2(n_264),
.B1(n_255),
.B2(n_238),
.Y(n_333)
);

OAI22x1_ASAP7_75t_L g285 ( 
.A1(n_241),
.A2(n_210),
.B1(n_233),
.B2(n_207),
.Y(n_285)
);

OA21x2_ASAP7_75t_L g351 ( 
.A1(n_285),
.A2(n_284),
.B(n_310),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_241),
.A2(n_213),
.B(n_221),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_301),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_204),
.B(n_219),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_309),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_225),
.B(n_223),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_305),
.B(n_218),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_244),
.B(n_242),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_244),
.B(n_240),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_309),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_259),
.A2(n_266),
.B1(n_261),
.B2(n_241),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_290),
.Y(n_319)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_319),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_321),
.B(n_332),
.C(n_306),
.Y(n_358)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_292),
.Y(n_322)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_322),
.Y(n_382)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_290),
.Y(n_323)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_323),
.Y(n_369)
);

INVx5_ASAP7_75t_L g324 ( 
.A(n_288),
.Y(n_324)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_324),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_325),
.B(n_333),
.Y(n_362)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_296),
.Y(n_326)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_326),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_310),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_327),
.B(n_349),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_298),
.B(n_227),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_328),
.B(n_342),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_329),
.A2(n_352),
.B1(n_280),
.B2(n_311),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_301),
.A2(n_216),
.B1(n_260),
.B2(n_251),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g387 ( 
.A1(n_330),
.A2(n_349),
.B1(n_344),
.B2(n_323),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_298),
.B(n_237),
.C(n_226),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_331),
.B(n_348),
.C(n_300),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_282),
.B(n_229),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_334),
.B(n_338),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_287),
.A2(n_211),
.B1(n_257),
.B2(n_215),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_335),
.A2(n_337),
.B1(n_341),
.B2(n_347),
.Y(n_378)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_296),
.Y(n_336)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_336),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_276),
.A2(n_211),
.B1(n_243),
.B2(n_222),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_303),
.B(n_263),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_302),
.B(n_239),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_340),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_276),
.A2(n_235),
.B1(n_230),
.B2(n_212),
.Y(n_341)
);

AO22x1_ASAP7_75t_SL g342 ( 
.A1(n_276),
.A2(n_315),
.B1(n_274),
.B2(n_281),
.Y(n_342)
);

AO22x1_ASAP7_75t_L g343 ( 
.A1(n_269),
.A2(n_285),
.B1(n_275),
.B2(n_304),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_343),
.A2(n_291),
.B(n_311),
.Y(n_373)
);

NAND2x1p5_ASAP7_75t_L g345 ( 
.A(n_314),
.B(n_295),
.Y(n_345)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_345),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_275),
.A2(n_273),
.B1(n_279),
.B2(n_283),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_346),
.A2(n_350),
.B1(n_355),
.B2(n_297),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_279),
.A2(n_270),
.B1(n_317),
.B2(n_286),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_305),
.B(n_299),
.C(n_294),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_284),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_278),
.A2(n_294),
.B1(n_307),
.B2(n_316),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_351),
.B(n_312),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_307),
.B(n_302),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_353),
.B(n_354),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_271),
.B(n_277),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_300),
.A2(n_293),
.B1(n_292),
.B2(n_271),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_277),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_356),
.B(n_289),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_354),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_357),
.B(n_377),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_358),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_359),
.B(n_344),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_360),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_332),
.B(n_291),
.C(n_289),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_364),
.B(n_348),
.C(n_356),
.Y(n_403)
);

A2O1A1Ixp33_ASAP7_75t_L g366 ( 
.A1(n_339),
.A2(n_328),
.B(n_320),
.C(n_345),
.Y(n_366)
);

OA21x2_ASAP7_75t_L g407 ( 
.A1(n_366),
.A2(n_365),
.B(n_361),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_367),
.A2(n_373),
.B(n_385),
.Y(n_412)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_371),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_343),
.A2(n_297),
.B1(n_313),
.B2(n_308),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_376),
.A2(n_385),
.B1(n_341),
.B2(n_335),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_350),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_355),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_379),
.B(n_380),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_326),
.B(n_313),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_383),
.A2(n_351),
.B(n_347),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_343),
.A2(n_288),
.B1(n_308),
.B2(n_312),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_336),
.B(n_319),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_386),
.B(n_387),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_388),
.B(n_396),
.C(n_403),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_389),
.A2(n_393),
.B1(n_404),
.B2(n_378),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_391),
.A2(n_397),
.B(n_400),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_368),
.A2(n_339),
.B1(n_342),
.B2(n_320),
.Y(n_393)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_371),
.Y(n_395)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_395),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_366),
.B(n_331),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_383),
.A2(n_351),
.B(n_345),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_368),
.A2(n_346),
.B1(n_342),
.B2(n_325),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_398),
.A2(n_406),
.B1(n_413),
.B2(n_381),
.Y(n_415)
);

AO21x1_ASAP7_75t_SL g400 ( 
.A1(n_383),
.A2(n_333),
.B(n_337),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_380),
.Y(n_401)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_401),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_357),
.A2(n_322),
.B1(n_324),
.B2(n_387),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_370),
.B(n_386),
.Y(n_405)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_405),
.Y(n_423)
);

AOI322xp5_ASAP7_75t_L g406 ( 
.A1(n_375),
.A2(n_362),
.A3(n_366),
.B1(n_361),
.B2(n_369),
.C1(n_363),
.C2(n_384),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_407),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_365),
.B(n_359),
.C(n_358),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_408),
.B(n_388),
.C(n_403),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_373),
.A2(n_360),
.B(n_377),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_409),
.Y(n_427)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_363),
.Y(n_411)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_411),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_412),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_378),
.A2(n_384),
.B1(n_381),
.B2(n_369),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_415),
.A2(n_421),
.B1(n_432),
.B2(n_399),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_417),
.B(n_433),
.C(n_437),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_388),
.B(n_359),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_418),
.B(n_419),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_408),
.B(n_364),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_396),
.B(n_364),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_420),
.B(n_426),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_408),
.B(n_375),
.Y(n_426)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_411),
.Y(n_428)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_428),
.Y(n_444)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_410),
.Y(n_429)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_429),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_403),
.B(n_370),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_430),
.B(n_402),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_399),
.A2(n_379),
.B1(n_367),
.B2(n_376),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_392),
.B(n_372),
.C(n_362),
.Y(n_433)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_410),
.Y(n_435)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_435),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_391),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_436),
.B(n_409),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_396),
.B(n_374),
.C(n_382),
.Y(n_437)
);

A2O1A1Ixp33_ASAP7_75t_SL g468 ( 
.A1(n_440),
.A2(n_427),
.B(n_431),
.C(n_436),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_418),
.B(n_391),
.C(n_397),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_442),
.B(n_445),
.C(n_456),
.Y(n_459)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_414),
.Y(n_443)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_443),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_416),
.B(n_397),
.C(n_407),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_422),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_446),
.B(n_447),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_423),
.B(n_413),
.Y(n_447)
);

NOR2x1_ASAP7_75t_R g450 ( 
.A(n_431),
.B(n_393),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_450),
.Y(n_464)
);

INVxp67_ASAP7_75t_SL g451 ( 
.A(n_433),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_405),
.Y(n_470)
);

OAI22xp33_ASAP7_75t_SL g452 ( 
.A1(n_421),
.A2(n_390),
.B1(n_398),
.B2(n_401),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_452),
.A2(n_453),
.B1(n_398),
.B2(n_390),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_425),
.B(n_404),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_454),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_455),
.B(n_419),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_416),
.B(n_407),
.C(n_402),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_439),
.B(n_417),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_457),
.B(n_461),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_438),
.B(n_437),
.C(n_426),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_462),
.B(n_465),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_463),
.A2(n_447),
.B1(n_454),
.B2(n_441),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_439),
.B(n_438),
.C(n_445),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_456),
.B(n_430),
.C(n_420),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_467),
.B(n_468),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_449),
.A2(n_434),
.B(n_427),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_469),
.A2(n_441),
.B(n_440),
.Y(n_474)
);

NAND3xp33_ASAP7_75t_L g482 ( 
.A(n_470),
.B(n_446),
.C(n_443),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_459),
.B(n_442),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_471),
.B(n_481),
.Y(n_483)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_460),
.Y(n_472)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_472),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_473),
.A2(n_479),
.B1(n_468),
.B2(n_394),
.Y(n_490)
);

AOI21x1_ASAP7_75t_L g491 ( 
.A1(n_474),
.A2(n_412),
.B(n_466),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_457),
.B(n_448),
.C(n_455),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_478),
.B(n_480),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_458),
.A2(n_454),
.B1(n_434),
.B2(n_407),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_459),
.B(n_374),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_465),
.B(n_448),
.C(n_450),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_481),
.B(n_464),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_482),
.Y(n_485)
);

NOR2xp67_ASAP7_75t_SL g494 ( 
.A(n_483),
.B(n_484),
.Y(n_494)
);

NAND2xp33_ASAP7_75t_R g486 ( 
.A(n_477),
.B(n_464),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_486),
.A2(n_491),
.B(n_492),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_479),
.A2(n_468),
.B(n_406),
.Y(n_487)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_487),
.B(n_490),
.Y(n_496)
);

NOR2x1_ASAP7_75t_L g492 ( 
.A(n_471),
.B(n_394),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_485),
.B(n_476),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_495),
.B(n_497),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_488),
.B(n_473),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_489),
.B(n_492),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_498),
.B(n_500),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_484),
.A2(n_475),
.B(n_468),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_499),
.A2(n_487),
.B(n_491),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_483),
.B(n_475),
.C(n_478),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_502),
.B(n_505),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_496),
.A2(n_490),
.B1(n_389),
.B2(n_444),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_503),
.B(n_504),
.Y(n_507)
);

INVx6_ASAP7_75t_L g504 ( 
.A(n_494),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_500),
.B(n_395),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_505),
.B(n_496),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_509),
.B(n_510),
.C(n_501),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_506),
.B(n_493),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_511),
.A2(n_512),
.B(n_508),
.Y(n_513)
);

AO21x2_ASAP7_75t_L g512 ( 
.A1(n_507),
.A2(n_503),
.B(n_504),
.Y(n_512)
);

BUFx24_ASAP7_75t_SL g514 ( 
.A(n_513),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_514),
.A2(n_508),
.B(n_424),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_515),
.A2(n_382),
.B(n_400),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_400),
.Y(n_517)
);


endmodule