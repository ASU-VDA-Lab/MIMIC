module fake_ariane_1114_n_1918 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1918);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1918;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_699;
wire n_590;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g185 ( 
.A(n_99),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_22),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_79),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_106),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_46),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_6),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_71),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_65),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_0),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_132),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_76),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_56),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_75),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_62),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_112),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_180),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_173),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_154),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_80),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_7),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_56),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_14),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_57),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_171),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_145),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_51),
.Y(n_210)
);

BUFx2_ASAP7_75t_SL g211 ( 
.A(n_152),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_14),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_92),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_134),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_38),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_121),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_96),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_84),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_7),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_2),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_128),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_139),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_63),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_16),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_12),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_71),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_120),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_28),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_135),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_162),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_20),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_10),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_90),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_115),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_55),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_101),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_86),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_142),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_117),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_49),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_21),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_40),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_10),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_37),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_64),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_44),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_45),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_64),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_104),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_158),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_22),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_34),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_131),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_49),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_53),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_11),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_118),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_32),
.Y(n_260)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_165),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_21),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_33),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_1),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_77),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_50),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_13),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_3),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_36),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_127),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_94),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_170),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_167),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_58),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_184),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_141),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_111),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_175),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_52),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_89),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_55),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_114),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_140),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_144),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_164),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_45),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_93),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_72),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_137),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_126),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_78),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_107),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_85),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_13),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_172),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_83),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_136),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_155),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_159),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_0),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_169),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_9),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_35),
.Y(n_303)
);

BUFx2_ASAP7_75t_SL g304 ( 
.A(n_123),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_153),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_52),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_183),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_174),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_138),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_61),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_46),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_8),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_129),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_57),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_133),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_73),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_59),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_48),
.Y(n_318)
);

BUFx2_ASAP7_75t_SL g319 ( 
.A(n_98),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_95),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_38),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_70),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_151),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_28),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_25),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_54),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_67),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_16),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_74),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_157),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_31),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_37),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_36),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_176),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_27),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_103),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_59),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_43),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_108),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_182),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_50),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_116),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_150),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_87),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_35),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_102),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_43),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_17),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_119),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_113),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_105),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_23),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_65),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_178),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_42),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_60),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_88),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_48),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_41),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_156),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_23),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_58),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_24),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_110),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_143),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_124),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_125),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_130),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_91),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_68),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_181),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_168),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_1),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_31),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_194),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_251),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_185),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_185),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_191),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_231),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_199),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_277),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_199),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_285),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_191),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_216),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_209),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_209),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_342),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_214),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_227),
.B(n_2),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_216),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_214),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_215),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_322),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_354),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_212),
.B(n_3),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_267),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_267),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_186),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_230),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_215),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_212),
.B(n_4),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_190),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_192),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_186),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_218),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_360),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_218),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_204),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_360),
.Y(n_411)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_189),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_322),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_219),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_210),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_250),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_237),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_269),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_206),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_221),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_222),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_219),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_327),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_237),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_241),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_241),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_189),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_367),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_270),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_362),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_374),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_R g432 ( 
.A(n_217),
.B(n_122),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_270),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_226),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_228),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_282),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_233),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_367),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_282),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_283),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_243),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_280),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_193),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_280),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_283),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_245),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_329),
.B(n_4),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_284),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_248),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_254),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_284),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_210),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_256),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_257),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_287),
.Y(n_455)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_231),
.Y(n_456)
);

INVxp67_ASAP7_75t_SL g457 ( 
.A(n_205),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_258),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_287),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_262),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_263),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_225),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_225),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_289),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_289),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_341),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_332),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_264),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_329),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_377),
.B(n_378),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_377),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_399),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_378),
.B(n_292),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_401),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_381),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_417),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_381),
.B(n_292),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_417),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_417),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_383),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_424),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_383),
.B(n_332),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_387),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_424),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_424),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_387),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_388),
.Y(n_487)
);

NAND2xp33_ASAP7_75t_R g488 ( 
.A(n_398),
.B(n_404),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_388),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_390),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_399),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_390),
.B(n_297),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_393),
.B(n_193),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_393),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_394),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_466),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_391),
.A2(n_373),
.B1(n_205),
.B2(n_213),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_394),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_380),
.B(n_196),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_402),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_408),
.B(n_275),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_402),
.Y(n_502)
);

INVx5_ASAP7_75t_L g503 ( 
.A(n_380),
.Y(n_503)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_380),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_407),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_407),
.B(n_196),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_409),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_409),
.B(n_414),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_414),
.B(n_297),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_422),
.Y(n_510)
);

OA21x2_ASAP7_75t_L g511 ( 
.A1(n_422),
.A2(n_308),
.B(n_305),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_425),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_425),
.B(n_426),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_466),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_426),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_429),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_429),
.B(n_207),
.Y(n_517)
);

INVx2_ASAP7_75t_SL g518 ( 
.A(n_432),
.Y(n_518)
);

CKINVDCx8_ASAP7_75t_R g519 ( 
.A(n_408),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_433),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_433),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_436),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_442),
.A2(n_352),
.B1(n_328),
.B2(n_370),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_436),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_439),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_444),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_439),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_440),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_440),
.B(n_305),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_385),
.A2(n_373),
.B1(n_213),
.B2(n_234),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_392),
.Y(n_531)
);

BUFx8_ASAP7_75t_L g532 ( 
.A(n_379),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_445),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_416),
.B(n_268),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_445),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_448),
.Y(n_536)
);

INVx6_ASAP7_75t_L g537 ( 
.A(n_456),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_456),
.B(n_308),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_448),
.B(n_207),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_451),
.B(n_242),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_392),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_451),
.Y(n_542)
);

BUFx8_ASAP7_75t_L g543 ( 
.A(n_379),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_455),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_455),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_452),
.B(n_339),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_375),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_459),
.Y(n_548)
);

AND2x2_ASAP7_75t_SL g549 ( 
.A(n_511),
.B(n_447),
.Y(n_549)
);

INVx5_ASAP7_75t_L g550 ( 
.A(n_502),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_502),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_538),
.A2(n_397),
.B1(n_403),
.B2(n_447),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_476),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_476),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_476),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_518),
.B(n_411),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_502),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_484),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_502),
.Y(n_559)
);

NAND3xp33_ASAP7_75t_L g560 ( 
.A(n_546),
.B(n_518),
.C(n_410),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_484),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_503),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_484),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_518),
.B(n_411),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_502),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_504),
.B(n_428),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_479),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_508),
.B(n_428),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_503),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_508),
.B(n_438),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_504),
.B(n_438),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_502),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_508),
.B(n_400),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_L g574 ( 
.A(n_502),
.B(n_261),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_479),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_514),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_508),
.B(n_405),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_514),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_504),
.B(n_419),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_512),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_504),
.B(n_420),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_546),
.A2(n_385),
.B1(n_413),
.B2(n_469),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_512),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_537),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_530),
.A2(n_413),
.B1(n_395),
.B2(n_386),
.Y(n_585)
);

BUFx10_ASAP7_75t_L g586 ( 
.A(n_537),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_512),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_512),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_508),
.B(n_400),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_512),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_512),
.Y(n_591)
);

AND2x6_ASAP7_75t_L g592 ( 
.A(n_513),
.B(n_339),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_513),
.B(n_459),
.Y(n_593)
);

AO22x2_ASAP7_75t_L g594 ( 
.A1(n_530),
.A2(n_391),
.B1(n_412),
.B2(n_406),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_513),
.B(n_421),
.Y(n_595)
);

INVxp33_ASAP7_75t_L g596 ( 
.A(n_491),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_512),
.Y(n_597)
);

NAND3xp33_ASAP7_75t_SL g598 ( 
.A(n_523),
.B(n_435),
.C(n_434),
.Y(n_598)
);

INVxp33_ASAP7_75t_SL g599 ( 
.A(n_547),
.Y(n_599)
);

NAND2xp33_ASAP7_75t_L g600 ( 
.A(n_516),
.B(n_261),
.Y(n_600)
);

INVx5_ASAP7_75t_L g601 ( 
.A(n_516),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_479),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_516),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_479),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_537),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_481),
.Y(n_606)
);

OAI22xp33_ASAP7_75t_L g607 ( 
.A1(n_523),
.A2(n_441),
.B1(n_446),
.B2(n_437),
.Y(n_607)
);

OR2x6_ASAP7_75t_L g608 ( 
.A(n_537),
.B(n_452),
.Y(n_608)
);

OAI22xp33_ASAP7_75t_L g609 ( 
.A1(n_496),
.A2(n_450),
.B1(n_453),
.B2(n_449),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_503),
.Y(n_610)
);

BUFx4f_ASAP7_75t_L g611 ( 
.A(n_516),
.Y(n_611)
);

INVx1_ASAP7_75t_SL g612 ( 
.A(n_472),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_L g613 ( 
.A(n_516),
.B(n_261),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_537),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_503),
.Y(n_615)
);

BUFx10_ASAP7_75t_L g616 ( 
.A(n_513),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_516),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_513),
.B(n_406),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_516),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_472),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_496),
.Y(n_621)
);

NOR3xp33_ASAP7_75t_L g622 ( 
.A(n_497),
.B(n_458),
.C(n_454),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_507),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_501),
.B(n_460),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_507),
.Y(n_625)
);

INVxp33_ASAP7_75t_L g626 ( 
.A(n_491),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_471),
.B(n_461),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_519),
.B(n_468),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_493),
.B(n_412),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_507),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_507),
.B(n_464),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_481),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_519),
.B(n_376),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_471),
.B(n_463),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_490),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_490),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_475),
.B(n_464),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_531),
.Y(n_638)
);

CKINVDCx6p67_ASAP7_75t_R g639 ( 
.A(n_474),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_499),
.A2(n_465),
.B1(n_457),
.B2(n_427),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_475),
.B(n_465),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_519),
.B(n_382),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_481),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_526),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_482),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_490),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_481),
.Y(n_647)
);

NOR2x1p5_ASAP7_75t_L g648 ( 
.A(n_488),
.B(n_427),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_531),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_480),
.B(n_483),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_480),
.B(n_457),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_497),
.A2(n_311),
.B1(n_321),
.B2(n_310),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_493),
.B(n_463),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_494),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_483),
.B(n_443),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_503),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_499),
.A2(n_324),
.B1(n_274),
.B2(n_303),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_485),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_485),
.Y(n_659)
);

AND2x6_ASAP7_75t_L g660 ( 
.A(n_494),
.B(n_344),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_486),
.B(n_443),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_499),
.B(n_415),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_486),
.B(n_384),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_487),
.B(n_299),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_494),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_482),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_500),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_487),
.B(n_365),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_489),
.B(n_396),
.Y(n_669)
);

INVx4_ASAP7_75t_L g670 ( 
.A(n_503),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_500),
.Y(n_671)
);

AND2x2_ASAP7_75t_SL g672 ( 
.A(n_511),
.B(n_275),
.Y(n_672)
);

NAND3xp33_ASAP7_75t_L g673 ( 
.A(n_470),
.B(n_314),
.C(n_312),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_485),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_500),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_489),
.B(n_495),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_515),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_495),
.B(n_498),
.Y(n_678)
);

OAI22xp33_ASAP7_75t_L g679 ( 
.A1(n_541),
.A2(n_325),
.B1(n_335),
.B2(n_361),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_498),
.B(n_462),
.Y(n_680)
);

OAI22xp33_ASAP7_75t_SL g681 ( 
.A1(n_473),
.A2(n_331),
.B1(n_338),
.B2(n_345),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_532),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_515),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_541),
.B(n_467),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_499),
.B(n_234),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_515),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_485),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_478),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_520),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_520),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_520),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_522),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_478),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_503),
.Y(n_694)
);

AND3x1_ASAP7_75t_L g695 ( 
.A(n_470),
.B(n_246),
.C(n_244),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_522),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_478),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_482),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_505),
.B(n_344),
.Y(n_699)
);

NAND3xp33_ASAP7_75t_L g700 ( 
.A(n_505),
.B(n_355),
.C(n_348),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_478),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_552),
.A2(n_521),
.B1(n_545),
.B2(n_544),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_L g703 ( 
.A1(n_552),
.A2(n_510),
.B1(n_545),
.B2(n_544),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_616),
.B(n_510),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_L g705 ( 
.A(n_592),
.B(n_521),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_596),
.B(n_626),
.Y(n_706)
);

INVxp33_ASAP7_75t_L g707 ( 
.A(n_621),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_621),
.B(n_526),
.Y(n_708)
);

BUFx6f_ASAP7_75t_SL g709 ( 
.A(n_608),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_556),
.B(n_389),
.Y(n_710)
);

OR2x2_ASAP7_75t_L g711 ( 
.A(n_612),
.B(n_534),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_623),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_586),
.Y(n_713)
);

A2O1A1Ixp33_ASAP7_75t_L g714 ( 
.A1(n_573),
.A2(n_477),
.B(n_473),
.C(n_509),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_627),
.B(n_573),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_553),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_616),
.B(n_525),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_623),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_573),
.A2(n_525),
.B1(n_542),
.B2(n_536),
.Y(n_719)
);

INVxp67_ASAP7_75t_SL g720 ( 
.A(n_584),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_589),
.B(n_527),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_616),
.B(n_527),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_589),
.B(n_528),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_549),
.B(n_528),
.Y(n_724)
);

AND2x2_ASAP7_75t_SL g725 ( 
.A(n_549),
.B(n_511),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_584),
.B(n_493),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_618),
.B(n_629),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_618),
.B(n_533),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_553),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_549),
.B(n_533),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_L g731 ( 
.A1(n_560),
.A2(n_536),
.B1(n_542),
.B2(n_509),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_554),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_629),
.B(n_522),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_620),
.B(n_532),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_586),
.B(n_524),
.Y(n_735)
);

OAI22xp33_ASAP7_75t_L g736 ( 
.A1(n_652),
.A2(n_492),
.B1(n_529),
.B2(n_477),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_645),
.B(n_524),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_620),
.B(n_532),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_648),
.A2(n_532),
.B1(n_543),
.B2(n_499),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_576),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_554),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_586),
.B(n_524),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_SL g743 ( 
.A(n_599),
.B(n_532),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_623),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_624),
.B(n_543),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_605),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_645),
.B(n_535),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_666),
.B(n_535),
.Y(n_748)
);

INVxp67_ASAP7_75t_L g749 ( 
.A(n_578),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_648),
.A2(n_548),
.B1(n_535),
.B2(n_540),
.Y(n_750)
);

INVx8_ASAP7_75t_L g751 ( 
.A(n_592),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_644),
.Y(n_752)
);

INVxp33_ASAP7_75t_L g753 ( 
.A(n_649),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_625),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_555),
.Y(n_755)
);

OAI22xp33_ASAP7_75t_L g756 ( 
.A1(n_652),
.A2(n_529),
.B1(n_492),
.B2(n_548),
.Y(n_756)
);

INVx8_ASAP7_75t_L g757 ( 
.A(n_592),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_564),
.B(n_543),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_609),
.B(n_548),
.Y(n_759)
);

OAI21xp5_ASAP7_75t_L g760 ( 
.A1(n_672),
.A2(n_511),
.B(n_506),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_666),
.B(n_698),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_555),
.Y(n_762)
);

OAI22xp5_ASAP7_75t_L g763 ( 
.A1(n_593),
.A2(n_356),
.B1(n_358),
.B2(n_300),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_625),
.B(n_539),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_625),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_558),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_605),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_558),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_698),
.B(n_506),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_579),
.B(n_506),
.Y(n_770)
);

OR2x2_ASAP7_75t_SL g771 ( 
.A(n_598),
.B(n_543),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_630),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_649),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_663),
.B(n_543),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_684),
.B(n_534),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_669),
.B(n_418),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_608),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_672),
.A2(n_511),
.B1(n_539),
.B2(n_540),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_581),
.B(n_517),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_630),
.B(n_672),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_630),
.B(n_539),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_651),
.B(n_517),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_664),
.B(n_668),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_582),
.B(n_517),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_690),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_561),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_634),
.B(n_539),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_638),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_676),
.Y(n_789)
);

XOR2xp5_ASAP7_75t_L g790 ( 
.A(n_599),
.B(n_423),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_653),
.B(n_539),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_577),
.B(n_430),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_650),
.B(n_540),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_635),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_678),
.B(n_540),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_592),
.A2(n_540),
.B1(n_237),
.B2(n_242),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_580),
.B(n_346),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_684),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_568),
.A2(n_306),
.B1(n_253),
.B2(n_317),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_561),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_571),
.B(n_680),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_653),
.B(n_431),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_640),
.B(n_614),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_595),
.B(n_244),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_580),
.B(n_346),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_563),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_563),
.Y(n_807)
);

INVx4_ASAP7_75t_L g808 ( 
.A(n_592),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_635),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_614),
.B(n_260),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_690),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_568),
.B(n_260),
.Y(n_812)
);

A2O1A1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_631),
.A2(n_306),
.B(n_266),
.C(n_281),
.Y(n_813)
);

OAI221xp5_ASAP7_75t_L g814 ( 
.A1(n_657),
.A2(n_249),
.B1(n_302),
.B2(n_247),
.C(n_317),
.Y(n_814)
);

AND2x2_ASAP7_75t_SL g815 ( 
.A(n_622),
.B(n_369),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_580),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_566),
.B(n_279),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_690),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_692),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_692),
.Y(n_820)
);

NAND3xp33_ASAP7_75t_L g821 ( 
.A(n_657),
.B(n_372),
.C(n_357),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_580),
.B(n_357),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_655),
.B(n_279),
.Y(n_823)
);

O2A1O1Ixp5_ASAP7_75t_L g824 ( 
.A1(n_611),
.A2(n_372),
.B(n_266),
.C(n_246),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_580),
.B(n_369),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_661),
.B(n_247),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_608),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_692),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_592),
.B(n_249),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_636),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_592),
.B(n_253),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_591),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_637),
.B(n_281),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_591),
.B(n_261),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_608),
.B(n_570),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_636),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_591),
.B(n_261),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_662),
.B(n_286),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_572),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_646),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_662),
.B(n_286),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_572),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_641),
.B(n_294),
.Y(n_843)
);

NAND2xp33_ASAP7_75t_SL g844 ( 
.A(n_628),
.B(n_294),
.Y(n_844)
);

NAND2x1p5_ASAP7_75t_L g845 ( 
.A(n_685),
.B(n_351),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_685),
.A2(n_211),
.B1(n_304),
.B2(n_319),
.Y(n_846)
);

INVx8_ASAP7_75t_L g847 ( 
.A(n_660),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_607),
.B(n_300),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_SL g849 ( 
.A(n_682),
.B(n_351),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_662),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_685),
.Y(n_851)
);

A2O1A1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_646),
.A2(n_326),
.B(n_363),
.C(n_359),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_633),
.B(n_302),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_642),
.B(n_318),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_654),
.B(n_318),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_594),
.B(n_326),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_673),
.B(n_333),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_654),
.B(n_665),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_591),
.B(n_261),
.Y(n_859)
);

INVx5_ASAP7_75t_L g860 ( 
.A(n_591),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_611),
.A2(n_478),
.B(n_200),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_665),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_679),
.B(n_700),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_681),
.B(n_333),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_667),
.B(n_337),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_611),
.B(n_261),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_671),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_695),
.B(n_337),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_671),
.B(n_347),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_572),
.B(n_347),
.Y(n_870)
);

NAND2xp33_ASAP7_75t_L g871 ( 
.A(n_550),
.B(n_261),
.Y(n_871)
);

AOI22xp5_ASAP7_75t_L g872 ( 
.A1(n_675),
.A2(n_211),
.B1(n_304),
.B2(n_319),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_801),
.B(n_675),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_724),
.A2(n_557),
.B(n_551),
.Y(n_874)
);

OR2x6_ASAP7_75t_L g875 ( 
.A(n_751),
.B(n_594),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_715),
.B(n_677),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_774),
.A2(n_594),
.B1(n_686),
.B2(n_691),
.Y(n_877)
);

BUFx8_ASAP7_75t_L g878 ( 
.A(n_708),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_808),
.B(n_550),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_727),
.B(n_677),
.Y(n_880)
);

AO21x1_ASAP7_75t_L g881 ( 
.A1(n_730),
.A2(n_699),
.B(n_686),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_736),
.B(n_683),
.Y(n_882)
);

NOR2x2_ASAP7_75t_L g883 ( 
.A(n_790),
.B(n_594),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_808),
.A2(n_603),
.B1(n_683),
.B2(n_696),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_730),
.A2(n_565),
.B(n_559),
.Y(n_885)
);

AOI21x1_ASAP7_75t_L g886 ( 
.A1(n_866),
.A2(n_691),
.B(n_689),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_780),
.A2(n_565),
.B(n_559),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_783),
.B(n_689),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_789),
.B(n_696),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_760),
.A2(n_587),
.B(n_583),
.Y(n_890)
);

NAND2x1p5_ASAP7_75t_L g891 ( 
.A(n_808),
.B(n_550),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_716),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_713),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_780),
.A2(n_587),
.B(n_583),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_858),
.A2(n_590),
.B(n_588),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_863),
.A2(n_363),
.B(n_353),
.C(n_359),
.Y(n_896)
);

BUFx12f_ASAP7_75t_L g897 ( 
.A(n_752),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_770),
.B(n_585),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_713),
.B(n_550),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_704),
.A2(n_590),
.B(n_588),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_704),
.A2(n_722),
.B(n_717),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_729),
.Y(n_902)
);

INVx1_ASAP7_75t_SL g903 ( 
.A(n_711),
.Y(n_903)
);

OAI21xp5_ASAP7_75t_L g904 ( 
.A1(n_725),
.A2(n_617),
.B(n_597),
.Y(n_904)
);

NAND2xp33_ASAP7_75t_L g905 ( 
.A(n_751),
.B(n_603),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_717),
.A2(n_617),
.B(n_597),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_745),
.B(n_603),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_SL g908 ( 
.A1(n_856),
.A2(n_353),
.B1(n_660),
.B2(n_198),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_791),
.B(n_567),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_722),
.A2(n_779),
.B(n_793),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_725),
.A2(n_619),
.B(n_688),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_795),
.A2(n_619),
.B(n_688),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_705),
.A2(n_697),
.B(n_693),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_756),
.B(n_575),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_734),
.B(n_602),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_705),
.A2(n_697),
.B(n_693),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_794),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_787),
.B(n_602),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_714),
.A2(n_701),
.B(n_606),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_733),
.A2(n_701),
.B(n_600),
.Y(n_920)
);

BUFx2_ASAP7_75t_L g921 ( 
.A(n_773),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_811),
.A2(n_600),
.B(n_574),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_782),
.B(n_604),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_809),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_811),
.A2(n_819),
.B(n_818),
.Y(n_925)
);

OR2x6_ASAP7_75t_L g926 ( 
.A(n_751),
.B(n_639),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_818),
.A2(n_613),
.B(n_574),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_713),
.B(n_550),
.Y(n_928)
);

AOI21xp33_ASAP7_75t_L g929 ( 
.A1(n_776),
.A2(n_606),
.B(n_604),
.Y(n_929)
);

AO21x1_ASAP7_75t_L g930 ( 
.A1(n_848),
.A2(n_613),
.B(n_632),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_819),
.A2(n_601),
.B(n_550),
.Y(n_931)
);

OR2x2_ASAP7_75t_L g932 ( 
.A(n_775),
.B(n_639),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_746),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_721),
.B(n_632),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_723),
.A2(n_658),
.B1(n_687),
.B2(n_674),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_728),
.B(n_738),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_836),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_SL g938 ( 
.A1(n_703),
.A2(n_643),
.B(n_647),
.C(n_658),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_729),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_719),
.A2(n_687),
.B1(n_659),
.B2(n_647),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_798),
.B(n_643),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_820),
.A2(n_601),
.B(n_659),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_726),
.B(n_660),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_SL g944 ( 
.A(n_743),
.B(n_660),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_820),
.A2(n_601),
.B(n_670),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_828),
.A2(n_601),
.B(n_670),
.Y(n_946)
);

NAND2xp33_ASAP7_75t_L g947 ( 
.A(n_751),
.B(n_601),
.Y(n_947)
);

O2A1O1Ixp5_ASAP7_75t_L g948 ( 
.A1(n_759),
.A2(n_569),
.B(n_670),
.C(n_610),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_866),
.A2(n_601),
.B(n_660),
.Y(n_949)
);

INVx1_ASAP7_75t_SL g950 ( 
.A(n_740),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_746),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_828),
.A2(n_610),
.B(n_569),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_713),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_726),
.B(n_660),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_737),
.Y(n_955)
);

AND2x2_ASAP7_75t_SL g956 ( 
.A(n_815),
.B(n_237),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_726),
.B(n_660),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_732),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_816),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_757),
.B(n_562),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_769),
.B(n_198),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_747),
.A2(n_610),
.B(n_569),
.Y(n_962)
);

HB1xp67_ASAP7_75t_L g963 ( 
.A(n_850),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_812),
.B(n_198),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_761),
.B(n_198),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_732),
.Y(n_966)
);

O2A1O1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_764),
.A2(n_694),
.B(n_656),
.C(n_615),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_748),
.A2(n_562),
.B(n_656),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_851),
.B(n_198),
.Y(n_969)
);

OR2x6_ASAP7_75t_L g970 ( 
.A(n_757),
.B(n_615),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_802),
.Y(n_971)
);

INVx4_ASAP7_75t_L g972 ( 
.A(n_757),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_702),
.B(n_237),
.Y(n_973)
);

OAI321xp33_ASAP7_75t_L g974 ( 
.A1(n_814),
.A2(n_237),
.A3(n_478),
.B1(n_320),
.B2(n_9),
.C(n_11),
.Y(n_974)
);

NOR2xp67_ASAP7_75t_L g975 ( 
.A(n_706),
.B(n_710),
.Y(n_975)
);

OAI321xp33_ASAP7_75t_L g976 ( 
.A1(n_821),
.A2(n_478),
.A3(n_320),
.B1(n_8),
.B2(n_12),
.C(n_15),
.Y(n_976)
);

INVx2_ASAP7_75t_SL g977 ( 
.A(n_788),
.Y(n_977)
);

OAI21xp33_ASAP7_75t_L g978 ( 
.A1(n_753),
.A2(n_371),
.B(n_187),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_735),
.A2(n_368),
.B(n_366),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_757),
.A2(n_364),
.B1(n_350),
.B2(n_349),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_835),
.B(n_188),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_707),
.B(n_5),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_815),
.B(n_261),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_817),
.B(n_838),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_735),
.A2(n_343),
.B(n_340),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_841),
.B(n_195),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_764),
.A2(n_5),
.B(n_6),
.C(n_15),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_804),
.B(n_197),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_742),
.A2(n_336),
.B(n_334),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_742),
.A2(n_330),
.B(n_323),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_830),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_830),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_839),
.A2(n_271),
.B(n_316),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_840),
.Y(n_994)
);

AOI222xp33_ASAP7_75t_L g995 ( 
.A1(n_784),
.A2(n_265),
.B1(n_315),
.B2(n_313),
.C1(n_309),
.C2(n_307),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_839),
.A2(n_252),
.B(n_301),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_777),
.B(n_201),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_839),
.A2(n_255),
.B(n_298),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_707),
.B(n_17),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_827),
.B(n_202),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_741),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_753),
.B(n_18),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_816),
.B(n_320),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_842),
.A2(n_240),
.B(n_296),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_712),
.A2(n_239),
.B(n_295),
.Y(n_1005)
);

AO21x1_ASAP7_75t_L g1006 ( 
.A1(n_759),
.A2(n_825),
.B(n_834),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_857),
.B(n_203),
.Y(n_1007)
);

NOR2xp67_ASAP7_75t_L g1008 ( 
.A(n_749),
.B(n_208),
.Y(n_1008)
);

BUFx3_ASAP7_75t_L g1009 ( 
.A(n_767),
.Y(n_1009)
);

INVx1_ASAP7_75t_SL g1010 ( 
.A(n_849),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_750),
.B(n_823),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_718),
.A2(n_259),
.B(n_293),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_803),
.B(n_220),
.Y(n_1013)
);

AOI21xp33_ASAP7_75t_L g1014 ( 
.A1(n_853),
.A2(n_272),
.B(n_291),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_842),
.A2(n_754),
.B(n_772),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_778),
.A2(n_238),
.B1(n_290),
.B2(n_288),
.Y(n_1016)
);

OAI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_744),
.A2(n_235),
.B(n_278),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_842),
.A2(n_232),
.B(n_276),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_758),
.B(n_273),
.Y(n_1019)
);

INVx1_ASAP7_75t_SL g1020 ( 
.A(n_844),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_792),
.B(n_18),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_854),
.B(n_236),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_846),
.A2(n_765),
.B1(n_785),
.B2(n_781),
.Y(n_1023)
);

NAND2x1_ASAP7_75t_L g1024 ( 
.A(n_785),
.B(n_320),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_868),
.B(n_19),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_840),
.A2(n_229),
.B(n_224),
.Y(n_1026)
);

AOI21xp33_ASAP7_75t_L g1027 ( 
.A1(n_799),
.A2(n_223),
.B(n_320),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_862),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_862),
.A2(n_867),
.B(n_781),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_826),
.B(n_19),
.Y(n_1030)
);

OAI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_837),
.A2(n_320),
.B(n_179),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_833),
.B(n_20),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_843),
.B(n_24),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_785),
.A2(n_720),
.B(n_731),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_SL g1035 ( 
.A(n_709),
.B(n_25),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_855),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_816),
.Y(n_1037)
);

INVx4_ASAP7_75t_L g1038 ( 
.A(n_767),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_816),
.A2(n_166),
.B(n_161),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_741),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_832),
.A2(n_160),
.B(n_149),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_755),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_832),
.A2(n_148),
.B(n_147),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_829),
.B(n_831),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_864),
.A2(n_870),
.B(n_872),
.C(n_813),
.Y(n_1045)
);

OR2x2_ASAP7_75t_L g1046 ( 
.A(n_763),
.B(n_26),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_832),
.B(n_26),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_832),
.A2(n_146),
.B(n_109),
.Y(n_1048)
);

INVxp67_ASAP7_75t_L g1049 ( 
.A(n_709),
.Y(n_1049)
);

NAND3xp33_ASAP7_75t_SL g1050 ( 
.A(n_813),
.B(n_739),
.C(n_844),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_709),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_762),
.A2(n_100),
.B(n_97),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_868),
.Y(n_1053)
);

NOR3xp33_ASAP7_75t_L g1054 ( 
.A(n_852),
.B(n_27),
.C(n_29),
.Y(n_1054)
);

INVx4_ASAP7_75t_L g1055 ( 
.A(n_847),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_865),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_762),
.A2(n_82),
.B(n_81),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_950),
.B(n_845),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_917),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_936),
.A2(n_871),
.B(n_859),
.Y(n_1060)
);

INVx5_ASAP7_75t_L g1061 ( 
.A(n_970),
.Y(n_1061)
);

NOR3xp33_ASAP7_75t_L g1062 ( 
.A(n_1021),
.B(n_852),
.C(n_824),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_898),
.B(n_845),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_975),
.A2(n_868),
.B1(n_796),
.B2(n_810),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_921),
.B(n_860),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_878),
.Y(n_1066)
);

NOR3xp33_ASAP7_75t_L g1067 ( 
.A(n_1050),
.B(n_869),
.C(n_797),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_873),
.A2(n_882),
.B(n_907),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_878),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_892),
.Y(n_1070)
);

AOI21xp33_ASAP7_75t_L g1071 ( 
.A1(n_877),
.A2(n_805),
.B(n_797),
.Y(n_1071)
);

NOR3xp33_ASAP7_75t_SL g1072 ( 
.A(n_1002),
.B(n_822),
.C(n_805),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_880),
.A2(n_860),
.B1(n_847),
.B2(n_771),
.Y(n_1073)
);

AO21x1_ASAP7_75t_L g1074 ( 
.A1(n_983),
.A2(n_825),
.B(n_822),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_888),
.B(n_806),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_977),
.B(n_860),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_955),
.B(n_806),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_924),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_1020),
.B(n_956),
.Y(n_1079)
);

O2A1O1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_1046),
.A2(n_807),
.B(n_800),
.C(n_786),
.Y(n_1080)
);

O2A1O1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_896),
.A2(n_807),
.B(n_800),
.C(n_786),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_902),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_959),
.Y(n_1083)
);

AO32x2_ASAP7_75t_L g1084 ( 
.A1(n_1023),
.A2(n_768),
.A3(n_766),
.B1(n_847),
.B2(n_33),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1036),
.B(n_768),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1056),
.B(n_766),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_937),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_926),
.B(n_847),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_889),
.A2(n_861),
.B1(n_30),
.B2(n_32),
.Y(n_1089)
);

AO32x2_ASAP7_75t_L g1090 ( 
.A1(n_935),
.A2(n_29),
.A3(n_30),
.B1(n_34),
.B2(n_39),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_956),
.B(n_39),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_896),
.A2(n_40),
.B(n_41),
.C(n_42),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_947),
.A2(n_44),
.B(n_47),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_905),
.A2(n_47),
.B(n_51),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_1053),
.B(n_53),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_926),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_910),
.B(n_54),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_SL g1098 ( 
.A1(n_1005),
.A2(n_60),
.B(n_61),
.C(n_62),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_1045),
.A2(n_63),
.B(n_66),
.C(n_67),
.Y(n_1099)
);

O2A1O1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_1045),
.A2(n_1030),
.B(n_982),
.C(n_1032),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_876),
.B(n_66),
.Y(n_1101)
);

OAI21xp33_ASAP7_75t_SL g1102 ( 
.A1(n_1033),
.A2(n_68),
.B(n_69),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_971),
.A2(n_69),
.B1(n_70),
.B2(n_1050),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_915),
.A2(n_914),
.B1(n_988),
.B2(n_1007),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_939),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_915),
.A2(n_901),
.B(n_982),
.C(n_974),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_R g1107 ( 
.A(n_1035),
.B(n_1009),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_1002),
.A2(n_1022),
.B(n_1011),
.C(n_984),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_971),
.B(n_963),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_938),
.A2(n_1034),
.B(n_934),
.Y(n_1110)
);

INVx1_ASAP7_75t_SL g1111 ( 
.A(n_903),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_941),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_958),
.Y(n_1113)
);

NOR3xp33_ASAP7_75t_SL g1114 ( 
.A(n_978),
.B(n_1047),
.C(n_987),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_991),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_893),
.B(n_953),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_932),
.B(n_963),
.Y(n_1117)
);

INVx2_ASAP7_75t_SL g1118 ( 
.A(n_1051),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_1047),
.A2(n_1014),
.B(n_1054),
.C(n_983),
.Y(n_1119)
);

O2A1O1Ixp5_ASAP7_75t_SL g1120 ( 
.A1(n_1003),
.A2(n_929),
.B(n_964),
.C(n_1027),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_919),
.A2(n_886),
.B(n_874),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1019),
.A2(n_972),
.B1(n_909),
.B2(n_1055),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_976),
.A2(n_1029),
.B(n_1031),
.C(n_1026),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_972),
.A2(n_909),
.B1(n_1055),
.B2(n_904),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_943),
.A2(n_954),
.B1(n_957),
.B2(n_918),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_992),
.B(n_994),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_R g1127 ( 
.A(n_1009),
.B(n_944),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_945),
.A2(n_946),
.B(n_913),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_926),
.Y(n_1129)
);

AO21x1_ASAP7_75t_L g1130 ( 
.A1(n_973),
.A2(n_911),
.B(n_1003),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_875),
.A2(n_995),
.B1(n_908),
.B2(n_1025),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1010),
.A2(n_981),
.B1(n_1008),
.B2(n_999),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_966),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_959),
.Y(n_1134)
);

INVx4_ASAP7_75t_L g1135 ( 
.A(n_893),
.Y(n_1135)
);

AOI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_986),
.A2(n_1016),
.B1(n_875),
.B2(n_1054),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1028),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_997),
.B(n_1000),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_1049),
.B(n_1038),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_SL g1140 ( 
.A1(n_875),
.A2(n_908),
.B1(n_1049),
.B2(n_883),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_923),
.B(n_1044),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_916),
.A2(n_962),
.B(n_912),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_884),
.A2(n_951),
.B1(n_933),
.B2(n_1038),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1001),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_890),
.A2(n_895),
.B(n_925),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_1040),
.A2(n_1042),
.B1(n_1051),
.B2(n_1013),
.Y(n_1146)
);

INVx2_ASAP7_75t_SL g1147 ( 
.A(n_933),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_1012),
.A2(n_1017),
.B1(n_980),
.B2(n_951),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_959),
.B(n_1037),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_922),
.A2(n_927),
.B(n_1015),
.C(n_967),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_893),
.B(n_953),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_893),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_R g1153 ( 
.A(n_953),
.B(n_959),
.Y(n_1153)
);

NOR2xp67_ASAP7_75t_L g1154 ( 
.A(n_979),
.B(n_985),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_953),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_1037),
.Y(n_1156)
);

AOI221x1_ASAP7_75t_L g1157 ( 
.A1(n_885),
.A2(n_887),
.B1(n_894),
.B2(n_920),
.C(n_961),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_1037),
.B(n_989),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_SL g1159 ( 
.A1(n_879),
.A2(n_928),
.B(n_899),
.C(n_960),
.Y(n_1159)
);

BUFx12f_ASAP7_75t_L g1160 ( 
.A(n_1037),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_969),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_938),
.A2(n_942),
.B(n_931),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_952),
.A2(n_968),
.B(n_906),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_948),
.A2(n_900),
.B(n_940),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_965),
.A2(n_996),
.B(n_993),
.C(n_1018),
.Y(n_1165)
);

OAI21xp33_ASAP7_75t_L g1166 ( 
.A1(n_998),
.A2(n_1004),
.B(n_990),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_970),
.B(n_899),
.Y(n_1167)
);

NAND3xp33_ASAP7_75t_SL g1168 ( 
.A(n_1039),
.B(n_1041),
.C(n_1043),
.Y(n_1168)
);

INVx6_ASAP7_75t_L g1169 ( 
.A(n_970),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_879),
.A2(n_928),
.B(n_948),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_949),
.A2(n_960),
.B(n_1024),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_891),
.A2(n_1057),
.B(n_1052),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_891),
.B(n_1048),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_910),
.A2(n_936),
.B(n_801),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_975),
.B(n_950),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_888),
.B(n_873),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_888),
.B(n_873),
.Y(n_1177)
);

NAND3xp33_ASAP7_75t_SL g1178 ( 
.A(n_1021),
.B(n_547),
.C(n_776),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_936),
.A2(n_873),
.B(n_715),
.Y(n_1179)
);

O2A1O1Ixp5_ASAP7_75t_SL g1180 ( 
.A1(n_1047),
.A2(n_983),
.B(n_1003),
.C(n_759),
.Y(n_1180)
);

BUFx10_ASAP7_75t_L g1181 ( 
.A(n_982),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_888),
.B(n_873),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_888),
.B(n_873),
.Y(n_1183)
);

INVx4_ASAP7_75t_L g1184 ( 
.A(n_926),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_950),
.B(n_599),
.Y(n_1185)
);

OR2x2_ASAP7_75t_L g1186 ( 
.A(n_903),
.B(n_612),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_897),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_888),
.B(n_873),
.Y(n_1188)
);

OR2x2_ASAP7_75t_L g1189 ( 
.A(n_903),
.B(n_612),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_936),
.A2(n_873),
.B(n_715),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_936),
.A2(n_873),
.B(n_715),
.Y(n_1191)
);

BUFx12f_ASAP7_75t_L g1192 ( 
.A(n_897),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_950),
.B(n_599),
.Y(n_1193)
);

BUFx3_ASAP7_75t_L g1194 ( 
.A(n_897),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_888),
.B(n_873),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_888),
.B(n_873),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_936),
.A2(n_715),
.B1(n_801),
.B2(n_552),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_917),
.Y(n_1198)
);

AOI21x1_ASAP7_75t_L g1199 ( 
.A1(n_930),
.A2(n_881),
.B(n_961),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_936),
.A2(n_873),
.B(n_715),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_917),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_936),
.A2(n_715),
.B1(n_801),
.B2(n_552),
.Y(n_1202)
);

INVx3_ASAP7_75t_L g1203 ( 
.A(n_1055),
.Y(n_1203)
);

O2A1O1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_936),
.A2(n_801),
.B(n_715),
.C(n_776),
.Y(n_1204)
);

OA22x2_ASAP7_75t_L g1205 ( 
.A1(n_875),
.A2(n_652),
.B1(n_497),
.B2(n_391),
.Y(n_1205)
);

O2A1O1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_936),
.A2(n_801),
.B(n_715),
.C(n_776),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_975),
.B(n_950),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_975),
.B(n_950),
.Y(n_1208)
);

INVx4_ASAP7_75t_L g1209 ( 
.A(n_926),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_950),
.B(n_599),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_897),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_888),
.B(n_873),
.Y(n_1212)
);

INVx2_ASAP7_75t_SL g1213 ( 
.A(n_1187),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1176),
.B(n_1177),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1128),
.A2(n_1142),
.B(n_1163),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1068),
.A2(n_1174),
.B(n_1190),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1059),
.Y(n_1217)
);

O2A1O1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_1197),
.A2(n_1202),
.B(n_1204),
.C(n_1206),
.Y(n_1218)
);

INVx3_ASAP7_75t_SL g1219 ( 
.A(n_1211),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1191),
.A2(n_1200),
.B(n_1179),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_1192),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1078),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1106),
.A2(n_1100),
.B(n_1123),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1121),
.A2(n_1162),
.B(n_1145),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1194),
.Y(n_1225)
);

OA21x2_ASAP7_75t_L g1226 ( 
.A1(n_1110),
.A2(n_1157),
.B(n_1164),
.Y(n_1226)
);

OAI22x1_ASAP7_75t_L g1227 ( 
.A1(n_1103),
.A2(n_1136),
.B1(n_1132),
.B2(n_1058),
.Y(n_1227)
);

AOI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1170),
.A2(n_1097),
.B(n_1172),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1108),
.A2(n_1119),
.B(n_1138),
.C(n_1063),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1176),
.B(n_1177),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1182),
.B(n_1183),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1087),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1109),
.B(n_1117),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1114),
.A2(n_1179),
.B(n_1104),
.C(n_1072),
.Y(n_1234)
);

OAI22x1_ASAP7_75t_L g1235 ( 
.A1(n_1095),
.A2(n_1205),
.B1(n_1118),
.B2(n_1091),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1171),
.A2(n_1173),
.B(n_1180),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1182),
.A2(n_1212),
.B(n_1196),
.Y(n_1237)
);

BUFx10_ASAP7_75t_L g1238 ( 
.A(n_1185),
.Y(n_1238)
);

BUFx12f_ASAP7_75t_L g1239 ( 
.A(n_1069),
.Y(n_1239)
);

INVx4_ASAP7_75t_L g1240 ( 
.A(n_1160),
.Y(n_1240)
);

BUFx10_ASAP7_75t_L g1241 ( 
.A(n_1193),
.Y(n_1241)
);

CKINVDCx8_ASAP7_75t_R g1242 ( 
.A(n_1210),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1183),
.A2(n_1212),
.B(n_1196),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1168),
.A2(n_1097),
.B(n_1120),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1082),
.Y(n_1245)
);

AOI221xp5_ASAP7_75t_L g1246 ( 
.A1(n_1092),
.A2(n_1178),
.B1(n_1099),
.B2(n_1102),
.C(n_1131),
.Y(n_1246)
);

INVx4_ASAP7_75t_L g1247 ( 
.A(n_1152),
.Y(n_1247)
);

AOI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1205),
.A2(n_1181),
.B1(n_1175),
.B2(n_1207),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1112),
.B(n_1186),
.Y(n_1249)
);

O2A1O1Ixp33_ASAP7_75t_SL g1250 ( 
.A1(n_1188),
.A2(n_1195),
.B(n_1101),
.C(n_1098),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1189),
.B(n_1181),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1198),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1188),
.B(n_1195),
.Y(n_1253)
);

AO32x2_ASAP7_75t_L g1254 ( 
.A1(n_1140),
.A2(n_1089),
.A3(n_1125),
.B1(n_1073),
.B2(n_1143),
.Y(n_1254)
);

AOI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1158),
.A2(n_1060),
.B(n_1154),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1141),
.B(n_1075),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1141),
.B(n_1075),
.Y(n_1257)
);

AO32x2_ASAP7_75t_L g1258 ( 
.A1(n_1096),
.A2(n_1209),
.A3(n_1184),
.B1(n_1124),
.B2(n_1084),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1150),
.A2(n_1165),
.B(n_1159),
.Y(n_1259)
);

AOI221xp5_ASAP7_75t_SL g1260 ( 
.A1(n_1101),
.A2(n_1094),
.B1(n_1093),
.B2(n_1148),
.C(n_1166),
.Y(n_1260)
);

OA21x2_ASAP7_75t_L g1261 ( 
.A1(n_1071),
.A2(n_1161),
.B(n_1067),
.Y(n_1261)
);

INVx3_ASAP7_75t_L g1262 ( 
.A(n_1088),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1149),
.A2(n_1122),
.B(n_1077),
.Y(n_1263)
);

AOI31xp67_ASAP7_75t_L g1264 ( 
.A1(n_1116),
.A2(n_1149),
.A3(n_1079),
.B(n_1126),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1071),
.A2(n_1111),
.B1(n_1062),
.B2(n_1133),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1081),
.A2(n_1080),
.B(n_1126),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1064),
.A2(n_1146),
.B(n_1201),
.C(n_1139),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1085),
.A2(n_1086),
.B(n_1077),
.Y(n_1268)
);

AOI21xp33_ASAP7_75t_L g1269 ( 
.A1(n_1085),
.A2(n_1086),
.B(n_1115),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1151),
.A2(n_1203),
.B(n_1076),
.Y(n_1270)
);

OR2x2_ASAP7_75t_L g1271 ( 
.A(n_1208),
.B(n_1137),
.Y(n_1271)
);

INVx6_ASAP7_75t_L g1272 ( 
.A(n_1096),
.Y(n_1272)
);

OAI22x1_ASAP7_75t_L g1273 ( 
.A1(n_1129),
.A2(n_1209),
.B1(n_1184),
.B2(n_1065),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1105),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1113),
.B(n_1144),
.Y(n_1275)
);

INVxp67_ASAP7_75t_SL g1276 ( 
.A(n_1083),
.Y(n_1276)
);

AO31x2_ASAP7_75t_L g1277 ( 
.A1(n_1084),
.A2(n_1156),
.A3(n_1135),
.B(n_1090),
.Y(n_1277)
);

INVx1_ASAP7_75t_SL g1278 ( 
.A(n_1127),
.Y(n_1278)
);

BUFx10_ASAP7_75t_L g1279 ( 
.A(n_1083),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1083),
.A2(n_1134),
.B(n_1088),
.Y(n_1280)
);

O2A1O1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_1147),
.A2(n_1066),
.B(n_1155),
.C(n_1090),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1061),
.A2(n_1153),
.B(n_1134),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1169),
.Y(n_1283)
);

AO31x2_ASAP7_75t_L g1284 ( 
.A1(n_1135),
.A2(n_1090),
.A3(n_1061),
.B(n_1134),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1061),
.A2(n_1169),
.B(n_1107),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1169),
.A2(n_1068),
.B(n_1174),
.Y(n_1286)
);

OA21x2_ASAP7_75t_L g1287 ( 
.A1(n_1110),
.A2(n_1142),
.B(n_1157),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1106),
.A2(n_1100),
.B(n_1123),
.Y(n_1288)
);

INVx3_ASAP7_75t_L g1289 ( 
.A(n_1088),
.Y(n_1289)
);

INVx2_ASAP7_75t_SL g1290 ( 
.A(n_1187),
.Y(n_1290)
);

CKINVDCx16_ASAP7_75t_R g1291 ( 
.A(n_1066),
.Y(n_1291)
);

O2A1O1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1197),
.A2(n_801),
.B(n_1202),
.C(n_1204),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1059),
.Y(n_1293)
);

AND2x6_ASAP7_75t_L g1294 ( 
.A(n_1088),
.B(n_1167),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1109),
.B(n_621),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1070),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1059),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1176),
.B(n_1177),
.Y(n_1298)
);

CKINVDCx11_ASAP7_75t_R g1299 ( 
.A(n_1066),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1176),
.B(n_1177),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1128),
.A2(n_1142),
.B(n_1163),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1160),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1185),
.B(n_599),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_SL g1304 ( 
.A1(n_1205),
.A2(n_774),
.B1(n_532),
.B2(n_543),
.Y(n_1304)
);

HB1xp67_ASAP7_75t_L g1305 ( 
.A(n_1109),
.Y(n_1305)
);

AOI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1185),
.A2(n_776),
.B1(n_774),
.B2(n_745),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1088),
.B(n_926),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1070),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1068),
.A2(n_1174),
.B(n_1190),
.Y(n_1309)
);

BUFx10_ASAP7_75t_L g1310 ( 
.A(n_1185),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1070),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1068),
.A2(n_1174),
.B(n_1190),
.Y(n_1312)
);

O2A1O1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1197),
.A2(n_801),
.B(n_1202),
.C(n_1204),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1128),
.A2(n_1142),
.B(n_1163),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1128),
.A2(n_1142),
.B(n_1163),
.Y(n_1315)
);

BUFx10_ASAP7_75t_L g1316 ( 
.A(n_1185),
.Y(n_1316)
);

AOI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1199),
.A2(n_1110),
.B(n_1162),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1106),
.A2(n_1100),
.B(n_1123),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1068),
.A2(n_1174),
.B(n_1190),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1106),
.A2(n_1100),
.B(n_1123),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1128),
.A2(n_1142),
.B(n_1163),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_1111),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1068),
.A2(n_1174),
.B(n_1190),
.Y(n_1323)
);

A2O1A1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1204),
.A2(n_1206),
.B(n_774),
.C(n_1100),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1160),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1176),
.B(n_1177),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1059),
.Y(n_1327)
);

AO32x2_ASAP7_75t_L g1328 ( 
.A1(n_1140),
.A2(n_1202),
.A3(n_1197),
.B1(n_1104),
.B2(n_703),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1070),
.Y(n_1329)
);

A2O1A1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1204),
.A2(n_1206),
.B(n_774),
.C(n_1100),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1128),
.A2(n_1142),
.B(n_1163),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1068),
.A2(n_1174),
.B(n_1190),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1068),
.A2(n_1174),
.B(n_1190),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1088),
.Y(n_1334)
);

BUFx2_ASAP7_75t_L g1335 ( 
.A(n_1107),
.Y(n_1335)
);

A2O1A1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1204),
.A2(n_1206),
.B(n_774),
.C(n_1100),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1068),
.A2(n_1174),
.B(n_1190),
.Y(n_1337)
);

INVxp67_ASAP7_75t_SL g1338 ( 
.A(n_1109),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1068),
.A2(n_1174),
.B(n_1190),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1070),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1109),
.B(n_621),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1128),
.A2(n_1142),
.B(n_1163),
.Y(n_1342)
);

OA21x2_ASAP7_75t_L g1343 ( 
.A1(n_1110),
.A2(n_1142),
.B(n_1157),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1068),
.A2(n_1174),
.B(n_1190),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_1160),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1128),
.A2(n_1142),
.B(n_1163),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1068),
.A2(n_1174),
.B(n_1190),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1068),
.A2(n_1174),
.B(n_1190),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1192),
.Y(n_1349)
);

NOR3xp33_ASAP7_75t_L g1350 ( 
.A(n_1178),
.B(n_776),
.C(n_774),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1197),
.A2(n_1202),
.B1(n_1176),
.B2(n_1182),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1205),
.A2(n_776),
.B1(n_594),
.B2(n_774),
.Y(n_1352)
);

NAND2x1_ASAP7_75t_L g1353 ( 
.A(n_1203),
.B(n_1135),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1068),
.A2(n_1174),
.B(n_1190),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1106),
.A2(n_1100),
.B(n_1123),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1176),
.B(n_1177),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1128),
.A2(n_1142),
.B(n_1163),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1128),
.A2(n_1142),
.B(n_1163),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1110),
.A2(n_1142),
.B(n_1157),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1176),
.B(n_1177),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1059),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1186),
.B(n_1189),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1128),
.A2(n_1142),
.B(n_1163),
.Y(n_1363)
);

OAI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1106),
.A2(n_1100),
.B(n_1123),
.Y(n_1364)
);

OAI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1106),
.A2(n_1100),
.B(n_1123),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1176),
.B(n_1177),
.Y(n_1366)
);

O2A1O1Ixp33_ASAP7_75t_SL g1367 ( 
.A1(n_1197),
.A2(n_1202),
.B(n_1106),
.C(n_1177),
.Y(n_1367)
);

AO31x2_ASAP7_75t_L g1368 ( 
.A1(n_1130),
.A2(n_881),
.A3(n_1074),
.B(n_1006),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1109),
.B(n_621),
.Y(n_1369)
);

CKINVDCx8_ASAP7_75t_R g1370 ( 
.A(n_1291),
.Y(n_1370)
);

CKINVDCx11_ASAP7_75t_R g1371 ( 
.A(n_1299),
.Y(n_1371)
);

INVx4_ASAP7_75t_L g1372 ( 
.A(n_1302),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1351),
.B(n_1237),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1217),
.Y(n_1374)
);

INVx8_ASAP7_75t_L g1375 ( 
.A(n_1239),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1338),
.Y(n_1376)
);

BUFx2_ASAP7_75t_L g1377 ( 
.A(n_1305),
.Y(n_1377)
);

OAI22xp33_ASAP7_75t_SL g1378 ( 
.A1(n_1306),
.A2(n_1351),
.B1(n_1214),
.B2(n_1298),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_SL g1379 ( 
.A1(n_1242),
.A2(n_1352),
.B1(n_1304),
.B2(n_1303),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1235),
.A2(n_1246),
.B1(n_1227),
.B2(n_1350),
.Y(n_1380)
);

AOI22xp5_ASAP7_75t_SL g1381 ( 
.A1(n_1328),
.A2(n_1294),
.B1(n_1320),
.B2(n_1318),
.Y(n_1381)
);

BUFx10_ASAP7_75t_L g1382 ( 
.A(n_1221),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1222),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1349),
.Y(n_1384)
);

INVx3_ASAP7_75t_SL g1385 ( 
.A(n_1219),
.Y(n_1385)
);

BUFx8_ASAP7_75t_SL g1386 ( 
.A(n_1225),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1246),
.A2(n_1265),
.B1(n_1237),
.B2(n_1243),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1232),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1233),
.B(n_1362),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1230),
.A2(n_1300),
.B1(n_1366),
.B2(n_1253),
.Y(n_1390)
);

CKINVDCx6p67_ASAP7_75t_R g1391 ( 
.A(n_1238),
.Y(n_1391)
);

BUFx6f_ASAP7_75t_SL g1392 ( 
.A(n_1302),
.Y(n_1392)
);

INVx5_ASAP7_75t_L g1393 ( 
.A(n_1294),
.Y(n_1393)
);

BUFx4_ASAP7_75t_R g1394 ( 
.A(n_1238),
.Y(n_1394)
);

AOI22xp5_ASAP7_75t_SL g1395 ( 
.A1(n_1328),
.A2(n_1294),
.B1(n_1365),
.B2(n_1364),
.Y(n_1395)
);

BUFx12f_ASAP7_75t_L g1396 ( 
.A(n_1335),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_SL g1397 ( 
.A1(n_1248),
.A2(n_1278),
.B1(n_1213),
.B2(n_1290),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1241),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1230),
.A2(n_1300),
.B1(n_1326),
.B2(n_1253),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1292),
.A2(n_1313),
.B1(n_1234),
.B2(n_1218),
.Y(n_1400)
);

BUFx8_ASAP7_75t_L g1401 ( 
.A(n_1302),
.Y(n_1401)
);

INVx6_ASAP7_75t_L g1402 ( 
.A(n_1325),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1252),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1256),
.B(n_1257),
.Y(n_1404)
);

BUFx10_ASAP7_75t_L g1405 ( 
.A(n_1325),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1231),
.A2(n_1326),
.B1(n_1356),
.B2(n_1360),
.Y(n_1406)
);

OAI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1231),
.A2(n_1356),
.B1(n_1360),
.B2(n_1278),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_1241),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1324),
.A2(n_1336),
.B1(n_1330),
.B2(n_1229),
.Y(n_1409)
);

OAI22xp33_ASAP7_75t_SL g1410 ( 
.A1(n_1328),
.A2(n_1256),
.B1(n_1257),
.B2(n_1320),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1293),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1245),
.A2(n_1311),
.B1(n_1308),
.B2(n_1296),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1295),
.B(n_1341),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1297),
.Y(n_1414)
);

CKINVDCx11_ASAP7_75t_R g1415 ( 
.A(n_1310),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1329),
.A2(n_1340),
.B1(n_1274),
.B2(n_1249),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_SL g1417 ( 
.A1(n_1223),
.A2(n_1288),
.B1(n_1365),
.B2(n_1364),
.Y(n_1417)
);

INVx6_ASAP7_75t_L g1418 ( 
.A(n_1345),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1327),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1223),
.A2(n_1288),
.B1(n_1355),
.B2(n_1318),
.Y(n_1420)
);

INVx2_ASAP7_75t_SL g1421 ( 
.A(n_1345),
.Y(n_1421)
);

INVx4_ASAP7_75t_L g1422 ( 
.A(n_1345),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1310),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1361),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1275),
.Y(n_1425)
);

OAI22xp33_ASAP7_75t_R g1426 ( 
.A1(n_1271),
.A2(n_1322),
.B1(n_1316),
.B2(n_1367),
.Y(n_1426)
);

CKINVDCx20_ASAP7_75t_R g1427 ( 
.A(n_1316),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1355),
.A2(n_1261),
.B1(n_1369),
.B2(n_1294),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1275),
.Y(n_1429)
);

BUFx4_ASAP7_75t_R g1430 ( 
.A(n_1279),
.Y(n_1430)
);

CKINVDCx11_ASAP7_75t_R g1431 ( 
.A(n_1247),
.Y(n_1431)
);

BUFx12f_ASAP7_75t_L g1432 ( 
.A(n_1240),
.Y(n_1432)
);

BUFx10_ASAP7_75t_L g1433 ( 
.A(n_1272),
.Y(n_1433)
);

INVx2_ASAP7_75t_SL g1434 ( 
.A(n_1240),
.Y(n_1434)
);

BUFx12f_ASAP7_75t_L g1435 ( 
.A(n_1251),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1264),
.Y(n_1436)
);

CKINVDCx11_ASAP7_75t_R g1437 ( 
.A(n_1283),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1250),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1268),
.B(n_1269),
.Y(n_1439)
);

INVx4_ASAP7_75t_L g1440 ( 
.A(n_1272),
.Y(n_1440)
);

AOI22xp5_ASAP7_75t_SL g1441 ( 
.A1(n_1307),
.A2(n_1273),
.B1(n_1285),
.B2(n_1261),
.Y(n_1441)
);

NAND2x1p5_ASAP7_75t_L g1442 ( 
.A(n_1282),
.B(n_1285),
.Y(n_1442)
);

BUFx2_ASAP7_75t_SL g1443 ( 
.A(n_1262),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1269),
.A2(n_1268),
.B1(n_1262),
.B2(n_1289),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1267),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1309),
.A2(n_1332),
.B1(n_1347),
.B2(n_1312),
.Y(n_1446)
);

OAI21xp5_ASAP7_75t_SL g1447 ( 
.A1(n_1281),
.A2(n_1259),
.B(n_1332),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1309),
.A2(n_1354),
.B1(n_1347),
.B2(n_1333),
.Y(n_1448)
);

AOI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1334),
.A2(n_1260),
.B1(n_1276),
.B2(n_1286),
.Y(n_1449)
);

BUFx2_ASAP7_75t_SL g1450 ( 
.A(n_1280),
.Y(n_1450)
);

INVx6_ASAP7_75t_L g1451 ( 
.A(n_1280),
.Y(n_1451)
);

INVx3_ASAP7_75t_L g1452 ( 
.A(n_1353),
.Y(n_1452)
);

INVx6_ASAP7_75t_L g1453 ( 
.A(n_1270),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1312),
.B(n_1333),
.Y(n_1454)
);

INVx1_ASAP7_75t_SL g1455 ( 
.A(n_1270),
.Y(n_1455)
);

INVx6_ASAP7_75t_L g1456 ( 
.A(n_1254),
.Y(n_1456)
);

OAI21xp5_ASAP7_75t_SL g1457 ( 
.A1(n_1319),
.A2(n_1339),
.B(n_1354),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1277),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1284),
.B(n_1254),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1254),
.Y(n_1460)
);

BUFx10_ASAP7_75t_L g1461 ( 
.A(n_1260),
.Y(n_1461)
);

OAI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1263),
.A2(n_1348),
.B1(n_1216),
.B2(n_1337),
.Y(n_1462)
);

CKINVDCx20_ASAP7_75t_R g1463 ( 
.A(n_1226),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1258),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1258),
.Y(n_1465)
);

BUFx4f_ASAP7_75t_SL g1466 ( 
.A(n_1258),
.Y(n_1466)
);

CKINVDCx6p67_ASAP7_75t_R g1467 ( 
.A(n_1244),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_SL g1468 ( 
.A1(n_1319),
.A2(n_1339),
.B1(n_1323),
.B2(n_1344),
.Y(n_1468)
);

INVx6_ASAP7_75t_L g1469 ( 
.A(n_1255),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1266),
.A2(n_1220),
.B1(n_1226),
.B2(n_1236),
.Y(n_1470)
);

BUFx2_ASAP7_75t_SL g1471 ( 
.A(n_1287),
.Y(n_1471)
);

CKINVDCx11_ASAP7_75t_R g1472 ( 
.A(n_1368),
.Y(n_1472)
);

OAI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1228),
.A2(n_1359),
.B1(n_1287),
.B2(n_1343),
.Y(n_1473)
);

CKINVDCx11_ASAP7_75t_R g1474 ( 
.A(n_1317),
.Y(n_1474)
);

OAI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1343),
.A2(n_1359),
.B1(n_1224),
.B2(n_1301),
.Y(n_1475)
);

INVx6_ASAP7_75t_L g1476 ( 
.A(n_1215),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1314),
.A2(n_1315),
.B1(n_1321),
.B2(n_1331),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1342),
.A2(n_1346),
.B1(n_1357),
.B2(n_1358),
.Y(n_1478)
);

AOI22xp5_ASAP7_75t_SL g1479 ( 
.A1(n_1363),
.A2(n_774),
.B1(n_1235),
.B2(n_1227),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_SL g1480 ( 
.A1(n_1351),
.A2(n_1205),
.B1(n_774),
.B2(n_1140),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1351),
.B(n_1237),
.Y(n_1481)
);

INVxp67_ASAP7_75t_SL g1482 ( 
.A(n_1226),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1217),
.Y(n_1483)
);

CKINVDCx20_ASAP7_75t_R g1484 ( 
.A(n_1299),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1305),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1338),
.Y(n_1486)
);

INVx1_ASAP7_75t_SL g1487 ( 
.A(n_1322),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_1225),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1352),
.A2(n_1205),
.B1(n_776),
.B2(n_774),
.Y(n_1489)
);

OAI22xp5_ASAP7_75t_SL g1490 ( 
.A1(n_1242),
.A2(n_790),
.B1(n_776),
.B2(n_1352),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_SL g1491 ( 
.A1(n_1351),
.A2(n_1205),
.B1(n_774),
.B2(n_1140),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1217),
.Y(n_1492)
);

CKINVDCx11_ASAP7_75t_R g1493 ( 
.A(n_1299),
.Y(n_1493)
);

CKINVDCx20_ASAP7_75t_R g1494 ( 
.A(n_1299),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1351),
.A2(n_1205),
.B1(n_774),
.B2(n_1140),
.Y(n_1495)
);

INVx6_ASAP7_75t_L g1496 ( 
.A(n_1302),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1475),
.A2(n_1478),
.B(n_1477),
.Y(n_1497)
);

BUFx3_ASAP7_75t_L g1498 ( 
.A(n_1376),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1459),
.B(n_1381),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1417),
.A2(n_1495),
.B1(n_1491),
.B2(n_1480),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1373),
.Y(n_1501)
);

NOR2x1_ASAP7_75t_L g1502 ( 
.A(n_1447),
.B(n_1420),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1480),
.A2(n_1495),
.B1(n_1491),
.B2(n_1489),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1373),
.Y(n_1504)
);

INVxp67_ASAP7_75t_SL g1505 ( 
.A(n_1486),
.Y(n_1505)
);

BUFx2_ASAP7_75t_L g1506 ( 
.A(n_1467),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1481),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1485),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1481),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1439),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1439),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1381),
.B(n_1395),
.Y(n_1512)
);

CKINVDCx6p67_ASAP7_75t_R g1513 ( 
.A(n_1392),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1377),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1395),
.B(n_1460),
.Y(n_1515)
);

BUFx5_ASAP7_75t_L g1516 ( 
.A(n_1461),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1374),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1454),
.Y(n_1518)
);

BUFx12f_ASAP7_75t_L g1519 ( 
.A(n_1371),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1383),
.Y(n_1520)
);

OAI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1417),
.A2(n_1420),
.B(n_1409),
.Y(n_1521)
);

INVx4_ASAP7_75t_SL g1522 ( 
.A(n_1451),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1454),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1436),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1388),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1403),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1411),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1414),
.Y(n_1528)
);

NAND2x1_ASAP7_75t_L g1529 ( 
.A(n_1453),
.B(n_1469),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1419),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1487),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1424),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1460),
.B(n_1456),
.Y(n_1533)
);

CKINVDCx20_ASAP7_75t_R g1534 ( 
.A(n_1484),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1483),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1492),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1455),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_SL g1538 ( 
.A1(n_1409),
.A2(n_1400),
.B(n_1447),
.Y(n_1538)
);

INVx3_ASAP7_75t_L g1539 ( 
.A(n_1476),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1455),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1390),
.B(n_1399),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1425),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1429),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1389),
.Y(n_1544)
);

BUFx6f_ASAP7_75t_L g1545 ( 
.A(n_1393),
.Y(n_1545)
);

INVxp67_ASAP7_75t_L g1546 ( 
.A(n_1413),
.Y(n_1546)
);

NAND2x1p5_ASAP7_75t_L g1547 ( 
.A(n_1393),
.B(n_1441),
.Y(n_1547)
);

AOI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1490),
.A2(n_1426),
.B1(n_1379),
.B2(n_1380),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1458),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1475),
.A2(n_1446),
.B(n_1448),
.Y(n_1550)
);

OAI21x1_ASAP7_75t_L g1551 ( 
.A1(n_1446),
.A2(n_1448),
.B(n_1470),
.Y(n_1551)
);

OAI21x1_ASAP7_75t_L g1552 ( 
.A1(n_1457),
.A2(n_1438),
.B(n_1482),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1482),
.Y(n_1553)
);

A2O1A1Ixp33_ASAP7_75t_L g1554 ( 
.A1(n_1479),
.A2(n_1445),
.B(n_1387),
.C(n_1400),
.Y(n_1554)
);

BUFx2_ASAP7_75t_L g1555 ( 
.A(n_1463),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1393),
.Y(n_1556)
);

OAI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1457),
.A2(n_1449),
.B(n_1442),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1464),
.B(n_1465),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1406),
.B(n_1404),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1410),
.Y(n_1560)
);

OAI21x1_ASAP7_75t_L g1561 ( 
.A1(n_1442),
.A2(n_1444),
.B(n_1452),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1410),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1471),
.Y(n_1563)
);

BUFx6f_ASAP7_75t_L g1564 ( 
.A(n_1474),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1472),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1466),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1450),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1462),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1407),
.B(n_1378),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1441),
.B(n_1452),
.Y(n_1570)
);

OAI21x1_ASAP7_75t_L g1571 ( 
.A1(n_1468),
.A2(n_1473),
.B(n_1412),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1468),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1378),
.Y(n_1573)
);

BUFx2_ASAP7_75t_L g1574 ( 
.A(n_1435),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1428),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1428),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1479),
.Y(n_1577)
);

OAI21x1_ASAP7_75t_L g1578 ( 
.A1(n_1416),
.A2(n_1443),
.B(n_1430),
.Y(n_1578)
);

BUFx4f_ASAP7_75t_SL g1579 ( 
.A(n_1494),
.Y(n_1579)
);

INVx4_ASAP7_75t_SL g1580 ( 
.A(n_1397),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1440),
.Y(n_1581)
);

CKINVDCx6p67_ASAP7_75t_R g1582 ( 
.A(n_1493),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1440),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1391),
.B(n_1423),
.Y(n_1584)
);

INVx6_ASAP7_75t_L g1585 ( 
.A(n_1401),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1398),
.B(n_1408),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1508),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1499),
.B(n_1515),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1499),
.B(n_1415),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1555),
.B(n_1437),
.Y(n_1590)
);

AO32x2_ASAP7_75t_L g1591 ( 
.A1(n_1500),
.A2(n_1421),
.A3(n_1372),
.B1(n_1422),
.B2(n_1434),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1535),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1525),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1525),
.Y(n_1594)
);

INVx3_ASAP7_75t_L g1595 ( 
.A(n_1539),
.Y(n_1595)
);

NOR2x1p5_ASAP7_75t_L g1596 ( 
.A(n_1582),
.B(n_1396),
.Y(n_1596)
);

AOI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1521),
.A2(n_1427),
.B(n_1422),
.Y(n_1597)
);

AO32x2_ASAP7_75t_L g1598 ( 
.A1(n_1560),
.A2(n_1394),
.A3(n_1370),
.B1(n_1431),
.B2(n_1496),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1570),
.B(n_1488),
.Y(n_1599)
);

A2O1A1Ixp33_ASAP7_75t_L g1600 ( 
.A1(n_1548),
.A2(n_1375),
.B(n_1384),
.C(n_1402),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1544),
.B(n_1385),
.Y(n_1601)
);

O2A1O1Ixp33_ASAP7_75t_L g1602 ( 
.A1(n_1538),
.A2(n_1401),
.B(n_1433),
.C(n_1418),
.Y(n_1602)
);

OA21x2_ASAP7_75t_L g1603 ( 
.A1(n_1550),
.A2(n_1433),
.B(n_1405),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1502),
.B(n_1496),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1502),
.B(n_1402),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1510),
.B(n_1382),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1510),
.B(n_1382),
.Y(n_1607)
);

AOI221xp5_ASAP7_75t_L g1608 ( 
.A1(n_1569),
.A2(n_1375),
.B1(n_1386),
.B2(n_1432),
.C(n_1573),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1505),
.B(n_1514),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1531),
.B(n_1546),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1559),
.B(n_1511),
.Y(n_1611)
);

AO21x2_ASAP7_75t_L g1612 ( 
.A1(n_1577),
.A2(n_1538),
.B(n_1562),
.Y(n_1612)
);

AND2x4_ASAP7_75t_L g1613 ( 
.A(n_1570),
.B(n_1522),
.Y(n_1613)
);

OA21x2_ASAP7_75t_L g1614 ( 
.A1(n_1550),
.A2(n_1551),
.B(n_1552),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1503),
.A2(n_1512),
.B1(n_1554),
.B2(n_1580),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1533),
.B(n_1501),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1574),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1570),
.B(n_1522),
.Y(n_1618)
);

A2O1A1Ixp33_ASAP7_75t_L g1619 ( 
.A1(n_1575),
.A2(n_1576),
.B(n_1541),
.C(n_1570),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1501),
.B(n_1504),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1504),
.B(n_1507),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1526),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1498),
.B(n_1581),
.Y(n_1623)
);

OAI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1572),
.A2(n_1568),
.B(n_1571),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1575),
.A2(n_1576),
.B1(n_1585),
.B2(n_1564),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1533),
.B(n_1507),
.Y(n_1626)
);

OAI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1571),
.A2(n_1551),
.B(n_1537),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1509),
.B(n_1498),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1526),
.Y(n_1629)
);

A2O1A1Ixp33_ASAP7_75t_L g1630 ( 
.A1(n_1578),
.A2(n_1557),
.B(n_1566),
.C(n_1564),
.Y(n_1630)
);

OAI21x1_ASAP7_75t_L g1631 ( 
.A1(n_1552),
.A2(n_1497),
.B(n_1557),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1564),
.B(n_1565),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1583),
.B(n_1564),
.Y(n_1633)
);

OAI21x1_ASAP7_75t_L g1634 ( 
.A1(n_1497),
.A2(n_1561),
.B(n_1529),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1517),
.B(n_1520),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1518),
.B(n_1523),
.Y(n_1636)
);

A2O1A1Ixp33_ASAP7_75t_L g1637 ( 
.A1(n_1578),
.A2(n_1561),
.B(n_1506),
.C(n_1556),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1517),
.B(n_1520),
.Y(n_1638)
);

AOI211xp5_ASAP7_75t_L g1639 ( 
.A1(n_1506),
.A2(n_1563),
.B(n_1530),
.C(n_1536),
.Y(n_1639)
);

NOR2x1_ASAP7_75t_SL g1640 ( 
.A(n_1545),
.B(n_1556),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1542),
.B(n_1543),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1527),
.B(n_1528),
.Y(n_1642)
);

CKINVDCx14_ASAP7_75t_R g1643 ( 
.A(n_1582),
.Y(n_1643)
);

OAI21xp5_ASAP7_75t_L g1644 ( 
.A1(n_1537),
.A2(n_1540),
.B(n_1567),
.Y(n_1644)
);

OAI221xp5_ASAP7_75t_SL g1645 ( 
.A1(n_1615),
.A2(n_1523),
.B1(n_1540),
.B2(n_1536),
.C(n_1532),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1593),
.Y(n_1646)
);

BUFx2_ASAP7_75t_L g1647 ( 
.A(n_1644),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1587),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1594),
.Y(n_1649)
);

INVxp67_ASAP7_75t_L g1650 ( 
.A(n_1609),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_SL g1651 ( 
.A1(n_1624),
.A2(n_1547),
.B1(n_1516),
.B2(n_1580),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1611),
.B(n_1532),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_1643),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1616),
.B(n_1553),
.Y(n_1654)
);

INVx3_ASAP7_75t_L g1655 ( 
.A(n_1603),
.Y(n_1655)
);

NOR2x1p5_ASAP7_75t_L g1656 ( 
.A(n_1589),
.B(n_1519),
.Y(n_1656)
);

NOR2x1_ASAP7_75t_L g1657 ( 
.A(n_1620),
.B(n_1621),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1626),
.B(n_1553),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1628),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1622),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1629),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1626),
.B(n_1558),
.Y(n_1662)
);

INVx3_ASAP7_75t_L g1663 ( 
.A(n_1603),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1610),
.B(n_1558),
.Y(n_1664)
);

BUFx2_ASAP7_75t_L g1665 ( 
.A(n_1603),
.Y(n_1665)
);

INVxp67_ASAP7_75t_L g1666 ( 
.A(n_1601),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1636),
.B(n_1516),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1592),
.Y(n_1668)
);

INVx3_ASAP7_75t_L g1669 ( 
.A(n_1595),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1642),
.B(n_1549),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_SL g1671 ( 
.A1(n_1589),
.A2(n_1547),
.B1(n_1534),
.B2(n_1574),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1641),
.Y(n_1672)
);

INVx1_ASAP7_75t_SL g1673 ( 
.A(n_1617),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1612),
.B(n_1549),
.Y(n_1674)
);

AOI222xp33_ASAP7_75t_L g1675 ( 
.A1(n_1619),
.A2(n_1625),
.B1(n_1608),
.B2(n_1627),
.C1(n_1588),
.C2(n_1600),
.Y(n_1675)
);

INVxp67_ASAP7_75t_L g1676 ( 
.A(n_1606),
.Y(n_1676)
);

AOI21xp5_ASAP7_75t_SL g1677 ( 
.A1(n_1656),
.A2(n_1630),
.B(n_1637),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1646),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1654),
.B(n_1614),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_SL g1680 ( 
.A1(n_1653),
.A2(n_1643),
.B1(n_1519),
.B2(n_1585),
.Y(n_1680)
);

AOI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1675),
.A2(n_1619),
.B1(n_1600),
.B2(n_1605),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1664),
.B(n_1635),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1664),
.B(n_1638),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1646),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1657),
.Y(n_1685)
);

BUFx2_ASAP7_75t_L g1686 ( 
.A(n_1655),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1654),
.B(n_1614),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1658),
.B(n_1614),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1649),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1647),
.B(n_1630),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1647),
.B(n_1631),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1649),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1658),
.B(n_1631),
.Y(n_1693)
);

BUFx6f_ASAP7_75t_L g1694 ( 
.A(n_1663),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1662),
.B(n_1607),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1662),
.B(n_1623),
.Y(n_1696)
);

INVxp67_ASAP7_75t_SL g1697 ( 
.A(n_1657),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1651),
.A2(n_1599),
.B1(n_1597),
.B2(n_1516),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_SL g1699 ( 
.A1(n_1671),
.A2(n_1590),
.B1(n_1598),
.B2(n_1618),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1665),
.B(n_1595),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1665),
.B(n_1672),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1669),
.B(n_1613),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1670),
.B(n_1634),
.Y(n_1703)
);

OA21x2_ASAP7_75t_L g1704 ( 
.A1(n_1674),
.A2(n_1634),
.B(n_1637),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1673),
.B(n_1604),
.Y(n_1705)
);

AOI221xp5_ASAP7_75t_SL g1706 ( 
.A1(n_1650),
.A2(n_1639),
.B1(n_1604),
.B2(n_1605),
.C(n_1602),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1648),
.B(n_1524),
.Y(n_1707)
);

OAI221xp5_ASAP7_75t_L g1708 ( 
.A1(n_1645),
.A2(n_1598),
.B1(n_1591),
.B2(n_1585),
.C(n_1633),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1697),
.B(n_1660),
.Y(n_1709)
);

NOR2x1_ASAP7_75t_L g1710 ( 
.A(n_1677),
.B(n_1656),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1679),
.B(n_1659),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1678),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1702),
.B(n_1671),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1697),
.B(n_1685),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1679),
.B(n_1676),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1682),
.B(n_1668),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1678),
.Y(n_1717)
);

INVxp67_ASAP7_75t_SL g1718 ( 
.A(n_1685),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1684),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1682),
.B(n_1652),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1684),
.Y(n_1721)
);

NOR2x1_ASAP7_75t_L g1722 ( 
.A(n_1691),
.B(n_1596),
.Y(n_1722)
);

INVx5_ASAP7_75t_L g1723 ( 
.A(n_1694),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1701),
.B(n_1689),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1702),
.B(n_1640),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1701),
.B(n_1661),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1702),
.B(n_1666),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1692),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1692),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1686),
.Y(n_1730)
);

AND2x4_ASAP7_75t_L g1731 ( 
.A(n_1702),
.B(n_1613),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1687),
.B(n_1688),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1693),
.B(n_1667),
.Y(n_1733)
);

INVxp67_ASAP7_75t_L g1734 ( 
.A(n_1708),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1682),
.B(n_1683),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1699),
.B(n_1632),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1712),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1734),
.B(n_1706),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1734),
.B(n_1706),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1735),
.B(n_1703),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1712),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1717),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1735),
.B(n_1703),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1717),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1719),
.Y(n_1745)
);

INVx1_ASAP7_75t_SL g1746 ( 
.A(n_1710),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1720),
.B(n_1701),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1713),
.B(n_1699),
.Y(n_1748)
);

A2O1A1Ixp33_ASAP7_75t_L g1749 ( 
.A1(n_1710),
.A2(n_1681),
.B(n_1708),
.C(n_1690),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1720),
.B(n_1695),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1713),
.B(n_1731),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1719),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1730),
.Y(n_1753)
);

INVxp67_ASAP7_75t_L g1754 ( 
.A(n_1722),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1721),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1731),
.B(n_1696),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1716),
.B(n_1695),
.Y(n_1757)
);

BUFx2_ASAP7_75t_L g1758 ( 
.A(n_1722),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1731),
.B(n_1696),
.Y(n_1759)
);

OR2x2_ASAP7_75t_L g1760 ( 
.A(n_1716),
.B(n_1703),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1731),
.B(n_1696),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1730),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1731),
.B(n_1700),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1726),
.B(n_1691),
.Y(n_1764)
);

O2A1O1Ixp33_ASAP7_75t_L g1765 ( 
.A1(n_1718),
.A2(n_1690),
.B(n_1691),
.C(n_1705),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1718),
.B(n_1695),
.Y(n_1766)
);

O2A1O1Ixp33_ASAP7_75t_L g1767 ( 
.A1(n_1714),
.A2(n_1690),
.B(n_1705),
.C(n_1686),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1725),
.B(n_1700),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1726),
.B(n_1707),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1709),
.Y(n_1770)
);

HB1xp67_ASAP7_75t_L g1771 ( 
.A(n_1709),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1728),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1728),
.Y(n_1773)
);

INVx3_ASAP7_75t_L g1774 ( 
.A(n_1725),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1729),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1737),
.Y(n_1776)
);

BUFx2_ASAP7_75t_L g1777 ( 
.A(n_1758),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1737),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1738),
.B(n_1711),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1751),
.B(n_1727),
.Y(n_1780)
);

INVxp67_ASAP7_75t_SL g1781 ( 
.A(n_1739),
.Y(n_1781)
);

NAND2x1p5_ASAP7_75t_L g1782 ( 
.A(n_1758),
.B(n_1681),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1741),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1741),
.Y(n_1784)
);

NOR2xp33_ASAP7_75t_L g1785 ( 
.A(n_1746),
.B(n_1680),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1742),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1753),
.Y(n_1787)
);

NAND3xp33_ASAP7_75t_SL g1788 ( 
.A(n_1749),
.B(n_1714),
.C(n_1736),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1742),
.Y(n_1789)
);

AOI21x1_ASAP7_75t_L g1790 ( 
.A1(n_1748),
.A2(n_1730),
.B(n_1686),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_SL g1791 ( 
.A(n_1748),
.B(n_1680),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1753),
.Y(n_1792)
);

INVx2_ASAP7_75t_SL g1793 ( 
.A(n_1751),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1756),
.B(n_1727),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1756),
.B(n_1725),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_SL g1796 ( 
.A(n_1754),
.B(n_1725),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1770),
.B(n_1711),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1750),
.B(n_1724),
.Y(n_1798)
);

INVxp67_ASAP7_75t_L g1799 ( 
.A(n_1771),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1759),
.B(n_1733),
.Y(n_1800)
);

NAND2x1p5_ASAP7_75t_L g1801 ( 
.A(n_1774),
.B(n_1723),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1757),
.B(n_1724),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1744),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1759),
.B(n_1733),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1740),
.B(n_1729),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1765),
.B(n_1715),
.Y(n_1806)
);

INVx1_ASAP7_75t_SL g1807 ( 
.A(n_1762),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1761),
.B(n_1733),
.Y(n_1808)
);

NOR2x1_ASAP7_75t_L g1809 ( 
.A(n_1767),
.B(n_1584),
.Y(n_1809)
);

OAI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1766),
.A2(n_1736),
.B(n_1698),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1762),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1744),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1788),
.A2(n_1704),
.B1(n_1732),
.B2(n_1772),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1779),
.B(n_1747),
.Y(n_1814)
);

AOI21xp33_ASAP7_75t_L g1815 ( 
.A1(n_1782),
.A2(n_1752),
.B(n_1745),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1803),
.Y(n_1816)
);

BUFx3_ASAP7_75t_L g1817 ( 
.A(n_1777),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1781),
.B(n_1761),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1776),
.Y(n_1819)
);

INVx1_ASAP7_75t_SL g1820 ( 
.A(n_1791),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_L g1821 ( 
.A(n_1791),
.B(n_1653),
.Y(n_1821)
);

OAI21xp33_ASAP7_75t_L g1822 ( 
.A1(n_1806),
.A2(n_1743),
.B(n_1740),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1776),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1778),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1780),
.B(n_1763),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1782),
.Y(n_1826)
);

OAI322xp33_ASAP7_75t_L g1827 ( 
.A1(n_1782),
.A2(n_1764),
.A3(n_1760),
.B1(n_1743),
.B2(n_1769),
.C1(n_1775),
.C2(n_1755),
.Y(n_1827)
);

AOI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1809),
.A2(n_1704),
.B1(n_1732),
.B2(n_1599),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1778),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1780),
.B(n_1794),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1783),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1798),
.B(n_1769),
.Y(n_1832)
);

OAI31xp33_ASAP7_75t_SL g1833 ( 
.A1(n_1809),
.A2(n_1763),
.A3(n_1768),
.B(n_1732),
.Y(n_1833)
);

AND2x2_ASAP7_75t_SL g1834 ( 
.A(n_1777),
.B(n_1698),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1783),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1798),
.B(n_1760),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1802),
.B(n_1745),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1784),
.Y(n_1838)
);

OAI311xp33_ASAP7_75t_L g1839 ( 
.A1(n_1813),
.A2(n_1822),
.A3(n_1818),
.B1(n_1828),
.C1(n_1810),
.Y(n_1839)
);

INVx1_ASAP7_75t_SL g1840 ( 
.A(n_1820),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1817),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1830),
.B(n_1799),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1819),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1817),
.Y(n_1844)
);

INVxp67_ASAP7_75t_L g1845 ( 
.A(n_1821),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1823),
.Y(n_1846)
);

AOI221xp5_ASAP7_75t_L g1847 ( 
.A1(n_1813),
.A2(n_1810),
.B1(n_1807),
.B2(n_1787),
.C(n_1792),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1824),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1830),
.B(n_1793),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1825),
.B(n_1793),
.Y(n_1850)
);

NOR2xp33_ASAP7_75t_L g1851 ( 
.A(n_1821),
.B(n_1785),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1825),
.B(n_1794),
.Y(n_1852)
);

INVx1_ASAP7_75t_SL g1853 ( 
.A(n_1826),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1815),
.B(n_1800),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1826),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1833),
.B(n_1800),
.Y(n_1856)
);

A2O1A1Ixp33_ASAP7_75t_L g1857 ( 
.A1(n_1834),
.A2(n_1807),
.B(n_1811),
.C(n_1787),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1829),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1852),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1850),
.Y(n_1860)
);

NAND2xp33_ASAP7_75t_SL g1861 ( 
.A(n_1841),
.B(n_1816),
.Y(n_1861)
);

NAND3xp33_ASAP7_75t_L g1862 ( 
.A(n_1857),
.B(n_1834),
.C(n_1831),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1852),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1841),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1844),
.Y(n_1865)
);

OAI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1840),
.A2(n_1836),
.B1(n_1814),
.B2(n_1832),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1844),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1850),
.B(n_1832),
.Y(n_1868)
);

AOI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1839),
.A2(n_1827),
.B(n_1796),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_SL g1870 ( 
.A(n_1851),
.B(n_1579),
.Y(n_1870)
);

OAI221xp5_ASAP7_75t_L g1871 ( 
.A1(n_1847),
.A2(n_1790),
.B1(n_1836),
.B2(n_1787),
.C(n_1792),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1860),
.B(n_1849),
.Y(n_1872)
);

OAI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1869),
.A2(n_1856),
.B1(n_1845),
.B2(n_1854),
.Y(n_1873)
);

NAND3xp33_ASAP7_75t_L g1874 ( 
.A(n_1862),
.B(n_1842),
.C(n_1843),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1860),
.B(n_1853),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1868),
.B(n_1853),
.Y(n_1876)
);

NAND3xp33_ASAP7_75t_L g1877 ( 
.A(n_1861),
.B(n_1871),
.C(n_1865),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1859),
.Y(n_1878)
);

NAND2xp33_ASAP7_75t_SL g1879 ( 
.A(n_1866),
.B(n_1856),
.Y(n_1879)
);

OAI221xp5_ASAP7_75t_L g1880 ( 
.A1(n_1861),
.A2(n_1839),
.B1(n_1790),
.B2(n_1855),
.C(n_1811),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1863),
.B(n_1843),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1864),
.B(n_1846),
.Y(n_1882)
);

AND2x4_ASAP7_75t_L g1883 ( 
.A(n_1867),
.B(n_1846),
.Y(n_1883)
);

INVx1_ASAP7_75t_SL g1884 ( 
.A(n_1876),
.Y(n_1884)
);

AOI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1880),
.A2(n_1870),
.B1(n_1855),
.B2(n_1792),
.Y(n_1885)
);

AOI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1879),
.A2(n_1811),
.B1(n_1848),
.B2(n_1858),
.Y(n_1886)
);

O2A1O1Ixp33_ASAP7_75t_L g1887 ( 
.A1(n_1873),
.A2(n_1848),
.B(n_1858),
.C(n_1838),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1875),
.Y(n_1888)
);

NAND3xp33_ASAP7_75t_SL g1889 ( 
.A(n_1877),
.B(n_1801),
.C(n_1837),
.Y(n_1889)
);

HB1xp67_ASAP7_75t_L g1890 ( 
.A(n_1884),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1886),
.B(n_1883),
.Y(n_1891)
);

OAI22xp33_ASAP7_75t_SL g1892 ( 
.A1(n_1885),
.A2(n_1882),
.B1(n_1881),
.B2(n_1872),
.Y(n_1892)
);

AOI221xp5_ASAP7_75t_L g1893 ( 
.A1(n_1887),
.A2(n_1874),
.B1(n_1883),
.B2(n_1878),
.C(n_1835),
.Y(n_1893)
);

OAI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1888),
.A2(n_1837),
.B1(n_1797),
.B2(n_1801),
.Y(n_1894)
);

AOI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1889),
.A2(n_1812),
.B1(n_1784),
.B2(n_1786),
.Y(n_1895)
);

CKINVDCx16_ASAP7_75t_R g1896 ( 
.A(n_1884),
.Y(n_1896)
);

INVx1_ASAP7_75t_SL g1897 ( 
.A(n_1896),
.Y(n_1897)
);

AND2x4_ASAP7_75t_L g1898 ( 
.A(n_1890),
.B(n_1795),
.Y(n_1898)
);

INVx1_ASAP7_75t_SL g1899 ( 
.A(n_1891),
.Y(n_1899)
);

AOI22xp5_ASAP7_75t_L g1900 ( 
.A1(n_1892),
.A2(n_1812),
.B1(n_1786),
.B2(n_1789),
.Y(n_1900)
);

INVx1_ASAP7_75t_SL g1901 ( 
.A(n_1895),
.Y(n_1901)
);

INVx2_ASAP7_75t_SL g1902 ( 
.A(n_1894),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_SL g1903 ( 
.A(n_1897),
.B(n_1899),
.Y(n_1903)
);

NOR2x1p5_ASAP7_75t_L g1904 ( 
.A(n_1898),
.B(n_1893),
.Y(n_1904)
);

AOI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1901),
.A2(n_1789),
.B(n_1801),
.Y(n_1905)
);

BUFx6f_ASAP7_75t_L g1906 ( 
.A(n_1903),
.Y(n_1906)
);

AOI22x1_ASAP7_75t_L g1907 ( 
.A1(n_1906),
.A2(n_1904),
.B1(n_1902),
.B2(n_1905),
.Y(n_1907)
);

AOI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1907),
.A2(n_1906),
.B1(n_1900),
.B2(n_1774),
.Y(n_1908)
);

OAI22x1_ASAP7_75t_L g1909 ( 
.A1(n_1907),
.A2(n_1906),
.B1(n_1586),
.B2(n_1774),
.Y(n_1909)
);

XNOR2xp5_ASAP7_75t_L g1910 ( 
.A(n_1909),
.B(n_1908),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1908),
.Y(n_1911)
);

OAI21xp33_ASAP7_75t_L g1912 ( 
.A1(n_1910),
.A2(n_1906),
.B(n_1795),
.Y(n_1912)
);

AO22x2_ASAP7_75t_L g1913 ( 
.A1(n_1911),
.A2(n_1805),
.B1(n_1808),
.B2(n_1804),
.Y(n_1913)
);

AOI22xp33_ASAP7_75t_L g1914 ( 
.A1(n_1913),
.A2(n_1805),
.B1(n_1808),
.B2(n_1804),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1914),
.B(n_1912),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1915),
.Y(n_1916)
);

AOI221xp5_ASAP7_75t_L g1917 ( 
.A1(n_1916),
.A2(n_1752),
.B1(n_1775),
.B2(n_1773),
.C(n_1772),
.Y(n_1917)
);

AOI211xp5_ASAP7_75t_L g1918 ( 
.A1(n_1917),
.A2(n_1802),
.B(n_1513),
.C(n_1764),
.Y(n_1918)
);


endmodule