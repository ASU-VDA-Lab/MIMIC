module fake_jpeg_10460_n_41 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_41);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_41;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_21),
.Y(n_30)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_11),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_15),
.B(n_0),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_17),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_16),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_19),
.B1(n_18),
.B2(n_4),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_26),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_20),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_22),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_28),
.Y(n_33)
);

AO22x1_ASAP7_75t_SL g28 ( 
.A1(n_24),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_22),
.Y(n_31)
);

FAx1_ASAP7_75t_SL g36 ( 
.A(n_33),
.B(n_31),
.CI(n_32),
.CON(n_36),
.SN(n_36)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_SL g37 ( 
.A(n_35),
.B(n_32),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_38),
.A2(n_36),
.B(n_37),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_39),
.A2(n_38),
.B(n_34),
.Y(n_40)
);

AO21x1_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_28),
.B(n_30),
.Y(n_41)
);


endmodule