module fake_jpeg_30383_n_317 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_317);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_20),
.B(n_10),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_20),
.B(n_10),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_24),
.B(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_57),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_10),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_56),
.B(n_58),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_0),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_0),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_42),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_23),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_65),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_24),
.B(n_9),
.Y(n_64)
);

NAND3xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_22),
.C(n_25),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_37),
.B1(n_28),
.B2(n_40),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_80),
.A2(n_82),
.B1(n_98),
.B2(n_70),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_47),
.A2(n_29),
.B1(n_41),
.B2(n_34),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_91),
.B1(n_101),
.B2(n_111),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_60),
.A2(n_40),
.B1(n_39),
.B2(n_28),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_93),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_89),
.B(n_96),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_63),
.A2(n_41),
.B1(n_21),
.B2(n_30),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_39),
.Y(n_93)
);

INVx6_ASAP7_75t_SL g95 ( 
.A(n_67),
.Y(n_95)
);

INVx4_ASAP7_75t_SL g128 ( 
.A(n_95),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_69),
.A2(n_22),
.B1(n_25),
.B2(n_27),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_49),
.A2(n_25),
.B1(n_27),
.B2(n_41),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_48),
.B(n_27),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_102),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_68),
.A2(n_21),
.B1(n_33),
.B2(n_38),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_51),
.B(n_43),
.Y(n_102)
);

NOR3xp33_ASAP7_75t_L g106 ( 
.A(n_57),
.B(n_43),
.C(n_19),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_42),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_57),
.A2(n_43),
.B(n_19),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_109),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_71),
.A2(n_73),
.B1(n_46),
.B2(n_59),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_115),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_113),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_116),
.Y(n_183)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_120),
.Y(n_174)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_19),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_123),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_26),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_99),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_124),
.B(n_142),
.Y(n_176)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_26),
.C(n_38),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_66),
.C(n_100),
.Y(n_155)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_129),
.Y(n_166)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_134),
.Y(n_161)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_132),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_78),
.B(n_26),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_133),
.B(n_145),
.Y(n_180)
);

AOI32xp33_ASAP7_75t_L g134 ( 
.A1(n_84),
.A2(n_52),
.A3(n_33),
.B1(n_36),
.B2(n_30),
.Y(n_134)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_136),
.Y(n_175)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_138),
.Y(n_165)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_109),
.A2(n_42),
.B(n_65),
.C(n_61),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_139),
.A2(n_101),
.B1(n_91),
.B2(n_81),
.Y(n_156)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_143),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g178 ( 
.A1(n_141),
.A2(n_88),
.B(n_1),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_87),
.B(n_30),
.Y(n_142)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_77),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_79),
.B(n_33),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_150),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_85),
.B(n_38),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_147),
.B(n_148),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_104),
.B(n_36),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_86),
.B(n_36),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_149),
.B(n_151),
.Y(n_184)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

AO22x2_ASAP7_75t_SL g152 ( 
.A1(n_111),
.A2(n_72),
.B1(n_54),
.B2(n_65),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_152),
.A2(n_75),
.B1(n_108),
.B2(n_107),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_155),
.B(n_156),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_144),
.A2(n_114),
.B1(n_94),
.B2(n_105),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_159),
.A2(n_171),
.B1(n_177),
.B2(n_179),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_123),
.C(n_135),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_162),
.B(n_169),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_119),
.A2(n_135),
.B1(n_139),
.B2(n_152),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_168),
.A2(n_182),
.B1(n_142),
.B2(n_128),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_126),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_124),
.B(n_15),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_172),
.A2(n_12),
.B(n_4),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_118),
.B(n_15),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_18),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_151),
.A2(n_105),
.B1(n_94),
.B2(n_108),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_178),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_152),
.A2(n_107),
.B1(n_53),
.B2(n_88),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_125),
.B(n_62),
.C(n_2),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_181),
.B(n_17),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_149),
.A2(n_11),
.B1(n_2),
.B2(n_4),
.Y(n_182)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_186),
.A2(n_196),
.B1(n_213),
.B2(n_171),
.Y(n_218)
);

AND2x4_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_128),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_189),
.Y(n_214)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_156),
.B(n_184),
.Y(n_189)
);

AND2x2_ASAP7_75t_SL g190 ( 
.A(n_157),
.B(n_121),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_190),
.B(n_208),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_191),
.B(n_210),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_132),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_197),
.Y(n_226)
);

NAND3xp33_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_176),
.C(n_180),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_184),
.A2(n_146),
.B1(n_136),
.B2(n_129),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_157),
.B(n_127),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_162),
.B(n_120),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_205),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_201),
.Y(n_217)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_200),
.Y(n_237)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_206),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_155),
.B(n_140),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_204),
.A2(n_174),
.B(n_183),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_176),
.B(n_143),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_159),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_169),
.B(n_153),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_212),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_115),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_116),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_211),
.B(n_14),
.Y(n_233)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_177),
.A2(n_131),
.B1(n_4),
.B2(n_5),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_215),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_218),
.A2(n_221),
.B1(n_223),
.B2(n_227),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_172),
.C(n_167),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_224),
.C(n_190),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_186),
.A2(n_179),
.B1(n_166),
.B2(n_154),
.Y(n_221)
);

AOI322xp5_ASAP7_75t_L g222 ( 
.A1(n_189),
.A2(n_194),
.A3(n_205),
.B1(n_198),
.B2(n_187),
.C1(n_202),
.C2(n_207),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_222),
.B(n_233),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_202),
.A2(n_166),
.B1(n_154),
.B2(n_175),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_164),
.C(n_158),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_209),
.A2(n_182),
.B1(n_131),
.B2(n_175),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_209),
.A2(n_158),
.B1(n_174),
.B2(n_183),
.Y(n_230)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_232),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_187),
.A2(n_160),
.B(n_0),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_235),
.A2(n_188),
.B(n_185),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_196),
.A2(n_160),
.B1(n_8),
.B2(n_9),
.Y(n_236)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_204),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_241),
.C(n_243),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_225),
.B(n_191),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_240),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_204),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_197),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_226),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_192),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_248),
.C(n_255),
.Y(n_269)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_229),
.Y(n_249)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_200),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_250),
.A2(n_226),
.B(n_234),
.Y(n_270)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_217),
.Y(n_252)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_234),
.B(n_211),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_219),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_190),
.C(n_187),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_217),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_256),
.B(n_228),
.Y(n_258)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_258),
.Y(n_273)
);

AOI322xp5_ASAP7_75t_L g259 ( 
.A1(n_253),
.A2(n_228),
.A3(n_227),
.B1(n_235),
.B2(n_230),
.C1(n_187),
.C2(n_237),
.Y(n_259)
);

AOI322xp5_ASAP7_75t_L g274 ( 
.A1(n_259),
.A2(n_247),
.A3(n_249),
.B1(n_252),
.B2(n_256),
.C1(n_244),
.C2(n_239),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_263),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_245),
.A2(n_218),
.B1(n_220),
.B2(n_216),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_261),
.A2(n_262),
.B1(n_250),
.B2(n_239),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_242),
.A2(n_237),
.B1(n_216),
.B2(n_220),
.Y(n_262)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_270),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_242),
.A2(n_221),
.B1(n_223),
.B2(n_193),
.Y(n_271)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_271),
.Y(n_283)
);

OAI322xp33_ASAP7_75t_L g272 ( 
.A1(n_254),
.A2(n_225),
.A3(n_233),
.B1(n_190),
.B2(n_232),
.C1(n_195),
.C2(n_212),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_243),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_276),
.C(n_282),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_248),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_268),
.B(n_257),
.Y(n_277)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_277),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_278),
.B(n_279),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_264),
.B(n_241),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_246),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_284),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_267),
.C(n_263),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_261),
.A2(n_251),
.B1(n_255),
.B2(n_213),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_285),
.B(n_260),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_294),
.C(n_295),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_269),
.C(n_238),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_289),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_266),
.C(n_265),
.Y(n_289)
);

NOR3xp33_ASAP7_75t_SL g290 ( 
.A(n_273),
.B(n_272),
.C(n_258),
.Y(n_290)
);

OA21x2_ASAP7_75t_SL g296 ( 
.A1(n_290),
.A2(n_273),
.B(n_270),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_285),
.C(n_281),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_266),
.C(n_265),
.Y(n_295)
);

OAI21x1_ASAP7_75t_L g304 ( 
.A1(n_296),
.A2(n_302),
.B(n_293),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_286),
.A2(n_275),
.B(n_283),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_297),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_292),
.A2(n_275),
.B(n_283),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_301),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_291),
.A2(n_278),
.B(n_271),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_292),
.A2(n_262),
.B(n_203),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_298),
.A2(n_293),
.B1(n_201),
.B2(n_12),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_303),
.A2(n_304),
.B1(n_14),
.B2(n_15),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_7),
.C(n_11),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_306),
.A2(n_18),
.B(n_16),
.Y(n_312)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_299),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_307),
.B(n_7),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_310),
.Y(n_314)
);

BUFx24_ASAP7_75t_SL g310 ( 
.A(n_305),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_311),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_308),
.C(n_303),
.Y(n_315)
);

OAI22xp33_ASAP7_75t_R g316 ( 
.A1(n_315),
.A2(n_306),
.B1(n_314),
.B2(n_312),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_16),
.Y(n_317)
);


endmodule