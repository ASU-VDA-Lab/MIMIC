module fake_jpeg_26690_n_225 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_225);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_3),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_21),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_18),
.B1(n_26),
.B2(n_25),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_45),
.A2(n_47),
.B1(n_48),
.B2(n_55),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_18),
.B1(n_26),
.B2(n_16),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_44),
.A2(n_18),
.B1(n_26),
.B2(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_36),
.B(n_23),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_54),
.B(n_57),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_23),
.B1(n_21),
.B2(n_24),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_33),
.B1(n_19),
.B2(n_22),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_56),
.A2(n_48),
.B1(n_46),
.B2(n_50),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_27),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

OR2x2_ASAP7_75t_SL g68 ( 
.A(n_58),
.B(n_64),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_35),
.A2(n_33),
.B1(n_22),
.B2(n_28),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_63),
.B1(n_27),
.B2(n_32),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_27),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_62),
.A2(n_24),
.B(n_28),
.C(n_17),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_35),
.A2(n_28),
.B1(n_17),
.B2(n_33),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_60),
.A2(n_29),
.B1(n_32),
.B2(n_20),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_66),
.A2(n_83),
.B(n_63),
.Y(n_97)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_69),
.Y(n_91)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_71),
.Y(n_100)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_77),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_75),
.Y(n_103)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_80),
.B1(n_88),
.B2(n_51),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_30),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_81),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_32),
.B1(n_20),
.B2(n_29),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_63),
.A2(n_29),
.B1(n_20),
.B2(n_24),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_31),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_87),
.B(n_22),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_51),
.A2(n_33),
.B1(n_22),
.B2(n_30),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_89),
.A2(n_97),
.B(n_106),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_67),
.B(n_59),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_92),
.B(n_94),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_81),
.A2(n_53),
.B1(n_51),
.B2(n_58),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_93),
.A2(n_108),
.B1(n_49),
.B2(n_1),
.Y(n_127)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_68),
.B1(n_69),
.B2(n_84),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_59),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_101),
.Y(n_120)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_83),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_102),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_65),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_105),
.B(n_110),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_73),
.A2(n_31),
.B(n_30),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_53),
.B1(n_52),
.B2(n_65),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_65),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_111),
.A2(n_84),
.B(n_1),
.Y(n_121)
);

OAI32xp33_ASAP7_75t_L g112 ( 
.A1(n_71),
.A2(n_53),
.A3(n_31),
.B1(n_2),
.B2(n_3),
.Y(n_112)
);

A2O1A1O1Ixp25_ASAP7_75t_L g116 ( 
.A1(n_112),
.A2(n_68),
.B(n_66),
.C(n_76),
.D(n_3),
.Y(n_116)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_110),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_113),
.B(n_117),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_82),
.C(n_72),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_109),
.C(n_91),
.Y(n_145)
);

OAI32xp33_ASAP7_75t_L g146 ( 
.A1(n_116),
.A2(n_109),
.A3(n_112),
.B1(n_105),
.B2(n_91),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_128),
.B1(n_111),
.B2(n_94),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_125),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_9),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_126),
.Y(n_139)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_9),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_127),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_89),
.A2(n_49),
.B1(n_1),
.B2(n_0),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_103),
.B(n_8),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_10),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_102),
.A2(n_8),
.B1(n_14),
.B2(n_2),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_90),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_100),
.B(n_8),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_133),
.B(n_104),
.Y(n_143)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_96),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_120),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_135),
.Y(n_166)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_136),
.B(n_142),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_138),
.A2(n_7),
.B1(n_4),
.B2(n_5),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_89),
.B1(n_95),
.B2(n_104),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_140),
.A2(n_134),
.B1(n_117),
.B2(n_125),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_106),
.B(n_97),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_141),
.A2(n_123),
.B(n_1),
.Y(n_163)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_147),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_148),
.Y(n_160)
);

AOI322xp5_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_116),
.A3(n_121),
.B1(n_131),
.B2(n_126),
.C1(n_129),
.C2(n_130),
.Y(n_157)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_101),
.C(n_90),
.Y(n_148)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_96),
.C(n_99),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_152),
.B(n_154),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_99),
.Y(n_155)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_157),
.B(n_139),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_169),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_137),
.A2(n_114),
.B(n_122),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_161),
.A2(n_163),
.B(n_137),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_140),
.A2(n_114),
.B1(n_122),
.B2(n_99),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_162),
.A2(n_170),
.B1(n_136),
.B2(n_153),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_165),
.Y(n_173)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_151),
.A2(n_11),
.B1(n_4),
.B2(n_5),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_171),
.A2(n_143),
.B1(n_144),
.B2(n_151),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_156),
.C(n_164),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_145),
.C(n_148),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_179),
.C(n_156),
.Y(n_188)
);

XNOR2x2_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_141),
.Y(n_176)
);

XNOR2x1_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_163),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_177),
.A2(n_169),
.B(n_135),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_166),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_180),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_147),
.C(n_142),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_183),
.Y(n_192)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_159),
.A2(n_138),
.B(n_144),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_184),
.A2(n_168),
.B(n_172),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_185),
.A2(n_184),
.B1(n_168),
.B2(n_170),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_180),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_187),
.B(n_196),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_189),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_191),
.A2(n_193),
.B(n_194),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_146),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_195),
.A2(n_193),
.B(n_186),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_139),
.C(n_167),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_179),
.C(n_174),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_190),
.A2(n_182),
.B1(n_181),
.B2(n_177),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_198),
.A2(n_6),
.B1(n_12),
.B2(n_13),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_182),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_201),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_183),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_204),
.B(n_173),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_205),
.B(n_188),
.C(n_173),
.Y(n_208)
);

NOR2xp67_ASAP7_75t_SL g206 ( 
.A(n_202),
.B(n_197),
.Y(n_206)
);

NOR2xp67_ASAP7_75t_SL g215 ( 
.A(n_206),
.B(n_203),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_209),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_208),
.B(n_203),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_200),
.A2(n_154),
.B(n_4),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_212),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_6),
.C(n_14),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_213),
.A2(n_215),
.B(n_216),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_210),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_214),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_212),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_219),
.B(n_207),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_220),
.B(n_205),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_221),
.A2(n_222),
.B1(n_218),
.B2(n_15),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_15),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_0),
.Y(n_225)
);


endmodule