module fake_netlist_1_12195_n_873 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_237, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_242, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_873);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_237;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_242;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_873;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_462;
wire n_316;
wire n_545;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_476;
wire n_617;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_724;
wire n_857;
wire n_786;
wire n_345;
wire n_360;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_567;
wire n_809;
wire n_580;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_533;
wire n_506;
wire n_393;
wire n_490;
wire n_247;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_666;
wire n_621;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_573;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_837;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_126), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_131), .Y(n_245) );
BUFx2_ASAP7_75t_L g246 ( .A(n_192), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_236), .Y(n_247) );
BUFx10_ASAP7_75t_L g248 ( .A(n_99), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_75), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_124), .Y(n_250) );
INVxp67_ASAP7_75t_L g251 ( .A(n_199), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g252 ( .A(n_242), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_39), .Y(n_253) );
CKINVDCx20_ASAP7_75t_R g254 ( .A(n_88), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_163), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_170), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_68), .Y(n_257) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_182), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_237), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_210), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_13), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_40), .Y(n_262) );
INVxp67_ASAP7_75t_L g263 ( .A(n_147), .Y(n_263) );
BUFx10_ASAP7_75t_L g264 ( .A(n_191), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_203), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g266 ( .A(n_230), .Y(n_266) );
INVx3_ASAP7_75t_L g267 ( .A(n_204), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_202), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_130), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_33), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_3), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_188), .Y(n_272) );
INVxp33_ASAP7_75t_SL g273 ( .A(n_102), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_34), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_181), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_93), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_10), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_171), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_103), .Y(n_279) );
CKINVDCx20_ASAP7_75t_R g280 ( .A(n_226), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_114), .Y(n_281) );
BUFx8_ASAP7_75t_SL g282 ( .A(n_137), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_145), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_29), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_57), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_217), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_216), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_166), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_59), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_24), .Y(n_290) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_81), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_43), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_127), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_89), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_118), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_87), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_26), .Y(n_297) );
CKINVDCx20_ASAP7_75t_R g298 ( .A(n_231), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_44), .Y(n_299) );
INVx1_ASAP7_75t_SL g300 ( .A(n_21), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_121), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_142), .Y(n_302) );
INVxp67_ASAP7_75t_L g303 ( .A(n_151), .Y(n_303) );
BUFx10_ASAP7_75t_L g304 ( .A(n_47), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_45), .Y(n_305) );
CKINVDCx14_ASAP7_75t_R g306 ( .A(n_28), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_157), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_101), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_113), .Y(n_309) );
BUFx10_ASAP7_75t_L g310 ( .A(n_243), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_227), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_164), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_235), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_5), .Y(n_314) );
INVx2_ASAP7_75t_SL g315 ( .A(n_122), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_129), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_154), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_32), .Y(n_318) );
CKINVDCx20_ASAP7_75t_R g319 ( .A(n_209), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_167), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_38), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_66), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_1), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_15), .Y(n_324) );
INVx1_ASAP7_75t_SL g325 ( .A(n_115), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_92), .Y(n_326) );
INVxp67_ASAP7_75t_L g327 ( .A(n_187), .Y(n_327) );
INVxp33_ASAP7_75t_SL g328 ( .A(n_42), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_72), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_225), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_76), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_197), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_19), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_22), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_90), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_98), .Y(n_336) );
CKINVDCx16_ASAP7_75t_R g337 ( .A(n_159), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_132), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_67), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_6), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_117), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_51), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_105), .Y(n_343) );
CKINVDCx20_ASAP7_75t_R g344 ( .A(n_222), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_85), .Y(n_345) );
INVx1_ASAP7_75t_SL g346 ( .A(n_84), .Y(n_346) );
CKINVDCx20_ASAP7_75t_R g347 ( .A(n_54), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_10), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_165), .Y(n_349) );
INVx1_ASAP7_75t_SL g350 ( .A(n_111), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_229), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_37), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_207), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_139), .Y(n_354) );
BUFx3_ASAP7_75t_L g355 ( .A(n_48), .Y(n_355) );
INVx2_ASAP7_75t_SL g356 ( .A(n_240), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_49), .Y(n_357) );
INVx1_ASAP7_75t_SL g358 ( .A(n_31), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_100), .Y(n_359) );
CKINVDCx16_ASAP7_75t_R g360 ( .A(n_97), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_106), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_110), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_9), .Y(n_363) );
INVx1_ASAP7_75t_SL g364 ( .A(n_172), .Y(n_364) );
BUFx3_ASAP7_75t_L g365 ( .A(n_233), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_41), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_21), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_11), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_140), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_345), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_345), .B(n_0), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_252), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_261), .Y(n_373) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_262), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_246), .B(n_2), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_337), .B(n_3), .Y(n_376) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_262), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_290), .Y(n_378) );
NAND2xp5_ASAP7_75t_SL g379 ( .A(n_267), .B(n_4), .Y(n_379) );
CKINVDCx8_ASAP7_75t_R g380 ( .A(n_360), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_315), .B(n_4), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_271), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_267), .Y(n_383) );
INVx6_ASAP7_75t_L g384 ( .A(n_248), .Y(n_384) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_262), .Y(n_385) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_262), .Y(n_386) );
CKINVDCx20_ASAP7_75t_R g387 ( .A(n_282), .Y(n_387) );
AND2x4_ASAP7_75t_L g388 ( .A(n_277), .B(n_5), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_282), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_314), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_333), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_306), .B(n_6), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_334), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_393) );
INVx2_ASAP7_75t_SL g394 ( .A(n_248), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_340), .B(n_7), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_306), .B(n_8), .Y(n_396) );
OAI21x1_ASAP7_75t_L g397 ( .A1(n_285), .A2(n_27), .B(n_25), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_348), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_398) );
CKINVDCx6p67_ASAP7_75t_R g399 ( .A(n_387), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_374), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_383), .Y(n_401) );
INVx3_ASAP7_75t_L g402 ( .A(n_388), .Y(n_402) );
OAI22xp33_ASAP7_75t_L g403 ( .A1(n_372), .A2(n_300), .B1(n_324), .B2(n_323), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_389), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_370), .A2(n_367), .B1(n_368), .B2(n_363), .Y(n_405) );
NOR2x1p5_ASAP7_75t_L g406 ( .A(n_378), .B(n_355), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_374), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_374), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_388), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_382), .Y(n_410) );
NOR2x1p5_ASAP7_75t_L g411 ( .A(n_390), .B(n_365), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_395), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_374), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_391), .Y(n_414) );
INVx3_ASAP7_75t_L g415 ( .A(n_395), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_384), .B(n_356), .Y(n_416) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_381), .B(n_286), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_381), .B(n_287), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_379), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_394), .B(n_301), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_397), .B(n_305), .Y(n_421) );
NAND3xp33_ASAP7_75t_L g422 ( .A(n_371), .B(n_375), .C(n_373), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_377), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_379), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_385), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_385), .Y(n_426) );
INVxp67_ASAP7_75t_L g427 ( .A(n_373), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_419), .B(n_392), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_401), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g430 ( .A1(n_421), .A2(n_396), .B(n_250), .Y(n_430) );
NOR2x1p5_ASAP7_75t_L g431 ( .A(n_399), .B(n_380), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_427), .B(n_376), .Y(n_432) );
INVx8_ASAP7_75t_L g433 ( .A(n_402), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_427), .B(n_371), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_410), .B(n_384), .Y(n_435) );
NOR2xp67_ASAP7_75t_L g436 ( .A(n_404), .B(n_375), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_422), .B(n_384), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_414), .B(n_251), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_405), .A2(n_372), .B1(n_258), .B2(n_266), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_409), .B(n_273), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_424), .B(n_328), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g442 ( .A(n_412), .B(n_244), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_411), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_403), .B(n_398), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_403), .A2(n_254), .B1(n_291), .B2(n_280), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_420), .Y(n_446) );
AND2x4_ASAP7_75t_L g447 ( .A(n_406), .B(n_393), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_415), .A2(n_247), .B1(n_259), .B2(n_256), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_416), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_417), .B(n_251), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_417), .A2(n_418), .B1(n_298), .B2(n_332), .Y(n_451) );
NOR2x1p5_ASAP7_75t_L g452 ( .A(n_418), .B(n_319), .Y(n_452) );
INVx2_ASAP7_75t_SL g453 ( .A(n_426), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_425), .B(n_263), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_400), .B(n_264), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_400), .B(n_303), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_407), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_407), .B(n_327), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_408), .B(n_269), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_408), .B(n_245), .Y(n_460) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_444), .A2(n_272), .B(n_279), .C(n_276), .Y(n_461) );
AOI21xp33_ASAP7_75t_L g462 ( .A1(n_434), .A2(n_347), .B(n_344), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_449), .B(n_249), .Y(n_463) );
AOI21x1_ASAP7_75t_L g464 ( .A1(n_430), .A2(n_423), .B(n_413), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_441), .A2(n_284), .B(n_281), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_441), .A2(n_299), .B(n_293), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_428), .A2(n_308), .B(n_302), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_451), .A2(n_312), .B1(n_316), .B2(n_309), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_432), .B(n_264), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_431), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_428), .A2(n_318), .B(n_317), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_450), .A2(n_321), .B(n_320), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_429), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_437), .A2(n_335), .B(n_339), .C(n_331), .Y(n_474) );
CKINVDCx10_ASAP7_75t_R g475 ( .A(n_452), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_442), .A2(n_343), .B(n_341), .Y(n_476) );
INVx6_ASAP7_75t_L g477 ( .A(n_433), .Y(n_477) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_440), .A2(n_351), .B(n_359), .C(n_361), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_439), .A2(n_362), .B1(n_369), .B2(n_253), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g480 ( .A1(n_438), .A2(n_346), .B(n_350), .C(n_358), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_435), .A2(n_330), .B(n_311), .Y(n_481) );
OAI21xp33_ASAP7_75t_L g482 ( .A1(n_448), .A2(n_257), .B(n_255), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_446), .B(n_304), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_458), .A2(n_364), .B(n_325), .Y(n_484) );
CKINVDCx8_ASAP7_75t_R g485 ( .A(n_447), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_458), .A2(n_265), .B(n_260), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_459), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_447), .A2(n_307), .B1(n_268), .B2(n_270), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_443), .B(n_304), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_445), .A2(n_313), .B1(n_274), .B2(n_275), .Y(n_490) );
INVx4_ASAP7_75t_L g491 ( .A(n_433), .Y(n_491) );
OAI21xp33_ASAP7_75t_L g492 ( .A1(n_456), .A2(n_283), .B(n_278), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_460), .A2(n_454), .B(n_457), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_436), .B(n_288), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_455), .A2(n_336), .B1(n_292), .B2(n_294), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_493), .A2(n_453), .B(n_295), .Y(n_496) );
NAND3xp33_ASAP7_75t_L g497 ( .A(n_480), .B(n_366), .C(n_296), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_469), .B(n_289), .Y(n_498) );
AO31x2_ASAP7_75t_L g499 ( .A1(n_474), .A2(n_377), .A3(n_385), .B(n_386), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_473), .Y(n_500) );
AND2x2_ASAP7_75t_SL g501 ( .A(n_491), .B(n_366), .Y(n_501) );
OAI21x1_ASAP7_75t_L g502 ( .A1(n_464), .A2(n_366), .B(n_30), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_465), .B(n_297), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_487), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_466), .B(n_322), .Y(n_505) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_467), .A2(n_329), .B(n_326), .Y(n_506) );
AO32x2_ASAP7_75t_L g507 ( .A1(n_468), .A2(n_377), .A3(n_386), .B1(n_310), .B2(n_16), .Y(n_507) );
AOI221xp5_ASAP7_75t_L g508 ( .A1(n_479), .A2(n_352), .B1(n_357), .B2(n_354), .C(n_353), .Y(n_508) );
INVxp67_ASAP7_75t_SL g509 ( .A(n_491), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_478), .B(n_338), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_462), .B(n_310), .Y(n_511) );
NAND2x1p5_ASAP7_75t_L g512 ( .A(n_477), .B(n_12), .Y(n_512) );
BUFx2_ASAP7_75t_L g513 ( .A(n_477), .Y(n_513) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_463), .Y(n_514) );
OAI21x1_ASAP7_75t_SL g515 ( .A1(n_484), .A2(n_14), .B(n_15), .Y(n_515) );
AO32x2_ASAP7_75t_L g516 ( .A1(n_490), .A2(n_386), .A3(n_16), .B1(n_17), .B2(n_18), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_461), .B(n_342), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_471), .A2(n_349), .B(n_149), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_486), .A2(n_148), .B(n_241), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_488), .B(n_14), .Y(n_520) );
NAND2x1p5_ASAP7_75t_L g521 ( .A(n_483), .B(n_17), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_472), .B(n_18), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_494), .A2(n_150), .B(n_239), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g524 ( .A1(n_476), .A2(n_146), .B(n_238), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_485), .B(n_19), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_489), .B(n_20), .Y(n_526) );
OAI21x1_ASAP7_75t_SL g527 ( .A1(n_481), .A2(n_20), .B(n_22), .Y(n_527) );
OAI21xp5_ASAP7_75t_L g528 ( .A1(n_492), .A2(n_153), .B(n_234), .Y(n_528) );
AO31x2_ASAP7_75t_L g529 ( .A1(n_495), .A2(n_23), .A3(n_24), .B(n_35), .Y(n_529) );
OAI21x1_ASAP7_75t_L g530 ( .A1(n_482), .A2(n_155), .B(n_36), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_470), .B(n_23), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_475), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_475), .A2(n_46), .B(n_50), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_485), .B(n_52), .Y(n_534) );
INVxp67_ASAP7_75t_SL g535 ( .A(n_501), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_504), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_504), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_500), .Y(n_538) );
OAI21x1_ASAP7_75t_L g539 ( .A1(n_502), .A2(n_53), .B(n_55), .Y(n_539) );
OAI21xp5_ASAP7_75t_L g540 ( .A1(n_519), .A2(n_56), .B(n_58), .Y(n_540) );
AO21x2_ASAP7_75t_L g541 ( .A1(n_528), .A2(n_60), .B(n_61), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_509), .B(n_62), .Y(n_542) );
OA21x2_ASAP7_75t_L g543 ( .A1(n_530), .A2(n_63), .B(n_64), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_512), .Y(n_544) );
NOR2x1_ASAP7_75t_SL g545 ( .A(n_514), .B(n_65), .Y(n_545) );
CKINVDCx11_ASAP7_75t_R g546 ( .A(n_532), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_511), .B(n_69), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_514), .Y(n_548) );
BUFx10_ASAP7_75t_L g549 ( .A(n_534), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_515), .Y(n_550) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_513), .Y(n_551) );
OAI21x1_ASAP7_75t_L g552 ( .A1(n_496), .A2(n_70), .B(n_71), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_514), .A2(n_73), .B1(n_74), .B2(n_77), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_520), .A2(n_78), .B1(n_79), .B2(n_80), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_525), .B(n_82), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_499), .Y(n_556) );
A2O1A1Ixp33_ASAP7_75t_L g557 ( .A1(n_522), .A2(n_83), .B(n_86), .C(n_91), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_499), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_527), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_498), .B(n_94), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_521), .B(n_95), .Y(n_561) );
OR2x6_ASAP7_75t_L g562 ( .A(n_533), .B(n_96), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_526), .B(n_104), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_517), .B(n_107), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_510), .A2(n_108), .B1(n_109), .B2(n_112), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_531), .B(n_116), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_503), .B(n_119), .Y(n_567) );
O2A1O1Ixp33_ASAP7_75t_SL g568 ( .A1(n_524), .A2(n_120), .B(n_123), .C(n_125), .Y(n_568) );
INVx1_ASAP7_75t_SL g569 ( .A(n_505), .Y(n_569) );
AO31x2_ASAP7_75t_L g570 ( .A1(n_523), .A2(n_128), .A3(n_133), .B(n_134), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_506), .B(n_135), .Y(n_571) );
OAI21xp5_ASAP7_75t_L g572 ( .A1(n_518), .A2(n_136), .B(n_138), .Y(n_572) );
AO21x2_ASAP7_75t_L g573 ( .A1(n_497), .A2(n_141), .B(n_143), .Y(n_573) );
OR2x6_ASAP7_75t_L g574 ( .A(n_507), .B(n_144), .Y(n_574) );
OA21x2_ASAP7_75t_L g575 ( .A1(n_499), .A2(n_152), .B(n_156), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_508), .B(n_232), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_529), .B(n_158), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_507), .A2(n_160), .B1(n_161), .B2(n_162), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_507), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_516), .B(n_168), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_516), .A2(n_169), .B1(n_173), .B2(n_174), .Y(n_581) );
OAI21xp5_ASAP7_75t_L g582 ( .A1(n_516), .A2(n_175), .B(n_176), .Y(n_582) );
OAI21x1_ASAP7_75t_L g583 ( .A1(n_529), .A2(n_177), .B(n_178), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_500), .Y(n_584) );
OAI21x1_ASAP7_75t_L g585 ( .A1(n_502), .A2(n_179), .B(n_180), .Y(n_585) );
OAI21x1_ASAP7_75t_L g586 ( .A1(n_502), .A2(n_183), .B(n_184), .Y(n_586) );
O2A1O1Ixp33_ASAP7_75t_SL g587 ( .A1(n_504), .A2(n_185), .B(n_186), .C(n_189), .Y(n_587) );
AO21x2_ASAP7_75t_L g588 ( .A1(n_502), .A2(n_190), .B(n_193), .Y(n_588) );
O2A1O1Ixp33_ASAP7_75t_SL g589 ( .A1(n_504), .A2(n_194), .B(n_195), .C(n_196), .Y(n_589) );
BUFx2_ASAP7_75t_L g590 ( .A(n_509), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_500), .Y(n_591) );
OAI21x1_ASAP7_75t_L g592 ( .A1(n_502), .A2(n_198), .B(n_200), .Y(n_592) );
AO32x2_ASAP7_75t_L g593 ( .A1(n_507), .A2(n_201), .A3(n_205), .B1(n_206), .B2(n_208), .Y(n_593) );
INVx2_ASAP7_75t_SL g594 ( .A(n_590), .Y(n_594) );
INVx2_ASAP7_75t_SL g595 ( .A(n_551), .Y(n_595) );
INVx2_ASAP7_75t_SL g596 ( .A(n_544), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_536), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_584), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_591), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_575), .Y(n_600) );
OA21x2_ASAP7_75t_L g601 ( .A1(n_583), .A2(n_211), .B(n_212), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_588), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_548), .Y(n_603) );
INVxp67_ASAP7_75t_L g604 ( .A(n_535), .Y(n_604) );
INVx3_ASAP7_75t_L g605 ( .A(n_562), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_588), .Y(n_606) );
AO21x2_ASAP7_75t_L g607 ( .A1(n_582), .A2(n_213), .B(n_214), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_569), .B(n_215), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_539), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_561), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_550), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_559), .Y(n_612) );
OAI21x1_ASAP7_75t_L g613 ( .A1(n_585), .A2(n_218), .B(n_219), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_549), .B(n_220), .Y(n_614) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_574), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_549), .B(n_221), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_586), .Y(n_617) );
BUFx3_ASAP7_75t_L g618 ( .A(n_546), .Y(n_618) );
INVx2_ASAP7_75t_SL g619 ( .A(n_562), .Y(n_619) );
BUFx2_ASAP7_75t_L g620 ( .A(n_562), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_542), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_574), .Y(n_622) );
OAI21x1_ASAP7_75t_L g623 ( .A1(n_592), .A2(n_223), .B(n_224), .Y(n_623) );
INVx2_ASAP7_75t_SL g624 ( .A(n_566), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_571), .B(n_228), .Y(n_625) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_552), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_574), .Y(n_627) );
NAND4xp25_ASAP7_75t_L g628 ( .A(n_547), .B(n_582), .C(n_578), .D(n_581), .Y(n_628) );
OAI21x1_ASAP7_75t_L g629 ( .A1(n_543), .A2(n_577), .B(n_540), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_578), .A2(n_581), .B1(n_580), .B2(n_563), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_560), .B(n_593), .Y(n_631) );
AO21x2_ASAP7_75t_L g632 ( .A1(n_541), .A2(n_540), .B(n_572), .Y(n_632) );
INVx3_ASAP7_75t_L g633 ( .A(n_567), .Y(n_633) );
OAI21x1_ASAP7_75t_L g634 ( .A1(n_572), .A2(n_565), .B(n_553), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_570), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_576), .B(n_555), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_570), .Y(n_637) );
INVx3_ASAP7_75t_L g638 ( .A(n_573), .Y(n_638) );
BUFx3_ASAP7_75t_L g639 ( .A(n_570), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_545), .Y(n_640) );
BUFx2_ASAP7_75t_L g641 ( .A(n_557), .Y(n_641) );
OAI21x1_ASAP7_75t_L g642 ( .A1(n_554), .A2(n_564), .B(n_568), .Y(n_642) );
AOI22xp33_ASAP7_75t_SL g643 ( .A1(n_541), .A2(n_573), .B1(n_587), .B2(n_589), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_538), .Y(n_644) );
INVx2_ASAP7_75t_SL g645 ( .A(n_590), .Y(n_645) );
CKINVDCx5p33_ASAP7_75t_R g646 ( .A(n_546), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_536), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_538), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_538), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_537), .B(n_590), .Y(n_650) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_537), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_536), .Y(n_652) );
OA21x2_ASAP7_75t_L g653 ( .A1(n_556), .A2(n_558), .B(n_583), .Y(n_653) );
BUFx12f_ASAP7_75t_L g654 ( .A(n_546), .Y(n_654) );
AND2x4_ASAP7_75t_L g655 ( .A(n_536), .B(n_537), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_536), .B(n_584), .Y(n_656) );
OAI22xp33_ASAP7_75t_L g657 ( .A1(n_574), .A2(n_535), .B1(n_537), .B2(n_445), .Y(n_657) );
O2A1O1Ixp33_ASAP7_75t_L g658 ( .A1(n_569), .A2(n_403), .B(n_372), .C(n_478), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_537), .B(n_590), .Y(n_659) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_548), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_538), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_536), .Y(n_662) );
AND2x4_ASAP7_75t_L g663 ( .A(n_536), .B(n_537), .Y(n_663) );
AO31x2_ASAP7_75t_L g664 ( .A1(n_556), .A2(n_558), .A3(n_579), .B(n_581), .Y(n_664) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_537), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_536), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_569), .B(n_485), .Y(n_667) );
INVx3_ASAP7_75t_L g668 ( .A(n_590), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_536), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_669), .B(n_647), .Y(n_670) );
AND2x2_ASAP7_75t_SL g671 ( .A(n_620), .B(n_615), .Y(n_671) );
AND2x4_ASAP7_75t_L g672 ( .A(n_605), .B(n_619), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_650), .B(n_659), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_598), .Y(n_674) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_651), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_599), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_644), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_655), .B(n_663), .Y(n_678) );
AO31x2_ASAP7_75t_L g679 ( .A1(n_637), .A2(n_635), .A3(n_630), .B(n_606), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_655), .B(n_663), .Y(n_680) );
OAI21xp5_ASAP7_75t_SL g681 ( .A1(n_657), .A2(n_605), .B(n_615), .Y(n_681) );
BUFx6f_ASAP7_75t_L g682 ( .A(n_660), .Y(n_682) );
INVx3_ASAP7_75t_L g683 ( .A(n_660), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_648), .B(n_649), .Y(n_684) );
INVx2_ASAP7_75t_R g685 ( .A(n_639), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_661), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_594), .B(n_645), .Y(n_687) );
INVxp67_ASAP7_75t_L g688 ( .A(n_651), .Y(n_688) );
AND2x4_ASAP7_75t_L g689 ( .A(n_622), .B(n_627), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_668), .B(n_665), .Y(n_690) );
BUFx3_ASAP7_75t_L g691 ( .A(n_596), .Y(n_691) );
AND2x4_ASAP7_75t_SL g692 ( .A(n_652), .B(n_669), .Y(n_692) );
INVxp67_ASAP7_75t_L g693 ( .A(n_611), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_667), .B(n_595), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_656), .B(n_597), .Y(n_695) );
BUFx2_ASAP7_75t_L g696 ( .A(n_604), .Y(n_696) );
INVxp67_ASAP7_75t_SL g697 ( .A(n_630), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_667), .B(n_610), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_662), .B(n_666), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_666), .B(n_604), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_603), .Y(n_701) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_612), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_624), .B(n_633), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_614), .B(n_616), .Y(n_704) );
OR2x2_ASAP7_75t_L g705 ( .A(n_608), .B(n_657), .Y(n_705) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_664), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_608), .Y(n_707) );
INVx4_ASAP7_75t_L g708 ( .A(n_660), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_616), .B(n_621), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_664), .Y(n_710) );
AND2x2_ASAP7_75t_L g711 ( .A(n_618), .B(n_658), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_664), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_658), .B(n_636), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_631), .B(n_625), .Y(n_714) );
AOI22xp33_ASAP7_75t_SL g715 ( .A1(n_641), .A2(n_607), .B1(n_639), .B2(n_632), .Y(n_715) );
BUFx3_ASAP7_75t_L g716 ( .A(n_654), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_640), .Y(n_717) );
AND2x2_ASAP7_75t_L g718 ( .A(n_646), .B(n_637), .Y(n_718) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_653), .Y(n_719) );
INVx3_ASAP7_75t_L g720 ( .A(n_626), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_602), .B(n_634), .Y(n_721) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_602), .Y(n_722) );
OR2x2_ASAP7_75t_L g723 ( .A(n_628), .B(n_632), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_613), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_623), .B(n_601), .Y(n_725) );
AND2x2_ASAP7_75t_L g726 ( .A(n_601), .B(n_629), .Y(n_726) );
AND2x4_ASAP7_75t_L g727 ( .A(n_609), .B(n_617), .Y(n_727) );
INVx5_ASAP7_75t_SL g728 ( .A(n_626), .Y(n_728) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_617), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_642), .B(n_600), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_626), .Y(n_731) );
INVxp67_ASAP7_75t_L g732 ( .A(n_638), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_638), .B(n_626), .Y(n_733) );
NOR2x1_ASAP7_75t_R g734 ( .A(n_643), .B(n_654), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_643), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_669), .B(n_647), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_657), .A2(n_620), .B1(n_574), .B2(n_628), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_650), .B(n_659), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_650), .B(n_659), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_689), .B(n_697), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_673), .B(n_738), .Y(n_741) );
AND2x2_ASAP7_75t_L g742 ( .A(n_678), .B(n_680), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_711), .B(n_709), .Y(n_743) );
AND2x2_ASAP7_75t_L g744 ( .A(n_739), .B(n_698), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_694), .B(n_687), .Y(n_745) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_675), .Y(n_746) );
INVx2_ASAP7_75t_SL g747 ( .A(n_692), .Y(n_747) );
OR2x2_ASAP7_75t_L g748 ( .A(n_675), .B(n_688), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_689), .B(n_697), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_690), .B(n_703), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_674), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_737), .A2(n_681), .B1(n_671), .B2(n_691), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_676), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_677), .Y(n_754) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_688), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_686), .Y(n_756) );
AND2x4_ASAP7_75t_L g757 ( .A(n_672), .B(n_733), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_713), .B(n_717), .Y(n_758) );
INVx2_ASAP7_75t_SL g759 ( .A(n_692), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_670), .B(n_736), .Y(n_760) );
AND2x2_ASAP7_75t_L g761 ( .A(n_670), .B(n_736), .Y(n_761) );
AND2x2_ASAP7_75t_L g762 ( .A(n_718), .B(n_700), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_684), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_702), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_701), .B(n_699), .Y(n_765) );
OR2x2_ASAP7_75t_L g766 ( .A(n_696), .B(n_695), .Y(n_766) );
INVx3_ASAP7_75t_L g767 ( .A(n_708), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_693), .B(n_737), .Y(n_768) );
AND2x2_ASAP7_75t_L g769 ( .A(n_671), .B(n_704), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_707), .B(n_714), .Y(n_770) );
BUFx4_ASAP7_75t_SL g771 ( .A(n_716), .Y(n_771) );
AND2x2_ASAP7_75t_L g772 ( .A(n_705), .B(n_735), .Y(n_772) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_722), .Y(n_773) );
AND2x4_ASAP7_75t_L g774 ( .A(n_720), .B(n_721), .Y(n_774) );
AND2x2_ASAP7_75t_L g775 ( .A(n_723), .B(n_708), .Y(n_775) );
BUFx2_ASAP7_75t_L g776 ( .A(n_734), .Y(n_776) );
INVx4_ASAP7_75t_L g777 ( .A(n_767), .Y(n_777) );
OR2x2_ASAP7_75t_SL g778 ( .A(n_771), .B(n_716), .Y(n_778) );
NAND2x1_ASAP7_75t_L g779 ( .A(n_776), .B(n_725), .Y(n_779) );
AND2x4_ASAP7_75t_L g780 ( .A(n_775), .B(n_732), .Y(n_780) );
OR2x2_ASAP7_75t_L g781 ( .A(n_760), .B(n_706), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_772), .B(n_712), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_750), .B(n_683), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_764), .B(n_712), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_751), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_763), .B(n_710), .Y(n_786) );
OR2x2_ASAP7_75t_L g787 ( .A(n_760), .B(n_679), .Y(n_787) );
OR2x2_ASAP7_75t_L g788 ( .A(n_761), .B(n_679), .Y(n_788) );
NOR2xp33_ASAP7_75t_L g789 ( .A(n_758), .B(n_732), .Y(n_789) );
NAND4xp25_ASAP7_75t_L g790 ( .A(n_758), .B(n_715), .C(n_730), .D(n_726), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_770), .B(n_679), .Y(n_791) );
INVx3_ASAP7_75t_L g792 ( .A(n_767), .Y(n_792) );
AND2x2_ASAP7_75t_L g793 ( .A(n_762), .B(n_685), .Y(n_793) );
AND2x2_ASAP7_75t_L g794 ( .A(n_741), .B(n_685), .Y(n_794) );
AND2x2_ASAP7_75t_L g795 ( .A(n_742), .B(n_682), .Y(n_795) );
OR2x2_ASAP7_75t_L g796 ( .A(n_761), .B(n_679), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_753), .Y(n_797) );
AND2x4_ASAP7_75t_L g798 ( .A(n_757), .B(n_731), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_746), .B(n_719), .Y(n_799) );
AND2x4_ASAP7_75t_L g800 ( .A(n_757), .B(n_727), .Y(n_800) );
INVx2_ASAP7_75t_SL g801 ( .A(n_771), .Y(n_801) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_773), .Y(n_802) );
AND2x2_ASAP7_75t_L g803 ( .A(n_745), .B(n_719), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_754), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_743), .B(n_724), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_756), .Y(n_806) );
AND2x2_ASAP7_75t_L g807 ( .A(n_743), .B(n_728), .Y(n_807) );
OR2x2_ASAP7_75t_L g808 ( .A(n_766), .B(n_729), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_744), .B(n_728), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_785), .Y(n_810) );
INVx2_ASAP7_75t_SL g811 ( .A(n_777), .Y(n_811) );
AND2x4_ASAP7_75t_L g812 ( .A(n_777), .B(n_774), .Y(n_812) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_805), .A2(n_752), .B1(n_768), .B2(n_769), .Y(n_813) );
OR2x2_ASAP7_75t_L g814 ( .A(n_781), .B(n_748), .Y(n_814) );
NOR2xp33_ASAP7_75t_L g815 ( .A(n_789), .B(n_755), .Y(n_815) );
HB1xp67_ASAP7_75t_L g816 ( .A(n_802), .Y(n_816) );
BUFx3_ASAP7_75t_L g817 ( .A(n_778), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_797), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_804), .Y(n_819) );
INVx2_ASAP7_75t_L g820 ( .A(n_784), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_806), .Y(n_821) );
AND2x2_ASAP7_75t_L g822 ( .A(n_803), .B(n_757), .Y(n_822) );
HB1xp67_ASAP7_75t_L g823 ( .A(n_802), .Y(n_823) );
AND2x2_ASAP7_75t_L g824 ( .A(n_787), .B(n_740), .Y(n_824) );
NOR2xp33_ASAP7_75t_SL g825 ( .A(n_801), .B(n_759), .Y(n_825) );
AND2x2_ASAP7_75t_L g826 ( .A(n_794), .B(n_749), .Y(n_826) );
AND2x4_ASAP7_75t_L g827 ( .A(n_780), .B(n_774), .Y(n_827) );
AND2x2_ASAP7_75t_L g828 ( .A(n_793), .B(n_740), .Y(n_828) );
INVxp67_ASAP7_75t_SL g829 ( .A(n_799), .Y(n_829) );
INVxp67_ASAP7_75t_L g830 ( .A(n_805), .Y(n_830) );
AND2x2_ASAP7_75t_L g831 ( .A(n_827), .B(n_800), .Y(n_831) );
OR2x2_ASAP7_75t_L g832 ( .A(n_829), .B(n_788), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_810), .Y(n_833) );
OR2x2_ASAP7_75t_L g834 ( .A(n_814), .B(n_796), .Y(n_834) );
INVx2_ASAP7_75t_L g835 ( .A(n_811), .Y(n_835) );
AND2x2_ASAP7_75t_L g836 ( .A(n_827), .B(n_800), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_820), .B(n_791), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_818), .Y(n_838) );
AND2x2_ASAP7_75t_L g839 ( .A(n_827), .B(n_795), .Y(n_839) );
OAI221xp5_ASAP7_75t_L g840 ( .A1(n_813), .A2(n_790), .B1(n_779), .B2(n_789), .C(n_791), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_819), .Y(n_841) );
OR2x2_ASAP7_75t_L g842 ( .A(n_820), .B(n_782), .Y(n_842) );
AOI22xp5_ASAP7_75t_L g843 ( .A1(n_825), .A2(n_790), .B1(n_807), .B2(n_759), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_837), .B(n_830), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_837), .B(n_824), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_834), .Y(n_846) );
OAI32xp33_ASAP7_75t_L g847 ( .A1(n_840), .A2(n_817), .A3(n_815), .B1(n_823), .B2(n_816), .Y(n_847) );
OR2x2_ASAP7_75t_L g848 ( .A(n_832), .B(n_816), .Y(n_848) );
INVxp67_ASAP7_75t_L g849 ( .A(n_835), .Y(n_849) );
AOI21xp33_ASAP7_75t_L g850 ( .A1(n_843), .A2(n_817), .B(n_815), .Y(n_850) );
AOI311xp33_ASAP7_75t_L g851 ( .A1(n_850), .A2(n_833), .A3(n_838), .B(n_841), .C(n_821), .Y(n_851) );
OAI22xp33_ASAP7_75t_L g852 ( .A1(n_850), .A2(n_843), .B1(n_747), .B2(n_792), .Y(n_852) );
AOI21xp5_ASAP7_75t_L g853 ( .A1(n_847), .A2(n_823), .B(n_812), .Y(n_853) );
OAI21xp33_ASAP7_75t_L g854 ( .A1(n_844), .A2(n_824), .B(n_842), .Y(n_854) );
AOI22xp5_ASAP7_75t_L g855 ( .A1(n_846), .A2(n_780), .B1(n_809), .B2(n_812), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_855), .Y(n_856) );
XNOR2xp5_ASAP7_75t_L g857 ( .A(n_852), .B(n_812), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_854), .Y(n_858) );
NAND3xp33_ASAP7_75t_L g859 ( .A(n_858), .B(n_851), .C(n_853), .Y(n_859) );
NOR4xp25_ASAP7_75t_L g860 ( .A(n_856), .B(n_849), .C(n_848), .D(n_845), .Y(n_860) );
NOR2x1_ASAP7_75t_L g861 ( .A(n_857), .B(n_792), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_859), .Y(n_862) );
NOR2xp67_ASAP7_75t_L g863 ( .A(n_860), .B(n_831), .Y(n_863) );
BUFx6f_ASAP7_75t_L g864 ( .A(n_862), .Y(n_864) );
NAND4xp75_ASAP7_75t_L g865 ( .A(n_863), .B(n_861), .C(n_836), .D(n_839), .Y(n_865) );
INVx2_ASAP7_75t_L g866 ( .A(n_864), .Y(n_866) );
AOI21xp5_ASAP7_75t_L g867 ( .A1(n_866), .A2(n_864), .B(n_865), .Y(n_867) );
AND2x2_ASAP7_75t_L g868 ( .A(n_867), .B(n_822), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_868), .Y(n_869) );
NAND3x2_ASAP7_75t_L g870 ( .A(n_869), .B(n_808), .C(n_798), .Y(n_870) );
OA21x2_ASAP7_75t_L g871 ( .A1(n_870), .A2(n_765), .B(n_786), .Y(n_871) );
INVxp67_ASAP7_75t_SL g872 ( .A(n_871), .Y(n_872) );
AOI22xp5_ASAP7_75t_L g873 ( .A1(n_872), .A2(n_828), .B1(n_826), .B2(n_783), .Y(n_873) );
endmodule