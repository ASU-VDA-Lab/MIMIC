module fake_ariane_3210_n_918 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_918);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_918;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_584;
wire n_528;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_349;
wire n_391;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_207;
wire n_857;
wire n_898;
wire n_790;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_193;
wire n_761;
wire n_733;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_754;
wire n_731;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_481;
wire n_433;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_839;
wire n_821;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_899;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_889;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_747;
wire n_772;
wire n_741;
wire n_847;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_916;
wire n_254;
wire n_596;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_915;
wire n_215;
wire n_252;
wire n_664;
wire n_629;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_882;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_184;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_353;
wire n_767;
wire n_736;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

INVx2_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_16),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_44),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g189 ( 
.A(n_62),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_143),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_103),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_47),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_65),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_79),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_152),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_70),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_90),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_13),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_149),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_3),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_41),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_180),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_127),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_88),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_67),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_145),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_139),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_106),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

BUFx10_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_110),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_133),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_36),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_21),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_181),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_43),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_102),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_86),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_128),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_89),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_156),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_95),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_87),
.Y(n_224)
);

BUFx10_ASAP7_75t_L g225 ( 
.A(n_24),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_138),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_66),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_183),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_2),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_21),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_92),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_6),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_98),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_129),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_136),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_82),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_115),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_142),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_2),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_148),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_68),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_59),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_3),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_15),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_83),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_23),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_153),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_18),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_155),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_80),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_119),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_130),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_94),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_33),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_50),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_101),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_251),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_185),
.Y(n_258)
);

INVxp33_ASAP7_75t_L g259 ( 
.A(n_214),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_251),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_253),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_0),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_206),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_229),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_199),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_186),
.B(n_0),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_244),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_201),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_206),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_191),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_239),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_191),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_191),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_211),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_248),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_246),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_211),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_211),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_225),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_225),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_190),
.Y(n_283)
);

INVxp67_ASAP7_75t_SL g284 ( 
.A(n_184),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_187),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_225),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_190),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_188),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_192),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_194),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_215),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_230),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_223),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_232),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_208),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_223),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_250),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_250),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_209),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_210),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_254),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_217),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_220),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_221),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_193),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_256),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_258),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_285),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_285),
.Y(n_309)
);

AND2x4_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_184),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_305),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_306),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_264),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_257),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_289),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_289),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_265),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_264),
.B(n_222),
.Y(n_318)
);

CKINVDCx9p33_ASAP7_75t_R g319 ( 
.A(n_260),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_270),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_268),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_305),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_278),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_283),
.Y(n_324)
);

NAND2x1_ASAP7_75t_L g325 ( 
.A(n_288),
.B(n_198),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_262),
.Y(n_326)
);

AND2x4_ASAP7_75t_L g327 ( 
.A(n_300),
.B(n_231),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_283),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_259),
.B(n_200),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_272),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_276),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_287),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_287),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_296),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_296),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_277),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_262),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_262),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_290),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_295),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_304),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_R g342 ( 
.A(n_297),
.B(n_195),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_299),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_297),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_298),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_266),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_284),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_302),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_298),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_303),
.B(n_213),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_304),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_267),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_291),
.Y(n_353)
);

BUFx8_ASAP7_75t_L g354 ( 
.A(n_281),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_271),
.B(n_234),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_269),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_263),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_293),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_293),
.Y(n_359)
);

CKINVDCx11_ASAP7_75t_R g360 ( 
.A(n_292),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_301),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_271),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_293),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_261),
.Y(n_364)
);

AO22x2_ASAP7_75t_L g365 ( 
.A1(n_329),
.A2(n_282),
.B1(n_286),
.B2(n_235),
.Y(n_365)
);

INVx5_ASAP7_75t_L g366 ( 
.A(n_309),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_341),
.Y(n_367)
);

NAND2xp33_ASAP7_75t_L g368 ( 
.A(n_357),
.B(n_189),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_357),
.B(n_273),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_341),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_357),
.B(n_347),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_329),
.B(n_261),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_309),
.Y(n_373)
);

INVx5_ASAP7_75t_L g374 ( 
.A(n_309),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_350),
.B(n_273),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_357),
.B(n_274),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g377 ( 
.A(n_341),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_309),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_358),
.A2(n_294),
.B1(n_274),
.B2(n_279),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_307),
.Y(n_380)
);

CKINVDCx8_ASAP7_75t_R g381 ( 
.A(n_312),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_351),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_357),
.B(n_240),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_309),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_364),
.B(n_275),
.Y(n_385)
);

INVx2_ASAP7_75t_SL g386 ( 
.A(n_351),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_308),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_317),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_308),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_330),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_327),
.B(n_241),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_323),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_352),
.B(n_196),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_323),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_315),
.Y(n_395)
);

BUFx10_ASAP7_75t_L g396 ( 
.A(n_358),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_353),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_315),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_331),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_355),
.B(n_197),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_311),
.Y(n_401)
);

AND2x2_ASAP7_75t_SL g402 ( 
.A(n_310),
.B(n_245),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_316),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_346),
.B(n_280),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_316),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_318),
.B(n_202),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g407 ( 
.A(n_353),
.B(n_1),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_336),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_339),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_316),
.Y(n_410)
);

OR2x2_ASAP7_75t_L g411 ( 
.A(n_361),
.B(n_4),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_340),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_343),
.Y(n_413)
);

OR2x6_ASAP7_75t_L g414 ( 
.A(n_361),
.B(n_247),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_327),
.B(n_249),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_325),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_362),
.B(n_313),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_311),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_325),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_327),
.B(n_252),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_310),
.B(n_4),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_310),
.B(n_203),
.Y(n_422)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_326),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_321),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_313),
.B(n_204),
.Y(n_425)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_326),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_342),
.B(n_198),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_337),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_348),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_337),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_314),
.Y(n_431)
);

OAI22xp33_ASAP7_75t_L g432 ( 
.A1(n_324),
.A2(n_226),
.B1(n_242),
.B2(n_238),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_338),
.Y(n_433)
);

AND2x6_ASAP7_75t_L g434 ( 
.A(n_338),
.B(n_198),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_324),
.B(n_5),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_359),
.B(n_205),
.Y(n_436)
);

OR2x2_ASAP7_75t_L g437 ( 
.A(n_328),
.B(n_5),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_356),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_401),
.B(n_322),
.Y(n_439)
);

NOR3xp33_ASAP7_75t_L g440 ( 
.A(n_432),
.B(n_333),
.C(n_332),
.Y(n_440)
);

INVx2_ASAP7_75t_SL g441 ( 
.A(n_401),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_369),
.B(n_332),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_402),
.A2(n_349),
.B1(n_335),
.B2(n_344),
.Y(n_443)
);

NAND2x1_ASAP7_75t_L g444 ( 
.A(n_423),
.B(n_198),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_375),
.B(n_333),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_428),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g447 ( 
.A(n_418),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_371),
.B(n_359),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_371),
.B(n_363),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_428),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_402),
.A2(n_354),
.B1(n_334),
.B2(n_345),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_370),
.B(n_363),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_400),
.B(n_334),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_369),
.B(n_376),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_406),
.B(n_344),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_418),
.B(n_189),
.Y(n_456)
);

NAND3xp33_ASAP7_75t_L g457 ( 
.A(n_436),
.B(n_354),
.C(n_320),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_377),
.B(n_403),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_L g459 ( 
.A1(n_365),
.A2(n_354),
.B1(n_224),
.B2(n_320),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_387),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_393),
.B(n_6),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_391),
.B(n_319),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_377),
.B(n_207),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_367),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_367),
.B(n_7),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_372),
.B(n_360),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_417),
.B(n_7),
.Y(n_467)
);

OR2x6_ASAP7_75t_L g468 ( 
.A(n_414),
.B(n_224),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_403),
.B(n_212),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_387),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_421),
.B(n_189),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_404),
.B(n_8),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_386),
.B(n_216),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_405),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_391),
.B(n_8),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_397),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g477 ( 
.A1(n_365),
.A2(n_421),
.B1(n_391),
.B2(n_420),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_386),
.B(n_218),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_425),
.B(n_9),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_389),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_389),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_436),
.B(n_219),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_431),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_382),
.B(n_9),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_382),
.B(n_227),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_L g486 ( 
.A1(n_365),
.A2(n_224),
.B1(n_189),
.B2(n_236),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_405),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_383),
.A2(n_255),
.B1(n_237),
.B2(n_228),
.Y(n_488)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_419),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_383),
.A2(n_189),
.B1(n_224),
.B2(n_12),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_380),
.B(n_189),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_388),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_423),
.B(n_10),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_390),
.B(n_189),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_424),
.B(n_11),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_397),
.Y(n_496)
);

OAI221xp5_ASAP7_75t_L g497 ( 
.A1(n_435),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.C(n_16),
.Y(n_497)
);

INVxp33_ASAP7_75t_L g498 ( 
.A(n_385),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_399),
.B(n_14),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_408),
.B(n_409),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_410),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_438),
.B(n_17),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_381),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_503)
);

AND2x6_ASAP7_75t_SL g504 ( 
.A(n_414),
.B(n_20),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_398),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_412),
.B(n_20),
.Y(n_506)
);

AND2x6_ASAP7_75t_SL g507 ( 
.A(n_414),
.B(n_22),
.Y(n_507)
);

CKINVDCx11_ASAP7_75t_R g508 ( 
.A(n_381),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_413),
.B(n_22),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_396),
.B(n_23),
.Y(n_510)
);

AO221x1_ASAP7_75t_L g511 ( 
.A1(n_432),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.C(n_27),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_379),
.Y(n_512)
);

NAND3xp33_ASAP7_75t_L g513 ( 
.A(n_423),
.B(n_25),
.C(n_26),
.Y(n_513)
);

AO22x1_ASAP7_75t_L g514 ( 
.A1(n_421),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_429),
.B(n_28),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_415),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_516)
);

INVx4_ASAP7_75t_L g517 ( 
.A(n_489),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_448),
.B(n_415),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_489),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_500),
.Y(n_520)
);

AND2x6_ASAP7_75t_L g521 ( 
.A(n_475),
.B(n_416),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_460),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_508),
.Y(n_523)
);

BUFx12f_ASAP7_75t_L g524 ( 
.A(n_508),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_462),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_R g526 ( 
.A(n_483),
.B(n_396),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_454),
.B(n_419),
.Y(n_527)
);

CKINVDCx8_ASAP7_75t_R g528 ( 
.A(n_462),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_443),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_447),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_449),
.B(n_415),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_453),
.B(n_420),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_512),
.A2(n_437),
.B1(n_420),
.B2(n_416),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_455),
.B(n_442),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_442),
.B(n_396),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_482),
.B(n_410),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_476),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_496),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_474),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_464),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_487),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_464),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_445),
.B(n_407),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_460),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_501),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_440),
.A2(n_427),
.B1(n_416),
.B2(n_422),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_454),
.B(n_419),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_441),
.B(n_419),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_470),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_466),
.Y(n_550)
);

INVx4_ASAP7_75t_L g551 ( 
.A(n_468),
.Y(n_551)
);

AO221x1_ASAP7_75t_L g552 ( 
.A1(n_503),
.A2(n_394),
.B1(n_392),
.B2(n_395),
.C(n_384),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_468),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_R g554 ( 
.A(n_451),
.B(n_411),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_470),
.Y(n_555)
);

AND2x6_ASAP7_75t_L g556 ( 
.A(n_475),
.B(n_373),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_446),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_480),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_450),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_468),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_480),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_467),
.B(n_427),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_481),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_481),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_505),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_505),
.Y(n_566)
);

NAND2x1p5_ASAP7_75t_L g567 ( 
.A(n_471),
.B(n_426),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_491),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_495),
.Y(n_569)
);

NAND3xp33_ASAP7_75t_L g570 ( 
.A(n_461),
.B(n_368),
.C(n_426),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_461),
.B(n_452),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_479),
.B(n_430),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_439),
.B(n_426),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_499),
.Y(n_574)
);

NOR3xp33_ASAP7_75t_SL g575 ( 
.A(n_497),
.B(n_433),
.C(n_31),
.Y(n_575)
);

AO31x2_ASAP7_75t_L g576 ( 
.A1(n_568),
.A2(n_493),
.A3(n_494),
.B(n_484),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g577 ( 
.A1(n_571),
.A2(n_439),
.B(n_471),
.Y(n_577)
);

NOR2x1_ASAP7_75t_L g578 ( 
.A(n_517),
.B(n_457),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_538),
.B(n_477),
.Y(n_579)
);

A2O1A1Ixp33_ASAP7_75t_L g580 ( 
.A1(n_534),
.A2(n_531),
.B(n_518),
.C(n_532),
.Y(n_580)
);

AOI211x1_ASAP7_75t_L g581 ( 
.A1(n_533),
.A2(n_514),
.B(n_492),
.C(n_515),
.Y(n_581)
);

OAI21x1_ASAP7_75t_L g582 ( 
.A1(n_527),
.A2(n_456),
.B(n_373),
.Y(n_582)
);

OAI21x1_ASAP7_75t_L g583 ( 
.A1(n_527),
.A2(n_456),
.B(n_458),
.Y(n_583)
);

AO21x1_ASAP7_75t_L g584 ( 
.A1(n_547),
.A2(n_493),
.B(n_484),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_535),
.B(n_477),
.Y(n_585)
);

OAI21x1_ASAP7_75t_L g586 ( 
.A1(n_547),
.A2(n_444),
.B(n_395),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_543),
.B(n_498),
.Y(n_587)
);

O2A1O1Ixp5_ASAP7_75t_L g588 ( 
.A1(n_571),
.A2(n_465),
.B(n_509),
.C(n_506),
.Y(n_588)
);

AOI221xp5_ASAP7_75t_L g589 ( 
.A1(n_529),
.A2(n_472),
.B1(n_516),
.B2(n_459),
.C(n_502),
.Y(n_589)
);

OA22x2_ASAP7_75t_L g590 ( 
.A1(n_550),
.A2(n_511),
.B1(n_510),
.B2(n_507),
.Y(n_590)
);

AO22x1_ASAP7_75t_L g591 ( 
.A1(n_521),
.A2(n_504),
.B1(n_459),
.B2(n_465),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_520),
.B(n_395),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_521),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g594 ( 
.A1(n_536),
.A2(n_463),
.B(n_469),
.Y(n_594)
);

AOI21x1_ASAP7_75t_L g595 ( 
.A1(n_574),
.A2(n_473),
.B(n_478),
.Y(n_595)
);

A2O1A1Ixp33_ASAP7_75t_L g596 ( 
.A1(n_573),
.A2(n_486),
.B(n_490),
.C(n_513),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_L g597 ( 
.A1(n_570),
.A2(n_368),
.B(n_486),
.Y(n_597)
);

OAI21x1_ASAP7_75t_L g598 ( 
.A1(n_568),
.A2(n_398),
.B(n_485),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_L g599 ( 
.A1(n_572),
.A2(n_488),
.B(n_366),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_525),
.B(n_392),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_521),
.B(n_392),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_525),
.B(n_392),
.Y(n_602)
);

CKINVDCx11_ASAP7_75t_R g603 ( 
.A(n_524),
.Y(n_603)
);

CKINVDCx8_ASAP7_75t_R g604 ( 
.A(n_523),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_573),
.A2(n_562),
.B(n_546),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_537),
.B(n_394),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_521),
.B(n_394),
.Y(n_607)
);

AOI221x1_ASAP7_75t_L g608 ( 
.A1(n_561),
.A2(n_394),
.B1(n_384),
.B2(n_378),
.C(n_374),
.Y(n_608)
);

AOI21x1_ASAP7_75t_L g609 ( 
.A1(n_539),
.A2(n_384),
.B(n_378),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_521),
.B(n_378),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_519),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_556),
.B(n_378),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_519),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_567),
.A2(n_384),
.B(n_366),
.Y(n_614)
);

OR2x6_ASAP7_75t_L g615 ( 
.A(n_551),
.B(n_366),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_541),
.Y(n_616)
);

OAI21x1_ASAP7_75t_L g617 ( 
.A1(n_567),
.A2(n_374),
.B(n_366),
.Y(n_617)
);

OR2x6_ASAP7_75t_L g618 ( 
.A(n_551),
.B(n_374),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_575),
.A2(n_374),
.B1(n_32),
.B2(n_33),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_L g620 ( 
.A1(n_545),
.A2(n_434),
.B(n_32),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_548),
.A2(n_109),
.B(n_179),
.Y(n_621)
);

OAI21x1_ASAP7_75t_L g622 ( 
.A1(n_522),
.A2(n_434),
.B(n_108),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_557),
.Y(n_623)
);

AOI21x1_ASAP7_75t_L g624 ( 
.A1(n_609),
.A2(n_559),
.B(n_565),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_616),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_587),
.B(n_537),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_585),
.B(n_553),
.Y(n_627)
);

OAI21x1_ASAP7_75t_L g628 ( 
.A1(n_598),
.A2(n_583),
.B(n_582),
.Y(n_628)
);

OAI21x1_ASAP7_75t_SL g629 ( 
.A1(n_577),
.A2(n_560),
.B(n_552),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_L g630 ( 
.A1(n_580),
.A2(n_575),
.B(n_548),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_623),
.Y(n_631)
);

AOI21xp33_ASAP7_75t_L g632 ( 
.A1(n_589),
.A2(n_569),
.B(n_563),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_L g633 ( 
.A1(n_605),
.A2(n_556),
.B(n_530),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_579),
.B(n_554),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_606),
.Y(n_635)
);

OAI21x1_ASAP7_75t_L g636 ( 
.A1(n_586),
.A2(n_544),
.B(n_558),
.Y(n_636)
);

OAI21x1_ASAP7_75t_L g637 ( 
.A1(n_622),
.A2(n_544),
.B(n_558),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_594),
.A2(n_542),
.B(n_540),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_592),
.Y(n_639)
);

OAI21x1_ASAP7_75t_SL g640 ( 
.A1(n_584),
.A2(n_522),
.B(n_556),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_592),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_591),
.B(n_528),
.Y(n_642)
);

OAI21x1_ASAP7_75t_L g643 ( 
.A1(n_595),
.A2(n_564),
.B(n_555),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_593),
.Y(n_644)
);

OAI21x1_ASAP7_75t_L g645 ( 
.A1(n_588),
.A2(n_564),
.B(n_555),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_602),
.Y(n_646)
);

OAI21xp5_ASAP7_75t_L g647 ( 
.A1(n_596),
.A2(n_434),
.B(n_526),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_600),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_593),
.B(n_519),
.Y(n_649)
);

OAI21x1_ASAP7_75t_SL g650 ( 
.A1(n_597),
.A2(n_599),
.B(n_620),
.Y(n_650)
);

A2O1A1Ixp33_ASAP7_75t_L g651 ( 
.A1(n_597),
.A2(n_542),
.B(n_540),
.C(n_566),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_L g652 ( 
.A1(n_599),
.A2(n_434),
.B(n_526),
.Y(n_652)
);

OR2x6_ASAP7_75t_SL g653 ( 
.A(n_619),
.B(n_540),
.Y(n_653)
);

INVx3_ASAP7_75t_SL g654 ( 
.A(n_590),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_578),
.Y(n_655)
);

AOI221xp5_ASAP7_75t_L g656 ( 
.A1(n_581),
.A2(n_566),
.B1(n_549),
.B2(n_542),
.C(n_540),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_576),
.B(n_542),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_611),
.B(n_549),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_619),
.B(n_549),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_611),
.B(n_549),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_608),
.A2(n_566),
.B(n_111),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_576),
.Y(n_662)
);

AO21x2_ASAP7_75t_L g663 ( 
.A1(n_612),
.A2(n_566),
.B(n_434),
.Y(n_663)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_576),
.B(n_30),
.Y(n_664)
);

INVxp67_ASAP7_75t_SL g665 ( 
.A(n_601),
.Y(n_665)
);

AOI21x1_ASAP7_75t_L g666 ( 
.A1(n_614),
.A2(n_107),
.B(n_176),
.Y(n_666)
);

OAI22xp33_ASAP7_75t_L g667 ( 
.A1(n_620),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_667)
);

OAI21x1_ASAP7_75t_L g668 ( 
.A1(n_617),
.A2(n_105),
.B(n_175),
.Y(n_668)
);

A2O1A1Ixp33_ASAP7_75t_L g669 ( 
.A1(n_621),
.A2(n_34),
.B(n_35),
.C(n_37),
.Y(n_669)
);

OAI21x1_ASAP7_75t_L g670 ( 
.A1(n_612),
.A2(n_112),
.B(n_174),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_626),
.Y(n_671)
);

O2A1O1Ixp33_ASAP7_75t_SL g672 ( 
.A1(n_669),
.A2(n_610),
.B(n_607),
.C(n_613),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_625),
.Y(n_673)
);

OAI21x1_ASAP7_75t_L g674 ( 
.A1(n_628),
.A2(n_613),
.B(n_618),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_SL g675 ( 
.A1(n_634),
.A2(n_618),
.B1(n_615),
.B2(n_603),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_631),
.Y(n_676)
);

CKINVDCx11_ASAP7_75t_R g677 ( 
.A(n_654),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_657),
.Y(n_678)
);

NAND2x1p5_ASAP7_75t_L g679 ( 
.A(n_644),
.B(n_615),
.Y(n_679)
);

AOI222xp33_ASAP7_75t_L g680 ( 
.A1(n_654),
.A2(n_37),
.B1(n_38),
.B2(n_604),
.C1(n_618),
.C2(n_615),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_653),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_681)
);

BUFx2_ASAP7_75t_L g682 ( 
.A(n_635),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_649),
.B(n_42),
.Y(n_683)
);

OAI221xp5_ASAP7_75t_L g684 ( 
.A1(n_630),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.C(n_49),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_646),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_642),
.B(n_51),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_627),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_649),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_627),
.Y(n_689)
);

NAND2xp33_ASAP7_75t_L g690 ( 
.A(n_669),
.B(n_52),
.Y(n_690)
);

NOR3xp33_ASAP7_75t_SL g691 ( 
.A(n_667),
.B(n_53),
.C(n_54),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_639),
.Y(n_692)
);

AOI21xp33_ASAP7_75t_L g693 ( 
.A1(n_650),
.A2(n_55),
.B(n_56),
.Y(n_693)
);

AND2x2_ASAP7_75t_SL g694 ( 
.A(n_664),
.B(n_57),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_648),
.B(n_655),
.Y(n_695)
);

A2O1A1Ixp33_ASAP7_75t_L g696 ( 
.A1(n_647),
.A2(n_58),
.B(n_60),
.C(n_61),
.Y(n_696)
);

NAND2xp33_ASAP7_75t_SL g697 ( 
.A(n_644),
.B(n_63),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_664),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_641),
.B(n_64),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_649),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_658),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_644),
.B(n_69),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_633),
.B(n_71),
.Y(n_703)
);

OAI21xp5_ASAP7_75t_L g704 ( 
.A1(n_651),
.A2(n_72),
.B(n_73),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_659),
.Y(n_705)
);

NAND2x1_ASAP7_75t_L g706 ( 
.A(n_629),
.B(n_74),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_660),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_653),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_632),
.A2(n_78),
.B1(n_81),
.B2(n_84),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_665),
.B(n_85),
.Y(n_710)
);

NOR2xp67_ASAP7_75t_L g711 ( 
.A(n_638),
.B(n_91),
.Y(n_711)
);

BUFx2_ASAP7_75t_SL g712 ( 
.A(n_662),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_651),
.B(n_93),
.Y(n_713)
);

NAND3xp33_ASAP7_75t_L g714 ( 
.A(n_656),
.B(n_96),
.C(n_97),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_645),
.Y(n_715)
);

INVx5_ASAP7_75t_L g716 ( 
.A(n_662),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_652),
.B(n_99),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_SL g718 ( 
.A1(n_640),
.A2(n_100),
.B1(n_104),
.B2(n_113),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_643),
.B(n_114),
.Y(n_719)
);

CKINVDCx16_ASAP7_75t_R g720 ( 
.A(n_663),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_643),
.Y(n_721)
);

OAI22xp33_ASAP7_75t_L g722 ( 
.A1(n_661),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_645),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_624),
.Y(n_724)
);

OAI22xp33_ASAP7_75t_L g725 ( 
.A1(n_681),
.A2(n_708),
.B1(n_684),
.B2(n_671),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_682),
.B(n_636),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_687),
.B(n_689),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_673),
.Y(n_728)
);

AOI221xp5_ASAP7_75t_L g729 ( 
.A1(n_681),
.A2(n_663),
.B1(n_670),
.B2(n_666),
.C(n_636),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_694),
.A2(n_670),
.B1(n_637),
.B2(n_668),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_680),
.A2(n_637),
.B1(n_668),
.B2(n_628),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_707),
.B(n_120),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_676),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_708),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_734)
);

OAI22xp33_ASAP7_75t_L g735 ( 
.A1(n_684),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_735)
);

AOI21xp33_ASAP7_75t_L g736 ( 
.A1(n_690),
.A2(n_131),
.B(n_132),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_677),
.A2(n_134),
.B1(n_135),
.B2(n_137),
.Y(n_737)
);

OAI22xp33_ASAP7_75t_SL g738 ( 
.A1(n_698),
.A2(n_140),
.B1(n_141),
.B2(n_144),
.Y(n_738)
);

AOI221xp5_ASAP7_75t_L g739 ( 
.A1(n_685),
.A2(n_691),
.B1(n_693),
.B2(n_686),
.C(n_672),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_675),
.A2(n_146),
.B1(n_147),
.B2(n_150),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_SL g741 ( 
.A1(n_713),
.A2(n_151),
.B1(n_154),
.B2(n_157),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_701),
.A2(n_158),
.B1(n_160),
.B2(n_162),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_692),
.Y(n_743)
);

AOI222xp33_ASAP7_75t_L g744 ( 
.A1(n_704),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.C1(n_166),
.C2(n_168),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_713),
.A2(n_169),
.B1(n_170),
.B2(n_172),
.Y(n_745)
);

OAI211xp5_ASAP7_75t_SL g746 ( 
.A1(n_691),
.A2(n_173),
.B(n_177),
.C(n_693),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_705),
.B(n_695),
.Y(n_747)
);

AND2x6_ASAP7_75t_SL g748 ( 
.A(n_683),
.B(n_699),
.Y(n_748)
);

OAI22xp33_ASAP7_75t_L g749 ( 
.A1(n_705),
.A2(n_714),
.B1(n_699),
.B2(n_710),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_703),
.A2(n_675),
.B1(n_697),
.B2(n_717),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_678),
.A2(n_709),
.B1(n_720),
.B2(n_710),
.Y(n_751)
);

OAI21x1_ASAP7_75t_L g752 ( 
.A1(n_674),
.A2(n_706),
.B(n_724),
.Y(n_752)
);

BUFx4f_ASAP7_75t_SL g753 ( 
.A(n_700),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_678),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_696),
.A2(n_718),
.B1(n_702),
.B2(n_679),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_712),
.Y(n_756)
);

BUFx4f_ASAP7_75t_L g757 ( 
.A(n_683),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_718),
.A2(n_688),
.B1(n_716),
.B2(n_722),
.Y(n_758)
);

AOI221xp5_ASAP7_75t_L g759 ( 
.A1(n_723),
.A2(n_702),
.B1(n_719),
.B2(n_721),
.C(n_688),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_716),
.A2(n_711),
.B1(n_679),
.B2(n_715),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_715),
.Y(n_761)
);

OA21x2_ASAP7_75t_L g762 ( 
.A1(n_716),
.A2(n_628),
.B(n_724),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_716),
.Y(n_763)
);

OAI22xp5_ASAP7_75t_L g764 ( 
.A1(n_691),
.A2(n_653),
.B1(n_451),
.B2(n_529),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_L g765 ( 
.A1(n_691),
.A2(n_653),
.B1(n_451),
.B2(n_529),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_682),
.B(n_671),
.Y(n_766)
);

AO22x1_ASAP7_75t_L g767 ( 
.A1(n_681),
.A2(n_708),
.B1(n_654),
.B2(n_671),
.Y(n_767)
);

OAI22xp33_ASAP7_75t_SL g768 ( 
.A1(n_681),
.A2(n_654),
.B1(n_653),
.B2(n_708),
.Y(n_768)
);

AOI221xp5_ASAP7_75t_L g769 ( 
.A1(n_681),
.A2(n_512),
.B1(n_451),
.B2(n_503),
.C(n_554),
.Y(n_769)
);

BUFx2_ASAP7_75t_L g770 ( 
.A(n_761),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_757),
.Y(n_771)
);

OAI22xp33_ASAP7_75t_L g772 ( 
.A1(n_764),
.A2(n_765),
.B1(n_757),
.B2(n_725),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_762),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_756),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_762),
.Y(n_775)
);

CKINVDCx6p67_ASAP7_75t_R g776 ( 
.A(n_766),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_747),
.B(n_762),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_726),
.B(n_754),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_763),
.B(n_752),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_728),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_733),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_743),
.Y(n_782)
);

OR2x2_ASAP7_75t_SL g783 ( 
.A(n_767),
.B(n_725),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_753),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_727),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_748),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_753),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_730),
.B(n_759),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_732),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_760),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_749),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_755),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_729),
.Y(n_793)
);

AND2x4_ASAP7_75t_L g794 ( 
.A(n_730),
.B(n_758),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_731),
.B(n_750),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_740),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_749),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_739),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_731),
.B(n_750),
.Y(n_799)
);

INVx2_ASAP7_75t_R g800 ( 
.A(n_768),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_738),
.Y(n_801)
);

INVx2_ASAP7_75t_R g802 ( 
.A(n_735),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_745),
.B(n_744),
.Y(n_803)
);

OAI31xp33_ASAP7_75t_SL g804 ( 
.A1(n_772),
.A2(n_735),
.A3(n_746),
.B(n_769),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_782),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_776),
.Y(n_806)
);

INVxp67_ASAP7_75t_SL g807 ( 
.A(n_773),
.Y(n_807)
);

OAI211xp5_ASAP7_75t_L g808 ( 
.A1(n_798),
.A2(n_745),
.B(n_734),
.C(n_741),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_773),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_782),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_782),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_776),
.B(n_737),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_777),
.B(n_751),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_803),
.A2(n_736),
.B1(n_742),
.B2(n_802),
.Y(n_814)
);

BUFx2_ASAP7_75t_SL g815 ( 
.A(n_787),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_777),
.B(n_779),
.Y(n_816)
);

AOI221xp5_ASAP7_75t_L g817 ( 
.A1(n_798),
.A2(n_793),
.B1(n_791),
.B2(n_797),
.C(n_795),
.Y(n_817)
);

NAND3xp33_ASAP7_75t_L g818 ( 
.A(n_791),
.B(n_797),
.C(n_803),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_780),
.Y(n_819)
);

AOI222xp33_ASAP7_75t_L g820 ( 
.A1(n_803),
.A2(n_795),
.B1(n_799),
.B2(n_794),
.C1(n_797),
.C2(n_796),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_780),
.Y(n_821)
);

BUFx2_ASAP7_75t_SL g822 ( 
.A(n_787),
.Y(n_822)
);

NOR5xp2_ASAP7_75t_SL g823 ( 
.A(n_783),
.B(n_802),
.C(n_772),
.D(n_776),
.E(n_800),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_777),
.B(n_778),
.Y(n_824)
);

NAND3xp33_ASAP7_75t_L g825 ( 
.A(n_793),
.B(n_792),
.C(n_799),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_816),
.B(n_824),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_805),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_824),
.B(n_785),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_816),
.B(n_774),
.Y(n_829)
);

NAND2x1_ASAP7_75t_SL g830 ( 
.A(n_816),
.B(n_786),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_816),
.B(n_774),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_825),
.B(n_785),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_825),
.B(n_778),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_813),
.B(n_774),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_813),
.B(n_778),
.Y(n_835)
);

OR2x2_ASAP7_75t_L g836 ( 
.A(n_805),
.B(n_793),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_815),
.B(n_770),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_810),
.B(n_779),
.Y(n_838)
);

OR2x2_ASAP7_75t_L g839 ( 
.A(n_811),
.B(n_793),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_811),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_809),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_826),
.B(n_815),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_832),
.B(n_820),
.Y(n_843)
);

AOI211xp5_ASAP7_75t_L g844 ( 
.A1(n_833),
.A2(n_818),
.B(n_804),
.C(n_812),
.Y(n_844)
);

OAI21xp33_ASAP7_75t_L g845 ( 
.A1(n_834),
.A2(n_788),
.B(n_795),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_826),
.B(n_831),
.Y(n_846)
);

OAI31xp33_ASAP7_75t_L g847 ( 
.A1(n_836),
.A2(n_818),
.A3(n_799),
.B(n_808),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_836),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_827),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_839),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_839),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_827),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_849),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_849),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_844),
.B(n_835),
.Y(n_855)
);

INVx1_ASAP7_75t_SL g856 ( 
.A(n_843),
.Y(n_856)
);

NAND4xp25_ASAP7_75t_L g857 ( 
.A(n_847),
.B(n_814),
.C(n_817),
.D(n_845),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_842),
.Y(n_858)
);

AOI221xp5_ASAP7_75t_L g859 ( 
.A1(n_848),
.A2(n_788),
.B1(n_794),
.B2(n_792),
.C(n_786),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_846),
.B(n_829),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_850),
.B(n_835),
.Y(n_861)
);

AOI221xp5_ASAP7_75t_L g862 ( 
.A1(n_851),
.A2(n_788),
.B1(n_794),
.B2(n_792),
.C(n_786),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_852),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_857),
.A2(n_786),
.B1(n_801),
.B2(n_794),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_854),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_853),
.Y(n_866)
);

AOI221xp5_ASAP7_75t_L g867 ( 
.A1(n_857),
.A2(n_794),
.B1(n_792),
.B2(n_786),
.C(n_801),
.Y(n_867)
);

NAND2xp33_ASAP7_75t_SL g868 ( 
.A(n_855),
.B(n_806),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_863),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_866),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_869),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_865),
.Y(n_872)
);

INVxp67_ASAP7_75t_L g873 ( 
.A(n_868),
.Y(n_873)
);

NAND2xp33_ASAP7_75t_SL g874 ( 
.A(n_872),
.B(n_860),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_870),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_871),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_873),
.B(n_864),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_875),
.B(n_856),
.Y(n_878)
);

NAND2x1_ASAP7_75t_L g879 ( 
.A(n_876),
.B(n_846),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_877),
.Y(n_880)
);

OAI21xp33_ASAP7_75t_L g881 ( 
.A1(n_874),
.A2(n_873),
.B(n_867),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_876),
.Y(n_882)
);

INVxp67_ASAP7_75t_L g883 ( 
.A(n_877),
.Y(n_883)
);

AOI211xp5_ASAP7_75t_SL g884 ( 
.A1(n_875),
.A2(n_862),
.B(n_859),
.C(n_861),
.Y(n_884)
);

AOI211xp5_ASAP7_75t_L g885 ( 
.A1(n_881),
.A2(n_858),
.B(n_784),
.C(n_801),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_880),
.Y(n_886)
);

NAND3xp33_ASAP7_75t_L g887 ( 
.A(n_883),
.B(n_801),
.C(n_852),
.Y(n_887)
);

AOI211xp5_ASAP7_75t_L g888 ( 
.A1(n_878),
.A2(n_784),
.B(n_796),
.C(n_787),
.Y(n_888)
);

XNOR2xp5_ASAP7_75t_L g889 ( 
.A(n_879),
.B(n_783),
.Y(n_889)
);

OAI221xp5_ASAP7_75t_L g890 ( 
.A1(n_884),
.A2(n_830),
.B1(n_796),
.B2(n_823),
.C(n_789),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_886),
.Y(n_891)
);

OAI211xp5_ASAP7_75t_SL g892 ( 
.A1(n_885),
.A2(n_882),
.B(n_784),
.C(n_828),
.Y(n_892)
);

XNOR2x1_ASAP7_75t_L g893 ( 
.A(n_889),
.B(n_823),
.Y(n_893)
);

NOR2xp67_ASAP7_75t_L g894 ( 
.A(n_887),
.B(n_842),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_890),
.A2(n_783),
.B1(n_834),
.B2(n_787),
.Y(n_895)
);

XNOR2xp5_ASAP7_75t_L g896 ( 
.A(n_888),
.B(n_789),
.Y(n_896)
);

NOR2x1_ASAP7_75t_L g897 ( 
.A(n_892),
.B(n_822),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_893),
.Y(n_898)
);

NOR2x1p5_ASAP7_75t_L g899 ( 
.A(n_891),
.B(n_837),
.Y(n_899)
);

AO22x1_ASAP7_75t_L g900 ( 
.A1(n_895),
.A2(n_837),
.B1(n_829),
.B2(n_831),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_894),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_898),
.A2(n_896),
.B1(n_796),
.B2(n_789),
.Y(n_902)
);

OR3x2_ASAP7_75t_L g903 ( 
.A(n_901),
.B(n_823),
.C(n_830),
.Y(n_903)
);

OAI322xp33_ASAP7_75t_L g904 ( 
.A1(n_899),
.A2(n_819),
.A3(n_821),
.B1(n_840),
.B2(n_781),
.C1(n_807),
.C2(n_775),
.Y(n_904)
);

NAND3xp33_ASAP7_75t_SL g905 ( 
.A(n_897),
.B(n_802),
.C(n_800),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_905),
.A2(n_900),
.B(n_819),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_903),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_907),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_906),
.Y(n_909)
);

AO22x2_ASAP7_75t_L g910 ( 
.A1(n_908),
.A2(n_902),
.B1(n_904),
.B2(n_822),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_909),
.A2(n_802),
.B1(n_800),
.B2(n_794),
.Y(n_911)
);

BUFx2_ASAP7_75t_L g912 ( 
.A(n_910),
.Y(n_912)
);

INVxp33_ASAP7_75t_SL g913 ( 
.A(n_911),
.Y(n_913)
);

OAI21x1_ASAP7_75t_SL g914 ( 
.A1(n_912),
.A2(n_821),
.B(n_800),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_914),
.A2(n_913),
.B1(n_838),
.B2(n_779),
.Y(n_915)
);

AOI322xp5_ASAP7_75t_L g916 ( 
.A1(n_915),
.A2(n_838),
.A3(n_790),
.B1(n_841),
.B2(n_773),
.C1(n_775),
.C2(n_809),
.Y(n_916)
);

AOI221xp5_ASAP7_75t_L g917 ( 
.A1(n_916),
.A2(n_838),
.B1(n_841),
.B2(n_779),
.C(n_790),
.Y(n_917)
);

AOI211xp5_ASAP7_75t_L g918 ( 
.A1(n_917),
.A2(n_771),
.B(n_779),
.C(n_781),
.Y(n_918)
);


endmodule