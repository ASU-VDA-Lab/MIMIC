module fake_netlist_1_353_n_26 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_26);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_26;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
INVx1_ASAP7_75t_L g11 ( .A(n_1), .Y(n_11) );
INVx3_ASAP7_75t_L g12 ( .A(n_9), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_3), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_10), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_12), .Y(n_16) );
AND2x4_ASAP7_75t_L g17 ( .A(n_12), .B(n_0), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_16), .B(n_13), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_18), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_19), .B(n_17), .Y(n_20) );
A2O1A1Ixp33_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_15), .B(n_14), .C(n_11), .Y(n_21) );
XNOR2x1_ASAP7_75t_L g22 ( .A(n_21), .B(n_0), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_21), .B(n_13), .Y(n_23) );
OAI221xp5_ASAP7_75t_L g24 ( .A1(n_22), .A2(n_2), .B1(n_4), .B2(n_5), .C(n_6), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
AOI22xp33_ASAP7_75t_SL g26 ( .A1(n_25), .A2(n_23), .B1(n_7), .B2(n_8), .Y(n_26) );
endmodule