module fake_netlist_1_330_n_638 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_638);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_638;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_SL g75 ( .A(n_65), .Y(n_75) );
BUFx6f_ASAP7_75t_L g76 ( .A(n_53), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_5), .Y(n_77) );
HB1xp67_ASAP7_75t_L g78 ( .A(n_34), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_61), .Y(n_79) );
INVx1_ASAP7_75t_SL g80 ( .A(n_18), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_0), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_31), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_1), .Y(n_83) );
INVx4_ASAP7_75t_R g84 ( .A(n_40), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_70), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_74), .Y(n_86) );
NOR2xp33_ASAP7_75t_L g87 ( .A(n_19), .B(n_22), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_13), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_49), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_71), .Y(n_90) );
CKINVDCx16_ASAP7_75t_R g91 ( .A(n_28), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_1), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_38), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_35), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_43), .Y(n_95) );
INVxp67_ASAP7_75t_L g96 ( .A(n_69), .Y(n_96) );
INVxp33_ASAP7_75t_SL g97 ( .A(n_12), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_48), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_62), .Y(n_99) );
INVx1_ASAP7_75t_SL g100 ( .A(n_50), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_13), .Y(n_101) );
CKINVDCx14_ASAP7_75t_R g102 ( .A(n_27), .Y(n_102) );
INVxp67_ASAP7_75t_SL g103 ( .A(n_11), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_52), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_41), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_54), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_56), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_15), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_4), .Y(n_109) );
BUFx3_ASAP7_75t_L g110 ( .A(n_29), .Y(n_110) );
BUFx2_ASAP7_75t_L g111 ( .A(n_26), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_36), .Y(n_112) );
INVxp33_ASAP7_75t_SL g113 ( .A(n_42), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_60), .Y(n_114) );
INVxp67_ASAP7_75t_L g115 ( .A(n_33), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_8), .Y(n_116) );
INVxp67_ASAP7_75t_SL g117 ( .A(n_17), .Y(n_117) );
CKINVDCx14_ASAP7_75t_R g118 ( .A(n_2), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_23), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_14), .Y(n_120) );
CKINVDCx16_ASAP7_75t_R g121 ( .A(n_91), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_111), .B(n_0), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_118), .Y(n_123) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_83), .Y(n_124) );
INVx3_ASAP7_75t_L g125 ( .A(n_108), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_108), .Y(n_126) );
NOR2xp33_ASAP7_75t_R g127 ( .A(n_102), .B(n_30), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_91), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_111), .B(n_2), .Y(n_129) );
AND2x4_ASAP7_75t_L g130 ( .A(n_108), .B(n_3), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_104), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_113), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_120), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_78), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_120), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_120), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_90), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_79), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_90), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_79), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_110), .B(n_3), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_85), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_97), .B(n_4), .Y(n_143) );
OR2x2_ASAP7_75t_L g144 ( .A(n_77), .B(n_5), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_85), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_90), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_86), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_76), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_76), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_86), .Y(n_150) );
XOR2xp5_ASAP7_75t_L g151 ( .A(n_103), .B(n_6), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_105), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_89), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_96), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_115), .Y(n_155) );
BUFx3_ASAP7_75t_L g156 ( .A(n_110), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_89), .B(n_6), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_105), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_110), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_105), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_77), .B(n_7), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_154), .B(n_119), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_155), .B(n_119), .Y(n_163) );
AND3x1_ASAP7_75t_L g164 ( .A(n_143), .B(n_101), .C(n_116), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_129), .B(n_88), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_138), .B(n_95), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_149), .Y(n_167) );
HB1xp67_ASAP7_75t_L g168 ( .A(n_121), .Y(n_168) );
BUFx3_ASAP7_75t_L g169 ( .A(n_156), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_137), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_156), .Y(n_171) );
BUFx3_ASAP7_75t_L g172 ( .A(n_156), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_130), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_149), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_137), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_138), .B(n_95), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_139), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_139), .Y(n_178) );
NAND2x1_ASAP7_75t_L g179 ( .A(n_141), .B(n_84), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_140), .B(n_99), .Y(n_180) );
NOR2x1p5_ASAP7_75t_L g181 ( .A(n_131), .B(n_117), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_148), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_130), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_148), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_130), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_130), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_129), .B(n_116), .Y(n_187) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_149), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_148), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_149), .Y(n_190) );
BUFx2_ASAP7_75t_L g191 ( .A(n_121), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_159), .A2(n_81), .B1(n_88), .B2(n_109), .Y(n_192) );
INVx8_ASAP7_75t_L g193 ( .A(n_141), .Y(n_193) );
AND2x4_ASAP7_75t_L g194 ( .A(n_141), .B(n_101), .Y(n_194) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_124), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_161), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_149), .Y(n_197) );
NAND2x1p5_ASAP7_75t_L g198 ( .A(n_141), .B(n_114), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_132), .B(n_114), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_161), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_128), .Y(n_201) );
BUFx2_ASAP7_75t_L g202 ( .A(n_134), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_140), .B(n_112), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_146), .Y(n_204) );
OR2x2_ASAP7_75t_L g205 ( .A(n_122), .B(n_109), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_148), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_142), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_142), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_145), .B(n_112), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_145), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_146), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_147), .B(n_99), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_193), .B(n_127), .Y(n_213) );
BUFx12f_ASAP7_75t_L g214 ( .A(n_191), .Y(n_214) );
BUFx2_ASAP7_75t_L g215 ( .A(n_195), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_171), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_202), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_171), .Y(n_218) );
OR2x2_ASAP7_75t_L g219 ( .A(n_191), .B(n_144), .Y(n_219) );
BUFx2_ASAP7_75t_L g220 ( .A(n_193), .Y(n_220) );
AND2x4_ASAP7_75t_L g221 ( .A(n_196), .B(n_144), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_165), .B(n_147), .Y(n_222) );
OR2x6_ASAP7_75t_L g223 ( .A(n_193), .B(n_198), .Y(n_223) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_202), .Y(n_224) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_201), .Y(n_225) );
INVx4_ASAP7_75t_L g226 ( .A(n_193), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_165), .B(n_150), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_173), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_173), .Y(n_229) );
INVx4_ASAP7_75t_L g230 ( .A(n_198), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_187), .B(n_150), .Y(n_231) );
OAI22xp5_ASAP7_75t_SL g232 ( .A1(n_201), .A2(n_151), .B1(n_164), .B2(n_123), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_194), .A2(n_153), .B1(n_157), .B2(n_81), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_187), .B(n_153), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_170), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_187), .B(n_80), .Y(n_236) );
BUFx2_ASAP7_75t_L g237 ( .A(n_168), .Y(n_237) );
INVx3_ASAP7_75t_L g238 ( .A(n_173), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_205), .B(n_125), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_170), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_175), .Y(n_241) );
BUFx10_ASAP7_75t_L g242 ( .A(n_199), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_175), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_177), .Y(n_244) );
INVxp67_ASAP7_75t_L g245 ( .A(n_162), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_200), .B(n_125), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_177), .Y(n_247) );
BUFx3_ASAP7_75t_L g248 ( .A(n_169), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_178), .Y(n_249) );
OR2x6_ASAP7_75t_L g250 ( .A(n_198), .B(n_92), .Y(n_250) );
NOR3xp33_ASAP7_75t_SL g251 ( .A(n_163), .B(n_203), .C(n_209), .Y(n_251) );
INVx4_ASAP7_75t_SL g252 ( .A(n_194), .Y(n_252) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_205), .Y(n_253) );
INVx2_ASAP7_75t_SL g254 ( .A(n_194), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_207), .B(n_125), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_178), .Y(n_256) );
AND2x4_ASAP7_75t_L g257 ( .A(n_183), .B(n_92), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_208), .B(n_80), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_204), .Y(n_259) );
AND2x4_ASAP7_75t_L g260 ( .A(n_185), .B(n_125), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_204), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_211), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_211), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_210), .B(n_126), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_186), .B(n_166), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_169), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_176), .Y(n_267) );
CKINVDCx20_ASAP7_75t_R g268 ( .A(n_192), .Y(n_268) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_179), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_180), .B(n_126), .Y(n_270) );
BUFx8_ASAP7_75t_L g271 ( .A(n_172), .Y(n_271) );
OAI22xp5_ASAP7_75t_SL g272 ( .A1(n_179), .A2(n_151), .B1(n_133), .B2(n_135), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_212), .Y(n_273) );
A2O1A1Ixp33_ASAP7_75t_L g274 ( .A1(n_267), .A2(n_152), .B(n_160), .C(n_158), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_245), .B(n_172), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_267), .B(n_181), .Y(n_276) );
INVx5_ASAP7_75t_L g277 ( .A(n_223), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_273), .A2(n_160), .B1(n_158), .B2(n_152), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_223), .Y(n_279) );
AOI22xp33_ASAP7_75t_SL g280 ( .A1(n_272), .A2(n_136), .B1(n_135), .B2(n_133), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_253), .B(n_136), .Y(n_281) );
A2O1A1Ixp33_ASAP7_75t_L g282 ( .A1(n_273), .A2(n_94), .B(n_107), .C(n_106), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_215), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_238), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_238), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_223), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_265), .A2(n_75), .B(n_82), .Y(n_287) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_223), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_238), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_235), .Y(n_290) );
INVx3_ASAP7_75t_L g291 ( .A(n_226), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_219), .B(n_7), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_222), .Y(n_293) );
INVx3_ASAP7_75t_L g294 ( .A(n_226), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_235), .Y(n_295) );
BUFx3_ASAP7_75t_L g296 ( .A(n_271), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_222), .B(n_100), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_227), .Y(n_298) );
NAND2x1p5_ASAP7_75t_L g299 ( .A(n_230), .B(n_100), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_226), .B(n_93), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_230), .B(n_98), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_230), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_227), .Y(n_303) );
INVxp67_ASAP7_75t_L g304 ( .A(n_220), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_260), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_250), .B(n_94), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_250), .Y(n_307) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_250), .Y(n_308) );
INVx3_ASAP7_75t_L g309 ( .A(n_250), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_228), .A2(n_106), .B(n_107), .Y(n_310) );
INVx2_ASAP7_75t_SL g311 ( .A(n_237), .Y(n_311) );
O2A1O1Ixp33_ASAP7_75t_L g312 ( .A1(n_234), .A2(n_107), .B(n_106), .C(n_87), .Y(n_312) );
OAI22xp33_ASAP7_75t_L g313 ( .A1(n_233), .A2(n_76), .B1(n_148), .B2(n_149), .Y(n_313) );
AND2x6_ASAP7_75t_L g314 ( .A(n_252), .B(n_76), .Y(n_314) );
NAND2x1_ASAP7_75t_L g315 ( .A(n_228), .B(n_84), .Y(n_315) );
AOI22x1_ASAP7_75t_L g316 ( .A1(n_229), .A2(n_206), .B1(n_182), .B2(n_184), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_241), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_237), .B(n_9), .Y(n_318) );
INVx6_ASAP7_75t_L g319 ( .A(n_271), .Y(n_319) );
AND2x2_ASAP7_75t_SL g320 ( .A(n_220), .B(n_76), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_260), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_271), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_241), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_233), .B(n_9), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_290), .Y(n_325) );
NAND2xp5_ASAP7_75t_SL g326 ( .A(n_308), .B(n_252), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_296), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_293), .B(n_221), .Y(n_328) );
NAND2x1_ASAP7_75t_L g329 ( .A(n_314), .B(n_243), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_296), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_322), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_290), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_277), .B(n_252), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_298), .B(n_221), .Y(n_334) );
A2O1A1Ixp33_ASAP7_75t_L g335 ( .A1(n_312), .A2(n_251), .B(n_254), .C(n_229), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_283), .A2(n_272), .B1(n_268), .B2(n_232), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_308), .A2(n_254), .B1(n_231), .B2(n_240), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_303), .B(n_221), .Y(n_338) );
OAI21x1_ASAP7_75t_L g339 ( .A1(n_316), .A2(n_264), .B(n_263), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_280), .A2(n_232), .B1(n_221), .B2(n_224), .Y(n_340) );
NAND2xp33_ASAP7_75t_SL g341 ( .A(n_308), .B(n_252), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_308), .B(n_243), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_295), .Y(n_343) );
INVxp67_ASAP7_75t_SL g344 ( .A(n_279), .Y(n_344) );
INVx4_ASAP7_75t_L g345 ( .A(n_277), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_295), .B(n_244), .Y(n_346) );
OAI221xp5_ASAP7_75t_L g347 ( .A1(n_280), .A2(n_217), .B1(n_236), .B2(n_239), .C(n_225), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_317), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_320), .A2(n_240), .B1(n_263), .B2(n_256), .Y(n_349) );
OAI221xp5_ASAP7_75t_L g350 ( .A1(n_276), .A2(n_217), .B1(n_225), .B2(n_269), .C(n_258), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_311), .A2(n_214), .B1(n_257), .B2(n_242), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_306), .A2(n_214), .B1(n_257), .B2(n_242), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_317), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_323), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_277), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_306), .A2(n_257), .B1(n_242), .B2(n_260), .Y(n_356) );
OR2x6_ASAP7_75t_L g357 ( .A(n_279), .B(n_257), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_306), .A2(n_213), .B1(n_260), .B2(n_246), .Y(n_358) );
INVx2_ASAP7_75t_SL g359 ( .A(n_333), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_332), .Y(n_360) );
OAI21x1_ASAP7_75t_L g361 ( .A1(n_339), .A2(n_310), .B(n_315), .Y(n_361) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_340), .A2(n_281), .B1(n_297), .B2(n_324), .C(n_246), .Y(n_362) );
INVx1_ASAP7_75t_SL g363 ( .A(n_342), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_325), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_336), .A2(n_319), .B1(n_322), .B2(n_320), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_347), .A2(n_319), .B1(n_292), .B2(n_307), .Y(n_366) );
AOI22xp33_ASAP7_75t_SL g367 ( .A1(n_349), .A2(n_319), .B1(n_277), .B2(n_299), .Y(n_367) );
AOI21xp33_ASAP7_75t_L g368 ( .A1(n_337), .A2(n_313), .B(n_282), .Y(n_368) );
OAI21x1_ASAP7_75t_L g369 ( .A1(n_339), .A2(n_323), .B(n_278), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_342), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_350), .A2(n_309), .B1(n_307), .B2(n_318), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_325), .Y(n_372) );
OR2x6_ASAP7_75t_L g373 ( .A(n_357), .B(n_279), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_353), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_332), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_343), .Y(n_376) );
AOI222xp33_ASAP7_75t_L g377 ( .A1(n_328), .A2(n_304), .B1(n_321), .B2(n_305), .C1(n_275), .C2(n_279), .Y(n_377) );
INVx2_ASAP7_75t_SL g378 ( .A(n_333), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_353), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_343), .Y(n_380) );
OAI22xp33_ASAP7_75t_L g381 ( .A1(n_327), .A2(n_299), .B1(n_304), .B2(n_286), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_334), .B(n_286), .Y(n_382) );
OAI21x1_ASAP7_75t_L g383 ( .A1(n_329), .A2(n_278), .B(n_309), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_338), .B(n_286), .Y(n_384) );
BUFx4f_ASAP7_75t_SL g385 ( .A(n_345), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_385), .Y(n_386) );
OAI221xp5_ASAP7_75t_L g387 ( .A1(n_362), .A2(n_352), .B1(n_356), .B2(n_351), .C(n_358), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_360), .B(n_348), .Y(n_388) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_363), .Y(n_389) );
BUFx2_ASAP7_75t_L g390 ( .A(n_373), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_360), .B(n_348), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_364), .Y(n_392) );
AO21x2_ASAP7_75t_L g393 ( .A1(n_369), .A2(n_282), .B(n_274), .Y(n_393) );
OAI211xp5_ASAP7_75t_SL g394 ( .A1(n_366), .A2(n_287), .B(n_335), .C(n_274), .Y(n_394) );
AO21x2_ASAP7_75t_L g395 ( .A1(n_369), .A2(n_313), .B(n_354), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_368), .A2(n_327), .B1(n_330), .B2(n_331), .C(n_275), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_375), .B(n_354), .Y(n_397) );
AOI222xp33_ASAP7_75t_L g398 ( .A1(n_365), .A2(n_330), .B1(n_331), .B2(n_288), .C1(n_355), .C2(n_346), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_375), .B(n_355), .Y(n_399) );
BUFx3_ASAP7_75t_L g400 ( .A(n_373), .Y(n_400) );
NOR3xp33_ASAP7_75t_SL g401 ( .A(n_381), .B(n_341), .C(n_326), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_377), .A2(n_357), .B1(n_288), .B2(n_301), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_364), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_364), .Y(n_404) );
OAI31xp33_ASAP7_75t_L g405 ( .A1(n_368), .A2(n_300), .A3(n_301), .B(n_333), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_376), .B(n_380), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_376), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_380), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_372), .B(n_346), .Y(n_409) );
NAND3xp33_ASAP7_75t_L g410 ( .A(n_377), .B(n_345), .C(n_76), .Y(n_410) );
AO21x2_ASAP7_75t_L g411 ( .A1(n_361), .A2(n_344), .B(n_255), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_372), .B(n_345), .Y(n_412) );
BUFx2_ASAP7_75t_L g413 ( .A(n_373), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_363), .B(n_370), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_372), .B(n_357), .Y(n_415) );
OR2x6_ASAP7_75t_L g416 ( .A(n_373), .B(n_357), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_374), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_409), .B(n_374), .Y(n_418) );
BUFx2_ASAP7_75t_SL g419 ( .A(n_386), .Y(n_419) );
INVx2_ASAP7_75t_SL g420 ( .A(n_412), .Y(n_420) );
INVx6_ASAP7_75t_L g421 ( .A(n_412), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_391), .B(n_370), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_399), .B(n_374), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_391), .B(n_379), .Y(n_424) );
INVx1_ASAP7_75t_SL g425 ( .A(n_409), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_417), .B(n_379), .Y(n_426) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_387), .A2(n_371), .B1(n_301), .B2(n_300), .C(n_384), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_392), .Y(n_428) );
INVx4_ASAP7_75t_L g429 ( .A(n_416), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_407), .Y(n_430) );
NAND3xp33_ASAP7_75t_L g431 ( .A(n_396), .B(n_367), .C(n_302), .Y(n_431) );
AND2x4_ASAP7_75t_L g432 ( .A(n_400), .B(n_379), .Y(n_432) );
AND2x4_ASAP7_75t_L g433 ( .A(n_400), .B(n_383), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_407), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_399), .B(n_373), .Y(n_435) );
AND2x4_ASAP7_75t_L g436 ( .A(n_400), .B(n_383), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_406), .B(n_382), .Y(n_437) );
OAI31xp33_ASAP7_75t_SL g438 ( .A1(n_410), .A2(n_396), .A3(n_387), .B(n_394), .Y(n_438) );
NOR3xp33_ASAP7_75t_L g439 ( .A(n_394), .B(n_378), .C(n_359), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_392), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_408), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_408), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_406), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g444 ( .A(n_410), .B(n_288), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_392), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_417), .B(n_378), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_388), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_403), .B(n_361), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_397), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_414), .B(n_288), .Y(n_450) );
NAND2x1_ASAP7_75t_L g451 ( .A(n_401), .B(n_314), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_397), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_403), .B(n_10), .Y(n_453) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_403), .Y(n_454) );
BUFx2_ASAP7_75t_L g455 ( .A(n_389), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_414), .Y(n_456) );
OAI221xp5_ASAP7_75t_L g457 ( .A1(n_405), .A2(n_270), .B1(n_302), .B2(n_285), .C(n_284), .Y(n_457) );
NAND3xp33_ASAP7_75t_L g458 ( .A(n_398), .B(n_302), .C(n_271), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_404), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_404), .Y(n_460) );
INVx3_ASAP7_75t_L g461 ( .A(n_404), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_425), .B(n_402), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_443), .B(n_390), .Y(n_463) );
INVx3_ASAP7_75t_L g464 ( .A(n_461), .Y(n_464) );
NAND3xp33_ASAP7_75t_SL g465 ( .A(n_458), .B(n_398), .C(n_405), .Y(n_465) );
AOI221x1_ASAP7_75t_L g466 ( .A1(n_439), .A2(n_415), .B1(n_300), .B2(n_411), .C(n_302), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_454), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_447), .B(n_390), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_430), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_454), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_461), .B(n_411), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_455), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_461), .B(n_411), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_434), .Y(n_474) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_420), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_441), .Y(n_476) );
INVx1_ASAP7_75t_SL g477 ( .A(n_419), .Y(n_477) );
INVx1_ASAP7_75t_SL g478 ( .A(n_421), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_442), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_418), .B(n_411), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_456), .B(n_413), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_420), .B(n_393), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_449), .B(n_415), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_452), .B(n_415), .Y(n_484) );
INVx2_ASAP7_75t_SL g485 ( .A(n_421), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_418), .B(n_415), .Y(n_486) );
OAI21xp5_ASAP7_75t_L g487 ( .A1(n_431), .A2(n_314), .B(n_416), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_448), .B(n_393), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_448), .B(n_393), .Y(n_489) );
AND2x2_ASAP7_75t_SL g490 ( .A(n_429), .B(n_416), .Y(n_490) );
NAND2xp33_ASAP7_75t_SL g491 ( .A(n_429), .B(n_395), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_459), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_453), .Y(n_493) );
INVxp67_ASAP7_75t_SL g494 ( .A(n_444), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_428), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_428), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_422), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_423), .B(n_416), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_440), .B(n_393), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_460), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_424), .B(n_416), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_437), .B(n_395), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_440), .B(n_395), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_445), .B(n_426), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_421), .B(n_395), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_445), .B(n_10), .Y(n_506) );
NAND2x1p5_ASAP7_75t_L g507 ( .A(n_444), .B(n_329), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_426), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_446), .B(n_11), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_446), .B(n_12), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_450), .B(n_14), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_433), .B(n_436), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_433), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_433), .B(n_15), .Y(n_514) );
INVxp67_ASAP7_75t_L g515 ( .A(n_432), .Y(n_515) );
AOI322xp5_ASAP7_75t_L g516 ( .A1(n_477), .A2(n_427), .A3(n_438), .B1(n_436), .B2(n_451), .C1(n_432), .C2(n_429), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_475), .B(n_432), .Y(n_517) );
OAI22xp33_ASAP7_75t_SL g518 ( .A1(n_485), .A2(n_457), .B1(n_435), .B2(n_450), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_469), .Y(n_519) );
OAI22xp33_ASAP7_75t_L g520 ( .A1(n_465), .A2(n_436), .B1(n_294), .B2(n_291), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_497), .B(n_16), .Y(n_521) );
NOR4xp25_ASAP7_75t_SL g522 ( .A(n_491), .B(n_16), .C(n_17), .D(n_314), .Y(n_522) );
OAI22xp5_ASAP7_75t_SL g523 ( .A1(n_490), .A2(n_294), .B1(n_291), .B2(n_289), .Y(n_523) );
NOR2x1_ASAP7_75t_L g524 ( .A(n_487), .B(n_247), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_490), .A2(n_249), .B(n_244), .C(n_262), .Y(n_525) );
BUFx2_ASAP7_75t_L g526 ( .A(n_485), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_474), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_478), .A2(n_249), .B1(n_262), .B2(n_261), .Y(n_528) );
AOI322xp5_ASAP7_75t_L g529 ( .A1(n_472), .A2(n_261), .A3(n_259), .B1(n_247), .B2(n_218), .C1(n_216), .C2(n_182), .Y(n_529) );
OR4x1_ASAP7_75t_L g530 ( .A(n_513), .B(n_20), .C(n_21), .D(n_24), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_476), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_514), .A2(n_314), .B1(n_259), .B2(n_266), .Y(n_532) );
NAND3xp33_ASAP7_75t_L g533 ( .A(n_466), .B(n_190), .C(n_174), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_462), .A2(n_266), .B1(n_218), .B2(n_216), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_476), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_512), .B(n_25), .Y(n_536) );
NOR2xp33_ASAP7_75t_SL g537 ( .A(n_494), .B(n_248), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_509), .B(n_32), .Y(n_538) );
OAI21xp33_ASAP7_75t_L g539 ( .A1(n_513), .A2(n_184), .B(n_189), .Y(n_539) );
AOI21xp33_ASAP7_75t_SL g540 ( .A1(n_506), .A2(n_37), .B(n_39), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_510), .A2(n_206), .B1(n_189), .B2(n_190), .Y(n_541) );
OAI22xp33_ASAP7_75t_L g542 ( .A1(n_506), .A2(n_44), .B1(n_45), .B2(n_46), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_479), .B(n_47), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_508), .B(n_51), .Y(n_544) );
INVxp67_ASAP7_75t_L g545 ( .A(n_511), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_492), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_500), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_508), .B(n_55), .Y(n_548) );
OAI21xp5_ASAP7_75t_SL g549 ( .A1(n_507), .A2(n_57), .B(n_58), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_512), .B(n_59), .Y(n_550) );
NOR2xp67_ASAP7_75t_SL g551 ( .A(n_464), .B(n_63), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_467), .Y(n_552) );
AOI22xp33_ASAP7_75t_SL g553 ( .A1(n_480), .A2(n_197), .B1(n_190), .B2(n_188), .Y(n_553) );
OAI33xp33_ASAP7_75t_L g554 ( .A1(n_502), .A2(n_64), .A3(n_66), .B1(n_67), .B2(n_68), .B3(n_72), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_501), .A2(n_73), .B1(n_167), .B2(n_174), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_501), .A2(n_197), .B1(n_174), .B2(n_188), .Y(n_556) );
AOI32xp33_ASAP7_75t_L g557 ( .A1(n_491), .A2(n_480), .A3(n_504), .B1(n_473), .B2(n_471), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_498), .A2(n_167), .B1(n_174), .B2(n_188), .Y(n_558) );
AOI21xp33_ASAP7_75t_SL g559 ( .A1(n_507), .A2(n_167), .B(n_174), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_468), .B(n_167), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_519), .Y(n_561) );
XNOR2xp5_ASAP7_75t_L g562 ( .A(n_526), .B(n_486), .Y(n_562) );
INVxp67_ASAP7_75t_L g563 ( .A(n_552), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_527), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_531), .Y(n_565) );
INVx3_ASAP7_75t_L g566 ( .A(n_517), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_535), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_537), .B(n_470), .Y(n_568) );
NOR3xp33_ASAP7_75t_SL g569 ( .A(n_520), .B(n_505), .C(n_484), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_537), .B(n_470), .Y(n_570) );
OAI22xp33_ASAP7_75t_L g571 ( .A1(n_549), .A2(n_515), .B1(n_507), .B2(n_481), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g572 ( .A(n_545), .Y(n_572) );
INVxp67_ASAP7_75t_L g573 ( .A(n_521), .Y(n_573) );
NOR2xp33_ASAP7_75t_SL g574 ( .A(n_549), .B(n_467), .Y(n_574) );
NAND4xp75_ASAP7_75t_L g575 ( .A(n_524), .B(n_489), .C(n_488), .D(n_483), .Y(n_575) );
OAI321xp33_ASAP7_75t_L g576 ( .A1(n_557), .A2(n_482), .A3(n_463), .B1(n_488), .B2(n_489), .C(n_493), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_518), .B(n_482), .Y(n_577) );
INVx2_ASAP7_75t_SL g578 ( .A(n_550), .Y(n_578) );
INVxp33_ASAP7_75t_L g579 ( .A(n_523), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_546), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_547), .B(n_471), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_536), .B(n_499), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_560), .Y(n_583) );
NOR3xp33_ASAP7_75t_SL g584 ( .A(n_554), .B(n_464), .C(n_503), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_543), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_516), .B(n_495), .Y(n_586) );
INVx1_ASAP7_75t_SL g587 ( .A(n_550), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_544), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_529), .B(n_496), .Y(n_589) );
AOI222xp33_ASAP7_75t_L g590 ( .A1(n_538), .A2(n_188), .B1(n_190), .B2(n_197), .C1(n_496), .C2(n_533), .Y(n_590) );
INVx1_ASAP7_75t_SL g591 ( .A(n_572), .Y(n_591) );
AND3x4_ASAP7_75t_L g592 ( .A(n_584), .B(n_569), .C(n_579), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_577), .A2(n_542), .B1(n_555), .B2(n_532), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_565), .Y(n_594) );
INVx1_ASAP7_75t_SL g595 ( .A(n_572), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_577), .B(n_548), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_561), .Y(n_597) );
AOI221x1_ASAP7_75t_L g598 ( .A1(n_586), .A2(n_540), .B1(n_539), .B2(n_556), .C(n_559), .Y(n_598) );
AOI211xp5_ASAP7_75t_SL g599 ( .A1(n_574), .A2(n_528), .B(n_525), .C(n_530), .Y(n_599) );
OAI21xp33_ASAP7_75t_L g600 ( .A1(n_579), .A2(n_553), .B(n_541), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_587), .Y(n_601) );
OAI32xp33_ASAP7_75t_L g602 ( .A1(n_566), .A2(n_522), .A3(n_551), .B1(n_558), .B2(n_534), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_564), .Y(n_603) );
INVxp67_ASAP7_75t_SL g604 ( .A(n_563), .Y(n_604) );
OAI21xp5_ASAP7_75t_SL g605 ( .A1(n_571), .A2(n_522), .B(n_190), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_573), .A2(n_188), .B1(n_197), .B2(n_585), .Y(n_606) );
XNOR2xp5_ASAP7_75t_L g607 ( .A(n_562), .B(n_197), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_567), .Y(n_608) );
NOR3x1_ASAP7_75t_L g609 ( .A(n_578), .B(n_575), .C(n_568), .Y(n_609) );
NOR3xp33_ASAP7_75t_L g610 ( .A(n_602), .B(n_576), .C(n_570), .Y(n_610) );
NOR2xp33_ASAP7_75t_R g611 ( .A(n_591), .B(n_588), .Y(n_611) );
OAI21xp5_ASAP7_75t_SL g612 ( .A1(n_599), .A2(n_590), .B(n_589), .Y(n_612) );
INVx1_ASAP7_75t_SL g613 ( .A(n_595), .Y(n_613) );
CKINVDCx16_ASAP7_75t_R g614 ( .A(n_601), .Y(n_614) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_604), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_592), .B(n_580), .Y(n_616) );
CKINVDCx14_ASAP7_75t_R g617 ( .A(n_607), .Y(n_617) );
AO22x2_ASAP7_75t_L g618 ( .A1(n_598), .A2(n_583), .B1(n_581), .B2(n_582), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_593), .A2(n_582), .B1(n_605), .B2(n_597), .Y(n_619) );
OAI22x1_ASAP7_75t_L g620 ( .A1(n_609), .A2(n_603), .B1(n_608), .B2(n_594), .Y(n_620) );
NAND4xp25_ASAP7_75t_L g621 ( .A(n_606), .B(n_599), .C(n_609), .D(n_598), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_592), .A2(n_577), .B1(n_596), .B2(n_600), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_604), .Y(n_623) );
AOI32xp33_ASAP7_75t_L g624 ( .A1(n_599), .A2(n_579), .A3(n_574), .B1(n_571), .B2(n_477), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_614), .Y(n_625) );
INVx1_ASAP7_75t_SL g626 ( .A(n_613), .Y(n_626) );
INVxp67_ASAP7_75t_SL g627 ( .A(n_615), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_623), .Y(n_628) );
BUFx4f_ASAP7_75t_SL g629 ( .A(n_613), .Y(n_629) );
XOR2xp5_ASAP7_75t_L g630 ( .A(n_625), .B(n_617), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_627), .Y(n_631) );
OAI211xp5_ASAP7_75t_SL g632 ( .A1(n_626), .A2(n_624), .B(n_622), .C(n_612), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_630), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_631), .Y(n_634) );
OAI221xp5_ASAP7_75t_L g635 ( .A1(n_633), .A2(n_632), .B1(n_621), .B2(n_610), .C(n_619), .Y(n_635) );
INVxp67_ASAP7_75t_SL g636 ( .A(n_634), .Y(n_636) );
AOI222xp33_ASAP7_75t_L g637 ( .A1(n_635), .A2(n_629), .B1(n_628), .B2(n_620), .C1(n_618), .C2(n_616), .Y(n_637) );
AO21x2_ASAP7_75t_L g638 ( .A1(n_637), .A2(n_636), .B(n_611), .Y(n_638) );
endmodule