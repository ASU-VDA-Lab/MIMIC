module fake_jpeg_16799_n_249 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_21),
.Y(n_35)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_32),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_37),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx4f_ASAP7_75t_SL g38 ( 
.A(n_19),
.Y(n_38)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_0),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_30),
.B1(n_27),
.B2(n_24),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_40),
.B1(n_23),
.B2(n_32),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_27),
.B1(n_24),
.B2(n_30),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_53),
.B1(n_17),
.B2(n_23),
.Y(n_72)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_52),
.Y(n_60)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_26),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_51),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_26),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_27),
.B1(n_24),
.B2(n_30),
.Y(n_53)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_68),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_31),
.B1(n_35),
.B2(n_36),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_59),
.A2(n_61),
.B1(n_83),
.B2(n_31),
.Y(n_92)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_43),
.B(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_64),
.B(n_21),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_66),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_37),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_22),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_22),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_75),
.Y(n_88)
);

CKINVDCx9p33_ASAP7_75t_R g70 ( 
.A(n_49),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_70),
.Y(n_87)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_72),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_16),
.B1(n_28),
.B2(n_20),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_73),
.A2(n_79),
.B1(n_84),
.B2(n_52),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_33),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_46),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_80),
.Y(n_95)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_78),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_42),
.A2(n_16),
.B1(n_28),
.B2(n_20),
.Y(n_79)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_41),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_82),
.Y(n_100)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_31),
.B1(n_20),
.B2(n_18),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_47),
.A2(n_52),
.B1(n_41),
.B2(n_29),
.Y(n_84)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_97),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_92),
.B(n_94),
.Y(n_129)
);

AND2x6_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_1),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_96),
.B(n_21),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_98),
.A2(n_109),
.B1(n_58),
.B2(n_29),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_67),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_57),
.B(n_83),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_106),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_25),
.B(n_18),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_62),
.B(n_33),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_101),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_21),
.Y(n_108)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_108),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_75),
.B1(n_62),
.B2(n_61),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_113),
.A2(n_117),
.B(n_133),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_115),
.B(n_118),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_101),
.A2(n_71),
.B1(n_82),
.B2(n_58),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_116),
.A2(n_124),
.B1(n_132),
.B2(n_102),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_119),
.B(n_121),
.Y(n_161)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_81),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_135),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_38),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_78),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_109),
.A2(n_65),
.B1(n_80),
.B2(n_38),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_85),
.B(n_15),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_127),
.B(n_15),
.Y(n_162)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_130),
.A2(n_89),
.B1(n_86),
.B2(n_18),
.Y(n_160)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_95),
.A2(n_38),
.B1(n_78),
.B2(n_66),
.Y(n_132)
);

AO21x1_ASAP7_75t_L g133 ( 
.A1(n_88),
.A2(n_96),
.B(n_92),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_134),
.A2(n_136),
.B(n_87),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_90),
.B(n_33),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_94),
.A2(n_21),
.B(n_26),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_128),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_137),
.B(n_139),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_98),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_138),
.B(n_140),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_97),
.Y(n_139)
);

AOI21xp33_ASAP7_75t_SL g140 ( 
.A1(n_123),
.A2(n_104),
.B(n_33),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_120),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_141),
.B(n_155),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_129),
.A2(n_122),
.B(n_132),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_154),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_162),
.Y(n_170)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_33),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_152),
.C(n_158),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_124),
.A2(n_114),
.B(n_115),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_126),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_156),
.B(n_157),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_112),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_113),
.A2(n_104),
.B(n_102),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_136),
.A2(n_89),
.B(n_106),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_26),
.C(n_19),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_160),
.A2(n_99),
.B1(n_29),
.B2(n_25),
.Y(n_180)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_118),
.B1(n_133),
.B2(n_134),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_177),
.C(n_158),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_125),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_171),
.B(n_181),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_147),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_178),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_99),
.C(n_26),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_180),
.B(n_139),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_99),
.Y(n_181)
);

OAI32xp33_ASAP7_75t_L g182 ( 
.A1(n_150),
.A2(n_25),
.A3(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_183),
.Y(n_199)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

XOR2x1_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_150),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_184),
.A2(n_154),
.B(n_182),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_190),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_142),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_138),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_191),
.B(n_196),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_192),
.A2(n_189),
.B1(n_166),
.B2(n_172),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_151),
.C(n_153),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_195),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_177),
.C(n_175),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_153),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_170),
.C(n_167),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_148),
.Y(n_206)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_207),
.Y(n_214)
);

BUFx12_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_205),
.Y(n_213)
);

BUFx24_ASAP7_75t_SL g205 ( 
.A(n_196),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_201),
.C(n_211),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_168),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_198),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_188),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_190),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_211),
.B(n_199),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_193),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_211),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_208),
.A2(n_173),
.B1(n_147),
.B2(n_148),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_215),
.A2(n_160),
.B1(n_159),
.B2(n_155),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_216),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_218),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_173),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_221),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_5),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_191),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_180),
.C(n_13),
.Y(n_228)
);

AOI21x1_ASAP7_75t_L g224 ( 
.A1(n_216),
.A2(n_204),
.B(n_189),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_224),
.A2(n_215),
.B(n_214),
.Y(n_232)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_225),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_230),
.C(n_231),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_1),
.C(n_2),
.Y(n_230)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_232),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_226),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_234),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_213),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_R g237 ( 
.A(n_230),
.B(n_223),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_237),
.A2(n_229),
.B(n_7),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_235),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_8),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_241),
.A2(n_6),
.B(n_7),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_236),
.C(n_7),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_243),
.Y(n_245)
);

AO21x1_ASAP7_75t_L g246 ( 
.A1(n_244),
.A2(n_239),
.B(n_9),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_246),
.Y(n_247)
);

AOI321xp33_ASAP7_75t_L g248 ( 
.A1(n_247),
.A2(n_8),
.A3(n_9),
.B1(n_11),
.B2(n_245),
.C(n_241),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_11),
.Y(n_249)
);


endmodule