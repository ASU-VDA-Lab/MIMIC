module fake_jpeg_10383_n_83 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_83);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_83;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_32),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_59)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_45),
.Y(n_54)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_0),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_7),
.Y(n_55)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_36),
.B(n_2),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_51),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_67)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_9),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_55),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_8),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_60),
.C(n_61),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_58),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_67),
.B1(n_30),
.B2(n_31),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_13),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_15),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_47),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_64),
.B(n_66),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_44),
.B(n_16),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_68),
.B1(n_64),
.B2(n_66),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_20),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_44),
.B(n_27),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_73),
.C(n_54),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_75),
.B(n_71),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_72),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_53),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_79),
.B(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_81),
.A2(n_74),
.B1(n_62),
.B2(n_70),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_56),
.Y(n_83)
);


endmodule