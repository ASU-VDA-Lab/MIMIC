module real_jpeg_9441_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_340, n_7, n_341, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_340;
input n_7;
input n_341;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_1),
.A2(n_68),
.B1(n_69),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_1),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_1),
.A2(n_48),
.B1(n_50),
.B2(n_98),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_98),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_1),
.A2(n_23),
.B1(n_25),
.B2(n_98),
.Y(n_239)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_3),
.A2(n_50),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_3),
.B(n_50),
.Y(n_103)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_3),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_3),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_3),
.B(n_26),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_L g191 ( 
.A1(n_3),
.A2(n_28),
.B(n_30),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_3),
.A2(n_23),
.B1(n_25),
.B2(n_114),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_4),
.A2(n_68),
.B1(n_69),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_4),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_4),
.A2(n_48),
.B1(n_50),
.B2(n_93),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_93),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_4),
.A2(n_23),
.B1(n_25),
.B2(n_93),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g95 ( 
.A(n_5),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_7),
.A2(n_23),
.B1(n_25),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_7),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_7),
.A2(n_60),
.B1(n_68),
.B2(n_69),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_7),
.A2(n_48),
.B1(n_50),
.B2(n_60),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_60),
.Y(n_266)
);

BUFx6f_ASAP7_75t_SL g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_11),
.A2(n_23),
.B1(n_25),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_11),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_11),
.A2(n_62),
.B1(n_68),
.B2(n_69),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_11),
.A2(n_48),
.B1(n_50),
.B2(n_62),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_62),
.Y(n_290)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_13),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_13),
.A2(n_24),
.B1(n_29),
.B2(n_30),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_13),
.A2(n_24),
.B1(n_48),
.B2(n_50),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_13),
.A2(n_24),
.B1(n_68),
.B2(n_69),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_14),
.A2(n_48),
.B1(n_50),
.B2(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_14),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_14),
.A2(n_68),
.B1(n_69),
.B2(n_105),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_105),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_14),
.A2(n_23),
.B1(n_25),
.B2(n_105),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_15),
.A2(n_23),
.B1(n_25),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_15),
.A2(n_34),
.B1(n_68),
.B2(n_69),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_15),
.A2(n_34),
.B1(n_48),
.B2(n_50),
.Y(n_204)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.C(n_338),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_80),
.B(n_336),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_38),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_20),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_32),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_21),
.A2(n_36),
.B(n_239),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_26),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_22),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_22),
.A2(n_26),
.B(n_35),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_23),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_23),
.A2(n_27),
.B(n_31),
.C(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_31),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_23),
.A2(n_31),
.B(n_114),
.C(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_26),
.B(n_33),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_26),
.A2(n_35),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_27),
.A2(n_36),
.B1(n_59),
.B2(n_61),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_27),
.A2(n_36),
.B1(n_211),
.B2(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_27),
.A2(n_36),
.B1(n_220),
.B2(n_239),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_27),
.A2(n_32),
.B(n_59),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_27)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

O2A1O1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_30),
.A2(n_45),
.B(n_46),
.C(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_46),
.Y(n_54)
);

HAxp5_ASAP7_75t_SL g144 ( 
.A(n_30),
.B(n_114),
.CON(n_144),
.SN(n_144)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_35),
.A2(n_75),
.B(n_76),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_36),
.A2(n_77),
.B(n_284),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_39),
.B(n_337),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_74),
.C(n_78),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_40),
.A2(n_41),
.B1(n_332),
.B2(n_334),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_57),
.C(n_63),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_42),
.A2(n_43),
.B1(n_63),
.B2(n_311),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_52),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_44),
.A2(n_163),
.B(n_207),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_51),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_51),
.B(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_45),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_45),
.A2(n_53),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_45),
.A2(n_53),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_46),
.B(n_50),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_48),
.A2(n_54),
.B1(n_144),
.B2(n_150),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_65),
.B(n_66),
.C(n_67),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_65),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_51),
.A2(n_53),
.B(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_52),
.A2(n_130),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_53),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_56),
.B(n_130),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_57),
.A2(n_58),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_63),
.A2(n_308),
.B1(n_311),
.B2(n_312),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_63),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_67),
.B(n_72),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_64),
.A2(n_67),
.B1(n_102),
.B2(n_104),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_64),
.A2(n_67),
.B1(n_104),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_64),
.A2(n_67),
.B1(n_132),
.B2(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_64),
.A2(n_142),
.B(n_179),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_64),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_64),
.A2(n_67),
.B1(n_226),
.B2(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_64),
.A2(n_246),
.B(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_65),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_65),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_67),
.B(n_114),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_67),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_67),
.B(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_67),
.A2(n_226),
.B(n_227),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_68),
.B(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_68),
.B(n_71),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_68),
.B(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_69),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_106)
);

BUFx24_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_73),
.B(n_180),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_73),
.A2(n_202),
.B(n_203),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_74),
.A2(n_78),
.B1(n_79),
.B2(n_333),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_74),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_329),
.B(n_335),
.Y(n_80)
);

OAI321xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_301),
.A3(n_322),
.B1(n_327),
.B2(n_328),
.C(n_340),
.Y(n_81)
);

AOI321xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_254),
.A3(n_276),
.B1(n_294),
.B2(n_300),
.C(n_341),
.Y(n_82)
);

NOR3xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_213),
.C(n_250),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_184),
.B(n_212),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_157),
.B(n_183),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_137),
.B(n_156),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_125),
.B(n_136),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_111),
.B(n_124),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_99),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_90),
.B(n_99),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_94),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_94),
.B(n_154),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_95),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_95),
.B(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_97),
.A2(n_117),
.B(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_106),
.B2(n_110),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_100),
.B(n_110),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_103),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_106),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_119),
.B(n_123),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_113),
.B(n_115),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_118),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_117),
.A2(n_152),
.B(n_153),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_117),
.A2(n_118),
.B1(n_169),
.B2(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_117),
.A2(n_153),
.B(n_194),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_117),
.A2(n_118),
.B(n_152),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_118),
.A2(n_169),
.B(n_170),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_126),
.B(n_127),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_128),
.B(n_138),
.Y(n_156)
);

FAx1_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_131),
.CI(n_133),
.CON(n_128),
.SN(n_128)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_130),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_130),
.A2(n_163),
.B1(n_165),
.B2(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_134),
.B(n_170),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_135),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_148),
.B2(n_155),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_143),
.B1(n_146),
.B2(n_147),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_141),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_143),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_147),
.C(n_155),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_145),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_148),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_151),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_158),
.B(n_159),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_175),
.B2(n_176),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_178),
.C(n_181),
.Y(n_185)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_166),
.B1(n_167),
.B2(n_174),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_162),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_163),
.A2(n_309),
.B(n_310),
.Y(n_308)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_168),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_171),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_172),
.C(n_174),
.Y(n_195)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_181),
.B2(n_182),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_177),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_178),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_179),
.B(n_227),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_185),
.B(n_186),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_198),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_188),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_188),
.B(n_197),
.C(n_198),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_193),
.Y(n_216)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_195),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_208),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_205),
.B2(n_206),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_205),
.C(n_208),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_228),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_203),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_213),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_232),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_214),
.B(n_232),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_223),
.C(n_230),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_215),
.B(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_218),
.C(n_222),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_222),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_221),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_223),
.A2(n_224),
.B1(n_230),
.B2(n_231),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_229),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_229),
.Y(n_235)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.Y(n_232)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_233),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_243),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_243),
.C(n_247),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_235),
.B(n_237),
.C(n_241),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_240),
.B2(n_241),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_242),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_245),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_251),
.B(n_252),
.Y(n_297)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_255),
.A2(n_295),
.B(n_299),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_256),
.B(n_257),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_275),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_268),
.B2(n_269),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_269),
.C(n_275),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_261),
.B(n_263),
.C(n_267),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_265),
.B2(n_267),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_265),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_266),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_274),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_270),
.A2(n_271),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_270),
.A2(n_283),
.B(n_286),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_272),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_272),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_277),
.B(n_278),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_278),
.Y(n_323)
);

FAx1_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_287),
.CI(n_293),
.CON(n_278),
.SN(n_278)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_285),
.B2(n_286),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_285),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_291),
.B(n_292),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_291),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_290),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_292),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_292),
.A2(n_303),
.B1(n_313),
.B2(n_326),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B(n_298),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_315),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_302),
.B(n_315),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_313),
.C(n_314),
.Y(n_302)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_303),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_304),
.A2(n_305),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_305),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_311),
.C(n_312),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_305),
.B(n_317),
.C(n_321),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_308),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_325),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_321),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_323),
.B(n_324),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_331),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_332),
.Y(n_334)
);


endmodule