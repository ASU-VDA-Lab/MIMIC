module fake_jpeg_7182_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx8_ASAP7_75t_SL g8 ( 
.A(n_3),
.Y(n_8)
);

INVxp67_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx6_ASAP7_75t_SL g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_2),
.B(n_6),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_19),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_13),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_11),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_32),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_18),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_16),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

O2A1O1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_25),
.B(n_10),
.C(n_9),
.Y(n_35)
);

AO21x1_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_39),
.B(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_40),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_9),
.B(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

OAI21xp33_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_28),
.B(n_15),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_18),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_26),
.C(n_19),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_27),
.C(n_12),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_45),
.A2(n_26),
.B1(n_28),
.B2(n_25),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_46),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_48),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_49),
.A2(n_41),
.B(n_43),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_49),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_50),
.A2(n_49),
.B(n_51),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_51),
.B1(n_26),
.B2(n_20),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_54),
.B(n_27),
.Y(n_56)
);

INVxp33_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_56),
.C(n_7),
.Y(n_58)
);

AOI221xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_7),
.B1(n_1),
.B2(n_0),
.C(n_12),
.Y(n_59)
);


endmodule