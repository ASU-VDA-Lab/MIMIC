module real_jpeg_27159_n_3 (n_1, n_0, n_2, n_3);

input n_1;
input n_0;
input n_2;

output n_3;

wire n_5;
wire n_8;
wire n_4;
wire n_6;
wire n_7;
wire n_10;
wire n_9;

HAxp5_ASAP7_75t_SL g7 ( 
.A(n_0),
.B(n_8),
.CON(n_7),
.SN(n_7)
);

NAND2xp5_ASAP7_75t_L g4 ( 
.A(n_1),
.B(n_5),
.Y(n_4)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_2),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g3 ( 
.A(n_4),
.B(n_9),
.Y(n_3)
);

CKINVDCx20_ASAP7_75t_R g5 ( 
.A(n_6),
.Y(n_5)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_6),
.B(n_10),
.Y(n_9)
);

CKINVDCx5p33_ASAP7_75t_R g6 ( 
.A(n_7),
.Y(n_6)
);

BUFx24_ASAP7_75t_SL g11 ( 
.A(n_7),
.Y(n_11)
);


endmodule