module fake_jpeg_1872_n_445 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_445);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_445;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_3),
.B(n_4),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_55),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_58),
.B(n_60),
.Y(n_120)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_59),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_23),
.B(n_9),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_63),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_64),
.Y(n_168)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_66),
.Y(n_158)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_68),
.Y(n_170)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_21),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_71),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_23),
.B(n_9),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_72),
.B(n_78),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_73),
.Y(n_171)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_74),
.Y(n_173)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_75),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

NOR3xp33_ASAP7_75t_L g77 ( 
.A(n_34),
.B(n_11),
.C(n_16),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_82),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_27),
.B(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_80),
.Y(n_174)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_81),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_21),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_27),
.B(n_11),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_83),
.B(n_84),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_28),
.B(n_16),
.Y(n_84)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_31),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_86),
.B(n_91),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_28),
.B(n_17),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_88),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_89),
.Y(n_184)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_29),
.B(n_15),
.Y(n_91)
);

BUFx16f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

BUFx12_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g121 ( 
.A(n_95),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_96),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_41),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_97),
.B(n_98),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_41),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_32),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_99),
.B(n_105),
.Y(n_136)
);

BUFx12_ASAP7_75t_L g100 ( 
.A(n_37),
.Y(n_100)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_101),
.Y(n_160)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_54),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_25),
.Y(n_106)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_19),
.Y(n_107)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_107),
.Y(n_159)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_19),
.Y(n_108)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_108),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_37),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_112),
.Y(n_119)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_43),
.Y(n_110)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_110),
.Y(n_176)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_18),
.Y(n_111)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_111),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g114 ( 
.A1(n_63),
.A2(n_53),
.B1(n_39),
.B2(n_38),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_114),
.A2(n_115),
.B1(n_124),
.B2(n_126),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_36),
.B1(n_18),
.B2(n_38),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_92),
.A2(n_106),
.B1(n_90),
.B2(n_55),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_89),
.A2(n_36),
.B1(n_50),
.B2(n_48),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_92),
.A2(n_20),
.B1(n_50),
.B2(n_48),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_128),
.A2(n_131),
.B1(n_132),
.B2(n_140),
.Y(n_235)
);

AOI21xp33_ASAP7_75t_L g130 ( 
.A1(n_74),
.A2(n_46),
.B(n_42),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_130),
.B(n_181),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_55),
.A2(n_46),
.B1(n_42),
.B2(n_53),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_56),
.A2(n_39),
.B1(n_34),
.B2(n_3),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_65),
.A2(n_37),
.B1(n_1),
.B2(n_3),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_59),
.A2(n_37),
.B1(n_3),
.B2(n_5),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_144),
.A2(n_149),
.B1(n_175),
.B2(n_178),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_62),
.A2(n_0),
.B1(n_5),
.B2(n_6),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_145),
.A2(n_165),
.B1(n_167),
.B2(n_169),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_71),
.A2(n_0),
.B1(n_6),
.B2(n_7),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_64),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_151),
.A2(n_146),
.B1(n_127),
.B2(n_141),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_73),
.A2(n_7),
.B1(n_13),
.B2(n_66),
.Y(n_157)
);

AO22x1_ASAP7_75t_L g196 ( 
.A1(n_157),
.A2(n_162),
.B1(n_119),
.B2(n_148),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_111),
.A2(n_112),
.B1(n_95),
.B2(n_103),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_107),
.A2(n_75),
.B1(n_96),
.B2(n_101),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_93),
.A2(n_104),
.B1(n_85),
.B2(n_108),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_102),
.A2(n_76),
.B1(n_74),
.B2(n_94),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_80),
.A2(n_109),
.B1(n_94),
.B2(n_100),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_109),
.A2(n_100),
.B1(n_92),
.B2(n_70),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_87),
.A2(n_70),
.B1(n_82),
.B2(n_35),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_L g210 ( 
.A1(n_180),
.A2(n_124),
.B1(n_184),
.B2(n_177),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_58),
.B(n_78),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_78),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_182),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_92),
.A2(n_70),
.B1(n_82),
.B2(n_19),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_183),
.A2(n_113),
.B1(n_147),
.B2(n_153),
.Y(n_220)
);

NAND2xp33_ASAP7_75t_SL g185 ( 
.A(n_119),
.B(n_142),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_185),
.B(n_225),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_136),
.B(n_138),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_188),
.B(n_195),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_143),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_189),
.B(n_193),
.Y(n_263)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_190),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_191),
.A2(n_220),
.B1(n_226),
.B2(n_238),
.Y(n_254)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_125),
.Y(n_192)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_192),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_173),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_134),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_194),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_120),
.B(n_172),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_196),
.A2(n_210),
.B1(n_204),
.B2(n_197),
.Y(n_284)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_148),
.Y(n_197)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_197),
.Y(n_267)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_134),
.Y(n_198)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_198),
.Y(n_257)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_155),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_199),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_154),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_200),
.B(n_201),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_117),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_139),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_202),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_133),
.B(n_163),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_203),
.B(n_204),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_155),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_118),
.B(n_122),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_205),
.B(n_214),
.Y(n_273)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_207),
.Y(n_258)
);

AND2x2_ASAP7_75t_SL g208 ( 
.A(n_176),
.B(n_129),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_208),
.B(n_224),
.C(n_203),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_131),
.A2(n_128),
.B(n_132),
.C(n_183),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_209),
.A2(n_244),
.B(n_227),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_173),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_211),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_212),
.Y(n_278)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_135),
.Y(n_213)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_213),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_154),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_156),
.Y(n_215)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_215),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_147),
.B(n_152),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_216),
.B(n_221),
.Y(n_283)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_217),
.Y(n_271)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_218),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_123),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_219),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_175),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_121),
.Y(n_222)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_222),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g224 ( 
.A(n_129),
.B(n_174),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_121),
.B(n_150),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_113),
.A2(n_158),
.B1(n_160),
.B2(n_164),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_152),
.B(n_160),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_227),
.B(n_233),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_153),
.B(n_158),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_229),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_161),
.B(n_166),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_239),
.Y(n_245)
);

OR2x4_ASAP7_75t_L g231 ( 
.A(n_145),
.B(n_178),
.Y(n_231)
);

NAND2xp67_ASAP7_75t_SL g286 ( 
.A(n_231),
.B(n_243),
.Y(n_286)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_166),
.Y(n_232)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_232),
.Y(n_289)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_123),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_137),
.B(n_171),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_234),
.Y(n_256)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_137),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_236),
.Y(n_266)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_168),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_237),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_116),
.A2(n_165),
.B1(n_144),
.B2(n_149),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_159),
.B(n_168),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_171),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_240),
.Y(n_277)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_140),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_241),
.B(n_242),
.Y(n_288)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_116),
.Y(n_242)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_134),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_179),
.Y(n_244)
);

AOI32xp33_ASAP7_75t_L g250 ( 
.A1(n_223),
.A2(n_185),
.A3(n_231),
.B1(n_221),
.B2(n_208),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_250),
.B(n_252),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_252),
.B(n_275),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_208),
.B(n_224),
.C(n_192),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_261),
.B(n_264),
.C(n_199),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_210),
.B(n_196),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_262),
.B(n_275),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_224),
.B(n_227),
.C(n_203),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_228),
.A2(n_235),
.B1(n_187),
.B2(n_206),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_269),
.A2(n_270),
.B1(n_274),
.B2(n_280),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_209),
.A2(n_233),
.B1(n_240),
.B2(n_207),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_217),
.A2(n_236),
.B1(n_232),
.B2(n_212),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_219),
.A2(n_244),
.B1(n_190),
.B2(n_218),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_284),
.A2(n_260),
.B1(n_285),
.B2(n_288),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_245),
.B(n_186),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_290),
.B(n_298),
.Y(n_324)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_291),
.Y(n_325)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_292),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_265),
.B(n_186),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_293),
.B(n_296),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_295),
.B(n_302),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_265),
.B(n_194),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_253),
.Y(n_297)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_297),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_245),
.B(n_242),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_271),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_284),
.A2(n_211),
.B1(n_243),
.B2(n_198),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_300),
.A2(n_315),
.B1(n_307),
.B2(n_292),
.Y(n_332)
);

NOR2x1_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_249),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_301),
.B(n_308),
.Y(n_343)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_258),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_303),
.B(n_305),
.Y(n_345)
);

OAI21xp33_ASAP7_75t_SL g338 ( 
.A1(n_304),
.A2(n_246),
.B(n_247),
.Y(n_338)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_257),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_282),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_307),
.B(n_309),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_255),
.B(n_263),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_255),
.B(n_256),
.Y(n_309)
);

O2A1O1Ixp33_ASAP7_75t_L g310 ( 
.A1(n_286),
.A2(n_288),
.B(n_262),
.C(n_254),
.Y(n_310)
);

O2A1O1Ixp33_ASAP7_75t_L g333 ( 
.A1(n_310),
.A2(n_279),
.B(n_289),
.C(n_251),
.Y(n_333)
);

NAND2x1p5_ASAP7_75t_L g311 ( 
.A(n_264),
.B(n_261),
.Y(n_311)
);

OA21x2_ASAP7_75t_L g323 ( 
.A1(n_311),
.A2(n_279),
.B(n_267),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_256),
.B(n_273),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_313),
.Y(n_326)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_271),
.Y(n_313)
);

INVx6_ASAP7_75t_L g314 ( 
.A(n_266),
.Y(n_314)
);

INVx11_ASAP7_75t_L g328 ( 
.A(n_314),
.Y(n_328)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_248),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_286),
.B(n_276),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_319),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_285),
.A2(n_260),
.B1(n_266),
.B2(n_276),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_318),
.A2(n_277),
.B1(n_278),
.B2(n_287),
.Y(n_340)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_281),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_260),
.A2(n_268),
.B(n_259),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_320),
.A2(n_291),
.B(n_301),
.Y(n_347)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_259),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_321),
.B(n_322),
.Y(n_335)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_268),
.Y(n_322)
);

XNOR2x1_ASAP7_75t_L g350 ( 
.A(n_323),
.B(n_347),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_332),
.B(n_334),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_333),
.Y(n_365)
);

OA21x2_ASAP7_75t_L g334 ( 
.A1(n_317),
.A2(n_289),
.B(n_267),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_310),
.A2(n_287),
.B1(n_278),
.B2(n_246),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_336),
.A2(n_344),
.B1(n_346),
.B2(n_320),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_338),
.B(n_302),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_295),
.B(n_247),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_294),
.C(n_311),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_340),
.A2(n_323),
.B1(n_334),
.B2(n_329),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_298),
.B(n_277),
.Y(n_341)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_341),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_306),
.A2(n_248),
.B1(n_257),
.B2(n_272),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_315),
.A2(n_248),
.B1(n_318),
.B2(n_290),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_343),
.B(n_312),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_348),
.B(n_359),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_327),
.B(n_294),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_349),
.B(n_351),
.C(n_358),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_327),
.B(n_294),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_353),
.A2(n_323),
.B1(n_330),
.B2(n_332),
.Y(n_378)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_342),
.Y(n_354)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_354),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_355),
.A2(n_337),
.B(n_326),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_346),
.Y(n_356)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_356),
.Y(n_383)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_328),
.Y(n_357)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_357),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_331),
.B(n_319),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_345),
.Y(n_360)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_360),
.Y(n_381)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_342),
.Y(n_361)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_361),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_344),
.A2(n_314),
.B1(n_322),
.B2(n_313),
.Y(n_362)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_362),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_339),
.B(n_311),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_363),
.B(n_366),
.C(n_323),
.Y(n_375)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_335),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_364),
.B(n_369),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_347),
.B(n_324),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_368),
.A2(n_330),
.B1(n_325),
.B2(n_326),
.Y(n_384)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_335),
.Y(n_369)
);

OA22x2_ASAP7_75t_L g370 ( 
.A1(n_336),
.A2(n_300),
.B1(n_299),
.B2(n_316),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_370),
.B(n_340),
.Y(n_374)
);

BUFx24_ASAP7_75t_SL g372 ( 
.A(n_366),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_372),
.Y(n_399)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_374),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_375),
.B(n_380),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_378),
.A2(n_374),
.B1(n_365),
.B2(n_367),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_349),
.B(n_329),
.C(n_325),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_379),
.B(n_350),
.C(n_363),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_384),
.Y(n_402)
);

XOR2x1_ASAP7_75t_L g385 ( 
.A(n_350),
.B(n_324),
.Y(n_385)
);

HAxp5_ASAP7_75t_SL g398 ( 
.A(n_385),
.B(n_358),
.CON(n_398),
.SN(n_398)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_365),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_387),
.B(n_388),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_368),
.A2(n_341),
.B1(n_337),
.B2(n_331),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_384),
.Y(n_390)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_390),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_388),
.B(n_352),
.Y(n_393)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_393),
.Y(n_407)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_376),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_394),
.A2(n_395),
.B1(n_396),
.B2(n_400),
.Y(n_411)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_376),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_371),
.B(n_367),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_397),
.Y(n_409)
);

HAxp5_ASAP7_75t_SL g412 ( 
.A(n_398),
.B(n_373),
.CON(n_412),
.SN(n_412)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_382),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_401),
.B(n_373),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_392),
.A2(n_367),
.B(n_380),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_405),
.A2(n_397),
.B(n_378),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_393),
.A2(n_381),
.B(n_392),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_406),
.B(n_414),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_408),
.B(n_413),
.Y(n_423)
);

A2O1A1Ixp33_ASAP7_75t_SL g410 ( 
.A1(n_403),
.A2(n_387),
.B(n_385),
.C(n_375),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_410),
.A2(n_412),
.B1(n_409),
.B2(n_402),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_395),
.A2(n_403),
.B1(n_402),
.B2(n_390),
.Y(n_413)
);

BUFx12_ASAP7_75t_L g414 ( 
.A(n_401),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_411),
.Y(n_415)
);

OR2x2_ASAP7_75t_L g424 ( 
.A(n_415),
.B(n_416),
.Y(n_424)
);

OAI211xp5_ASAP7_75t_L g425 ( 
.A1(n_417),
.A2(n_419),
.B(n_413),
.C(n_371),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_408),
.B(n_391),
.C(n_379),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_418),
.B(n_422),
.C(n_381),
.Y(n_426)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_407),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_404),
.B(n_389),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_421),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_405),
.B(n_391),
.C(n_351),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_425),
.B(n_426),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_420),
.A2(n_386),
.B1(n_383),
.B2(n_410),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_427),
.A2(n_422),
.B1(n_423),
.B2(n_410),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_416),
.A2(n_417),
.B1(n_386),
.B2(n_383),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_429),
.B(n_430),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_423),
.A2(n_334),
.B1(n_400),
.B2(n_394),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_433),
.A2(n_410),
.B1(n_427),
.B2(n_424),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_428),
.B(n_399),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_434),
.B(n_435),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_426),
.B(n_418),
.C(n_414),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_435),
.B(n_424),
.Y(n_436)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_436),
.Y(n_440)
);

AO221x1_ASAP7_75t_L g439 ( 
.A1(n_437),
.A2(n_432),
.B1(n_431),
.B2(n_412),
.C(n_438),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_439),
.B(n_440),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_441),
.B(n_377),
.C(n_396),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_442),
.B(n_377),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_443),
.B(n_382),
.Y(n_444)
);

HAxp5_ASAP7_75t_SL g445 ( 
.A(n_444),
.B(n_345),
.CON(n_445),
.SN(n_445)
);


endmodule