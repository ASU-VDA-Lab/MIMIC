module real_jpeg_7845_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_38;
wire n_33;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

INVx2_ASAP7_75t_SL g12 ( 
.A(n_0),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_0),
.B(n_17),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_3),
.A2(n_13),
.B1(n_19),
.B2(n_20),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_4),
.A2(n_13),
.B1(n_19),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

OAI21xp33_ASAP7_75t_L g10 ( 
.A1(n_5),
.A2(n_11),
.B(n_16),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_7),
.Y(n_6)
);

OAI22xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_9),
.B1(n_24),
.B2(n_38),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_9),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_10),
.B(n_21),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_11),
.B(n_18),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_13),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_23),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_12),
.A2(n_33),
.B(n_35),
.Y(n_32)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_13),
.A2(n_19),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

BUFx24_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_19),
.B(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_23),
.B(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_24),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_37),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_32),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_32),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);


endmodule