module real_jpeg_32852_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_578;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_605;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_599;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_608;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_588;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_568;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_0),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_0),
.Y(n_267)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_0),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_0),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_1),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_1),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_1),
.B(n_281),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_1),
.A2(n_8),
.B1(n_288),
.B2(n_290),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_1),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_1),
.B(n_469),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_1),
.B(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_1),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_2),
.B(n_605),
.Y(n_604)
);

CKINVDCx11_ASAP7_75t_R g606 ( 
.A(n_2),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_3),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_3),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_5),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_5),
.Y(n_232)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_5),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_6),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_6),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_6),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_6),
.B(n_300),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_6),
.B(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_6),
.B(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_6),
.B(n_452),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_6),
.Y(n_476)
);

INVxp33_ASAP7_75t_L g605 ( 
.A(n_7),
.Y(n_605)
);

NAND2x1_ASAP7_75t_SL g53 ( 
.A(n_8),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_8),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_8),
.B(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_8),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_8),
.B(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_8),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_8),
.B(n_278),
.Y(n_277)
);

NAND2x1_ASAP7_75t_SL g577 ( 
.A(n_8),
.B(n_578),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_9),
.Y(n_113)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_9),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_9),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_10),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_10),
.B(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_R g168 ( 
.A(n_10),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_10),
.B(n_249),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_10),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_10),
.B(n_345),
.Y(n_344)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_10),
.B(n_376),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_12),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_12),
.B(n_38),
.Y(n_37)
);

AND2x4_ASAP7_75t_SL g95 ( 
.A(n_12),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_12),
.B(n_62),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_12),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_12),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_12),
.B(n_199),
.Y(n_198)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_13),
.Y(n_93)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_13),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_14),
.B(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_14),
.B(n_317),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_14),
.B(n_331),
.Y(n_330)
);

NAND2x1_ASAP7_75t_L g340 ( 
.A(n_14),
.B(n_341),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_14),
.B(n_380),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_14),
.B(n_482),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_14),
.B(n_488),
.Y(n_487)
);

AND2x2_ASAP7_75t_SL g526 ( 
.A(n_14),
.B(n_527),
.Y(n_526)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_15),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_15),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_15),
.B(n_465),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_15),
.B(n_530),
.Y(n_529)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_16),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_16),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_16),
.Y(n_323)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_17),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_17),
.B(n_59),
.Y(n_58)
);

NAND2x1_ASAP7_75t_L g65 ( 
.A(n_17),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_17),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_17),
.Y(n_94)
);

NAND2x1p5_ASAP7_75t_L g116 ( 
.A(n_17),
.B(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_17),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_17),
.B(n_96),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_608),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_588),
.B1(n_606),
.B2(n_607),
.Y(n_19)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_20),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_569),
.Y(n_20)
);

OAI21x1_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_255),
.B(n_566),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_203),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_23),
.A2(n_567),
.B(n_568),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_171),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_24),
.B(n_171),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_107),
.C(n_132),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_25),
.B(n_107),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_71),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_26),
.B(n_86),
.C(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_46),
.C(n_57),
.Y(n_26)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_27),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_33),
.B(n_43),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_28),
.A2(n_44),
.B(n_45),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_28),
.A2(n_29),
.B1(n_116),
.B2(n_123),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_28),
.B(n_128),
.C(n_129),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_28),
.B(n_110),
.C(n_116),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_28),
.A2(n_29),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_29),
.B(n_325),
.C(n_330),
.Y(n_336)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_31),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_37),
.B(n_42),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_37),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_R g47 ( 
.A(n_34),
.B(n_48),
.C(n_52),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_34),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_34),
.A2(n_52),
.B1(n_53),
.B2(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_34),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_34),
.B(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_34),
.A2(n_137),
.B1(n_243),
.B2(n_264),
.Y(n_455)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_37),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_41),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_41),
.Y(n_190)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_41),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_41),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_41),
.Y(n_579)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_46),
.A2(n_47),
.B1(n_57),
.B2(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

XNOR2x1_ASAP7_75t_L g135 ( 
.A(n_48),
.B(n_136),
.Y(n_135)
);

XOR2x2_ASAP7_75t_L g195 ( 
.A(n_48),
.B(n_196),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_48),
.B(n_109),
.C(n_197),
.Y(n_580)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_51),
.Y(n_142)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_56),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_56),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_56),
.Y(n_523)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_57),
.Y(n_214)
);

XOR2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_63),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_58),
.B(n_67),
.C(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_58),
.Y(n_584)
);

MAJx2_ASAP7_75t_L g596 ( 
.A(n_58),
.B(n_139),
.C(n_197),
.Y(n_596)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_61),
.Y(n_186)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_61),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_62),
.Y(n_246)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_62),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_62),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_67),
.B2(n_70),
.Y(n_63)
);

MAJx2_ASAP7_75t_L g223 ( 
.A(n_64),
.B(n_224),
.C(n_227),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_64),
.A2(n_65),
.B1(n_225),
.B2(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_69),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_69),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_69),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_86),
.Y(n_71)
);

INVxp33_ASAP7_75t_SL g173 ( 
.A(n_72),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_73),
.B(n_85),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_73),
.B(n_85),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_81),
.B1(n_84),
.B2(n_85),
.Y(n_75)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_81),
.B(n_95),
.C(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_81),
.A2(n_85),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_83),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_84),
.A2(n_193),
.B(n_194),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_101),
.C(n_102),
.Y(n_86)
);

INVxp33_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_88),
.A2(n_89),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_95),
.C(n_97),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_90),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_90),
.A2(n_152),
.B1(n_299),
.B2(n_302),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_90),
.B(n_294),
.C(n_299),
.Y(n_355)
);

OR2x2_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_94),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_95),
.B(n_97),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_95),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_95),
.B(n_446),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_95),
.B(n_447),
.Y(n_519)
);

INVx4_ASAP7_75t_SL g279 ( 
.A(n_96),
.Y(n_279)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_101),
.A2(n_103),
.B1(n_104),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_101),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_101),
.B(n_162),
.C(n_166),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_101),
.A2(n_159),
.B1(n_166),
.B2(n_167),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g599 ( 
.A1(n_101),
.A2(n_139),
.B1(n_140),
.B2(n_159),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_106),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_124),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_108),
.A2(n_177),
.B(n_178),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_114),
.B2(n_115),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_109),
.A2(n_110),
.B1(n_197),
.B2(n_200),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_109),
.A2(n_110),
.B1(n_340),
.B2(n_343),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_109),
.B(n_340),
.C(n_344),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_116),
.A2(n_123),
.B1(n_598),
.B2(n_599),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_127),
.B1(n_130),
.B2(n_131),
.Y(n_124)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_127),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_130),
.B(n_131),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_130),
.B(n_131),
.Y(n_178)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_133),
.B(n_205),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_154),
.C(n_160),
.Y(n_133)
);

XNOR2x1_ASAP7_75t_L g208 ( 
.A(n_134),
.B(n_209),
.Y(n_208)
);

MAJx2_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.C(n_151),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_135),
.B(n_138),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.C(n_146),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g585 ( 
.A1(n_139),
.A2(n_140),
.B1(n_197),
.B2(n_200),
.Y(n_585)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2x1_ASAP7_75t_L g234 ( 
.A(n_140),
.B(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI22x1_ASAP7_75t_SL g235 ( 
.A1(n_143),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_235)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_149),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_149),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_150),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_150),
.Y(n_471)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_151),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_156),
.B(n_161),
.Y(n_209)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_162),
.B(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_163),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_163),
.A2(n_220),
.B1(n_307),
.B2(n_310),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_163),
.B(n_307),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx6_ASAP7_75t_L g450 ( 
.A(n_165),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_165),
.Y(n_503)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_174),
.B1(n_201),
.B2(n_202),
.Y(n_171)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_179),
.B2(n_180),
.Y(n_174)
);

INVxp67_ASAP7_75t_SL g175 ( 
.A(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_176),
.B(n_179),
.C(n_201),
.Y(n_571)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_191),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g587 ( 
.A(n_181),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_182),
.B(n_184),
.C(n_187),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.Y(n_183)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_192),
.B(n_195),
.C(n_587),
.Y(n_586)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_197),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_197),
.A2(n_200),
.B1(n_369),
.B2(n_370),
.Y(n_368)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_240),
.C(n_243),
.Y(n_239)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_199),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_204),
.B(n_206),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.C(n_215),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_208),
.B(n_211),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

INVxp33_ASAP7_75t_SL g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_216),
.B(n_430),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_236),
.C(n_252),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_217),
.B(n_417),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.C(n_233),
.Y(n_217)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_218),
.Y(n_402)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_219),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_223),
.B(n_234),
.Y(n_403)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_225),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_227),
.B(n_357),
.Y(n_356)
);

NOR2xp67_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_232),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_236),
.A2(n_237),
.B1(n_252),
.B2(n_253),
.Y(n_417)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_244),
.C(n_247),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2x1_ASAP7_75t_L g394 ( 
.A(n_239),
.B(n_395),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_240),
.A2(n_243),
.B1(n_264),
.B2(n_371),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_240),
.Y(n_371)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_245),
.B(n_248),
.Y(n_395)
);

INVxp33_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

OA21x2_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_406),
.B(n_557),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_384),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_347),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_259),
.B(n_347),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_303),
.C(n_333),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_260),
.B(n_434),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_275),
.Y(n_260)
);

MAJx2_ASAP7_75t_L g349 ( 
.A(n_261),
.B(n_276),
.C(n_293),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.C(n_268),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_262),
.A2(n_263),
.B1(n_441),
.B2(n_442),
.Y(n_440)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_265),
.A2(n_268),
.B1(n_269),
.B2(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_265),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_267),
.Y(n_289)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_272),
.Y(n_342)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_293),
.Y(n_275)
);

OA21x2_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_280),
.B(n_286),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_285),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_286),
.A2(n_287),
.B1(n_373),
.B2(n_374),
.Y(n_372)
);

INVxp33_ASAP7_75t_SL g286 ( 
.A(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_287),
.B(n_398),
.C(n_399),
.Y(n_397)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_292),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_298),
.Y(n_293)
);

NOR2x1_ASAP7_75t_R g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_308),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_295),
.B(n_502),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_295),
.B(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_299),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_301),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_304),
.B(n_334),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_311),
.C(n_324),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_305),
.A2(n_306),
.B1(n_311),
.B2(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_307),
.Y(n_310)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_311),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_316),
.C(n_319),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_312),
.A2(n_313),
.B1(n_319),
.B2(n_320),
.Y(n_542)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_316),
.B(n_542),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx8_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g437 ( 
.A(n_324),
.B(n_438),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_328),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_338),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_336),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_337),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_338),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_344),
.Y(n_338)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_340),
.Y(n_343)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_359),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_349),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_350),
.B(n_360),
.C(n_405),
.Y(n_404)
);

XNOR2x1_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_354),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

MAJx2_ASAP7_75t_L g392 ( 
.A(n_353),
.B(n_355),
.C(n_356),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_367),
.Y(n_360)
);

OA21x2_ASAP7_75t_L g386 ( 
.A1(n_361),
.A2(n_387),
.B(n_388),
.Y(n_386)
);

OAI21x1_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_365),
.B(n_366),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_363),
.B(n_364),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_372),
.B1(n_382),
.B2(n_383),
.Y(n_367)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_368),
.Y(n_383)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_372),
.Y(n_382)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_379),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_375),
.Y(n_398)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_379),
.Y(n_399)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_382),
.B(n_383),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_382),
.B(n_383),
.Y(n_388)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_384),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_404),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_385),
.B(n_404),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_389),
.Y(n_385)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_386),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_401),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_390),
.Y(n_412)
);

OAI22x1_ASAP7_75t_L g390 ( 
.A1(n_391),
.A2(n_392),
.B1(n_393),
.B2(n_400),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_392),
.B(n_423),
.C(n_424),
.Y(n_422)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_393),
.Y(n_400)
);

XNOR2x1_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_396),
.Y(n_393)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_394),
.Y(n_424)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_397),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_401),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_403),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_431),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_407),
.A2(n_558),
.B(n_562),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_408),
.A2(n_413),
.B1(n_425),
.B2(n_428),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_409),
.B(n_414),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_411),
.C(n_412),
.Y(n_409)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_418),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_416),
.B(n_422),
.C(n_427),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_422),
.Y(n_418)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_419),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_421),
.Y(n_419)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

NOR2x1_ASAP7_75t_L g563 ( 
.A(n_426),
.B(n_429),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_426),
.B(n_429),
.Y(n_565)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_429),
.Y(n_428)
);

AO21x1_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_456),
.B(n_556),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_433),
.B(n_435),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_433),
.B(n_435),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_440),
.C(n_444),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_436),
.A2(n_437),
.B1(n_553),
.B2(n_554),
.Y(n_552)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_440),
.B(n_444),
.Y(n_554)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_451),
.C(n_454),
.Y(n_444)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_445),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g448 ( 
.A(n_449),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_451),
.A2(n_454),
.B1(n_455),
.B2(n_546),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_451),
.Y(n_546)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_457),
.A2(n_550),
.B(n_555),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_458),
.A2(n_534),
.B(n_549),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_459),
.A2(n_512),
.B(n_533),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_460),
.A2(n_494),
.B(n_511),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_461),
.B(n_485),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_461),
.B(n_485),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_462),
.A2(n_463),
.B1(n_472),
.B2(n_473),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_464),
.B(n_468),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_464),
.B(n_468),
.C(n_472),
.Y(n_513)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx4_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_474),
.A2(n_475),
.B1(n_480),
.B2(n_481),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_475),
.B(n_480),
.Y(n_517)
);

NOR2x1_ASAP7_75t_SL g475 ( 
.A(n_476),
.B(n_477),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_479),
.Y(n_500)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_484),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_490),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_486),
.A2(n_487),
.B1(n_490),
.B2(n_491),
.Y(n_509)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

BUFx4f_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_495),
.A2(n_504),
.B(n_510),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_496),
.B(n_501),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_498),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_497),
.B(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_509),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_505),
.B(n_509),
.Y(n_510)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_514),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_513),
.B(n_514),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_520),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_516),
.A2(n_517),
.B1(n_518),
.B2(n_519),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_516),
.B(n_519),
.C(n_520),
.Y(n_535)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_524),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_521),
.B(n_526),
.C(n_528),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_523),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_525),
.A2(n_526),
.B1(n_528),
.B2(n_529),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx5_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx5_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_535),
.B(n_536),
.Y(n_534)
);

NOR2xp67_ASAP7_75t_L g549 ( 
.A(n_535),
.B(n_536),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_537),
.A2(n_543),
.B1(n_547),
.B2(n_548),
.Y(n_536)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_537),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_538),
.A2(n_539),
.B1(n_540),
.B2(n_541),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_539),
.B(n_540),
.C(n_548),
.Y(n_551)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_543),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_544),
.B(n_545),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_551),
.B(n_552),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_551),
.B(n_552),
.Y(n_555)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g558 ( 
.A1(n_559),
.A2(n_560),
.B(n_561),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_L g562 ( 
.A1(n_563),
.A2(n_564),
.B(n_565),
.Y(n_562)
);

INVxp33_ASAP7_75t_SL g569 ( 
.A(n_570),
.Y(n_569)
);

NOR2xp67_ASAP7_75t_L g570 ( 
.A(n_571),
.B(n_572),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_571),
.B(n_572),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_573),
.B(n_586),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_574),
.B(n_575),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_574),
.B(n_575),
.C(n_586),
.Y(n_602)
);

XOR2xp5_ASAP7_75t_L g575 ( 
.A(n_576),
.B(n_583),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_577),
.A2(n_580),
.B1(n_581),
.B2(n_582),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_577),
.Y(n_581)
);

BUFx4f_ASAP7_75t_SL g578 ( 
.A(n_579),
.Y(n_578)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_580),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_580),
.B(n_581),
.C(n_583),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_SL g583 ( 
.A(n_584),
.B(n_585),
.Y(n_583)
);

NOR3xp33_ASAP7_75t_L g588 ( 
.A(n_589),
.B(n_591),
.C(n_604),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_L g608 ( 
.A1(n_589),
.A2(n_609),
.B(n_610),
.Y(n_608)
);

INVxp67_ASAP7_75t_SL g589 ( 
.A(n_590),
.Y(n_589)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_592),
.B(n_604),
.Y(n_610)
);

AO21x1_ASAP7_75t_L g592 ( 
.A1(n_593),
.A2(n_602),
.B(n_603),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_593),
.B(n_602),
.Y(n_603)
);

XOR2xp5_ASAP7_75t_L g593 ( 
.A(n_594),
.B(n_601),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_595),
.A2(n_596),
.B1(n_597),
.B2(n_600),
.Y(n_594)
);

CKINVDCx14_ASAP7_75t_R g595 ( 
.A(n_596),
.Y(n_595)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_597),
.Y(n_600)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

INVxp33_ASAP7_75t_L g607 ( 
.A(n_604),
.Y(n_607)
);


endmodule