module fake_jpeg_25717_n_52 (n_3, n_2, n_1, n_0, n_4, n_5, n_52);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_52;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

INVx4_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

INVx11_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_13),
.A2(n_14),
.B1(n_11),
.B2(n_6),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_16),
.B(n_6),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

AO22x1_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_21),
.B1(n_15),
.B2(n_10),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_16),
.B(n_11),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_21),
.B(n_9),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_1),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_14),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_24),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_17),
.A2(n_13),
.B1(n_8),
.B2(n_15),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_12),
.Y(n_27)
);

OA21x2_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_24),
.B(n_12),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_9),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_30),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_29),
.A2(n_23),
.B1(n_15),
.B2(n_19),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_35),
.C(n_16),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_16),
.C(n_19),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_38),
.C(n_16),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_16),
.C(n_19),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

AOI21xp33_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_32),
.B(n_33),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_42),
.C(n_18),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_3),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_45),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_16),
.C(n_19),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_18),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

OAI211xp5_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_3),
.B(n_4),
.C(n_18),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_3),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_49),
.Y(n_52)
);


endmodule