module fake_netlist_1_9643_n_45 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_45);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_43;
wire n_40;
wire n_29;
wire n_39;
CKINVDCx20_ASAP7_75t_R g15 ( .A(n_10), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_2), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_11), .Y(n_17) );
HB1xp67_ASAP7_75t_L g18 ( .A(n_8), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_12), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_0), .Y(n_20) );
HB1xp67_ASAP7_75t_L g21 ( .A(n_6), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_1), .B(n_3), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_17), .Y(n_23) );
AOI22xp33_ASAP7_75t_L g24 ( .A1(n_16), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_24) );
NOR2xp33_ASAP7_75t_L g25 ( .A(n_18), .B(n_3), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_21), .B(n_4), .Y(n_26) );
OAI21x1_ASAP7_75t_L g27 ( .A1(n_23), .A2(n_17), .B(n_19), .Y(n_27) );
AO21x2_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_22), .B(n_20), .Y(n_28) );
AOI21xp5_ASAP7_75t_L g29 ( .A1(n_25), .A2(n_15), .B(n_9), .Y(n_29) );
OR2x2_ASAP7_75t_L g30 ( .A(n_28), .B(n_24), .Y(n_30) );
OR2x2_ASAP7_75t_L g31 ( .A(n_28), .B(n_24), .Y(n_31) );
INVx2_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
AND2x2_ASAP7_75t_L g33 ( .A(n_31), .B(n_29), .Y(n_33) );
INVxp67_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
INVx2_ASAP7_75t_L g35 ( .A(n_33), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_35), .Y(n_36) );
INVxp67_ASAP7_75t_L g37 ( .A(n_34), .Y(n_37) );
NAND2xp33_ASAP7_75t_L g38 ( .A(n_35), .B(n_15), .Y(n_38) );
NAND2xp5_ASAP7_75t_L g39 ( .A(n_36), .B(n_29), .Y(n_39) );
NOR2x1_ASAP7_75t_L g40 ( .A(n_38), .B(n_4), .Y(n_40) );
NOR3xp33_ASAP7_75t_SL g41 ( .A(n_36), .B(n_5), .C(n_6), .Y(n_41) );
NOR2xp33_ASAP7_75t_L g42 ( .A(n_40), .B(n_37), .Y(n_42) );
NAND3xp33_ASAP7_75t_L g43 ( .A(n_41), .B(n_5), .C(n_27), .Y(n_43) );
OAI22xp5_ASAP7_75t_SL g44 ( .A1(n_42), .A2(n_39), .B1(n_13), .B2(n_14), .Y(n_44) );
OAI21xp5_ASAP7_75t_L g45 ( .A1(n_44), .A2(n_43), .B(n_7), .Y(n_45) );
endmodule