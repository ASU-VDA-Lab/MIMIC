module fake_aes_1481_n_717 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_717);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_717;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_146;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_47), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_72), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_62), .Y(n_81) );
INVxp33_ASAP7_75t_L g82 ( .A(n_53), .Y(n_82) );
INVxp33_ASAP7_75t_L g83 ( .A(n_28), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_76), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_44), .Y(n_85) );
BUFx3_ASAP7_75t_L g86 ( .A(n_38), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_52), .Y(n_87) );
INVxp67_ASAP7_75t_L g88 ( .A(n_6), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_75), .Y(n_89) );
INVxp33_ASAP7_75t_L g90 ( .A(n_3), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_31), .Y(n_91) );
INVxp67_ASAP7_75t_L g92 ( .A(n_26), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_51), .Y(n_93) );
INVxp33_ASAP7_75t_SL g94 ( .A(n_10), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_36), .Y(n_95) );
INVxp33_ASAP7_75t_L g96 ( .A(n_10), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_54), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_2), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_67), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_5), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_37), .Y(n_101) );
INVxp67_ASAP7_75t_L g102 ( .A(n_23), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_59), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_19), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_66), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_4), .Y(n_106) );
INVxp67_ASAP7_75t_L g107 ( .A(n_42), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_61), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_15), .Y(n_110) );
BUFx3_ASAP7_75t_L g111 ( .A(n_3), .Y(n_111) );
INVxp33_ASAP7_75t_SL g112 ( .A(n_78), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_41), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_1), .Y(n_114) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_40), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_77), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_24), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_14), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_32), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_27), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_46), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_6), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_55), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_57), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_11), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_0), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_22), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_79), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_115), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_115), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_111), .B(n_0), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_79), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_98), .B(n_1), .Y(n_133) );
INVx1_ASAP7_75t_SL g134 ( .A(n_104), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_115), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_80), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_80), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_81), .Y(n_138) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_111), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_122), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_115), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_81), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_90), .B(n_4), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_85), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_85), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_115), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_87), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_120), .Y(n_148) );
AOI22xp5_ASAP7_75t_L g149 ( .A1(n_94), .A2(n_5), .B1(n_7), .B2(n_8), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_98), .B(n_7), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_120), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_125), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_87), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_91), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_120), .Y(n_155) );
OAI21x1_ASAP7_75t_L g156 ( .A1(n_84), .A2(n_35), .B(n_73), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_91), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_120), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_93), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_100), .B(n_8), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_100), .B(n_9), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_109), .B(n_9), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_120), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_96), .B(n_11), .Y(n_164) );
OAI21x1_ASAP7_75t_L g165 ( .A1(n_84), .A2(n_39), .B(n_71), .Y(n_165) );
INVxp33_ASAP7_75t_SL g166 ( .A(n_106), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_93), .Y(n_167) );
BUFx2_ASAP7_75t_L g168 ( .A(n_88), .Y(n_168) );
OAI21x1_ASAP7_75t_L g169 ( .A1(n_89), .A2(n_34), .B(n_70), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_97), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_97), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_139), .B(n_82), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_139), .B(n_83), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_145), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_145), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_135), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_135), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_145), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_128), .B(n_99), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_140), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_129), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_145), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_168), .B(n_127), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_145), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_134), .B(n_107), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_128), .B(n_102), .Y(n_186) );
NAND2x1p5_ASAP7_75t_L g187 ( .A(n_160), .B(n_119), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_160), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g189 ( .A1(n_160), .A2(n_126), .B1(n_109), .B2(n_110), .Y(n_189) );
OAI22xp5_ASAP7_75t_SL g190 ( .A1(n_149), .A2(n_127), .B1(n_126), .B2(n_110), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_129), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_160), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_135), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_168), .B(n_114), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_166), .B(n_92), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_134), .B(n_112), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_152), .B(n_103), .Y(n_197) );
BUFx2_ASAP7_75t_L g198 ( .A(n_143), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_160), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_161), .Y(n_200) );
BUFx2_ASAP7_75t_L g201 ( .A(n_143), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_161), .Y(n_202) );
AND2x6_ASAP7_75t_L g203 ( .A(n_161), .B(n_124), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_129), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_141), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_161), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_161), .Y(n_207) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_129), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_162), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_129), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_132), .B(n_116), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_143), .B(n_114), .Y(n_212) );
OAI21xp33_ASAP7_75t_L g213 ( .A1(n_132), .A2(n_118), .B(n_86), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_136), .B(n_105), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_162), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_162), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_162), .Y(n_217) );
OAI221xp5_ASAP7_75t_L g218 ( .A1(n_133), .A2(n_118), .B1(n_95), .B2(n_121), .C(n_119), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_162), .Y(n_219) );
BUFx4f_ASAP7_75t_L g220 ( .A(n_131), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_131), .Y(n_221) );
INVx2_ASAP7_75t_SL g222 ( .A(n_131), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_136), .B(n_89), .Y(n_223) );
AND2x4_ASAP7_75t_L g224 ( .A(n_131), .B(n_124), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_137), .B(n_123), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_131), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_141), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_137), .B(n_86), .Y(n_228) );
CKINVDCx16_ASAP7_75t_R g229 ( .A(n_164), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g230 ( .A1(n_164), .A2(n_123), .B1(n_121), .B2(n_117), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_141), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_138), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_138), .Y(n_233) );
INVxp67_ASAP7_75t_SL g234 ( .A(n_164), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_142), .B(n_117), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_142), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_144), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_220), .B(n_171), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_174), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_198), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_198), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_180), .Y(n_242) );
INVx2_ASAP7_75t_SL g243 ( .A(n_220), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_203), .A2(n_171), .B1(n_170), .B2(n_154), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_174), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_187), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_201), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_173), .B(n_170), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_201), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_234), .Y(n_250) );
AND2x6_ASAP7_75t_L g251 ( .A(n_188), .B(n_101), .Y(n_251) );
BUFx2_ASAP7_75t_L g252 ( .A(n_203), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_229), .A2(n_149), .B1(n_167), .B2(n_157), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_175), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_175), .Y(n_255) );
BUFx12f_ASAP7_75t_L g256 ( .A(n_180), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_195), .B(n_157), .Y(n_257) );
AOI221xp5_ASAP7_75t_L g258 ( .A1(n_190), .A2(n_154), .B1(n_159), .B2(n_167), .C(n_153), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_172), .Y(n_259) );
AND2x4_ASAP7_75t_L g260 ( .A(n_212), .B(n_133), .Y(n_260) );
BUFx12f_ASAP7_75t_L g261 ( .A(n_172), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_179), .B(n_153), .Y(n_262) );
BUFx12f_ASAP7_75t_L g263 ( .A(n_187), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_212), .B(n_147), .Y(n_264) );
INVx4_ASAP7_75t_L g265 ( .A(n_203), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_224), .B(n_150), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_186), .B(n_147), .Y(n_267) );
BUFx12f_ASAP7_75t_L g268 ( .A(n_187), .Y(n_268) );
BUFx3_ASAP7_75t_L g269 ( .A(n_203), .Y(n_269) );
INVxp67_ASAP7_75t_L g270 ( .A(n_183), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_232), .B(n_159), .Y(n_271) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_220), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_178), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_178), .Y(n_274) );
BUFx3_ASAP7_75t_L g275 ( .A(n_203), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_182), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_232), .B(n_144), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_196), .B(n_150), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_183), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_185), .B(n_113), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_203), .A2(n_101), .B1(n_108), .B2(n_113), .Y(n_281) );
INVx3_ASAP7_75t_L g282 ( .A(n_207), .Y(n_282) );
AO21x2_ASAP7_75t_L g283 ( .A1(n_188), .A2(n_169), .B(n_165), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_224), .B(n_169), .Y(n_284) );
INVx4_ASAP7_75t_L g285 ( .A(n_203), .Y(n_285) );
O2A1O1Ixp33_ASAP7_75t_L g286 ( .A1(n_218), .A2(n_108), .B(n_116), .C(n_163), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_182), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_194), .A2(n_169), .B1(n_165), .B2(n_156), .Y(n_288) );
CKINVDCx6p67_ASAP7_75t_R g289 ( .A(n_197), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_233), .Y(n_290) );
INVx5_ASAP7_75t_L g291 ( .A(n_207), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_233), .B(n_165), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_224), .B(n_156), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_236), .B(n_156), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_236), .B(n_163), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_222), .Y(n_296) );
INVx4_ASAP7_75t_L g297 ( .A(n_207), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_194), .A2(n_230), .B1(n_189), .B2(n_192), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_184), .Y(n_299) );
NAND2x1p5_ASAP7_75t_L g300 ( .A(n_209), .B(n_163), .Y(n_300) );
INVx4_ASAP7_75t_L g301 ( .A(n_209), .Y(n_301) );
INVx5_ASAP7_75t_L g302 ( .A(n_209), .Y(n_302) );
BUFx2_ASAP7_75t_L g303 ( .A(n_192), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_237), .B(n_158), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_237), .Y(n_305) );
BUFx12f_ASAP7_75t_L g306 ( .A(n_222), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_199), .B(n_49), .Y(n_307) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_246), .Y(n_308) );
INVx5_ASAP7_75t_L g309 ( .A(n_263), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_250), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_265), .B(n_217), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_263), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_239), .Y(n_313) );
INVx4_ASAP7_75t_L g314 ( .A(n_268), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_284), .A2(n_215), .B(n_216), .Y(n_315) );
INVx2_ASAP7_75t_SL g316 ( .A(n_268), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_260), .B(n_216), .Y(n_317) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_246), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_265), .B(n_217), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_246), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_260), .B(n_215), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_282), .Y(n_322) );
INVx5_ASAP7_75t_L g323 ( .A(n_246), .Y(n_323) );
NAND2x1_ASAP7_75t_L g324 ( .A(n_265), .B(n_217), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_282), .Y(n_325) );
INVx5_ASAP7_75t_L g326 ( .A(n_285), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_252), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_282), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_269), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_260), .A2(n_202), .B1(n_206), .B2(n_219), .Y(n_330) );
BUFx4_ASAP7_75t_SL g331 ( .A(n_242), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_264), .Y(n_332) );
INVx5_ASAP7_75t_L g333 ( .A(n_285), .Y(n_333) );
A2O1A1Ixp33_ASAP7_75t_L g334 ( .A1(n_257), .A2(n_206), .B(n_202), .C(n_219), .Y(n_334) );
CKINVDCx16_ASAP7_75t_R g335 ( .A(n_256), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_266), .B(n_200), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_239), .Y(n_337) );
INVx6_ASAP7_75t_L g338 ( .A(n_306), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_285), .B(n_226), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_271), .Y(n_340) );
INVx4_ASAP7_75t_L g341 ( .A(n_272), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g342 ( .A1(n_259), .A2(n_226), .B1(n_221), .B2(n_214), .Y(n_342) );
INVx4_ASAP7_75t_L g343 ( .A(n_272), .Y(n_343) );
OR2x6_ASAP7_75t_SL g344 ( .A(n_242), .B(n_211), .Y(n_344) );
BUFx3_ASAP7_75t_L g345 ( .A(n_269), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_245), .Y(n_346) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_252), .Y(n_347) );
O2A1O1Ixp33_ASAP7_75t_SL g348 ( .A1(n_292), .A2(n_221), .B(n_223), .C(n_225), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_277), .Y(n_349) );
BUFx3_ASAP7_75t_L g350 ( .A(n_275), .Y(n_350) );
AO32x2_ASAP7_75t_L g351 ( .A1(n_297), .A2(n_213), .A3(n_228), .B1(n_155), .B2(n_148), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_256), .Y(n_352) );
CKINVDCx20_ASAP7_75t_R g353 ( .A(n_259), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_266), .B(n_184), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_279), .B(n_235), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_270), .B(n_12), .Y(n_356) );
AOI21xp33_ASAP7_75t_L g357 ( .A1(n_243), .A2(n_231), .B(n_227), .Y(n_357) );
INVx2_ASAP7_75t_SL g358 ( .A(n_261), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_275), .B(n_12), .Y(n_359) );
BUFx2_ASAP7_75t_L g360 ( .A(n_261), .Y(n_360) );
BUFx10_ASAP7_75t_L g361 ( .A(n_266), .Y(n_361) );
AO31x2_ASAP7_75t_L g362 ( .A1(n_334), .A2(n_294), .A3(n_307), .B(n_305), .Y(n_362) );
AND2x6_ASAP7_75t_L g363 ( .A(n_359), .B(n_284), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_332), .B(n_298), .Y(n_364) );
OR2x6_ASAP7_75t_L g365 ( .A(n_314), .B(n_306), .Y(n_365) );
INVx3_ASAP7_75t_L g366 ( .A(n_309), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_340), .A2(n_303), .B1(n_293), .B2(n_284), .Y(n_367) );
OAI22xp33_ASAP7_75t_L g368 ( .A1(n_344), .A2(n_253), .B1(n_248), .B2(n_303), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_309), .A2(n_240), .B1(n_247), .B2(n_249), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_349), .B(n_267), .Y(n_370) );
AOI221xp5_ASAP7_75t_L g371 ( .A1(n_310), .A2(n_258), .B1(n_241), .B2(n_278), .C(n_355), .Y(n_371) );
OAI22xp33_ASAP7_75t_L g372 ( .A1(n_309), .A2(n_288), .B1(n_262), .B2(n_290), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_309), .A2(n_251), .B1(n_272), .B2(n_301), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_339), .A2(n_251), .B1(n_272), .B2(n_301), .Y(n_374) );
INVx2_ASAP7_75t_SL g375 ( .A(n_338), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_330), .A2(n_293), .B1(n_244), .B2(n_281), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_361), .B(n_280), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_312), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g379 ( .A1(n_348), .A2(n_293), .B(n_238), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_356), .Y(n_380) );
O2A1O1Ixp33_ASAP7_75t_L g381 ( .A1(n_334), .A2(n_286), .B(n_238), .C(n_243), .Y(n_381) );
INVx4_ASAP7_75t_L g382 ( .A(n_314), .Y(n_382) );
OAI21xp5_ASAP7_75t_L g383 ( .A1(n_315), .A2(n_273), .B(n_276), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_359), .A2(n_251), .B1(n_297), .B2(n_301), .Y(n_384) );
AOI22xp33_ASAP7_75t_SL g385 ( .A1(n_353), .A2(n_251), .B1(n_283), .B2(n_297), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_316), .B(n_289), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_361), .B(n_251), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_317), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_330), .B(n_251), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_313), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_359), .A2(n_273), .B1(n_274), .B2(n_245), .Y(n_391) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_353), .A2(n_254), .B1(n_255), .B2(n_274), .C(n_299), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_321), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_338), .A2(n_289), .B1(n_302), .B2(n_291), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_354), .Y(n_395) );
BUFx2_ASAP7_75t_L g396 ( .A(n_363), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_370), .B(n_313), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_390), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_388), .B(n_337), .Y(n_399) );
BUFx12f_ASAP7_75t_L g400 ( .A(n_382), .Y(n_400) );
BUFx2_ASAP7_75t_L g401 ( .A(n_363), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_368), .A2(n_339), .B1(n_358), .B2(n_360), .Y(n_402) );
INVx2_ASAP7_75t_SL g403 ( .A(n_366), .Y(n_403) );
OAI22xp33_ASAP7_75t_L g404 ( .A1(n_368), .A2(n_335), .B1(n_338), .B2(n_352), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_391), .A2(n_336), .B1(n_337), .B2(n_346), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_364), .B(n_352), .Y(n_406) );
INVx4_ASAP7_75t_L g407 ( .A(n_363), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_395), .Y(n_408) );
BUFx12f_ASAP7_75t_L g409 ( .A(n_382), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_391), .B(n_346), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_385), .A2(n_339), .B1(n_347), .B2(n_327), .Y(n_411) );
AOI22xp33_ASAP7_75t_SL g412 ( .A1(n_363), .A2(n_331), .B1(n_327), .B2(n_347), .Y(n_412) );
BUFx12f_ASAP7_75t_L g413 ( .A(n_365), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_384), .A2(n_323), .B1(n_342), .B2(n_318), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_385), .A2(n_311), .B1(n_319), .B2(n_296), .Y(n_415) );
A2O1A1Ixp33_ASAP7_75t_L g416 ( .A1(n_381), .A2(n_392), .B(n_367), .C(n_389), .Y(n_416) );
OAI22xp33_ASAP7_75t_L g417 ( .A1(n_365), .A2(n_331), .B1(n_326), .B2(n_333), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_384), .A2(n_323), .B1(n_318), .B2(n_308), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_363), .A2(n_311), .B1(n_319), .B2(n_296), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_371), .B(n_323), .Y(n_420) );
AOI21xp33_ASAP7_75t_L g421 ( .A1(n_372), .A2(n_341), .B(n_343), .Y(n_421) );
INVxp67_ASAP7_75t_L g422 ( .A(n_378), .Y(n_422) );
OAI22xp33_ASAP7_75t_L g423 ( .A1(n_365), .A2(n_326), .B1(n_333), .B2(n_323), .Y(n_423) );
OAI22xp33_ASAP7_75t_L g424 ( .A1(n_366), .A2(n_326), .B1(n_333), .B2(n_343), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_406), .B(n_386), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_398), .Y(n_426) );
AOI33xp33_ASAP7_75t_L g427 ( .A1(n_402), .A2(n_380), .A3(n_369), .B1(n_375), .B2(n_372), .B3(n_393), .Y(n_427) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_397), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_397), .Y(n_429) );
AOI222xp33_ASAP7_75t_L g430 ( .A1(n_404), .A2(n_376), .B1(n_377), .B2(n_383), .C1(n_373), .C2(n_387), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_398), .Y(n_431) );
AOI21xp33_ASAP7_75t_SL g432 ( .A1(n_417), .A2(n_394), .B(n_14), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_410), .Y(n_433) );
OR2x6_ASAP7_75t_L g434 ( .A(n_407), .B(n_308), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_399), .B(n_362), .Y(n_435) );
OAI222xp33_ASAP7_75t_L g436 ( .A1(n_412), .A2(n_379), .B1(n_374), .B2(n_341), .C1(n_320), .C2(n_322), .Y(n_436) );
BUFx2_ASAP7_75t_L g437 ( .A(n_418), .Y(n_437) );
NAND3xp33_ASAP7_75t_L g438 ( .A(n_415), .B(n_348), .C(n_148), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_410), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_408), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_413), .A2(n_325), .B1(n_328), .B2(n_296), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_408), .Y(n_442) );
OA21x2_ASAP7_75t_L g443 ( .A1(n_416), .A2(n_357), .B(n_151), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_399), .Y(n_444) );
OAI221xp5_ASAP7_75t_L g445 ( .A1(n_420), .A2(n_324), .B1(n_300), .B2(n_295), .C(n_304), .Y(n_445) );
OAI22xp33_ASAP7_75t_L g446 ( .A1(n_407), .A2(n_326), .B1(n_333), .B2(n_308), .Y(n_446) );
OAI221xp5_ASAP7_75t_L g447 ( .A1(n_422), .A2(n_300), .B1(n_320), .B2(n_302), .C(n_291), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_405), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_411), .A2(n_318), .B1(n_308), .B2(n_311), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_400), .Y(n_450) );
INVx2_ASAP7_75t_SL g451 ( .A(n_400), .Y(n_451) );
OAI22xp33_ASAP7_75t_L g452 ( .A1(n_407), .A2(n_318), .B1(n_329), .B2(n_350), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_396), .B(n_362), .Y(n_453) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_396), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_418), .Y(n_455) );
OAI221xp5_ASAP7_75t_L g456 ( .A1(n_419), .A2(n_291), .B1(n_302), .B2(n_299), .C(n_254), .Y(n_456) );
NAND2x1p5_ASAP7_75t_SL g457 ( .A(n_403), .B(n_362), .Y(n_457) );
OAI21x1_ASAP7_75t_L g458 ( .A1(n_405), .A2(n_146), .B(n_158), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_401), .B(n_403), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_409), .B(n_362), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_409), .B(n_255), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_430), .A2(n_413), .B1(n_401), .B2(n_423), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_435), .B(n_351), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_428), .B(n_414), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_435), .B(n_351), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_429), .B(n_421), .Y(n_466) );
INVxp67_ASAP7_75t_SL g467 ( .A(n_444), .Y(n_467) );
AOI221xp5_ASAP7_75t_L g468 ( .A1(n_425), .A2(n_146), .B1(n_158), .B2(n_151), .C(n_424), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_440), .B(n_13), .Y(n_469) );
OAI31xp33_ASAP7_75t_L g470 ( .A1(n_449), .A2(n_319), .A3(n_287), .B(n_276), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_444), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_440), .B(n_13), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_453), .B(n_351), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_453), .B(n_351), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_442), .B(n_15), .Y(n_475) );
OAI31xp33_ASAP7_75t_L g476 ( .A1(n_449), .A2(n_287), .A3(n_350), .B(n_345), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_432), .B(n_329), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_444), .B(n_151), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_442), .B(n_146), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_426), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_433), .B(n_16), .Y(n_481) );
AOI31xp33_ASAP7_75t_L g482 ( .A1(n_451), .A2(n_16), .A3(n_17), .B(n_18), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_426), .B(n_17), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_431), .Y(n_484) );
BUFx2_ASAP7_75t_L g485 ( .A(n_454), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_433), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_451), .B(n_18), .Y(n_487) );
AO22x1_ASAP7_75t_L g488 ( .A1(n_460), .A2(n_329), .B1(n_345), .B2(n_21), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_431), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_427), .B(n_19), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_433), .B(n_20), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_430), .B(n_20), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_439), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_448), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_439), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_432), .B(n_329), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_448), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_439), .B(n_21), .Y(n_498) );
BUFx3_ASAP7_75t_L g499 ( .A(n_454), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_461), .B(n_22), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_457), .Y(n_501) );
BUFx2_ASAP7_75t_L g502 ( .A(n_454), .Y(n_502) );
NAND4xp25_ASAP7_75t_L g503 ( .A(n_438), .B(n_177), .C(n_231), .D(n_227), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_443), .B(n_283), .Y(n_504) );
A2O1A1Ixp33_ASAP7_75t_SL g505 ( .A1(n_447), .A2(n_176), .B(n_205), .C(n_193), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_437), .A2(n_296), .B1(n_283), .B2(n_291), .Y(n_506) );
NOR3xp33_ASAP7_75t_SL g507 ( .A(n_436), .B(n_25), .C(n_29), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_457), .B(n_129), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_454), .B(n_30), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_459), .B(n_302), .Y(n_510) );
OAI33xp33_ASAP7_75t_L g511 ( .A1(n_459), .A2(n_176), .A3(n_205), .B1(n_193), .B2(n_177), .B3(n_129), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_457), .Y(n_512) );
NAND4xp25_ASAP7_75t_L g513 ( .A(n_438), .B(n_155), .C(n_148), .D(n_130), .Y(n_513) );
NOR3xp33_ASAP7_75t_L g514 ( .A(n_482), .B(n_450), .C(n_456), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_480), .Y(n_515) );
NAND4xp25_ASAP7_75t_SL g516 ( .A(n_462), .B(n_441), .C(n_455), .D(n_445), .Y(n_516) );
OAI21xp5_ASAP7_75t_L g517 ( .A1(n_492), .A2(n_458), .B(n_443), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_463), .B(n_437), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_484), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_489), .Y(n_520) );
INVx3_ASAP7_75t_L g521 ( .A(n_508), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_463), .B(n_455), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_489), .B(n_454), .Y(n_523) );
NAND4xp25_ASAP7_75t_SL g524 ( .A(n_462), .B(n_455), .C(n_434), .D(n_446), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_484), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_465), .B(n_443), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_481), .B(n_443), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_471), .Y(n_528) );
AND2x4_ASAP7_75t_L g529 ( .A(n_512), .B(n_434), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_465), .B(n_458), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_491), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_490), .A2(n_434), .B1(n_452), .B2(n_130), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_473), .B(n_434), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_473), .B(n_434), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_467), .B(n_155), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_491), .B(n_155), .Y(n_536) );
NAND2x1p5_ASAP7_75t_L g537 ( .A(n_509), .B(n_302), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_508), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_481), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_498), .Y(n_540) );
BUFx2_ASAP7_75t_L g541 ( .A(n_485), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_487), .A2(n_291), .B1(n_130), .B2(n_155), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_498), .B(n_155), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_479), .B(n_155), .Y(n_544) );
INVx1_ASAP7_75t_SL g545 ( .A(n_485), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_479), .Y(n_546) );
NAND3xp33_ASAP7_75t_L g547 ( .A(n_512), .B(n_148), .C(n_130), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_494), .B(n_148), .Y(n_548) );
BUFx2_ASAP7_75t_L g549 ( .A(n_502), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_464), .B(n_148), .Y(n_550) );
INVx1_ASAP7_75t_SL g551 ( .A(n_502), .Y(n_551) );
NAND2x1_ASAP7_75t_L g552 ( .A(n_509), .B(n_148), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_474), .B(n_130), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_469), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_466), .B(n_130), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_474), .B(n_130), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_477), .A2(n_208), .B1(n_204), .B2(n_191), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_472), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_475), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_494), .B(n_33), .Y(n_560) );
AND2x4_ASAP7_75t_L g561 ( .A(n_501), .B(n_43), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_486), .Y(n_562) );
NOR2x1_ASAP7_75t_L g563 ( .A(n_513), .B(n_210), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_466), .B(n_45), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_486), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_486), .B(n_48), .Y(n_566) );
NAND2x1p5_ASAP7_75t_L g567 ( .A(n_509), .B(n_50), .Y(n_567) );
AND2x4_ASAP7_75t_L g568 ( .A(n_501), .B(n_56), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_497), .B(n_58), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_483), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_493), .Y(n_571) );
NOR2x1_ASAP7_75t_L g572 ( .A(n_513), .B(n_210), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_497), .B(n_60), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_554), .B(n_495), .Y(n_574) );
AND2x4_ASAP7_75t_SL g575 ( .A(n_529), .B(n_509), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_515), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_558), .B(n_493), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_522), .B(n_501), .Y(n_578) );
INVxp67_ASAP7_75t_L g579 ( .A(n_541), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_559), .B(n_496), .Y(n_580) );
CKINVDCx16_ASAP7_75t_R g581 ( .A(n_533), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_528), .B(n_493), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_522), .B(n_495), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_520), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_570), .B(n_495), .Y(n_585) );
INVxp67_ASAP7_75t_L g586 ( .A(n_549), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_518), .B(n_499), .Y(n_587) );
NOR2x1_ASAP7_75t_L g588 ( .A(n_563), .B(n_572), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_525), .Y(n_589) );
AOI21xp33_ASAP7_75t_SL g590 ( .A1(n_514), .A2(n_488), .B(n_470), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_519), .Y(n_591) );
AOI221x1_ASAP7_75t_L g592 ( .A1(n_543), .A2(n_503), .B1(n_500), .B2(n_478), .C(n_504), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_518), .B(n_504), .Y(n_593) );
NAND2xp33_ASAP7_75t_SL g594 ( .A(n_552), .B(n_507), .Y(n_594) );
INVx1_ASAP7_75t_SL g595 ( .A(n_545), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_555), .Y(n_596) );
XOR2xp5_ASAP7_75t_L g597 ( .A(n_524), .B(n_488), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_550), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_546), .B(n_478), .Y(n_599) );
A2O1A1Ixp33_ASAP7_75t_L g600 ( .A1(n_561), .A2(n_470), .B(n_476), .C(n_503), .Y(n_600) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_538), .Y(n_601) );
NOR2x1_ASAP7_75t_L g602 ( .A(n_547), .B(n_499), .Y(n_602) );
INVxp67_ASAP7_75t_SL g603 ( .A(n_538), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_562), .Y(n_604) );
INVx2_ASAP7_75t_SL g605 ( .A(n_535), .Y(n_605) );
INVxp67_ASAP7_75t_L g606 ( .A(n_553), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_516), .A2(n_511), .B1(n_510), .B2(n_476), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_531), .B(n_506), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_539), .B(n_499), .Y(n_609) );
AND2x2_ASAP7_75t_SL g610 ( .A(n_561), .B(n_468), .Y(n_610) );
OR2x2_ASAP7_75t_L g611 ( .A(n_521), .B(n_551), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_526), .B(n_63), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_564), .B(n_64), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_526), .B(n_65), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_553), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_556), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_540), .B(n_505), .Y(n_617) );
OAI211xp5_ASAP7_75t_SL g618 ( .A1(n_542), .A2(n_68), .B(n_69), .C(n_74), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_530), .B(n_181), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_562), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_556), .Y(n_621) );
OAI21xp5_ASAP7_75t_L g622 ( .A1(n_573), .A2(n_181), .B(n_191), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_565), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_565), .B(n_181), .Y(n_624) );
NOR2x1p5_ASAP7_75t_L g625 ( .A(n_521), .B(n_210), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_574), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_601), .B(n_521), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_603), .B(n_530), .Y(n_628) );
NOR2xp67_ASAP7_75t_SL g629 ( .A(n_612), .B(n_573), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_581), .B(n_534), .Y(n_630) );
INVxp67_ASAP7_75t_L g631 ( .A(n_588), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_577), .Y(n_632) );
NAND4xp25_ASAP7_75t_L g633 ( .A(n_590), .B(n_532), .C(n_517), .D(n_529), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_578), .B(n_534), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_585), .Y(n_635) );
INVxp67_ASAP7_75t_SL g636 ( .A(n_625), .Y(n_636) );
OR2x2_ASAP7_75t_L g637 ( .A(n_593), .B(n_523), .Y(n_637) );
INVx3_ASAP7_75t_L g638 ( .A(n_575), .Y(n_638) );
AND2x4_ASAP7_75t_L g639 ( .A(n_605), .B(n_529), .Y(n_639) );
AOI221xp5_ASAP7_75t_L g640 ( .A1(n_580), .A2(n_532), .B1(n_533), .B2(n_527), .C(n_548), .Y(n_640) );
OAI211xp5_ASAP7_75t_L g641 ( .A1(n_597), .A2(n_557), .B(n_536), .C(n_560), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_595), .B(n_571), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_602), .B(n_568), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_576), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_584), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_579), .B(n_569), .Y(n_646) );
BUFx2_ASAP7_75t_L g647 ( .A(n_586), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_600), .A2(n_568), .B(n_561), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_589), .Y(n_649) );
XOR2xp5_ASAP7_75t_L g650 ( .A(n_587), .B(n_567), .Y(n_650) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_605), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_580), .B(n_544), .Y(n_652) );
NAND2x1_ASAP7_75t_L g653 ( .A(n_611), .B(n_568), .Y(n_653) );
OAI211xp5_ASAP7_75t_L g654 ( .A1(n_600), .A2(n_557), .B(n_566), .C(n_571), .Y(n_654) );
NOR2x1p5_ASAP7_75t_L g655 ( .A(n_617), .B(n_566), .Y(n_655) );
INVx2_ASAP7_75t_SL g656 ( .A(n_582), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_578), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_596), .B(n_537), .Y(n_658) );
AOI311xp33_ASAP7_75t_L g659 ( .A1(n_615), .A2(n_567), .A3(n_537), .B(n_204), .C(n_208), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_594), .A2(n_181), .B(n_191), .Y(n_660) );
INVxp67_ASAP7_75t_L g661 ( .A(n_591), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_604), .Y(n_662) );
INVx2_ASAP7_75t_SL g663 ( .A(n_575), .Y(n_663) );
XNOR2xp5_ASAP7_75t_L g664 ( .A(n_583), .B(n_181), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_583), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_610), .A2(n_191), .B1(n_204), .B2(n_208), .Y(n_666) );
AOI32xp33_ASAP7_75t_L g667 ( .A1(n_594), .A2(n_191), .A3(n_204), .B1(n_208), .B2(n_210), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_598), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_609), .Y(n_669) );
INVx1_ASAP7_75t_SL g670 ( .A(n_612), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_616), .B(n_204), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_621), .B(n_208), .Y(n_672) );
NAND4xp25_ASAP7_75t_L g673 ( .A(n_592), .B(n_607), .C(n_608), .D(n_613), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_606), .B(n_599), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_610), .B(n_622), .Y(n_675) );
INVxp67_ASAP7_75t_L g676 ( .A(n_619), .Y(n_676) );
XNOR2x1_ASAP7_75t_L g677 ( .A(n_614), .B(n_620), .Y(n_677) );
A2O1A1O1Ixp25_ASAP7_75t_L g678 ( .A1(n_613), .A2(n_607), .B(n_614), .C(n_624), .D(n_618), .Y(n_678) );
INVxp67_ASAP7_75t_L g679 ( .A(n_620), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_623), .B(n_595), .Y(n_680) );
OAI211xp5_ASAP7_75t_L g681 ( .A1(n_590), .A2(n_597), .B(n_600), .C(n_462), .Y(n_681) );
NOR4xp25_ASAP7_75t_L g682 ( .A(n_681), .B(n_631), .C(n_673), .D(n_654), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_633), .A2(n_675), .B1(n_631), .B2(n_641), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_626), .Y(n_684) );
OAI321xp33_ASAP7_75t_L g685 ( .A1(n_636), .A2(n_667), .A3(n_663), .B1(n_666), .B2(n_676), .C(n_647), .Y(n_685) );
O2A1O1Ixp33_ASAP7_75t_L g686 ( .A1(n_678), .A2(n_643), .B(n_651), .C(n_660), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_669), .B(n_651), .Y(n_687) );
AOI221x1_ASAP7_75t_SL g688 ( .A1(n_668), .A2(n_674), .B1(n_628), .B2(n_680), .C(n_627), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_635), .B(n_632), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g690 ( .A1(n_636), .A2(n_643), .B(n_648), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_646), .A2(n_655), .B1(n_677), .B2(n_652), .Y(n_691) );
A2O1A1Ixp33_ASAP7_75t_SL g692 ( .A1(n_666), .A2(n_646), .B(n_652), .C(n_629), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_645), .Y(n_693) );
INVx1_ASAP7_75t_SL g694 ( .A(n_642), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_670), .A2(n_639), .B1(n_676), .B2(n_640), .Y(n_695) );
AOI21xp33_ASAP7_75t_L g696 ( .A1(n_692), .A2(n_664), .B(n_672), .Y(n_696) );
O2A1O1Ixp33_ASAP7_75t_L g697 ( .A1(n_682), .A2(n_644), .B(n_661), .C(n_649), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_688), .A2(n_661), .B1(n_656), .B2(n_665), .C(n_657), .Y(n_698) );
OAI21xp5_ASAP7_75t_L g699 ( .A1(n_683), .A2(n_653), .B(n_650), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_684), .B(n_679), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_691), .B(n_634), .Y(n_701) );
OA22x2_ASAP7_75t_L g702 ( .A1(n_695), .A2(n_694), .B1(n_638), .B2(n_689), .Y(n_702) );
OAI211xp5_ASAP7_75t_L g703 ( .A1(n_686), .A2(n_659), .B(n_638), .C(n_658), .Y(n_703) );
INVx1_ASAP7_75t_SL g704 ( .A(n_700), .Y(n_704) );
OAI322xp33_ASAP7_75t_L g705 ( .A1(n_702), .A2(n_690), .A3(n_687), .B1(n_693), .B2(n_679), .C1(n_685), .C2(n_637), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_697), .Y(n_706) );
AND3x1_ASAP7_75t_L g707 ( .A(n_699), .B(n_687), .C(n_630), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_701), .B(n_639), .Y(n_708) );
XNOR2xp5_ASAP7_75t_L g709 ( .A(n_707), .B(n_703), .Y(n_709) );
NAND3x1_ASAP7_75t_L g710 ( .A(n_706), .B(n_698), .C(n_696), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_704), .Y(n_711) );
OAI221xp5_ASAP7_75t_L g712 ( .A1(n_709), .A2(n_706), .B1(n_711), .B2(n_708), .C(n_710), .Y(n_712) );
AND3x4_ASAP7_75t_L g713 ( .A(n_711), .B(n_705), .C(n_662), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_712), .Y(n_714) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_714), .Y(n_715) );
INVxp67_ASAP7_75t_L g716 ( .A(n_715), .Y(n_716) );
AOI21xp33_ASAP7_75t_L g717 ( .A1(n_716), .A2(n_713), .B(n_671), .Y(n_717) );
endmodule