module real_aes_8899_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g107 ( .A(n_0), .Y(n_107) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_1), .A2(n_136), .B(n_140), .C(n_221), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_2), .A2(n_170), .B(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g513 ( .A(n_3), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_4), .B(n_237), .Y(n_256) );
AOI21xp33_ASAP7_75t_L g478 ( .A1(n_5), .A2(n_170), .B(n_479), .Y(n_478) );
AND2x6_ASAP7_75t_L g136 ( .A(n_6), .B(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g211 ( .A(n_7), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_8), .B(n_113), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_8), .B(n_42), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_9), .A2(n_169), .B(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_10), .B(n_148), .Y(n_223) );
INVx1_ASAP7_75t_L g483 ( .A(n_11), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_12), .B(n_251), .Y(n_538) );
INVx1_ASAP7_75t_L g156 ( .A(n_13), .Y(n_156) );
INVx1_ASAP7_75t_L g550 ( .A(n_14), .Y(n_550) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_15), .A2(n_146), .B(n_233), .C(n_235), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_16), .B(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_17), .B(n_501), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_18), .B(n_170), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_19), .B(n_182), .Y(n_181) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_20), .A2(n_251), .B(n_266), .C(n_268), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_21), .B(n_237), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_22), .B(n_148), .Y(n_193) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_23), .A2(n_178), .B(n_235), .C(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_24), .B(n_148), .Y(n_147) );
CKINVDCx16_ASAP7_75t_R g187 ( .A(n_25), .Y(n_187) );
INVx1_ASAP7_75t_L g144 ( .A(n_26), .Y(n_144) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_27), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_28), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_29), .B(n_148), .Y(n_514) );
OAI22xp5_ASAP7_75t_SL g747 ( .A1(n_30), .A2(n_31), .B1(n_748), .B2(n_749), .Y(n_747) );
INVx1_ASAP7_75t_L g749 ( .A(n_30), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_31), .Y(n_748) );
INVx1_ASAP7_75t_L g176 ( .A(n_32), .Y(n_176) );
INVx1_ASAP7_75t_L g492 ( .A(n_33), .Y(n_492) );
INVx2_ASAP7_75t_L g134 ( .A(n_34), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_35), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_36), .A2(n_251), .B(n_252), .C(n_254), .Y(n_250) );
INVxp67_ASAP7_75t_L g177 ( .A(n_37), .Y(n_177) );
A2O1A1Ixp33_ASAP7_75t_L g139 ( .A1(n_38), .A2(n_140), .B(n_143), .C(n_151), .Y(n_139) );
CKINVDCx14_ASAP7_75t_R g249 ( .A(n_39), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_40), .A2(n_136), .B(n_140), .C(n_525), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_41), .A2(n_104), .B1(n_114), .B2(n_759), .Y(n_103) );
INVx1_ASAP7_75t_L g113 ( .A(n_42), .Y(n_113) );
INVx1_ASAP7_75t_L g491 ( .A(n_43), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_44), .A2(n_195), .B(n_209), .C(n_210), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_45), .B(n_148), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_46), .A2(n_746), .B1(n_747), .B2(n_750), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_46), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_47), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_48), .Y(n_172) );
INVx1_ASAP7_75t_L g264 ( .A(n_49), .Y(n_264) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_50), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_51), .B(n_170), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_52), .B(n_459), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_53), .A2(n_140), .B1(n_268), .B2(n_490), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_54), .Y(n_529) );
CKINVDCx16_ASAP7_75t_R g510 ( .A(n_55), .Y(n_510) );
CKINVDCx14_ASAP7_75t_R g207 ( .A(n_56), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_57), .A2(n_209), .B(n_254), .C(n_482), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_58), .Y(n_566) );
INVx1_ASAP7_75t_L g480 ( .A(n_59), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_60), .A2(n_89), .B1(n_450), .B2(n_451), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_60), .Y(n_451) );
INVx1_ASAP7_75t_L g137 ( .A(n_61), .Y(n_137) );
INVx1_ASAP7_75t_L g155 ( .A(n_62), .Y(n_155) );
INVx1_ASAP7_75t_SL g253 ( .A(n_63), .Y(n_253) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_64), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_65), .B(n_237), .Y(n_270) );
INVx1_ASAP7_75t_L g190 ( .A(n_66), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_SL g500 ( .A1(n_67), .A2(n_254), .B(n_501), .C(n_502), .Y(n_500) );
INVxp67_ASAP7_75t_L g503 ( .A(n_68), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g120 ( .A1(n_69), .A2(n_121), .B1(n_122), .B2(n_123), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_69), .Y(n_121) );
INVx1_ASAP7_75t_L g111 ( .A(n_70), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_71), .A2(n_170), .B(n_206), .Y(n_205) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_72), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_73), .A2(n_170), .B(n_230), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_74), .Y(n_495) );
INVx1_ASAP7_75t_L g560 ( .A(n_75), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_76), .A2(n_169), .B(n_171), .Y(n_168) );
CKINVDCx16_ASAP7_75t_R g138 ( .A(n_77), .Y(n_138) );
INVx1_ASAP7_75t_L g231 ( .A(n_78), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_L g561 ( .A1(n_79), .A2(n_136), .B(n_140), .C(n_562), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_80), .A2(n_170), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g234 ( .A(n_81), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_82), .B(n_145), .Y(n_526) );
INVx2_ASAP7_75t_L g153 ( .A(n_83), .Y(n_153) );
INVx1_ASAP7_75t_L g222 ( .A(n_84), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_85), .B(n_501), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_86), .A2(n_136), .B(n_140), .C(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g108 ( .A(n_87), .Y(n_108) );
OR2x2_ASAP7_75t_L g454 ( .A(n_87), .B(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g466 ( .A(n_87), .B(n_456), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g188 ( .A1(n_88), .A2(n_140), .B(n_189), .C(n_197), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_89), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_90), .B(n_152), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_91), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_92), .A2(n_136), .B(n_140), .C(n_536), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_93), .Y(n_542) );
INVx1_ASAP7_75t_L g499 ( .A(n_94), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g547 ( .A(n_95), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_96), .B(n_145), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_97), .B(n_160), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_98), .B(n_160), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_99), .B(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g267 ( .A(n_100), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_101), .A2(n_170), .B(n_498), .Y(n_497) );
AOI222xp33_ASAP7_75t_L g462 ( .A1(n_102), .A2(n_463), .B1(n_744), .B2(n_745), .C1(n_751), .C2(n_754), .Y(n_462) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_105), .Y(n_759) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_112), .Y(n_105) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_107), .B(n_108), .C(n_109), .Y(n_106) );
AND2x2_ASAP7_75t_L g456 ( .A(n_107), .B(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g469 ( .A(n_108), .B(n_456), .Y(n_469) );
NOR2x2_ASAP7_75t_L g756 ( .A(n_108), .B(n_455), .Y(n_756) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
AO21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_119), .B(n_461), .Y(n_114) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g758 ( .A(n_117), .Y(n_758) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI21xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_452), .B(n_458), .Y(n_119) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
XOR2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_449), .Y(n_123) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_124), .A2(n_464), .B1(n_467), .B2(n_470), .Y(n_463) );
INVx1_ASAP7_75t_L g752 ( .A(n_124), .Y(n_752) );
OR4x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_339), .C(n_386), .D(n_426), .Y(n_124) );
NAND3xp33_ASAP7_75t_SL g125 ( .A(n_126), .B(n_285), .C(n_314), .Y(n_125) );
AOI211xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_200), .B(n_238), .C(n_278), .Y(n_126) );
O2A1O1Ixp33_ASAP7_75t_L g314 ( .A1(n_127), .A2(n_298), .B(n_315), .C(n_319), .Y(n_314) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_162), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_129), .B(n_277), .Y(n_276) );
INVx3_ASAP7_75t_SL g281 ( .A(n_129), .Y(n_281) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_129), .Y(n_293) );
AND2x4_ASAP7_75t_L g297 ( .A(n_129), .B(n_245), .Y(n_297) );
AND2x2_ASAP7_75t_L g308 ( .A(n_129), .B(n_185), .Y(n_308) );
OR2x2_ASAP7_75t_L g332 ( .A(n_129), .B(n_241), .Y(n_332) );
AND2x2_ASAP7_75t_L g345 ( .A(n_129), .B(n_246), .Y(n_345) );
AND2x2_ASAP7_75t_L g385 ( .A(n_129), .B(n_371), .Y(n_385) );
AND2x2_ASAP7_75t_L g392 ( .A(n_129), .B(n_355), .Y(n_392) );
AND2x2_ASAP7_75t_L g422 ( .A(n_129), .B(n_163), .Y(n_422) );
OR2x6_ASAP7_75t_L g129 ( .A(n_130), .B(n_157), .Y(n_129) );
O2A1O1Ixp33_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_138), .B(n_139), .C(n_152), .Y(n_130) );
OAI21xp5_ASAP7_75t_L g186 ( .A1(n_131), .A2(n_187), .B(n_188), .Y(n_186) );
OAI21xp5_ASAP7_75t_L g218 ( .A1(n_131), .A2(n_219), .B(n_220), .Y(n_218) );
OAI22xp33_ASAP7_75t_L g488 ( .A1(n_131), .A2(n_180), .B1(n_489), .B2(n_493), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_131), .A2(n_510), .B(n_511), .Y(n_509) );
OAI21xp5_ASAP7_75t_L g559 ( .A1(n_131), .A2(n_560), .B(n_561), .Y(n_559) );
NAND2x1p5_ASAP7_75t_L g131 ( .A(n_132), .B(n_136), .Y(n_131) );
AND2x4_ASAP7_75t_L g170 ( .A(n_132), .B(n_136), .Y(n_170) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
INVx1_ASAP7_75t_L g150 ( .A(n_133), .Y(n_150) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g141 ( .A(n_134), .Y(n_141) );
INVx1_ASAP7_75t_L g269 ( .A(n_134), .Y(n_269) );
INVx1_ASAP7_75t_L g142 ( .A(n_135), .Y(n_142) );
INVx3_ASAP7_75t_L g146 ( .A(n_135), .Y(n_146) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_135), .Y(n_148) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_135), .Y(n_179) );
INVx1_ASAP7_75t_L g501 ( .A(n_135), .Y(n_501) );
BUFx3_ASAP7_75t_L g151 ( .A(n_136), .Y(n_151) );
INVx4_ASAP7_75t_SL g180 ( .A(n_136), .Y(n_180) );
INVx5_ASAP7_75t_L g173 ( .A(n_140), .Y(n_173) );
AND2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
BUFx3_ASAP7_75t_L g196 ( .A(n_141), .Y(n_196) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_141), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_145), .B(n_147), .C(n_149), .Y(n_143) );
OAI22xp33_ASAP7_75t_L g175 ( .A1(n_145), .A2(n_176), .B1(n_177), .B2(n_178), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_L g512 ( .A1(n_145), .A2(n_513), .B(n_514), .C(n_515), .Y(n_512) );
INVx5_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_146), .B(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_146), .B(n_483), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_146), .B(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g209 ( .A(n_148), .Y(n_209) );
INVx4_ASAP7_75t_L g251 ( .A(n_148), .Y(n_251) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_150), .B(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g183 ( .A(n_152), .Y(n_183) );
OA21x2_ASAP7_75t_L g204 ( .A1(n_152), .A2(n_205), .B(n_212), .Y(n_204) );
INVx1_ASAP7_75t_L g217 ( .A(n_152), .Y(n_217) );
OA21x2_ASAP7_75t_L g544 ( .A1(n_152), .A2(n_545), .B(n_551), .Y(n_544) );
AND2x2_ASAP7_75t_SL g152 ( .A(n_153), .B(n_154), .Y(n_152) );
AND2x2_ASAP7_75t_L g161 ( .A(n_153), .B(n_154), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
AO21x2_ASAP7_75t_L g185 ( .A1(n_159), .A2(n_186), .B(n_198), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_159), .B(n_225), .Y(n_224) );
INVx3_ASAP7_75t_L g237 ( .A(n_159), .Y(n_237) );
NOR2xp33_ASAP7_75t_SL g528 ( .A(n_159), .B(n_529), .Y(n_528) );
INVx4_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_160), .Y(n_228) );
OA21x2_ASAP7_75t_L g496 ( .A1(n_160), .A2(n_497), .B(n_504), .Y(n_496) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g167 ( .A(n_161), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_162), .B(n_349), .Y(n_361) );
AND2x2_ASAP7_75t_L g162 ( .A(n_163), .B(n_184), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_163), .B(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g299 ( .A(n_163), .B(n_184), .Y(n_299) );
BUFx3_ASAP7_75t_L g307 ( .A(n_163), .Y(n_307) );
OR2x2_ASAP7_75t_L g328 ( .A(n_163), .B(n_203), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_163), .B(n_349), .Y(n_439) );
OA21x2_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_168), .B(n_181), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AO21x2_ASAP7_75t_L g241 ( .A1(n_165), .A2(n_242), .B(n_243), .Y(n_241) );
AO21x2_ASAP7_75t_L g558 ( .A1(n_165), .A2(n_559), .B(n_565), .Y(n_558) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AOI21xp5_ASAP7_75t_SL g522 ( .A1(n_166), .A2(n_523), .B(n_524), .Y(n_522) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_167), .A2(n_488), .B(n_494), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_167), .B(n_495), .Y(n_494) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_167), .A2(n_509), .B(n_516), .Y(n_508) );
INVx1_ASAP7_75t_L g242 ( .A(n_168), .Y(n_242) );
BUFx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_SL g171 ( .A1(n_172), .A2(n_173), .B(n_174), .C(n_180), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_SL g206 ( .A1(n_173), .A2(n_180), .B(n_207), .C(n_208), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_SL g230 ( .A1(n_173), .A2(n_180), .B(n_231), .C(n_232), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g248 ( .A1(n_173), .A2(n_180), .B(n_249), .C(n_250), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_SL g263 ( .A1(n_173), .A2(n_180), .B(n_264), .C(n_265), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_173), .A2(n_180), .B(n_480), .C(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g498 ( .A1(n_173), .A2(n_180), .B(n_499), .C(n_500), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_L g546 ( .A1(n_173), .A2(n_180), .B(n_547), .C(n_548), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_178), .B(n_234), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_178), .B(n_267), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_178), .B(n_550), .Y(n_549) );
INVx4_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g192 ( .A(n_179), .Y(n_192) );
OAI22xp5_ASAP7_75t_SL g490 ( .A1(n_179), .A2(n_192), .B1(n_491), .B2(n_492), .Y(n_490) );
INVx1_ASAP7_75t_L g197 ( .A(n_180), .Y(n_197) );
INVx1_ASAP7_75t_L g243 ( .A(n_181), .Y(n_243) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_183), .B(n_199), .Y(n_198) );
AO21x2_ASAP7_75t_L g533 ( .A1(n_183), .A2(n_534), .B(n_541), .Y(n_533) );
AND2x2_ASAP7_75t_L g244 ( .A(n_184), .B(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g292 ( .A(n_184), .Y(n_292) );
AND2x2_ASAP7_75t_L g355 ( .A(n_184), .B(n_246), .Y(n_355) );
AOI221xp5_ASAP7_75t_L g357 ( .A1(n_184), .A2(n_358), .B1(n_360), .B2(n_362), .C(n_363), .Y(n_357) );
AND2x2_ASAP7_75t_L g371 ( .A(n_184), .B(n_241), .Y(n_371) );
AND2x2_ASAP7_75t_L g397 ( .A(n_184), .B(n_281), .Y(n_397) );
INVx2_ASAP7_75t_SL g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g277 ( .A(n_185), .B(n_246), .Y(n_277) );
BUFx2_ASAP7_75t_L g411 ( .A(n_185), .Y(n_411) );
O2A1O1Ixp33_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_193), .C(n_194), .Y(n_189) );
O2A1O1Ixp5_ASAP7_75t_L g221 ( .A1(n_191), .A2(n_194), .B(n_222), .C(n_223), .Y(n_221) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_194), .A2(n_526), .B(n_527), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_194), .A2(n_563), .B(n_564), .Y(n_562) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g235 ( .A(n_196), .Y(n_235) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
OAI32xp33_ASAP7_75t_L g377 ( .A1(n_201), .A2(n_338), .A3(n_352), .B1(n_378), .B2(n_379), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_202), .B(n_213), .Y(n_201) );
AND2x2_ASAP7_75t_L g318 ( .A(n_202), .B(n_260), .Y(n_318) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
OR2x2_ASAP7_75t_L g300 ( .A(n_203), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_203), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g372 ( .A(n_203), .B(n_260), .Y(n_372) );
AND2x2_ASAP7_75t_L g383 ( .A(n_203), .B(n_275), .Y(n_383) );
BUFx3_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
OR2x2_ASAP7_75t_L g284 ( .A(n_204), .B(n_261), .Y(n_284) );
AND2x2_ASAP7_75t_L g288 ( .A(n_204), .B(n_261), .Y(n_288) );
AND2x2_ASAP7_75t_L g323 ( .A(n_204), .B(n_274), .Y(n_323) );
AND2x2_ASAP7_75t_L g330 ( .A(n_204), .B(n_226), .Y(n_330) );
OAI211xp5_ASAP7_75t_L g335 ( .A1(n_204), .A2(n_281), .B(n_292), .C(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g389 ( .A(n_204), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_204), .B(n_215), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_213), .B(n_272), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_213), .B(n_288), .Y(n_378) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
OR2x2_ASAP7_75t_L g283 ( .A(n_214), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_226), .Y(n_214) );
AND2x2_ASAP7_75t_L g275 ( .A(n_215), .B(n_227), .Y(n_275) );
OR2x2_ASAP7_75t_L g290 ( .A(n_215), .B(n_227), .Y(n_290) );
AND2x2_ASAP7_75t_L g313 ( .A(n_215), .B(n_274), .Y(n_313) );
INVx1_ASAP7_75t_L g317 ( .A(n_215), .Y(n_317) );
AND2x2_ASAP7_75t_L g336 ( .A(n_215), .B(n_273), .Y(n_336) );
OAI22xp33_ASAP7_75t_L g346 ( .A1(n_215), .A2(n_301), .B1(n_347), .B2(n_348), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_215), .B(n_389), .Y(n_413) );
AND2x2_ASAP7_75t_L g428 ( .A(n_215), .B(n_288), .Y(n_428) );
INVx4_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
BUFx3_ASAP7_75t_L g258 ( .A(n_216), .Y(n_258) );
AND2x2_ASAP7_75t_L g302 ( .A(n_216), .B(n_227), .Y(n_302) );
AND2x2_ASAP7_75t_L g304 ( .A(n_216), .B(n_260), .Y(n_304) );
AND3x2_ASAP7_75t_L g366 ( .A(n_216), .B(n_330), .C(n_367), .Y(n_366) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_224), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_217), .B(n_517), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_217), .B(n_542), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_217), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g401 ( .A(n_226), .B(n_273), .Y(n_401) );
INVx1_ASAP7_75t_SL g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g260 ( .A(n_227), .B(n_261), .Y(n_260) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_227), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_227), .B(n_272), .Y(n_334) );
NAND3xp33_ASAP7_75t_L g441 ( .A(n_227), .B(n_313), .C(n_389), .Y(n_441) );
OA21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_236), .Y(n_227) );
OA21x2_ASAP7_75t_L g246 ( .A1(n_228), .A2(n_247), .B(n_256), .Y(n_246) );
OA21x2_ASAP7_75t_L g261 ( .A1(n_228), .A2(n_262), .B(n_270), .Y(n_261) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_237), .A2(n_478), .B(n_484), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_257), .B1(n_271), .B2(n_276), .Y(n_238) );
INVx1_ASAP7_75t_SL g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_244), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_241), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_SL g353 ( .A(n_241), .Y(n_353) );
OAI31xp33_ASAP7_75t_L g369 ( .A1(n_244), .A2(n_370), .A3(n_371), .B(n_372), .Y(n_369) );
AND2x2_ASAP7_75t_L g394 ( .A(n_244), .B(n_281), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_244), .B(n_307), .Y(n_440) );
AND2x2_ASAP7_75t_L g349 ( .A(n_245), .B(n_281), .Y(n_349) );
AND2x2_ASAP7_75t_L g410 ( .A(n_245), .B(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g280 ( .A(n_246), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g338 ( .A(n_246), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_251), .B(n_253), .Y(n_252) );
INVx3_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_255), .Y(n_539) );
OR2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
CKINVDCx16_ASAP7_75t_R g359 ( .A(n_258), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_259), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
AOI221x1_ASAP7_75t_SL g326 ( .A1(n_260), .A2(n_327), .B1(n_329), .B2(n_331), .C(n_333), .Y(n_326) );
INVx2_ASAP7_75t_L g274 ( .A(n_261), .Y(n_274) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_261), .Y(n_368) );
INVx2_ASAP7_75t_L g515 ( .A(n_268), .Y(n_515) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g356 ( .A(n_271), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_275), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_272), .B(n_289), .Y(n_381) );
INVx1_ASAP7_75t_SL g444 ( .A(n_272), .Y(n_444) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g362 ( .A(n_275), .B(n_288), .Y(n_362) );
INVx1_ASAP7_75t_L g430 ( .A(n_276), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_276), .B(n_359), .Y(n_443) );
INVx2_ASAP7_75t_SL g282 ( .A(n_277), .Y(n_282) );
AND2x2_ASAP7_75t_L g325 ( .A(n_277), .B(n_281), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_277), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_277), .B(n_352), .Y(n_379) );
AOI21xp33_ASAP7_75t_SL g278 ( .A1(n_279), .A2(n_282), .B(n_283), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_280), .B(n_352), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_280), .B(n_307), .Y(n_448) );
OR2x2_ASAP7_75t_L g320 ( .A(n_281), .B(n_299), .Y(n_320) );
AND2x2_ASAP7_75t_L g419 ( .A(n_281), .B(n_410), .Y(n_419) );
OAI22xp5_ASAP7_75t_SL g294 ( .A1(n_282), .A2(n_295), .B1(n_300), .B2(n_303), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_282), .B(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g342 ( .A(n_284), .B(n_290), .Y(n_342) );
INVx1_ASAP7_75t_L g406 ( .A(n_284), .Y(n_406) );
AOI311xp33_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_291), .A3(n_293), .B(n_294), .C(n_305), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
AOI221xp5_ASAP7_75t_L g432 ( .A1(n_289), .A2(n_421), .B1(n_433), .B2(n_436), .C(n_438), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_289), .B(n_444), .Y(n_446) );
INVx2_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g343 ( .A(n_291), .Y(n_343) );
AOI211xp5_ASAP7_75t_L g333 ( .A1(n_292), .A2(n_334), .B(n_335), .C(n_337), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
O2A1O1Ixp33_ASAP7_75t_SL g402 ( .A1(n_296), .A2(n_298), .B(n_403), .C(n_404), .Y(n_402) );
INVx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_297), .B(n_371), .Y(n_437) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
OAI221xp5_ASAP7_75t_L g319 ( .A1(n_300), .A2(n_320), .B1(n_321), .B2(n_324), .C(n_326), .Y(n_319) );
INVx1_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g322 ( .A(n_302), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g405 ( .A(n_302), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_306), .B(n_309), .Y(n_305) );
A2O1A1Ixp33_ASAP7_75t_L g363 ( .A1(n_306), .A2(n_364), .B(n_365), .C(n_369), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_307), .B(n_308), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_307), .B(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_307), .B(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVxp67_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g329 ( .A(n_313), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_317), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g431 ( .A(n_320), .Y(n_431) );
INVx1_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_323), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g358 ( .A(n_323), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_SL g435 ( .A(n_323), .Y(n_435) );
INVx1_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g376 ( .A(n_325), .B(n_352), .Y(n_376) );
INVx1_ASAP7_75t_SL g370 ( .A(n_332), .Y(n_370) );
INVx1_ASAP7_75t_L g347 ( .A(n_338), .Y(n_347) );
NAND3xp33_ASAP7_75t_SL g339 ( .A(n_340), .B(n_357), .C(n_373), .Y(n_339) );
AOI322xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_343), .A3(n_344), .B1(n_346), .B2(n_350), .C1(n_354), .C2(n_356), .Y(n_340) );
AOI211xp5_ASAP7_75t_L g393 ( .A1(n_341), .A2(n_394), .B(n_395), .C(n_402), .Y(n_393) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_344), .A2(n_365), .B1(n_396), .B2(n_398), .Y(n_395) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g354 ( .A(n_352), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g391 ( .A(n_352), .B(n_392), .Y(n_391) );
AOI32xp33_ASAP7_75t_L g442 ( .A1(n_352), .A2(n_443), .A3(n_444), .B1(n_445), .B2(n_447), .Y(n_442) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g364 ( .A(n_355), .Y(n_364) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_355), .A2(n_408), .B1(n_412), .B2(n_414), .C(n_417), .Y(n_407) );
AND2x2_ASAP7_75t_L g421 ( .A(n_355), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g424 ( .A(n_359), .B(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g434 ( .A(n_359), .B(n_435), .Y(n_434) );
INVxp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
INVxp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g425 ( .A(n_368), .B(n_389), .Y(n_425) );
AOI211xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_376), .B(n_377), .C(n_380), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AOI21xp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_382), .B(n_384), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OAI211xp5_ASAP7_75t_SL g386 ( .A1(n_387), .A2(n_390), .B(n_393), .C(n_407), .Y(n_386) );
INVxp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_401), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g416 ( .A(n_413), .Y(n_416) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AOI21xp33_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_420), .B(n_423), .Y(n_417) );
INVx1_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI211xp5_ASAP7_75t_SL g426 ( .A1(n_427), .A2(n_429), .B(n_432), .C(n_442), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_428), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
INVx1_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AOI21xp33_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_440), .B(n_441), .Y(n_438) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_454), .Y(n_460) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AOI21xp33_ASAP7_75t_L g461 ( .A1(n_458), .A2(n_462), .B(n_757), .Y(n_461) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OAI22x1_ASAP7_75t_L g751 ( .A1(n_464), .A2(n_467), .B1(n_752), .B2(n_753), .Y(n_751) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVxp67_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g753 ( .A(n_471), .Y(n_753) );
BUFx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND3x1_ASAP7_75t_L g472 ( .A(n_473), .B(n_666), .C(n_711), .Y(n_472) );
NOR4xp25_ASAP7_75t_L g473 ( .A(n_474), .B(n_589), .C(n_630), .D(n_647), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_505), .B(n_519), .C(n_552), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_485), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_476), .B(n_506), .Y(n_505) );
NOR4xp25_ASAP7_75t_L g613 ( .A(n_476), .B(n_607), .C(n_614), .D(n_620), .Y(n_613) );
AND2x2_ASAP7_75t_L g686 ( .A(n_476), .B(n_575), .Y(n_686) );
AND2x2_ASAP7_75t_L g705 ( .A(n_476), .B(n_651), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_476), .B(n_700), .Y(n_714) );
AND2x2_ASAP7_75t_L g727 ( .A(n_476), .B(n_518), .Y(n_727) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_SL g572 ( .A(n_477), .Y(n_572) );
AND2x2_ASAP7_75t_L g579 ( .A(n_477), .B(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g629 ( .A(n_477), .B(n_486), .Y(n_629) );
AND2x2_ASAP7_75t_SL g640 ( .A(n_477), .B(n_575), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_477), .B(n_486), .Y(n_644) );
AND2x2_ASAP7_75t_L g653 ( .A(n_477), .B(n_578), .Y(n_653) );
BUFx2_ASAP7_75t_L g676 ( .A(n_477), .Y(n_676) );
AND2x2_ASAP7_75t_L g680 ( .A(n_477), .B(n_496), .Y(n_680) );
OR2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_496), .Y(n_485) );
AND2x2_ASAP7_75t_L g518 ( .A(n_486), .B(n_496), .Y(n_518) );
BUFx2_ASAP7_75t_L g582 ( .A(n_486), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_486), .A2(n_615), .B1(n_617), .B2(n_618), .Y(n_614) );
OR2x2_ASAP7_75t_L g636 ( .A(n_486), .B(n_508), .Y(n_636) );
AND2x2_ASAP7_75t_L g700 ( .A(n_486), .B(n_578), .Y(n_700) );
INVx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g568 ( .A(n_487), .B(n_508), .Y(n_568) );
AND2x2_ASAP7_75t_L g575 ( .A(n_487), .B(n_496), .Y(n_575) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_487), .Y(n_617) );
OR2x2_ASAP7_75t_L g652 ( .A(n_487), .B(n_507), .Y(n_652) );
INVx1_ASAP7_75t_L g571 ( .A(n_496), .Y(n_571) );
INVx3_ASAP7_75t_L g580 ( .A(n_496), .Y(n_580) );
BUFx2_ASAP7_75t_L g604 ( .A(n_496), .Y(n_604) );
AND2x2_ASAP7_75t_L g637 ( .A(n_496), .B(n_572), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_505), .A2(n_723), .B1(n_724), .B2(n_725), .Y(n_722) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_518), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_507), .B(n_580), .Y(n_584) );
INVx1_ASAP7_75t_L g612 ( .A(n_507), .Y(n_612) );
INVx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx3_ASAP7_75t_L g578 ( .A(n_508), .Y(n_578) );
INVx1_ASAP7_75t_L g590 ( .A(n_518), .Y(n_590) );
NAND2x1_ASAP7_75t_SL g519 ( .A(n_520), .B(n_530), .Y(n_519) );
AND2x2_ASAP7_75t_L g588 ( .A(n_520), .B(n_543), .Y(n_588) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_520), .Y(n_662) );
AND2x2_ASAP7_75t_L g689 ( .A(n_520), .B(n_609), .Y(n_689) );
AND2x2_ASAP7_75t_L g697 ( .A(n_520), .B(n_659), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_520), .B(n_555), .Y(n_724) );
INVx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g556 ( .A(n_521), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g573 ( .A(n_521), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g594 ( .A(n_521), .Y(n_594) );
INVx1_ASAP7_75t_L g600 ( .A(n_521), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_521), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g633 ( .A(n_521), .B(n_558), .Y(n_633) );
OR2x2_ASAP7_75t_L g671 ( .A(n_521), .B(n_626), .Y(n_671) );
AOI32xp33_ASAP7_75t_L g683 ( .A1(n_521), .A2(n_684), .A3(n_687), .B1(n_688), .B2(n_689), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_521), .B(n_659), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_521), .B(n_619), .Y(n_734) );
OR2x6_ASAP7_75t_L g521 ( .A(n_522), .B(n_528), .Y(n_521) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OR2x2_ASAP7_75t_L g645 ( .A(n_531), .B(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_543), .Y(n_531) );
INVx1_ASAP7_75t_L g607 ( .A(n_532), .Y(n_607) );
AND2x2_ASAP7_75t_L g609 ( .A(n_532), .B(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_532), .B(n_557), .Y(n_626) );
AND2x2_ASAP7_75t_L g659 ( .A(n_532), .B(n_635), .Y(n_659) );
AND2x2_ASAP7_75t_L g696 ( .A(n_532), .B(n_558), .Y(n_696) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g555 ( .A(n_533), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_533), .B(n_557), .Y(n_586) );
AND2x2_ASAP7_75t_L g593 ( .A(n_533), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g634 ( .A(n_533), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_540), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_538), .B(n_539), .Y(n_536) );
INVx2_ASAP7_75t_L g610 ( .A(n_543), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_543), .B(n_557), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_543), .B(n_601), .Y(n_682) );
INVx1_ASAP7_75t_L g704 ( .A(n_543), .Y(n_704) );
INVx1_ASAP7_75t_L g721 ( .A(n_543), .Y(n_721) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g574 ( .A(n_544), .B(n_557), .Y(n_574) );
AND2x2_ASAP7_75t_L g596 ( .A(n_544), .B(n_558), .Y(n_596) );
INVx1_ASAP7_75t_L g635 ( .A(n_544), .Y(n_635) );
AOI221x1_ASAP7_75t_SL g552 ( .A1(n_553), .A2(n_567), .B1(n_573), .B2(n_575), .C(n_576), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_553), .A2(n_640), .B1(n_707), .B2(n_708), .Y(n_706) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_556), .Y(n_553) );
AND2x2_ASAP7_75t_L g598 ( .A(n_554), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g693 ( .A(n_554), .B(n_573), .Y(n_693) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g649 ( .A(n_555), .B(n_574), .Y(n_649) );
INVx1_ASAP7_75t_L g661 ( .A(n_556), .Y(n_661) );
AND2x2_ASAP7_75t_L g672 ( .A(n_556), .B(n_659), .Y(n_672) );
AND2x2_ASAP7_75t_L g739 ( .A(n_556), .B(n_634), .Y(n_739) );
INVx2_ASAP7_75t_L g601 ( .A(n_557), .Y(n_601) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_568), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g691 ( .A(n_568), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_569), .B(n_652), .Y(n_655) );
INVx3_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_570), .A2(n_691), .B(n_736), .Y(n_735) );
AND2x4_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
NOR2xp33_ASAP7_75t_SL g713 ( .A(n_573), .B(n_599), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_574), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g665 ( .A(n_574), .B(n_593), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_574), .B(n_600), .Y(n_742) );
AND2x2_ASAP7_75t_L g611 ( .A(n_575), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g678 ( .A(n_575), .Y(n_678) );
AOI21xp33_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_581), .B(n_585), .Y(n_576) );
NAND2x1_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_578), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g627 ( .A(n_578), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_SL g639 ( .A(n_578), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_578), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g663 ( .A(n_579), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_579), .B(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_579), .B(n_582), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
AOI211xp5_ASAP7_75t_L g650 ( .A1(n_582), .A2(n_621), .B(n_651), .C(n_653), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_582), .A2(n_669), .B1(n_672), .B2(n_673), .C(n_677), .Y(n_668) );
AND2x2_ASAP7_75t_L g664 ( .A(n_583), .B(n_617), .Y(n_664) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g624 ( .A(n_588), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g695 ( .A(n_588), .B(n_696), .Y(n_695) );
OAI211xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B(n_597), .C(n_622), .Y(n_589) );
NAND3xp33_ASAP7_75t_SL g708 ( .A(n_590), .B(n_709), .C(n_710), .Y(n_708) );
OR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_595), .Y(n_591) );
OR2x2_ASAP7_75t_L g681 ( .A(n_592), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AOI221xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_602), .B1(n_605), .B2(n_611), .C(n_613), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_599), .B(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_599), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g621 ( .A(n_604), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_604), .A2(n_661), .B1(n_662), .B2(n_663), .Y(n_660) );
OR2x2_ASAP7_75t_L g741 ( .A(n_604), .B(n_652), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_606), .B(n_608), .Y(n_605) );
INVxp67_ASAP7_75t_L g715 ( .A(n_607), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_609), .B(n_730), .Y(n_729) );
INVxp67_ASAP7_75t_L g616 ( .A(n_610), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_612), .B(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_612), .B(n_659), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_612), .B(n_679), .Y(n_718) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_616), .Y(n_642) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OR2x2_ASAP7_75t_L g732 ( .A(n_621), .B(n_652), .Y(n_732) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_627), .Y(n_623) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_SL g710 ( .A(n_627), .Y(n_710) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OAI322xp33_ASAP7_75t_SL g630 ( .A1(n_631), .A2(n_636), .A3(n_637), .B1(n_638), .B2(n_641), .C1(n_643), .C2(n_645), .Y(n_630) );
OAI322xp33_ASAP7_75t_L g712 ( .A1(n_631), .A2(n_713), .A3(n_714), .B1(n_715), .B2(n_716), .C1(n_717), .C2(n_719), .Y(n_712) );
CKINVDCx16_ASAP7_75t_R g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx4_ASAP7_75t_L g646 ( .A(n_633), .Y(n_646) );
AND2x2_ASAP7_75t_L g707 ( .A(n_633), .B(n_659), .Y(n_707) );
AND2x2_ASAP7_75t_L g720 ( .A(n_633), .B(n_721), .Y(n_720) );
CKINVDCx16_ASAP7_75t_R g731 ( .A(n_636), .Y(n_731) );
INVx1_ASAP7_75t_L g709 ( .A(n_637), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
OR2x2_ASAP7_75t_L g643 ( .A(n_639), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g726 ( .A(n_639), .B(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_639), .B(n_680), .Y(n_737) );
OR2x2_ASAP7_75t_L g670 ( .A(n_642), .B(n_671), .Y(n_670) );
INVxp33_ASAP7_75t_L g687 ( .A(n_642), .Y(n_687) );
OAI221xp5_ASAP7_75t_SL g647 ( .A1(n_646), .A2(n_648), .B1(n_650), .B2(n_654), .C(n_656), .Y(n_647) );
NOR2xp67_ASAP7_75t_L g703 ( .A(n_646), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g730 ( .A(n_646), .Y(n_730) );
INVx1_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
INVx3_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
AOI322xp5_ASAP7_75t_L g694 ( .A1(n_653), .A2(n_678), .A3(n_695), .B1(n_697), .B2(n_698), .C1(n_701), .C2(n_705), .Y(n_694) );
INVxp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_660), .B1(n_664), .B2(n_665), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_690), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_668), .B(n_683), .Y(n_667) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_671), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
NAND2xp33_ASAP7_75t_SL g688 ( .A(n_674), .B(n_685), .Y(n_688) );
INVx1_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
OAI322xp33_ASAP7_75t_L g728 ( .A1(n_676), .A2(n_729), .A3(n_731), .B1(n_732), .B2(n_733), .C1(n_735), .C2(n_738), .Y(n_728) );
AOI21xp33_ASAP7_75t_SL g677 ( .A1(n_678), .A2(n_679), .B(n_681), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_686), .B(n_734), .Y(n_743) );
OAI211xp5_ASAP7_75t_SL g690 ( .A1(n_691), .A2(n_692), .B(n_694), .C(n_706), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NOR4xp25_ASAP7_75t_L g711 ( .A(n_712), .B(n_722), .C(n_728), .D(n_740), .Y(n_711) );
INVxp67_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
INVxp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
CKINVDCx14_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
OAI21xp5_ASAP7_75t_SL g740 ( .A1(n_741), .A2(n_742), .B(n_743), .Y(n_740) );
CKINVDCx16_ASAP7_75t_R g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
INVx3_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
endmodule