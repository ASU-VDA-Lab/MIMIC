module fake_jpeg_29951_n_77 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_77);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_77;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_37),
.Y(n_42)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_34),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_28),
.A2(n_31),
.B1(n_27),
.B2(n_32),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_36),
.B1(n_38),
.B2(n_3),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_28),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_0),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_14),
.B1(n_22),
.B2(n_21),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_29),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_29),
.B1(n_32),
.B2(n_26),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_48),
.B1(n_5),
.B2(n_6),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_12),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_44),
.B(n_47),
.Y(n_50)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_3),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_4),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_49),
.Y(n_56)
);

OR2x6_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_16),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_10),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_45),
.B1(n_8),
.B2(n_9),
.Y(n_57)
);

AO22x1_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_53),
.B1(n_52),
.B2(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_56),
.B(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_58),
.B(n_59),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_11),
.C(n_19),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_62),
.C(n_61),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_51),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_51),
.A2(n_17),
.B(n_18),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_51),
.B(n_23),
.Y(n_65)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_68),
.C(n_59),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_61),
.B(n_62),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_64),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_71),
.B1(n_70),
.B2(n_69),
.Y(n_73)
);

AOI21x1_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_69),
.B(n_70),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_70),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_71),
.Y(n_77)
);


endmodule