module fake_jpeg_22447_n_230 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_230);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_37),
.B(n_40),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_0),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_44),
.Y(n_57)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_19),
.B(n_1),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_40),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_35),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_54),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_20),
.B1(n_19),
.B2(n_25),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_52),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_101)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_58),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_20),
.B1(n_19),
.B2(n_25),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_46),
.A2(n_25),
.B1(n_24),
.B2(n_30),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_24),
.B1(n_30),
.B2(n_29),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_69),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_24),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_70),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_41),
.A2(n_30),
.B1(n_23),
.B2(n_29),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_66),
.B1(n_71),
.B2(n_31),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_21),
.B1(n_23),
.B2(n_29),
.Y(n_66)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_32),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_41),
.A2(n_21),
.B1(n_23),
.B2(n_34),
.Y(n_71)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_74),
.B(n_81),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_41),
.B1(n_39),
.B2(n_38),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_75),
.A2(n_76),
.B1(n_49),
.B2(n_50),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_39),
.B1(n_38),
.B2(n_32),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_82),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_78),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_36),
.C(n_34),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_80),
.B(n_1),
.Y(n_123)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_33),
.Y(n_83)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_33),
.Y(n_84)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_86),
.Y(n_105)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_88),
.Y(n_115)
);

NAND2xp33_ASAP7_75t_SL g88 ( 
.A(n_58),
.B(n_32),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_31),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_93),
.Y(n_114)
);

NOR2x1_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_17),
.Y(n_90)
);

NOR3xp33_ASAP7_75t_SL g110 ( 
.A(n_90),
.B(n_27),
.C(n_18),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_64),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_28),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_95),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_28),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_97),
.Y(n_118)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_99),
.Y(n_120)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_36),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_72),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_107),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_93),
.B(n_27),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_106),
.B(n_18),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_17),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_91),
.B(n_50),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_100),
.C(n_88),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_116),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_111),
.A2(n_86),
.B1(n_77),
.B2(n_78),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_67),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_96),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_50),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_81),
.B(n_75),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_49),
.B1(n_55),
.B2(n_51),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_122),
.A2(n_101),
.B1(n_76),
.B2(n_49),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_103),
.Y(n_147)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_92),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_97),
.C(n_113),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_131),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_96),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_74),
.Y(n_132)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_90),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_133),
.B(n_146),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_144),
.B1(n_145),
.B2(n_118),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_135),
.A2(n_148),
.B(n_122),
.Y(n_157)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

BUFx24_ASAP7_75t_SL g137 ( 
.A(n_106),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_142),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_138),
.B(n_141),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_119),
.A2(n_75),
.B1(n_92),
.B2(n_80),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_143),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_115),
.A2(n_75),
.B1(n_85),
.B2(n_82),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_123),
.Y(n_155)
);

AND2x4_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_97),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_149),
.A2(n_112),
.B1(n_124),
.B2(n_125),
.Y(n_160)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_152),
.B(n_161),
.Y(n_179)
);

OAI32xp33_ASAP7_75t_L g153 ( 
.A1(n_131),
.A2(n_115),
.A3(n_102),
.B1(n_121),
.B2(n_111),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_139),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_169),
.C(n_127),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_157),
.A2(n_167),
.B(n_168),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_115),
.B1(n_112),
.B2(n_118),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_158),
.A2(n_159),
.B1(n_144),
.B2(n_148),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_160),
.A2(n_126),
.B(n_138),
.Y(n_180)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_SL g165 ( 
.A1(n_133),
.A2(n_110),
.A3(n_107),
.B1(n_125),
.B2(n_108),
.C1(n_116),
.C2(n_13),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_16),
.C(n_14),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_107),
.B(n_116),
.Y(n_167)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_129),
.A2(n_108),
.B(n_2),
.C(n_3),
.Y(n_168)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_181),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_172),
.A2(n_185),
.B1(n_154),
.B2(n_162),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_173),
.A2(n_177),
.B1(n_180),
.B2(n_163),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_128),
.Y(n_174)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_174),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_176),
.C(n_182),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_147),
.C(n_128),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_154),
.A2(n_134),
.B1(n_149),
.B2(n_130),
.Y(n_177)
);

OAI321xp33_ASAP7_75t_L g178 ( 
.A1(n_153),
.A2(n_159),
.A3(n_167),
.B1(n_152),
.B2(n_151),
.C(n_150),
.Y(n_178)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_168),
.Y(n_181)
);

A2O1A1O1Ixp25_ASAP7_75t_L g182 ( 
.A1(n_157),
.A2(n_143),
.B(n_142),
.C(n_141),
.D(n_6),
.Y(n_182)
);

NOR2x1_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_156),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_161),
.A2(n_126),
.B(n_113),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_16),
.C(n_13),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_12),
.C(n_2),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_185),
.Y(n_187)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_195),
.Y(n_200)
);

O2A1O1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_192),
.A2(n_193),
.B(n_8),
.C(n_9),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_172),
.A2(n_164),
.B1(n_163),
.B2(n_155),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_194),
.A2(n_179),
.B1(n_173),
.B2(n_183),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_166),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_8),
.Y(n_207)
);

NOR2x1_ASAP7_75t_R g198 ( 
.A(n_183),
.B(n_1),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_5),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_175),
.C(n_176),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_204),
.C(n_189),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_188),
.A2(n_181),
.B1(n_180),
.B2(n_171),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_201),
.A2(n_208),
.B1(n_197),
.B2(n_191),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_203),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_177),
.C(n_186),
.Y(n_204)
);

OAI21x1_ASAP7_75t_L g205 ( 
.A1(n_192),
.A2(n_182),
.B(n_12),
.Y(n_205)
);

A2O1A1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_205),
.A2(n_206),
.B(n_190),
.C(n_195),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_196),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_188),
.Y(n_209)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_209),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_210),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_202),
.A2(n_194),
.B(n_198),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_213),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_215),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_211),
.A2(n_208),
.B1(n_201),
.B2(n_199),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_209),
.C(n_204),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_223),
.C(n_224),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_212),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_219),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_220),
.A2(n_206),
.B(n_10),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_8),
.C(n_10),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_222),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_226),
.A2(n_227),
.B(n_11),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_225),
.A2(n_217),
.B1(n_10),
.B2(n_11),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_228),
.B(n_229),
.Y(n_230)
);


endmodule