module real_aes_9084_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g182 ( .A1(n_0), .A2(n_183), .B(n_184), .C(n_188), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_1), .B(n_177), .Y(n_190) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_2), .B(n_93), .C(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g126 ( .A(n_2), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_3), .B(n_162), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_4), .A2(n_171), .B(n_477), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_5), .A2(n_151), .B(n_168), .C(n_521), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_6), .A2(n_171), .B(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_7), .B(n_177), .Y(n_483) );
AO21x2_ASAP7_75t_L g264 ( .A1(n_8), .A2(n_143), .B(n_265), .Y(n_264) );
AND2x6_ASAP7_75t_L g168 ( .A(n_9), .B(n_169), .Y(n_168) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_10), .A2(n_151), .B(n_168), .C(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g574 ( .A(n_11), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_12), .B(n_108), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_12), .B(n_40), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_13), .B(n_187), .Y(n_523) );
INVx1_ASAP7_75t_L g148 ( .A(n_14), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_15), .B(n_162), .Y(n_271) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_16), .A2(n_163), .B(n_532), .C(n_534), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_17), .B(n_177), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_18), .B(n_205), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_19), .A2(n_151), .B(n_197), .C(n_204), .Y(n_196) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_20), .A2(n_186), .B(n_239), .C(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_21), .B(n_187), .Y(n_505) );
AOI222xp33_ASAP7_75t_L g452 ( .A1(n_22), .A2(n_453), .B1(n_723), .B2(n_724), .C1(n_733), .C2(n_737), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_23), .B(n_187), .Y(n_472) );
CKINVDCx16_ASAP7_75t_R g501 ( .A(n_24), .Y(n_501) );
INVx1_ASAP7_75t_L g471 ( .A(n_25), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_26), .A2(n_151), .B(n_204), .C(n_268), .Y(n_267) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_27), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_28), .Y(n_519) );
INVx1_ASAP7_75t_L g495 ( .A(n_29), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_30), .A2(n_171), .B(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_31), .B(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g153 ( .A(n_32), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_33), .A2(n_166), .B(n_220), .C(n_221), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_34), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_35), .A2(n_186), .B(n_480), .C(n_482), .Y(n_479) );
INVxp67_ASAP7_75t_L g496 ( .A(n_36), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_37), .B(n_270), .Y(n_269) );
CKINVDCx14_ASAP7_75t_R g478 ( .A(n_38), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_39), .A2(n_151), .B(n_204), .C(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g108 ( .A(n_40), .Y(n_108) );
A2O1A1Ixp33_ASAP7_75t_L g571 ( .A1(n_41), .A2(n_188), .B(n_572), .C(n_573), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_42), .B(n_195), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_43), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_44), .B(n_162), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_45), .B(n_171), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_46), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_47), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_48), .A2(n_166), .B(n_220), .C(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g185 ( .A(n_49), .Y(n_185) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_50), .A2(n_67), .B1(n_130), .B2(n_131), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_50), .Y(n_131) );
INVx1_ASAP7_75t_L g249 ( .A(n_51), .Y(n_249) );
INVx1_ASAP7_75t_L g539 ( .A(n_52), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_53), .B(n_171), .Y(n_246) );
OAI22xp5_ASAP7_75t_SL g133 ( .A1(n_54), .A2(n_72), .B1(n_134), .B2(n_135), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_54), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g209 ( .A(n_55), .Y(n_209) );
CKINVDCx14_ASAP7_75t_R g570 ( .A(n_56), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_57), .A2(n_105), .B1(n_113), .B2(n_740), .Y(n_104) );
INVx1_ASAP7_75t_L g169 ( .A(n_58), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_59), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_60), .B(n_177), .Y(n_262) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_61), .A2(n_158), .B(n_203), .C(n_260), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_62), .A2(n_71), .B1(n_730), .B2(n_731), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_62), .Y(n_730) );
INVx1_ASAP7_75t_L g147 ( .A(n_63), .Y(n_147) );
INVx1_ASAP7_75t_SL g481 ( .A(n_64), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_65), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_66), .B(n_162), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_67), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_67), .B(n_177), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_68), .B(n_163), .Y(n_236) );
INVx1_ASAP7_75t_L g504 ( .A(n_69), .Y(n_504) );
CKINVDCx16_ASAP7_75t_R g180 ( .A(n_70), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_71), .Y(n_731) );
INVx1_ASAP7_75t_L g135 ( .A(n_72), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_73), .B(n_199), .Y(n_198) );
A2O1A1Ixp33_ASAP7_75t_L g150 ( .A1(n_74), .A2(n_151), .B(n_156), .C(n_166), .Y(n_150) );
CKINVDCx16_ASAP7_75t_R g258 ( .A(n_75), .Y(n_258) );
INVx1_ASAP7_75t_L g112 ( .A(n_76), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_77), .A2(n_171), .B(n_569), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_78), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_79), .A2(n_171), .B(n_529), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_80), .A2(n_195), .B(n_491), .Y(n_490) );
CKINVDCx16_ASAP7_75t_R g468 ( .A(n_81), .Y(n_468) );
INVx1_ASAP7_75t_L g530 ( .A(n_82), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_83), .A2(n_727), .B1(n_728), .B2(n_729), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_83), .Y(n_727) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_84), .B(n_201), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_85), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_86), .A2(n_171), .B(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g533 ( .A(n_87), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g724 ( .A1(n_88), .A2(n_725), .B1(n_726), .B2(n_732), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_88), .Y(n_725) );
INVx2_ASAP7_75t_L g145 ( .A(n_89), .Y(n_145) );
INVx1_ASAP7_75t_L g522 ( .A(n_90), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_91), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_92), .B(n_187), .Y(n_237) );
OR2x2_ASAP7_75t_L g123 ( .A(n_93), .B(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g457 ( .A(n_93), .B(n_125), .Y(n_457) );
INVx2_ASAP7_75t_L g722 ( .A(n_93), .Y(n_722) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_94), .A2(n_151), .B(n_166), .C(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_95), .B(n_171), .Y(n_218) );
INVx1_ASAP7_75t_L g222 ( .A(n_96), .Y(n_222) );
INVxp67_ASAP7_75t_L g261 ( .A(n_97), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_98), .B(n_143), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_99), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g157 ( .A(n_100), .Y(n_157) );
INVx1_ASAP7_75t_L g232 ( .A(n_101), .Y(n_232) );
INVx2_ASAP7_75t_L g542 ( .A(n_102), .Y(n_542) );
AND2x2_ASAP7_75t_L g251 ( .A(n_103), .B(n_207), .Y(n_251) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx6p67_ASAP7_75t_R g741 ( .A(n_106), .Y(n_741) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OA21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_119), .B(n_451), .Y(n_113) );
BUFx2_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_115), .B(n_448), .C(n_452), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_128), .B(n_448), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_SL g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_123), .Y(n_450) );
NOR2x2_ASAP7_75t_L g739 ( .A(n_124), .B(n_722), .Y(n_739) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g721 ( .A(n_125), .B(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
AOI22xp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_132), .B1(n_446), .B2(n_447), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_129), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_132), .Y(n_447) );
XNOR2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_136), .Y(n_132) );
INVx1_ASAP7_75t_L g454 ( .A(n_136), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_136), .A2(n_459), .B1(n_734), .B2(n_735), .Y(n_733) );
OR3x1_ASAP7_75t_L g136 ( .A(n_137), .B(n_354), .C(n_403), .Y(n_136) );
NAND5xp2_ASAP7_75t_L g137 ( .A(n_138), .B(n_288), .C(n_317), .D(n_325), .E(n_340), .Y(n_137) );
O2A1O1Ixp33_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_211), .B(n_227), .C(n_272), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g139 ( .A(n_140), .B(n_191), .Y(n_139) );
AND2x2_ASAP7_75t_L g283 ( .A(n_140), .B(n_280), .Y(n_283) );
AND2x2_ASAP7_75t_L g316 ( .A(n_140), .B(n_192), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_140), .B(n_215), .Y(n_409) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_176), .Y(n_140) );
INVx2_ASAP7_75t_L g214 ( .A(n_141), .Y(n_214) );
BUFx2_ASAP7_75t_L g383 ( .A(n_141), .Y(n_383) );
AO21x2_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_149), .B(n_174), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_142), .B(n_175), .Y(n_174) );
INVx3_ASAP7_75t_L g177 ( .A(n_142), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_142), .B(n_226), .Y(n_225) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_142), .A2(n_231), .B(n_241), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_142), .B(n_474), .Y(n_473) );
AO21x2_ASAP7_75t_L g499 ( .A1(n_142), .A2(n_500), .B(n_507), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_142), .B(n_525), .Y(n_524) );
INVx4_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_143), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_143), .A2(n_266), .B(n_267), .Y(n_265) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g243 ( .A(n_144), .Y(n_243) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AND2x2_ASAP7_75t_SL g207 ( .A(n_145), .B(n_146), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_150), .B(n_170), .Y(n_149) );
INVx5_ASAP7_75t_L g181 ( .A(n_151), .Y(n_181) );
AND2x6_ASAP7_75t_L g151 ( .A(n_152), .B(n_154), .Y(n_151) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_152), .Y(n_165) );
BUFx3_ASAP7_75t_L g189 ( .A(n_152), .Y(n_189) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g173 ( .A(n_153), .Y(n_173) );
INVx1_ASAP7_75t_L g240 ( .A(n_153), .Y(n_240) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_155), .Y(n_160) );
INVx3_ASAP7_75t_L g163 ( .A(n_155), .Y(n_163) );
AND2x2_ASAP7_75t_L g172 ( .A(n_155), .B(n_173), .Y(n_172) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_155), .Y(n_187) );
INVx1_ASAP7_75t_L g270 ( .A(n_155), .Y(n_270) );
O2A1O1Ixp33_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_161), .C(n_164), .Y(n_156) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
OAI22xp33_ASAP7_75t_L g494 ( .A1(n_159), .A2(n_162), .B1(n_495), .B2(n_496), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_159), .B(n_533), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_159), .B(n_542), .Y(n_541) );
INVx4_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g199 ( .A(n_160), .Y(n_199) );
INVx2_ASAP7_75t_L g183 ( .A(n_162), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_162), .B(n_261), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_162), .A2(n_202), .B(n_471), .C(n_472), .Y(n_470) );
INVx5_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_163), .B(n_574), .Y(n_573) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx3_ASAP7_75t_L g482 ( .A(n_165), .Y(n_482) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
O2A1O1Ixp33_ASAP7_75t_SL g179 ( .A1(n_167), .A2(n_180), .B(n_181), .C(n_182), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_L g257 ( .A1(n_167), .A2(n_181), .B(n_258), .C(n_259), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g477 ( .A1(n_167), .A2(n_181), .B(n_478), .C(n_479), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_SL g491 ( .A1(n_167), .A2(n_181), .B(n_492), .C(n_493), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_SL g529 ( .A1(n_167), .A2(n_181), .B(n_530), .C(n_531), .Y(n_529) );
O2A1O1Ixp33_ASAP7_75t_SL g538 ( .A1(n_167), .A2(n_181), .B(n_539), .C(n_540), .Y(n_538) );
O2A1O1Ixp33_ASAP7_75t_SL g569 ( .A1(n_167), .A2(n_181), .B(n_570), .C(n_571), .Y(n_569) );
INVx4_ASAP7_75t_SL g167 ( .A(n_168), .Y(n_167) );
AND2x4_ASAP7_75t_L g171 ( .A(n_168), .B(n_172), .Y(n_171) );
BUFx3_ASAP7_75t_L g204 ( .A(n_168), .Y(n_204) );
NAND2x1p5_ASAP7_75t_L g233 ( .A(n_168), .B(n_172), .Y(n_233) );
BUFx2_ASAP7_75t_L g195 ( .A(n_171), .Y(n_195) );
INVx1_ASAP7_75t_L g203 ( .A(n_173), .Y(n_203) );
AND2x2_ASAP7_75t_L g191 ( .A(n_176), .B(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g281 ( .A(n_176), .Y(n_281) );
AND2x2_ASAP7_75t_L g367 ( .A(n_176), .B(n_280), .Y(n_367) );
AND2x2_ASAP7_75t_L g422 ( .A(n_176), .B(n_214), .Y(n_422) );
OA21x2_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_190), .Y(n_176) );
INVx2_ASAP7_75t_L g220 ( .A(n_181), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_186), .B(n_481), .Y(n_480) );
INVx4_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g572 ( .A(n_187), .Y(n_572) );
INVx2_ASAP7_75t_L g506 ( .A(n_188), .Y(n_506) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_189), .Y(n_224) );
INVx1_ASAP7_75t_L g534 ( .A(n_189), .Y(n_534) );
INVx1_ASAP7_75t_L g339 ( .A(n_191), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_191), .B(n_215), .Y(n_386) );
INVx5_ASAP7_75t_L g280 ( .A(n_192), .Y(n_280) );
AND2x4_ASAP7_75t_L g301 ( .A(n_192), .B(n_281), .Y(n_301) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_192), .Y(n_323) );
AND2x2_ASAP7_75t_L g398 ( .A(n_192), .B(n_383), .Y(n_398) );
AND2x2_ASAP7_75t_L g401 ( .A(n_192), .B(n_216), .Y(n_401) );
OR2x6_ASAP7_75t_L g192 ( .A(n_193), .B(n_208), .Y(n_192) );
AOI21xp5_ASAP7_75t_SL g193 ( .A1(n_194), .A2(n_196), .B(n_205), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_200), .B(n_202), .Y(n_197) );
INVx2_ASAP7_75t_L g201 ( .A(n_199), .Y(n_201) );
O2A1O1Ixp33_ASAP7_75t_L g221 ( .A1(n_201), .A2(n_222), .B(n_223), .C(n_224), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g248 ( .A1(n_201), .A2(n_224), .B(n_249), .C(n_250), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_L g503 ( .A1(n_201), .A2(n_504), .B(n_505), .C(n_506), .Y(n_503) );
O2A1O1Ixp5_ASAP7_75t_L g521 ( .A1(n_201), .A2(n_506), .B(n_522), .C(n_523), .Y(n_521) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_203), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_206), .B(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g210 ( .A(n_207), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_207), .A2(n_218), .B(n_219), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_207), .A2(n_246), .B(n_247), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g467 ( .A1(n_207), .A2(n_233), .B(n_468), .C(n_469), .Y(n_467) );
OA21x2_ASAP7_75t_L g567 ( .A1(n_207), .A2(n_568), .B(n_575), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
AO21x2_ASAP7_75t_L g517 ( .A1(n_210), .A2(n_518), .B(n_524), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_211), .B(n_281), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_211), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_SL g211 ( .A(n_212), .Y(n_211) );
OR2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_215), .Y(n_212) );
AND2x2_ASAP7_75t_L g306 ( .A(n_213), .B(n_281), .Y(n_306) );
AND2x2_ASAP7_75t_L g324 ( .A(n_213), .B(n_216), .Y(n_324) );
INVx1_ASAP7_75t_L g344 ( .A(n_213), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_213), .B(n_280), .Y(n_389) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_213), .Y(n_431) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_214), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_215), .B(n_279), .Y(n_278) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_215), .Y(n_333) );
O2A1O1Ixp33_ASAP7_75t_L g336 ( .A1(n_215), .A2(n_276), .B(n_337), .C(n_339), .Y(n_336) );
AND2x2_ASAP7_75t_L g343 ( .A(n_215), .B(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g352 ( .A(n_215), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g356 ( .A(n_215), .B(n_280), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_215), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g371 ( .A(n_215), .B(n_281), .Y(n_371) );
AND2x2_ASAP7_75t_L g421 ( .A(n_215), .B(n_422), .Y(n_421) );
INVx5_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
BUFx2_ASAP7_75t_L g285 ( .A(n_216), .Y(n_285) );
AND2x2_ASAP7_75t_L g326 ( .A(n_216), .B(n_279), .Y(n_326) );
AND2x2_ASAP7_75t_L g338 ( .A(n_216), .B(n_313), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_216), .B(n_367), .Y(n_385) );
OR2x6_ASAP7_75t_L g216 ( .A(n_217), .B(n_225), .Y(n_216) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_252), .Y(n_227) );
INVx1_ASAP7_75t_L g274 ( .A(n_228), .Y(n_274) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_244), .Y(n_228) );
OR2x2_ASAP7_75t_L g276 ( .A(n_229), .B(n_244), .Y(n_276) );
NAND3xp33_ASAP7_75t_L g282 ( .A(n_229), .B(n_283), .C(n_284), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_229), .B(n_254), .Y(n_293) );
OR2x2_ASAP7_75t_L g308 ( .A(n_229), .B(n_296), .Y(n_308) );
AND2x2_ASAP7_75t_L g314 ( .A(n_229), .B(n_263), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_229), .B(n_445), .Y(n_444) );
INVx5_ASAP7_75t_SL g229 ( .A(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_230), .B(n_254), .Y(n_311) );
AND2x2_ASAP7_75t_L g350 ( .A(n_230), .B(n_264), .Y(n_350) );
NAND2xp5_ASAP7_75t_SL g378 ( .A(n_230), .B(n_263), .Y(n_378) );
OR2x2_ASAP7_75t_L g381 ( .A(n_230), .B(n_263), .Y(n_381) );
OAI21xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_234), .Y(n_231) );
OAI21xp5_ASAP7_75t_L g500 ( .A1(n_233), .A2(n_501), .B(n_502), .Y(n_500) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_233), .A2(n_519), .B(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_238), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_238), .A2(n_269), .B(n_271), .Y(n_268) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
INVx2_ASAP7_75t_L g489 ( .A(n_243), .Y(n_489) );
INVx5_ASAP7_75t_SL g296 ( .A(n_244), .Y(n_296) );
OR2x2_ASAP7_75t_L g302 ( .A(n_244), .B(n_253), .Y(n_302) );
AND2x2_ASAP7_75t_L g318 ( .A(n_244), .B(n_319), .Y(n_318) );
AOI321xp33_ASAP7_75t_L g325 ( .A1(n_244), .A2(n_326), .A3(n_327), .B1(n_328), .B2(n_334), .C(n_336), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_244), .B(n_252), .Y(n_335) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_244), .Y(n_348) );
OR2x2_ASAP7_75t_L g395 ( .A(n_244), .B(n_293), .Y(n_395) );
AND2x2_ASAP7_75t_L g417 ( .A(n_244), .B(n_314), .Y(n_417) );
AND2x2_ASAP7_75t_L g436 ( .A(n_244), .B(n_254), .Y(n_436) );
OR2x6_ASAP7_75t_L g244 ( .A(n_245), .B(n_251), .Y(n_244) );
INVx1_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_263), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_254), .B(n_263), .Y(n_277) );
AND2x2_ASAP7_75t_L g286 ( .A(n_254), .B(n_287), .Y(n_286) );
INVx3_ASAP7_75t_L g313 ( .A(n_254), .Y(n_313) );
AND2x2_ASAP7_75t_L g319 ( .A(n_254), .B(n_314), .Y(n_319) );
INVxp67_ASAP7_75t_L g349 ( .A(n_254), .Y(n_349) );
OR2x2_ASAP7_75t_L g391 ( .A(n_254), .B(n_296), .Y(n_391) );
OA21x2_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_256), .B(n_262), .Y(n_254) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_255), .A2(n_476), .B(n_483), .Y(n_475) );
OA21x2_ASAP7_75t_L g527 ( .A1(n_255), .A2(n_528), .B(n_535), .Y(n_527) );
OA21x2_ASAP7_75t_L g536 ( .A1(n_255), .A2(n_537), .B(n_543), .Y(n_536) );
OR2x2_ASAP7_75t_L g273 ( .A(n_263), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_SL g287 ( .A(n_263), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_263), .B(n_276), .Y(n_320) );
AND2x2_ASAP7_75t_L g369 ( .A(n_263), .B(n_313), .Y(n_369) );
AND2x2_ASAP7_75t_L g407 ( .A(n_263), .B(n_296), .Y(n_407) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_264), .B(n_296), .Y(n_295) );
A2O1A1Ixp33_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_275), .B(n_278), .C(n_282), .Y(n_272) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_273), .A2(n_275), .B1(n_400), .B2(n_402), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_275), .A2(n_298), .B1(n_353), .B2(n_439), .Y(n_438) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
INVx1_ASAP7_75t_SL g427 ( .A(n_276), .Y(n_427) );
INVx1_ASAP7_75t_SL g327 ( .A(n_277), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_279), .B(n_299), .Y(n_329) );
AOI222xp33_ASAP7_75t_L g340 ( .A1(n_279), .A2(n_320), .B1(n_327), .B2(n_341), .C1(n_345), .C2(n_351), .Y(n_340) );
AND2x2_ASAP7_75t_L g430 ( .A(n_279), .B(n_431), .Y(n_430) );
AND2x4_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx2_ASAP7_75t_L g305 ( .A(n_280), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_280), .B(n_300), .Y(n_375) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_280), .Y(n_412) );
AND2x2_ASAP7_75t_L g415 ( .A(n_280), .B(n_324), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_280), .B(n_431), .Y(n_441) );
INVx1_ASAP7_75t_L g332 ( .A(n_281), .Y(n_332) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_281), .Y(n_360) );
O2A1O1Ixp33_ASAP7_75t_L g423 ( .A1(n_283), .A2(n_424), .B(n_425), .C(n_428), .Y(n_423) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
NAND3xp33_ASAP7_75t_L g346 ( .A(n_285), .B(n_347), .C(n_350), .Y(n_346) );
OR2x2_ASAP7_75t_L g374 ( .A(n_285), .B(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_285), .B(n_301), .Y(n_402) );
OR2x2_ASAP7_75t_L g307 ( .A(n_287), .B(n_308), .Y(n_307) );
AOI211xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_291), .B(n_297), .C(n_309), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_290), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g396 ( .A(n_291), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_292), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g310 ( .A(n_295), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_296), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g364 ( .A(n_296), .B(n_314), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_296), .B(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_296), .B(n_313), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_302), .B1(n_303), .B2(n_307), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_299), .B(n_371), .Y(n_370) );
BUFx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_301), .B(n_343), .Y(n_342) );
OAI221xp5_ASAP7_75t_SL g365 ( .A1(n_302), .A2(n_366), .B1(n_368), .B2(n_370), .C(n_372), .Y(n_365) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
AND2x2_ASAP7_75t_L g420 ( .A(n_305), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g433 ( .A(n_305), .B(n_422), .Y(n_433) );
INVx1_ASAP7_75t_L g353 ( .A(n_306), .Y(n_353) );
INVx1_ASAP7_75t_L g424 ( .A(n_307), .Y(n_424) );
AOI21xp5_ASAP7_75t_L g413 ( .A1(n_308), .A2(n_391), .B(n_414), .Y(n_413) );
AOI21xp33_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_312), .B(n_315), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OAI21xp5_ASAP7_75t_SL g317 ( .A1(n_318), .A2(n_320), .B(n_321), .Y(n_317) );
INVx1_ASAP7_75t_L g357 ( .A(n_318), .Y(n_357) );
AOI221xp5_ASAP7_75t_L g404 ( .A1(n_319), .A2(n_405), .B1(n_408), .B2(n_410), .C(n_413), .Y(n_404) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_327), .A2(n_417), .B1(n_418), .B2(n_420), .Y(n_416) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g393 ( .A(n_329), .Y(n_393) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NOR2xp67_ASAP7_75t_SL g331 ( .A(n_332), .B(n_333), .Y(n_331) );
AND2x2_ASAP7_75t_L g397 ( .A(n_333), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g362 ( .A(n_338), .Y(n_362) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_343), .B(n_367), .Y(n_419) );
INVxp67_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_349), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g435 ( .A(n_350), .B(n_436), .Y(n_435) );
AND2x4_ASAP7_75t_L g442 ( .A(n_350), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OAI211xp5_ASAP7_75t_SL g354 ( .A1(n_355), .A2(n_357), .B(n_358), .C(n_392), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AOI211xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_361), .B(n_365), .C(n_384), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_SL g445 ( .A(n_369), .Y(n_445) );
AND2x2_ASAP7_75t_L g382 ( .A(n_371), .B(n_383), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_376), .B1(n_380), .B2(n_382), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
OR2x2_ASAP7_75t_L g390 ( .A(n_378), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g443 ( .A(n_379), .Y(n_443) );
INVxp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AOI31xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_386), .A3(n_387), .B(n_390), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI211xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_394), .B(n_396), .C(n_399), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
CKINVDCx16_ASAP7_75t_R g400 ( .A(n_401), .Y(n_400) );
NAND5xp2_ASAP7_75t_L g403 ( .A(n_404), .B(n_416), .C(n_423), .D(n_437), .E(n_440), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_415), .A2(n_441), .B1(n_442), .B2(n_444), .Y(n_440) );
INVx1_ASAP7_75t_SL g439 ( .A(n_417), .Y(n_439) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AOI21xp33_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_432), .B(n_434), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVxp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OAI22xp5_ASAP7_75t_SL g453 ( .A1(n_454), .A2(n_455), .B1(n_458), .B2(n_721), .Y(n_453) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g734 ( .A(n_456), .Y(n_734) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OR3x1_ASAP7_75t_L g459 ( .A(n_460), .B(n_632), .C(n_679), .Y(n_459) );
NAND3xp33_ASAP7_75t_SL g460 ( .A(n_461), .B(n_578), .C(n_603), .Y(n_460) );
AOI221xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_516), .B1(n_544), .B2(n_547), .C(n_555), .Y(n_461) );
OAI21xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_484), .B(n_509), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_464), .B(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_464), .B(n_560), .Y(n_676) );
AND2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_475), .Y(n_464) );
AND2x2_ASAP7_75t_L g546 ( .A(n_465), .B(n_515), .Y(n_546) );
AND2x2_ASAP7_75t_L g596 ( .A(n_465), .B(n_514), .Y(n_596) );
AND2x2_ASAP7_75t_L g617 ( .A(n_465), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g622 ( .A(n_465), .B(n_589), .Y(n_622) );
OR2x2_ASAP7_75t_L g630 ( .A(n_465), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g702 ( .A(n_465), .B(n_498), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_465), .B(n_651), .Y(n_716) );
INVx3_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g561 ( .A(n_466), .B(n_475), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_466), .B(n_498), .Y(n_562) );
AND2x4_ASAP7_75t_L g584 ( .A(n_466), .B(n_515), .Y(n_584) );
AND2x2_ASAP7_75t_L g614 ( .A(n_466), .B(n_486), .Y(n_614) );
AND2x2_ASAP7_75t_L g623 ( .A(n_466), .B(n_613), .Y(n_623) );
AND2x2_ASAP7_75t_L g639 ( .A(n_466), .B(n_499), .Y(n_639) );
OR2x2_ASAP7_75t_L g648 ( .A(n_466), .B(n_631), .Y(n_648) );
AND2x2_ASAP7_75t_L g654 ( .A(n_466), .B(n_589), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_466), .B(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g668 ( .A(n_466), .B(n_511), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_466), .B(n_557), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g707 ( .A(n_466), .B(n_618), .Y(n_707) );
OR2x6_ASAP7_75t_L g466 ( .A(n_467), .B(n_473), .Y(n_466) );
INVx2_ASAP7_75t_L g515 ( .A(n_475), .Y(n_515) );
AND2x2_ASAP7_75t_L g613 ( .A(n_475), .B(n_498), .Y(n_613) );
AND2x2_ASAP7_75t_L g618 ( .A(n_475), .B(n_499), .Y(n_618) );
INVx1_ASAP7_75t_L g674 ( .A(n_475), .Y(n_674) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g583 ( .A(n_485), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_498), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_486), .B(n_546), .Y(n_545) );
BUFx3_ASAP7_75t_L g560 ( .A(n_486), .Y(n_560) );
OR2x2_ASAP7_75t_L g631 ( .A(n_486), .B(n_498), .Y(n_631) );
OR2x2_ASAP7_75t_L g692 ( .A(n_486), .B(n_599), .Y(n_692) );
OA21x2_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_490), .B(n_497), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_488), .A2(n_512), .B(n_513), .Y(n_511) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g512 ( .A(n_490), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_497), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_498), .B(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g651 ( .A(n_498), .B(n_511), .Y(n_651) );
INVx2_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g590 ( .A(n_499), .Y(n_590) );
INVx1_ASAP7_75t_SL g509 ( .A(n_510), .Y(n_509) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_510), .A2(n_696), .B1(n_700), .B2(n_703), .C(n_704), .Y(n_695) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_514), .Y(n_510) );
INVx1_ASAP7_75t_SL g558 ( .A(n_511), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_511), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g690 ( .A(n_511), .B(n_546), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_514), .B(n_560), .Y(n_682) );
AND2x2_ASAP7_75t_L g589 ( .A(n_515), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_SL g593 ( .A(n_516), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g629 ( .A(n_516), .B(n_599), .Y(n_629) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_526), .Y(n_516) );
AND2x2_ASAP7_75t_L g554 ( .A(n_517), .B(n_527), .Y(n_554) );
INVx4_ASAP7_75t_L g566 ( .A(n_517), .Y(n_566) );
BUFx3_ASAP7_75t_L g609 ( .A(n_517), .Y(n_609) );
AND3x2_ASAP7_75t_L g624 ( .A(n_517), .B(n_625), .C(n_626), .Y(n_624) );
AND2x2_ASAP7_75t_L g706 ( .A(n_526), .B(n_620), .Y(n_706) );
AND2x2_ASAP7_75t_L g714 ( .A(n_526), .B(n_599), .Y(n_714) );
INVx1_ASAP7_75t_SL g719 ( .A(n_526), .Y(n_719) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_536), .Y(n_526) );
INVx1_ASAP7_75t_SL g577 ( .A(n_527), .Y(n_577) );
AND2x2_ASAP7_75t_L g600 ( .A(n_527), .B(n_566), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_527), .B(n_550), .Y(n_602) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_527), .Y(n_642) );
OR2x2_ASAP7_75t_L g647 ( .A(n_527), .B(n_566), .Y(n_647) );
INVx2_ASAP7_75t_L g552 ( .A(n_536), .Y(n_552) );
AND2x2_ASAP7_75t_L g587 ( .A(n_536), .B(n_567), .Y(n_587) );
OR2x2_ASAP7_75t_L g607 ( .A(n_536), .B(n_567), .Y(n_607) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_536), .Y(n_627) );
INVx1_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
AOI21xp33_ASAP7_75t_L g677 ( .A1(n_545), .A2(n_586), .B(n_678), .Y(n_677) );
AOI322xp5_ASAP7_75t_L g713 ( .A1(n_547), .A2(n_557), .A3(n_584), .B1(n_714), .B2(n_715), .C1(n_717), .C2(n_720), .Y(n_713) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_553), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_549), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_550), .B(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g576 ( .A(n_551), .B(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g644 ( .A(n_552), .B(n_566), .Y(n_644) );
AND2x2_ASAP7_75t_L g711 ( .A(n_552), .B(n_567), .Y(n_711) );
INVx1_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g652 ( .A(n_554), .B(n_606), .Y(n_652) );
AOI31xp33_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_559), .A3(n_562), .B(n_563), .Y(n_555) );
AND2x2_ASAP7_75t_L g611 ( .A(n_557), .B(n_589), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_557), .B(n_581), .Y(n_693) );
AND2x2_ASAP7_75t_L g712 ( .A(n_557), .B(n_617), .Y(n_712) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_560), .B(n_589), .Y(n_601) );
NAND2x1p5_ASAP7_75t_L g635 ( .A(n_560), .B(n_618), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_560), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_560), .B(n_702), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_561), .B(n_618), .Y(n_650) );
INVx1_ASAP7_75t_L g694 ( .A(n_561), .Y(n_694) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_576), .Y(n_564) );
INVxp67_ASAP7_75t_L g646 ( .A(n_565), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_566), .B(n_577), .Y(n_582) );
INVx1_ASAP7_75t_L g688 ( .A(n_566), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_566), .B(n_665), .Y(n_699) );
BUFx3_ASAP7_75t_L g599 ( .A(n_567), .Y(n_599) );
AND2x2_ASAP7_75t_L g625 ( .A(n_567), .B(n_577), .Y(n_625) );
INVx2_ASAP7_75t_L g665 ( .A(n_567), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_576), .B(n_698), .Y(n_697) );
AOI211xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_583), .B(n_585), .C(n_594), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AOI21xp33_ASAP7_75t_L g628 ( .A1(n_580), .A2(n_629), .B(n_630), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_581), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_581), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g661 ( .A(n_582), .B(n_607), .Y(n_661) );
INVx3_ASAP7_75t_L g592 ( .A(n_584), .Y(n_592) );
OAI22xp5_ASAP7_75t_SL g585 ( .A1(n_586), .A2(n_588), .B1(n_591), .B2(n_593), .Y(n_585) );
OAI21xp5_ASAP7_75t_SL g610 ( .A1(n_587), .A2(n_611), .B(n_612), .Y(n_610) );
AND2x2_ASAP7_75t_L g636 ( .A(n_587), .B(n_600), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_587), .B(n_688), .Y(n_687) );
INVxp67_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g591 ( .A(n_590), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g660 ( .A(n_590), .Y(n_660) );
OAI21xp5_ASAP7_75t_SL g604 ( .A1(n_591), .A2(n_605), .B(n_610), .Y(n_604) );
OAI22xp33_ASAP7_75t_SL g594 ( .A1(n_595), .A2(n_597), .B1(n_601), .B2(n_602), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_596), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx1_ASAP7_75t_L g620 ( .A(n_599), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_599), .B(n_642), .Y(n_641) );
NOR3xp33_ASAP7_75t_L g603 ( .A(n_604), .B(n_615), .C(n_628), .Y(n_603) );
OAI22xp5_ASAP7_75t_SL g670 ( .A1(n_605), .A2(n_671), .B1(n_675), .B2(n_676), .Y(n_670) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_606), .B(n_608), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g675 ( .A(n_607), .B(n_608), .Y(n_675) );
AND2x2_ASAP7_75t_L g683 ( .A(n_608), .B(n_664), .Y(n_683) );
CKINVDCx16_ASAP7_75t_R g608 ( .A(n_609), .Y(n_608) );
O2A1O1Ixp33_ASAP7_75t_SL g691 ( .A1(n_609), .A2(n_692), .B(n_693), .C(n_694), .Y(n_691) );
OR2x2_ASAP7_75t_L g718 ( .A(n_609), .B(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
OAI21xp33_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_619), .B(n_621), .Y(n_615) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_L g653 ( .A1(n_617), .A2(n_654), .B(n_655), .C(n_658), .Y(n_653) );
OAI21xp33_ASAP7_75t_SL g621 ( .A1(n_622), .A2(n_623), .B(n_624), .Y(n_621) );
AND2x2_ASAP7_75t_L g686 ( .A(n_625), .B(n_644), .Y(n_686) );
INVxp67_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g664 ( .A(n_627), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g669 ( .A(n_629), .Y(n_669) );
NAND3xp33_ASAP7_75t_SL g632 ( .A(n_633), .B(n_653), .C(n_666), .Y(n_632) );
AOI211xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_636), .B(n_637), .C(n_645), .Y(n_633) );
INVx1_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
INVx1_ASAP7_75t_L g703 ( .A(n_640), .Y(n_703) );
OR2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
INVx1_ASAP7_75t_L g663 ( .A(n_642), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_642), .B(n_711), .Y(n_710) );
INVxp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
A2O1A1Ixp33_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_647), .B(n_648), .C(n_649), .Y(n_645) );
INVx2_ASAP7_75t_SL g657 ( .A(n_647), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_648), .A2(n_659), .B1(n_661), .B2(n_662), .Y(n_658) );
OAI21xp33_ASAP7_75t_SL g649 ( .A1(n_650), .A2(n_651), .B(n_652), .Y(n_649) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
AOI211xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_669), .B(n_670), .C(n_677), .Y(n_666) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
INVxp33_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g720 ( .A(n_674), .Y(n_720) );
NAND4xp25_ASAP7_75t_L g679 ( .A(n_680), .B(n_695), .C(n_708), .D(n_713), .Y(n_679) );
AOI211xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_683), .B(n_684), .C(n_691), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_687), .B(n_689), .Y(n_684) );
AOI21xp33_ASAP7_75t_L g704 ( .A1(n_685), .A2(n_705), .B(n_707), .Y(n_704) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_692), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_712), .Y(n_708) );
INVxp67_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g736 ( .A(n_721), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_724), .Y(n_723) );
CKINVDCx16_ASAP7_75t_R g732 ( .A(n_726), .Y(n_732) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx3_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
endmodule