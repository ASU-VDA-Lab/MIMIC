module fake_jpeg_13350_n_440 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_440);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_440;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_47),
.Y(n_104)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_53),
.Y(n_95)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_52),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_54),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_58),
.Y(n_100)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx5_ASAP7_75t_SL g116 ( 
.A(n_59),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_16),
.B(n_15),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_60),
.B(n_74),
.Y(n_115)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx2_ASAP7_75t_SL g120 ( 
.A(n_62),
.Y(n_120)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_70),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_69),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_34),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_71),
.Y(n_144)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_72),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_16),
.B(n_15),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_34),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_78),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_17),
.B(n_0),
.Y(n_78)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_79),
.B(n_83),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_40),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_87),
.Y(n_124)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_81),
.Y(n_129)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_86),
.Y(n_112)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_84),
.B(n_29),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_89),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

HAxp5_ASAP7_75t_SL g102 ( 
.A(n_90),
.B(n_29),
.CON(n_102),
.SN(n_102)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_21),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_42),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_90),
.A2(n_29),
.B1(n_45),
.B2(n_23),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_94),
.A2(n_103),
.B1(n_113),
.B2(n_118),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_97),
.B(n_4),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_23),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_99),
.B(n_106),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_102),
.B(n_73),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_68),
.A2(n_29),
.B1(n_43),
.B2(n_38),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_64),
.A2(n_20),
.B1(n_42),
.B2(n_39),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_SL g190 ( 
.A1(n_105),
.A2(n_106),
.B(n_130),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_45),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_51),
.A2(n_43),
.B1(n_38),
.B2(n_31),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_107),
.A2(n_131),
.B1(n_132),
.B2(n_136),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_75),
.A2(n_31),
.B1(n_30),
.B2(n_46),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_50),
.A2(n_30),
.B1(n_39),
.B2(n_36),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_76),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_55),
.A2(n_36),
.B1(n_35),
.B2(n_33),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_52),
.B(n_35),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_125),
.B(n_5),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_71),
.A2(n_33),
.B1(n_27),
.B2(n_25),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_85),
.A2(n_27),
.B1(n_25),
.B2(n_24),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_63),
.B(n_24),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_134),
.B(n_76),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_69),
.A2(n_83),
.B1(n_66),
.B2(n_65),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_54),
.B(n_20),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_138),
.B(n_140),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_89),
.B(n_17),
.Y(n_140)
);

NAND3xp33_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_59),
.C(n_1),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_145),
.B(n_149),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_146),
.Y(n_233)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_147),
.Y(n_206)
);

O2A1O1Ixp33_ASAP7_75t_SL g148 ( 
.A1(n_124),
.A2(n_81),
.B(n_47),
.C(n_89),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_148),
.A2(n_173),
.B(n_176),
.C(n_128),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_112),
.Y(n_149)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_150),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_151),
.B(n_156),
.Y(n_209)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_152),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_153),
.B(n_161),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_81),
.B1(n_73),
.B2(n_3),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_154),
.A2(n_167),
.B1(n_104),
.B2(n_139),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_155),
.A2(n_126),
.B(n_129),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_116),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_95),
.B(n_0),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_157),
.B(n_162),
.Y(n_204)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_93),
.Y(n_158)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_116),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_100),
.B(n_0),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_93),
.Y(n_163)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_101),
.B(n_1),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_166),
.B(n_169),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_189),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_116),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_170),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_138),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_171),
.B(n_181),
.Y(n_225)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_126),
.Y(n_172)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_172),
.Y(n_218)
);

O2A1O1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_124),
.A2(n_62),
.B(n_6),
.C(n_7),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_124),
.A2(n_62),
.B1(n_7),
.B2(n_8),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_174),
.A2(n_190),
.B1(n_104),
.B2(n_139),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_99),
.B(n_14),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_129),
.C(n_139),
.Y(n_207)
);

OA22x2_ASAP7_75t_L g176 ( 
.A1(n_102),
.A2(n_5),
.B1(n_8),
.B2(n_10),
.Y(n_176)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_96),
.Y(n_177)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

CKINVDCx9p33_ASAP7_75t_R g178 ( 
.A(n_130),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_178),
.Y(n_237)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_179),
.Y(n_232)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_126),
.Y(n_180)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_180),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_134),
.B(n_8),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_182),
.Y(n_235)
);

NAND2x1p5_ASAP7_75t_L g183 ( 
.A(n_97),
.B(n_115),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_183),
.A2(n_121),
.B(n_141),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_117),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_184),
.B(n_186),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_140),
.Y(n_186)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_187),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_136),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_191),
.Y(n_220)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_98),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_115),
.B(n_10),
.Y(n_191)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_96),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_104),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_171),
.A2(n_107),
.B1(n_143),
.B2(n_109),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_198),
.A2(n_199),
.B1(n_205),
.B2(n_228),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_159),
.A2(n_111),
.B1(n_143),
.B2(n_109),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_202),
.B(n_212),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g203 ( 
.A(n_159),
.B(n_115),
.C(n_111),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_203),
.B(n_168),
.C(n_176),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_188),
.A2(n_98),
.B1(n_137),
.B2(n_108),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_207),
.B(n_223),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_210),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_127),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_178),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_216),
.B(n_230),
.Y(n_270)
);

AO21x1_ASAP7_75t_L g258 ( 
.A1(n_221),
.A2(n_226),
.B(n_231),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_133),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_229),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_133),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_165),
.A2(n_121),
.B1(n_127),
.B2(n_122),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_194),
.A2(n_144),
.B1(n_137),
.B2(n_122),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_234),
.A2(n_164),
.B1(n_193),
.B2(n_182),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_185),
.A2(n_144),
.B1(n_128),
.B2(n_114),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_236),
.A2(n_170),
.B1(n_173),
.B2(n_146),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_238),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_225),
.B(n_149),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_239),
.B(n_241),
.Y(n_285)
);

BUFx12f_ASAP7_75t_L g240 ( 
.A(n_233),
.Y(n_240)
);

BUFx4f_ASAP7_75t_SL g297 ( 
.A(n_240),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_209),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_206),
.Y(n_242)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_242),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_220),
.A2(n_155),
.B1(n_165),
.B2(n_180),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_245),
.A2(n_246),
.B1(n_253),
.B2(n_255),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_220),
.A2(n_155),
.B1(n_183),
.B2(n_194),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_229),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_247),
.B(n_249),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_200),
.B(n_175),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_210),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_251),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_227),
.B(n_184),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_200),
.B(n_175),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_252),
.B(n_261),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_223),
.A2(n_183),
.B1(n_153),
.B2(n_148),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_254),
.B(n_264),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_226),
.A2(n_148),
.B1(n_176),
.B2(n_168),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_210),
.Y(n_256)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_256),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_211),
.B(n_156),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_257),
.B(n_267),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_205),
.A2(n_216),
.B1(n_198),
.B2(n_237),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_262),
.B1(n_271),
.B2(n_217),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_200),
.B(n_161),
.Y(n_261)
);

OA22x2_ASAP7_75t_L g263 ( 
.A1(n_221),
.A2(n_176),
.B1(n_163),
.B2(n_147),
.Y(n_263)
);

A2O1A1Ixp33_ASAP7_75t_SL g296 ( 
.A1(n_263),
.A2(n_212),
.B(n_114),
.C(n_208),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_207),
.B(n_152),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_203),
.B(n_158),
.C(n_189),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_219),
.C(n_218),
.Y(n_284)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_206),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_266),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_204),
.B(n_160),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_201),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_268),
.B(n_269),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_235),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_270),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_228),
.A2(n_150),
.B1(n_177),
.B2(n_146),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_272),
.A2(n_213),
.B1(n_233),
.B2(n_222),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_214),
.B(n_187),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_199),
.Y(n_291)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_196),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_275),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_276),
.A2(n_290),
.B1(n_300),
.B2(n_308),
.Y(n_311)
);

AO22x1_ASAP7_75t_L g277 ( 
.A1(n_263),
.A2(n_202),
.B1(n_219),
.B2(n_218),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_277),
.B(n_286),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_248),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_280),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_248),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_281),
.B(n_291),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_284),
.B(n_304),
.C(n_305),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_273),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_258),
.A2(n_201),
.B(n_195),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_287),
.A2(n_294),
.B(n_299),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_258),
.A2(n_236),
.B1(n_217),
.B2(n_215),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_248),
.A2(n_214),
.B(n_215),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_296),
.A2(n_306),
.B1(n_309),
.B2(n_256),
.Y(n_322)
);

A2O1A1Ixp33_ASAP7_75t_SL g299 ( 
.A1(n_253),
.A2(n_212),
.B(n_120),
.C(n_208),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_244),
.A2(n_213),
.B1(n_179),
.B2(n_232),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_264),
.B(n_196),
.C(n_197),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_274),
.B(n_197),
.C(n_232),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_274),
.B(n_222),
.C(n_11),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_299),
.C(n_288),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_243),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_243),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_282),
.Y(n_310)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_310),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_298),
.A2(n_244),
.B1(n_247),
.B2(n_262),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_312),
.A2(n_322),
.B1(n_326),
.B2(n_318),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_290),
.A2(n_255),
.B1(n_246),
.B2(n_245),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_313),
.A2(n_317),
.B1(n_321),
.B2(n_330),
.Y(n_361)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_300),
.Y(n_315)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_315),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_285),
.B(n_265),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_316),
.B(n_329),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_291),
.A2(n_254),
.B1(n_263),
.B2(n_266),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_303),
.B(n_288),
.Y(n_319)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_319),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_294),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_320),
.B(n_334),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_280),
.A2(n_263),
.B1(n_242),
.B2(n_256),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_289),
.B(n_249),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_323),
.B(n_335),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_302),
.A2(n_271),
.B1(n_261),
.B2(n_259),
.Y(n_325)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_325),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_298),
.A2(n_259),
.B1(n_252),
.B2(n_275),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_278),
.Y(n_327)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_327),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_283),
.B(n_269),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_281),
.A2(n_240),
.B1(n_12),
.B2(n_13),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_304),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_331),
.Y(n_342)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_301),
.Y(n_332)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_332),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_293),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_289),
.B(n_240),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_336),
.B(n_337),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_284),
.B(n_240),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_320),
.A2(n_279),
.B(n_277),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_338),
.A2(n_356),
.B(n_335),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_334),
.B(n_301),
.Y(n_341)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_341),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_313),
.A2(n_317),
.B1(n_311),
.B2(n_321),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_343),
.B(n_353),
.Y(n_377)
);

OA21x2_ASAP7_75t_L g347 ( 
.A1(n_315),
.A2(n_296),
.B(n_306),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_347),
.A2(n_349),
.B(n_318),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_314),
.B(n_279),
.Y(n_348)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_348),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_328),
.A2(n_296),
.B(n_295),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_312),
.B(n_295),
.Y(n_351)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_351),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_333),
.Y(n_353)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_354),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_328),
.A2(n_299),
.B(n_296),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_326),
.A2(n_305),
.B1(n_299),
.B2(n_307),
.Y(n_357)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_357),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_311),
.A2(n_292),
.B1(n_297),
.B2(n_13),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_360),
.B(n_330),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_355),
.B(n_342),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_374),
.Y(n_384)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_346),
.Y(n_366)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_366),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_368),
.A2(n_370),
.B(n_356),
.Y(n_393)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_341),
.Y(n_371)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_371),
.Y(n_389)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_350),
.Y(n_372)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_372),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_355),
.B(n_319),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_373),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_342),
.B(n_324),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_345),
.B(n_324),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_375),
.A2(n_381),
.B1(n_353),
.B2(n_358),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_352),
.B(n_337),
.C(n_336),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_376),
.B(n_352),
.C(n_379),
.Y(n_391)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_350),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_378),
.B(n_380),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_348),
.B(n_323),
.Y(n_379)
);

MAJx2_ASAP7_75t_L g382 ( 
.A(n_379),
.B(n_376),
.C(n_351),
.Y(n_382)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_339),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_386),
.C(n_391),
.Y(n_400)
);

AOI321xp33_ASAP7_75t_L g383 ( 
.A1(n_369),
.A2(n_340),
.A3(n_346),
.B1(n_349),
.B2(n_345),
.C(n_338),
.Y(n_383)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_383),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_367),
.A2(n_354),
.B1(n_357),
.B2(n_349),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_385),
.A2(n_396),
.B1(n_347),
.B2(n_377),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_370),
.B(n_359),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_367),
.A2(n_343),
.B1(n_361),
.B2(n_347),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_387),
.A2(n_362),
.B1(n_381),
.B2(n_344),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_390),
.B(n_394),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_393),
.A2(n_366),
.B1(n_368),
.B2(n_363),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_369),
.B(n_359),
.C(n_340),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_377),
.A2(n_344),
.B1(n_361),
.B2(n_347),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_399),
.B(n_401),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_394),
.B(n_359),
.C(n_365),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_402),
.B(n_403),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_391),
.B(n_365),
.C(n_371),
.Y(n_403)
);

AOI21x1_ASAP7_75t_L g404 ( 
.A1(n_384),
.A2(n_363),
.B(n_362),
.Y(n_404)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_404),
.Y(n_411)
);

BUFx24_ASAP7_75t_SL g405 ( 
.A(n_388),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_405),
.B(n_409),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_385),
.B(n_327),
.Y(n_406)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_406),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_408),
.Y(n_419)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_397),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_403),
.B(n_382),
.C(n_386),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_410),
.B(n_414),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_402),
.B(n_393),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_398),
.B(n_387),
.C(n_396),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_416),
.B(n_417),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_400),
.A2(n_395),
.B(n_389),
.Y(n_417)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_413),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_420),
.B(n_422),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_414),
.B(n_401),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_421),
.B(n_423),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_415),
.B(n_407),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_416),
.B(n_400),
.C(n_399),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_411),
.A2(n_395),
.B1(n_397),
.B2(n_392),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_426),
.A2(n_418),
.B(n_419),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_427),
.A2(n_428),
.B(n_429),
.Y(n_433)
);

AO21x2_ASAP7_75t_L g428 ( 
.A1(n_425),
.A2(n_412),
.B(n_383),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_424),
.A2(n_410),
.B(n_412),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_431),
.B(n_423),
.C(n_421),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_432),
.B(n_358),
.C(n_360),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_430),
.Y(n_434)
);

AOI21x1_ASAP7_75t_L g436 ( 
.A1(n_434),
.A2(n_372),
.B(n_378),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_435),
.A2(n_436),
.B1(n_380),
.B2(n_339),
.Y(n_437)
);

NAND2xp33_ASAP7_75t_SL g438 ( 
.A(n_437),
.B(n_433),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_438),
.A2(n_310),
.B(n_297),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_439),
.B(n_297),
.Y(n_440)
);


endmodule