module fake_jpeg_12723_n_562 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_562);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_562;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_15),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_54),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_20),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_55),
.B(n_63),
.Y(n_114)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_56),
.Y(n_122)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_57),
.Y(n_151)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_62),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_28),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_65),
.Y(n_145)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_28),
.Y(n_66)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_67),
.Y(n_137)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_68),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_28),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_69),
.B(n_78),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_70),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_71),
.Y(n_147)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g156 ( 
.A(n_72),
.Y(n_156)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_73),
.Y(n_152)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_75),
.Y(n_142)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_29),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_21),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_79),
.B(n_80),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_41),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_81),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_41),
.B(n_17),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_82),
.B(n_83),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_43),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_85),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx5_ASAP7_75t_SL g112 ( 
.A(n_87),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_43),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_88),
.B(n_89),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_33),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_36),
.B(n_17),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_90),
.B(n_100),
.Y(n_159)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_93),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_98),
.Y(n_155)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx3_ASAP7_75t_SL g174 ( 
.A(n_99),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_48),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_48),
.B(n_17),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_102),
.B(n_103),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_52),
.B(n_13),
.Y(n_103)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_21),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_107),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_52),
.B(n_30),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_108),
.B(n_37),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_81),
.A2(n_37),
.B1(n_30),
.B2(n_66),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_109),
.A2(n_74),
.B1(n_64),
.B2(n_107),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_55),
.B(n_25),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_118),
.B(n_128),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_58),
.A2(n_53),
.B1(n_20),
.B2(n_39),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_124),
.A2(n_44),
.B1(n_35),
.B2(n_45),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_76),
.B(n_25),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_54),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_132),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_59),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_138),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_87),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_146),
.B(n_165),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g148 ( 
.A(n_70),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_148),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_71),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_75),
.Y(n_161)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_161),
.Y(n_216)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_75),
.Y(n_162)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_162),
.Y(n_217)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_86),
.Y(n_164)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_164),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_93),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_167),
.B(n_171),
.Y(n_222)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_67),
.Y(n_168)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_168),
.Y(n_176)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_86),
.Y(n_170)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

AOI21xp33_ASAP7_75t_L g171 ( 
.A1(n_79),
.A2(n_34),
.B(n_51),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_79),
.B(n_51),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_172),
.B(n_32),
.Y(n_229)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_101),
.Y(n_175)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_131),
.Y(n_180)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_180),
.Y(n_272)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_121),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_181),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_182),
.Y(n_245)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_183),
.Y(n_274)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_122),
.Y(n_185)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_185),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_149),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_186),
.B(n_191),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_149),
.B(n_53),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_187),
.B(n_208),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_188),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_34),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_123),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_192),
.B(n_204),
.Y(n_246)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_127),
.Y(n_193)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_193),
.Y(n_289)
);

O2A1O1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_169),
.A2(n_104),
.B(n_93),
.C(n_65),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_L g292 ( 
.A1(n_194),
.A2(n_220),
.B(n_181),
.Y(n_292)
);

BUFx12f_ASAP7_75t_L g195 ( 
.A(n_154),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_195),
.Y(n_265)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_134),
.Y(n_196)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_196),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_123),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_197),
.Y(n_269)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_130),
.Y(n_198)
);

BUFx2_ASAP7_75t_SL g243 ( 
.A(n_198),
.Y(n_243)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_132),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_199),
.Y(n_260)
);

CKINVDCx9p33_ASAP7_75t_R g200 ( 
.A(n_112),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_200),
.Y(n_284)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_135),
.Y(n_201)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_201),
.Y(n_250)
);

AO22x1_ASAP7_75t_SL g202 ( 
.A1(n_114),
.A2(n_105),
.B1(n_72),
.B2(n_99),
.Y(n_202)
);

AO22x1_ASAP7_75t_L g249 ( 
.A1(n_202),
.A2(n_139),
.B1(n_143),
.B2(n_144),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_203),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_27),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_205),
.A2(n_220),
.B1(n_174),
.B2(n_119),
.Y(n_262)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_129),
.A2(n_172),
.B(n_114),
.C(n_167),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g266 ( 
.A1(n_207),
.A2(n_49),
.B(n_40),
.C(n_32),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_159),
.B(n_98),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_157),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_209),
.B(n_211),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_159),
.B(n_140),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_210),
.B(n_214),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_112),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_111),
.Y(n_212)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_212),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_129),
.B(n_60),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_213),
.B(n_225),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_140),
.B(n_160),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_137),
.Y(n_215)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_215),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_113),
.Y(n_218)
);

INVx5_ASAP7_75t_L g291 ( 
.A(n_218),
.Y(n_291)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_130),
.Y(n_219)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_219),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_174),
.A2(n_62),
.B1(n_95),
.B2(n_91),
.Y(n_220)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_126),
.Y(n_221)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_221),
.Y(n_248)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_150),
.Y(n_223)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_223),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_133),
.B(n_49),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_224),
.B(n_232),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_156),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_120),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_236),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_109),
.A2(n_106),
.B1(n_97),
.B2(n_92),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_228),
.A2(n_230),
.B1(n_233),
.B2(n_50),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_229),
.B(n_11),
.Y(n_287)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_138),
.Y(n_231)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_231),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_133),
.B(n_40),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_152),
.A2(n_73),
.B1(n_85),
.B2(n_84),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_116),
.Y(n_234)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_234),
.Y(n_285)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_125),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_117),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_237),
.B(n_136),
.Y(n_290)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_155),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_151),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_189),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_240),
.B(n_258),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_177),
.B(n_156),
.Y(n_247)
);

OAI21xp33_ASAP7_75t_L g319 ( 
.A1(n_247),
.A2(n_255),
.B(n_256),
.Y(n_319)
);

OA22x2_ASAP7_75t_L g337 ( 
.A1(n_249),
.A2(n_279),
.B1(n_35),
.B2(n_24),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_156),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_252),
.B(n_271),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_194),
.B(n_57),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_176),
.B(n_151),
.Y(n_256)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_222),
.B(n_145),
.CI(n_13),
.CON(n_258),
.SN(n_258)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_207),
.B(n_68),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_261),
.B(n_264),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_L g313 ( 
.A1(n_262),
.A2(n_179),
.B1(n_136),
.B2(n_231),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_266),
.B(n_22),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_190),
.B(n_158),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_267),
.B(n_268),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_197),
.B(n_126),
.Y(n_268)
);

AND2x2_ASAP7_75t_SL g271 ( 
.A(n_184),
.B(n_110),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_202),
.A2(n_115),
.B(n_1),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_275),
.B(n_277),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_216),
.B(n_152),
.C(n_147),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_228),
.A2(n_22),
.B1(n_50),
.B2(n_44),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_281),
.A2(n_295),
.B1(n_35),
.B2(n_44),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_217),
.B(n_147),
.C(n_141),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_282),
.B(n_292),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_181),
.B(n_13),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_286),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_11),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_205),
.A2(n_148),
.B(n_141),
.Y(n_288)
);

O2A1O1Ixp33_ASAP7_75t_L g329 ( 
.A1(n_288),
.A2(n_199),
.B(n_227),
.C(n_195),
.Y(n_329)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_290),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_182),
.A2(n_22),
.B1(n_50),
.B2(n_44),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_247),
.B(n_198),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_296),
.B(n_308),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_270),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_297),
.B(n_299),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_271),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_300),
.A2(n_330),
.B(n_341),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_284),
.A2(n_221),
.B1(n_219),
.B2(n_179),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_301),
.Y(n_362)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_273),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_303),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_304),
.B(n_312),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_271),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_305),
.B(n_310),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_244),
.B(n_178),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g375 ( 
.A(n_307),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_280),
.B(n_203),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_255),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_261),
.B(n_218),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_311),
.B(n_327),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_251),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_313),
.A2(n_316),
.B1(n_324),
.B2(n_335),
.Y(n_368)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_291),
.Y(n_314)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_314),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_256),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_315),
.B(n_321),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_279),
.A2(n_237),
.B1(n_39),
.B2(n_24),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_254),
.Y(n_317)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_317),
.Y(n_373)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_263),
.Y(n_318)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_318),
.Y(n_382)
);

INVx13_ASAP7_75t_L g320 ( 
.A(n_265),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_320),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_242),
.B(n_178),
.Y(n_321)
);

NAND2x1_ASAP7_75t_L g322 ( 
.A(n_252),
.B(n_206),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_322),
.A2(n_286),
.B(n_248),
.Y(n_364)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_273),
.Y(n_323)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_323),
.Y(n_383)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_276),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_325),
.B(n_328),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_246),
.B(n_206),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_274),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_329),
.A2(n_288),
.B(n_292),
.Y(n_345)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_258),
.B(n_239),
.Y(n_330)
);

AND2x6_ASAP7_75t_L g331 ( 
.A(n_258),
.B(n_11),
.Y(n_331)
);

AOI322xp5_ASAP7_75t_L g379 ( 
.A1(n_331),
.A2(n_257),
.A3(n_259),
.B1(n_188),
.B2(n_4),
.C1(n_6),
.C2(n_0),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_269),
.B(n_188),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_332),
.B(n_336),
.Y(n_372)
);

OAI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_275),
.A2(n_24),
.B1(n_39),
.B2(n_35),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_250),
.B(n_241),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_337),
.B(n_339),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_257),
.Y(n_339)
);

INVx13_ASAP7_75t_L g340 ( 
.A(n_265),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_340),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_283),
.B(n_195),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_281),
.A2(n_227),
.B1(n_239),
.B2(n_235),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_342),
.A2(n_260),
.B1(n_294),
.B2(n_248),
.Y(n_370)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_272),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_343),
.B(n_344),
.Y(n_367)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_285),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_345),
.A2(n_364),
.B(n_377),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_296),
.B(n_277),
.C(n_282),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_346),
.B(n_363),
.C(n_385),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_330),
.A2(n_322),
.B(n_333),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_347),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_302),
.A2(n_262),
.B1(n_249),
.B2(n_295),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g396 ( 
.A1(n_351),
.A2(n_355),
.B1(n_357),
.B2(n_369),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_297),
.A2(n_284),
.B1(n_291),
.B2(n_253),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_354),
.B(n_378),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_302),
.A2(n_266),
.B1(n_253),
.B2(n_245),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_311),
.A2(n_245),
.B1(n_243),
.B2(n_294),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_327),
.Y(n_358)
);

INVx13_ASAP7_75t_L g406 ( 
.A(n_358),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_308),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_361),
.B(n_379),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_334),
.B(n_309),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_300),
.A2(n_337),
.B1(n_326),
.B2(n_299),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_370),
.A2(n_376),
.B1(n_368),
.B2(n_383),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_326),
.A2(n_260),
.B1(n_289),
.B2(n_278),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_333),
.A2(n_326),
.B(n_322),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_337),
.A2(n_293),
.B1(n_235),
.B2(n_259),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_333),
.B(n_2),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_381),
.B(n_315),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_309),
.A2(n_3),
.B(n_4),
.Y(n_384)
);

AO22x1_ASAP7_75t_L g405 ( 
.A1(n_384),
.A2(n_386),
.B1(n_313),
.B2(n_344),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_309),
.B(n_319),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_298),
.A2(n_3),
.B(n_4),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_380),
.Y(n_387)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_387),
.Y(n_425)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_367),
.Y(n_389)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_389),
.Y(n_448)
);

AOI22x1_ASAP7_75t_L g390 ( 
.A1(n_360),
.A2(n_342),
.B1(n_316),
.B2(n_329),
.Y(n_390)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_390),
.Y(n_442)
);

AND2x6_ASAP7_75t_L g392 ( 
.A(n_377),
.B(n_331),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_392),
.A2(n_405),
.B(n_362),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_393),
.B(n_394),
.Y(n_445)
);

NOR2x1_ASAP7_75t_L g394 ( 
.A(n_381),
.B(n_341),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_361),
.A2(n_337),
.B1(n_310),
.B2(n_306),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_395),
.A2(n_413),
.B1(n_351),
.B2(n_378),
.Y(n_438)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_397),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_363),
.B(n_341),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_399),
.B(n_402),
.C(n_415),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_367),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_400),
.B(n_401),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_380),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_385),
.B(n_306),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_374),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_403),
.B(n_404),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_358),
.B(n_353),
.Y(n_404)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_374),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_407),
.B(n_416),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_372),
.B(n_312),
.Y(n_408)
);

CKINVDCx14_ASAP7_75t_R g426 ( 
.A(n_408),
.Y(n_426)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_373),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_409),
.B(n_410),
.Y(n_430)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_373),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_353),
.B(n_318),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_411),
.B(n_414),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_368),
.A2(n_360),
.B1(n_348),
.B2(n_347),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_348),
.B(n_317),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_352),
.B(n_338),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_382),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_352),
.B(n_325),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_417),
.B(n_421),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_371),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_418),
.Y(n_431)
);

OAI21xp33_ASAP7_75t_L g419 ( 
.A1(n_359),
.A2(n_343),
.B(n_328),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_419),
.A2(n_349),
.B1(n_365),
.B2(n_366),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_375),
.B(n_339),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_420),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_354),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_398),
.B(n_346),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_428),
.B(n_436),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_391),
.A2(n_350),
.B(n_345),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_433),
.A2(n_434),
.B(n_440),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_422),
.A2(n_362),
.B(n_364),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_398),
.B(n_359),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_399),
.B(n_376),
.C(n_369),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_437),
.B(n_395),
.C(n_391),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_438),
.A2(n_441),
.B1(n_390),
.B2(n_384),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_413),
.A2(n_355),
.B1(n_357),
.B2(n_324),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_404),
.B(n_350),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_443),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_422),
.A2(n_370),
.B(n_365),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_444),
.B(n_405),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_402),
.B(n_415),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_446),
.B(n_394),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_414),
.B(n_382),
.Y(n_447)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_447),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_411),
.B(n_383),
.Y(n_449)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_449),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_417),
.B(n_356),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_SL g468 ( 
.A(n_450),
.B(n_396),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_387),
.B(n_349),
.Y(n_451)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_451),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_453),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_454),
.B(n_457),
.C(n_466),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_431),
.B(n_403),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_455),
.B(n_458),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_428),
.B(n_393),
.C(n_406),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_431),
.B(n_386),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_442),
.A2(n_452),
.B1(n_432),
.B2(n_425),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_460),
.A2(n_473),
.B1(n_438),
.B2(n_443),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_462),
.B(n_423),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_426),
.B(n_412),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_465),
.B(n_467),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_436),
.B(n_406),
.C(n_366),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_435),
.B(n_450),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_468),
.B(n_314),
.Y(n_498)
);

CKINVDCx14_ASAP7_75t_R g469 ( 
.A(n_445),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_469),
.B(n_445),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_447),
.B(n_388),
.Y(n_470)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_470),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_429),
.B(n_388),
.Y(n_471)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_471),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_442),
.A2(n_390),
.B1(n_405),
.B2(n_392),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_474),
.A2(n_443),
.B(n_424),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_423),
.B(n_446),
.C(n_437),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_475),
.B(n_433),
.C(n_432),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_424),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_476),
.B(n_480),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_435),
.B(n_407),
.Y(n_477)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_477),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_SL g490 ( 
.A1(n_478),
.A2(n_452),
.B1(n_425),
.B2(n_448),
.Y(n_490)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_449),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_482),
.B(n_484),
.Y(n_503)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_483),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_485),
.B(n_492),
.C(n_481),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_487),
.A2(n_497),
.B(n_479),
.Y(n_512)
);

A2O1A1Ixp33_ASAP7_75t_SL g488 ( 
.A1(n_464),
.A2(n_434),
.B(n_440),
.C(n_444),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_488),
.B(n_463),
.C(n_478),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_490),
.B(n_484),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_473),
.A2(n_441),
.B1(n_427),
.B2(n_429),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_491),
.B(n_492),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_456),
.B(n_466),
.C(n_475),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_460),
.A2(n_448),
.B1(n_453),
.B2(n_451),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_493),
.B(n_495),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_457),
.B(n_439),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_494),
.B(n_496),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_470),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_462),
.B(n_439),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_464),
.A2(n_430),
.B(n_303),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_498),
.B(n_468),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_504),
.B(n_518),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_505),
.B(n_491),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_499),
.B(n_456),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_507),
.B(n_509),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_502),
.Y(n_511)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_511),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_512),
.A2(n_516),
.B(n_488),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_485),
.B(n_454),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_513),
.B(n_517),
.Y(n_529)
);

INVx5_ASAP7_75t_L g515 ( 
.A(n_501),
.Y(n_515)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_515),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_481),
.B(n_479),
.C(n_480),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_494),
.B(n_472),
.C(n_476),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_489),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_519),
.B(n_459),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_482),
.B(n_472),
.C(n_459),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_520),
.B(n_496),
.C(n_497),
.Y(n_525)
);

OR2x2_ASAP7_75t_L g542 ( 
.A(n_522),
.B(n_515),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_525),
.B(n_535),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_SL g526 ( 
.A(n_506),
.B(n_461),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_526),
.B(n_531),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_516),
.A2(n_461),
.B1(n_487),
.B2(n_486),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_527),
.A2(n_533),
.B1(n_505),
.B2(n_518),
.Y(n_536)
);

INVxp33_ASAP7_75t_L g540 ( 
.A(n_528),
.Y(n_540)
);

OAI321xp33_ASAP7_75t_L g530 ( 
.A1(n_508),
.A2(n_489),
.A3(n_500),
.B1(n_471),
.B2(n_488),
.C(n_493),
.Y(n_530)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_530),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_514),
.A2(n_488),
.B(n_498),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_532),
.A2(n_510),
.B(n_520),
.Y(n_537)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_511),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_503),
.B(n_323),
.C(n_340),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_536),
.A2(n_531),
.B1(n_532),
.B2(n_521),
.Y(n_549)
);

AOI21x1_ASAP7_75t_L g546 ( 
.A1(n_537),
.A2(n_542),
.B(n_525),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_534),
.B(n_517),
.C(n_503),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_539),
.B(n_543),
.C(n_544),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_529),
.B(n_320),
.C(n_4),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_523),
.B(n_9),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_546),
.A2(n_549),
.B1(n_540),
.B2(n_541),
.Y(n_552)
);

NOR3xp33_ASAP7_75t_SL g547 ( 
.A(n_538),
.B(n_522),
.C(n_524),
.Y(n_547)
);

NOR2x1_ASAP7_75t_L g554 ( 
.A(n_547),
.B(n_551),
.Y(n_554)
);

NAND2x1_ASAP7_75t_SL g548 ( 
.A(n_539),
.B(n_535),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g553 ( 
.A(n_548),
.B(n_540),
.Y(n_553)
);

AOI31xp67_ASAP7_75t_L g551 ( 
.A1(n_545),
.A2(n_526),
.A3(n_527),
.B(n_7),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_552),
.B(n_553),
.Y(n_555)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g556 ( 
.A1(n_553),
.A2(n_542),
.B(n_549),
.C(n_550),
.D(n_543),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_556),
.B(n_554),
.C(n_6),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_557),
.B(n_555),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_558),
.B(n_3),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_559),
.B(n_3),
.C(n_6),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_SL g561 ( 
.A1(n_560),
.A2(n_7),
.B(n_8),
.Y(n_561)
);

O2A1O1Ixp33_ASAP7_75t_SL g562 ( 
.A1(n_561),
.A2(n_7),
.B(n_8),
.C(n_426),
.Y(n_562)
);


endmodule