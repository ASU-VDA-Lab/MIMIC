module fake_jpeg_28379_n_165 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_165);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_24),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_14),
.Y(n_30)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_25),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_22),
.A2(n_11),
.B1(n_20),
.B2(n_10),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_10),
.B1(n_28),
.B2(n_18),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g32 ( 
.A1(n_24),
.A2(n_11),
.B1(n_14),
.B2(n_12),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_35),
.B1(n_28),
.B2(n_30),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_24),
.A2(n_11),
.B1(n_20),
.B2(n_14),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_34),
.A2(n_11),
.B1(n_24),
.B2(n_26),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_39),
.B1(n_29),
.B2(n_47),
.Y(n_54)
);

NAND3xp33_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_26),
.C(n_27),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_34),
.A2(n_26),
.B1(n_18),
.B2(n_17),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_32),
.A2(n_28),
.B1(n_20),
.B2(n_14),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_41),
.B1(n_45),
.B2(n_29),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_25),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_18),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_22),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_49),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_14),
.B1(n_25),
.B2(n_21),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_10),
.B1(n_13),
.B2(n_15),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_39),
.B1(n_29),
.B2(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_13),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_17),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_56),
.Y(n_64)
);

AND2x6_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_31),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_SL g71 ( 
.A(n_52),
.B(n_54),
.C(n_55),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_21),
.B1(n_15),
.B2(n_23),
.Y(n_75)
);

AND2x6_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_31),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_13),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_42),
.B(n_40),
.C(n_45),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_48),
.B(n_33),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_63),
.B1(n_21),
.B2(n_25),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_48),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_63),
.Y(n_82)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_66),
.B(n_69),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_55),
.A2(n_37),
.B1(n_42),
.B2(n_33),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_67),
.A2(n_74),
.B1(n_59),
.B2(n_55),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_68),
.A2(n_73),
.B(n_59),
.Y(n_78)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_76),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_51),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_72),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_57),
.A2(n_15),
.B1(n_29),
.B2(n_47),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_61),
.B1(n_56),
.B2(n_63),
.Y(n_86)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_80),
.A2(n_81),
.B1(n_71),
.B2(n_64),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_66),
.A2(n_61),
.B1(n_52),
.B2(n_58),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_64),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g83 ( 
.A(n_65),
.B(n_60),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_84),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_60),
.B(n_63),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_85),
.B(n_86),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_52),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_91),
.C(n_71),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_75),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_50),
.Y(n_90)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_21),
.C(n_23),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_78),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_95),
.A2(n_104),
.B1(n_101),
.B2(n_86),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_16),
.B1(n_12),
.B2(n_23),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_97),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_70),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_99),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_23),
.C(n_46),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_105),
.C(n_108),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_46),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_23),
.C(n_46),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_89),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_106),
.B(n_107),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_79),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_16),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_117),
.C(n_119),
.Y(n_122)
);

XNOR2x1_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_80),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_111),
.B(n_104),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_91),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_118),
.A2(n_94),
.B1(n_27),
.B2(n_16),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_23),
.C(n_27),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_27),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_117),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_128),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_95),
.B1(n_102),
.B2(n_97),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_124),
.A2(n_115),
.B1(n_114),
.B2(n_113),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_121),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_0),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_113),
.A2(n_98),
.B1(n_102),
.B2(n_92),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_126),
.A2(n_129),
.B1(n_125),
.B2(n_124),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_105),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_127),
.B(n_27),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_116),
.B(n_6),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_131),
.Y(n_134)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_136),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_109),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_137),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_126),
.A2(n_122),
.B1(n_16),
.B2(n_12),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_0),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_122),
.B(n_12),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_143),
.Y(n_151)
);

AO21x1_ASAP7_75t_L g141 ( 
.A1(n_132),
.A2(n_9),
.B(n_8),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_141),
.B(n_145),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_9),
.C(n_8),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_5),
.C(n_1),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_5),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_133),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_148),
.B(n_152),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_134),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_141),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_144),
.A2(n_5),
.B(n_1),
.Y(n_150)
);

AOI21xp33_ASAP7_75t_L g156 ( 
.A1(n_150),
.A2(n_1),
.B(n_2),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_155),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_147),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_155)
);

OAI221xp5_ASAP7_75t_L g158 ( 
.A1(n_156),
.A2(n_157),
.B1(n_147),
.B2(n_4),
.C(n_3),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_2),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_158),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_151),
.C(n_3),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_3),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_159),
.C(n_4),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_162),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_4),
.Y(n_165)
);


endmodule