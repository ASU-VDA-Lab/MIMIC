module real_aes_9895_n_9 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_1, n_9);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_1;
output n_9;
wire n_17;
wire n_22;
wire n_13;
wire n_24;
wire n_12;
wire n_19;
wire n_25;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_27;
wire n_23;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_10;
OAI221xp5_ASAP7_75t_L g20 ( .A1(n_0), .A2(n_7), .B1(n_21), .B2(n_22), .C(n_27), .Y(n_20) );
AOI221xp5_ASAP7_75t_L g9 ( .A1(n_1), .A2(n_10), .B1(n_16), .B2(n_17), .C(n_19), .Y(n_9) );
HB1xp67_ASAP7_75t_L g16 ( .A(n_2), .Y(n_16) );
OAI21xp33_ASAP7_75t_L g10 ( .A1(n_3), .A2(n_11), .B(n_12), .Y(n_10) );
HB1xp67_ASAP7_75t_L g11 ( .A(n_4), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_5), .B(n_14), .Y(n_18) );
INVx2_ASAP7_75t_L g15 ( .A(n_6), .Y(n_15) );
BUFx2_ASAP7_75t_L g26 ( .A(n_8), .Y(n_26) );
NOR2xp33_ASAP7_75t_L g12 ( .A(n_13), .B(n_16), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_14), .Y(n_13) );
NOR2xp33_ASAP7_75t_L g19 ( .A(n_14), .B(n_20), .Y(n_19) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_15), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g27 ( .A(n_16), .Y(n_27) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_18), .Y(n_17) );
INVx1_ASAP7_75t_SL g21 ( .A(n_22), .Y(n_21) );
INVx5_ASAP7_75t_L g22 ( .A(n_23), .Y(n_22) );
BUFx8_ASAP7_75t_SL g23 ( .A(n_24), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_25), .Y(n_24) );
BUFx2_ASAP7_75t_L g25 ( .A(n_26), .Y(n_25) );
endmodule