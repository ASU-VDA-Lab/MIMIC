module fake_jpeg_2024_n_190 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_190);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_12),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_0),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_14),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_2),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_25),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_27),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_28),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_69),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_0),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_67),
.B(n_51),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_77),
.B(n_49),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_62),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_82),
.B(n_83),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_59),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_50),
.B1(n_48),
.B2(n_72),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_60),
.Y(n_96)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_52),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_68),
.Y(n_95)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g89 ( 
.A1(n_86),
.A2(n_49),
.B(n_54),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_91),
.B(n_94),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_SL g91 ( 
.A1(n_84),
.A2(n_61),
.B(n_73),
.C(n_53),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_55),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_97),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_93),
.B(n_95),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_60),
.B(n_51),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_96),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_58),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_58),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_100),
.Y(n_114)
);

AOI21xp33_ASAP7_75t_SL g99 ( 
.A1(n_80),
.A2(n_55),
.B(n_53),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_75),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_54),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_75),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_85),
.Y(n_116)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_94),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_115),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_76),
.C(n_63),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_107),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_76),
.C(n_65),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_41),
.Y(n_142)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_64),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_120),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_24),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_101),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_121),
.B(n_21),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_91),
.A2(n_79),
.B1(n_46),
.B2(n_70),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_57),
.B1(n_23),
.B2(n_29),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_119),
.A2(n_91),
.B1(n_79),
.B2(n_85),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_124),
.B1(n_133),
.B2(n_136),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_104),
.A2(n_57),
.B1(n_2),
.B2(n_3),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_1),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_127),
.B(n_132),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_130),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_129),
.B(n_139),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_110),
.Y(n_130)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_1),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_19),
.B1(n_43),
.B2(n_42),
.Y(n_136)
);

AO22x1_ASAP7_75t_SL g138 ( 
.A1(n_122),
.A2(n_44),
.B1(n_17),
.B2(n_18),
.Y(n_138)
);

OA21x2_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_40),
.B(n_39),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_3),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_107),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_143),
.Y(n_147)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_141),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_142),
.A2(n_120),
.B(n_118),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_111),
.B(n_4),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_150),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_135),
.B(n_123),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_146),
.A2(n_155),
.B(n_157),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_113),
.Y(n_149)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_131),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_159),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_38),
.B(n_37),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_134),
.A2(n_4),
.B(n_5),
.Y(n_157)
);

OAI22x1_ASAP7_75t_SL g158 ( 
.A1(n_133),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_158)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_161),
.C(n_36),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_6),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_147),
.B(n_142),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_169),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_146),
.A2(n_124),
.B(n_138),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_166),
.A2(n_168),
.B(n_157),
.Y(n_175)
);

FAx1_ASAP7_75t_SL g169 ( 
.A(n_145),
.B(n_138),
.CI(n_9),
.CON(n_169),
.SN(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_170),
.Y(n_172)
);

AOI221xp5_ASAP7_75t_L g171 ( 
.A1(n_149),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.C(n_13),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_171),
.B(n_151),
.Y(n_176)
);

XOR2x2_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_144),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_173),
.A2(n_175),
.B(n_177),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_165),
.A2(n_163),
.B1(n_167),
.B2(n_144),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_158),
.B1(n_148),
.B2(n_151),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_176),
.A2(n_171),
.B(n_153),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_154),
.B(n_152),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_181),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_172),
.B(n_156),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_182),
.A2(n_176),
.B1(n_178),
.B2(n_162),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_179),
.B(n_155),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_185),
.A2(n_183),
.B(n_152),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_32),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_33),
.B(n_34),
.Y(n_188)
);

OAI321xp33_ASAP7_75t_L g189 ( 
.A1(n_188),
.A2(n_11),
.A3(n_13),
.B1(n_15),
.B2(n_16),
.C(n_155),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_15),
.Y(n_190)
);


endmodule