module fake_jpeg_6504_n_258 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_258);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_258;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_7),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_33),
.B(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_38),
.B1(n_41),
.B2(n_32),
.Y(n_51)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_7),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

CKINVDCx9p33_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_42),
.B(n_49),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_43),
.B(n_45),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_37),
.B1(n_28),
.B2(n_25),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_18),
.B1(n_27),
.B2(n_29),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_29),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_29),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_53),
.Y(n_79)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_0),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_26),
.B1(n_27),
.B2(n_20),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_58),
.A2(n_60),
.B1(n_18),
.B2(n_24),
.Y(n_84)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_38),
.A2(n_24),
.B1(n_23),
.B2(n_20),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_34),
.A2(n_19),
.B(n_16),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_61),
.A2(n_11),
.B1(n_8),
.B2(n_9),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_63),
.B(n_36),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_63),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_64),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_65),
.A2(n_54),
.B1(n_47),
.B2(n_42),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_67),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_62),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

BUFx2_ASAP7_75t_SL g107 ( 
.A(n_70),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_52),
.A2(n_36),
.B1(n_34),
.B2(n_12),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_78),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

NAND3xp33_ASAP7_75t_SL g78 ( 
.A(n_45),
.B(n_43),
.C(n_1),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_82),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_0),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_0),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_84),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_85),
.B(n_86),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_66),
.A2(n_48),
.B1(n_59),
.B2(n_46),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_87),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.Y(n_115)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_97),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_90),
.B(n_68),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_45),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_81),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_65),
.A2(n_46),
.B1(n_56),
.B2(n_54),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_75),
.A2(n_46),
.B1(n_56),
.B2(n_49),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_1),
.B(n_2),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_100),
.B(n_1),
.Y(n_131)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_104),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_78),
.A2(n_36),
.B1(n_23),
.B2(n_55),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_103),
.A2(n_71),
.B1(n_69),
.B2(n_72),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_74),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_77),
.A2(n_19),
.B1(n_2),
.B2(n_3),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_84),
.B1(n_70),
.B2(n_12),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_62),
.C(n_57),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_64),
.Y(n_114)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_83),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_112),
.B(n_113),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_120),
.B1(n_129),
.B2(n_130),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_126),
.Y(n_136)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_122),
.Y(n_155)
);

BUFx24_ASAP7_75t_SL g156 ( 
.A(n_118),
.Y(n_156)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_97),
.A2(n_67),
.B(n_68),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_134),
.B(n_100),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_89),
.B(n_83),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_128),
.B(n_131),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_62),
.Y(n_127)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_98),
.A2(n_72),
.B1(n_70),
.B2(n_62),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_91),
.A2(n_76),
.B1(n_82),
.B2(n_3),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_91),
.A2(n_76),
.B1(n_82),
.B2(n_3),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_92),
.B(n_110),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_111),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_2),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_133),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_94),
.A2(n_3),
.B(n_4),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_108),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_144),
.C(n_112),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_95),
.B1(n_93),
.B2(n_105),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_138),
.A2(n_115),
.B1(n_126),
.B2(n_128),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_125),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_142),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_115),
.A2(n_105),
.B1(n_103),
.B2(n_99),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_141),
.Y(n_158)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_123),
.A2(n_100),
.B1(n_129),
.B2(n_130),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_143),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_102),
.C(n_96),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_145),
.A2(n_147),
.B(n_154),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_110),
.B(n_106),
.Y(n_147)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_124),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_122),
.Y(n_162)
);

AND2x6_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_102),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_144),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_90),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_173),
.C(n_176),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_152),
.Y(n_160)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_162),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_132),
.Y(n_163)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_163),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_165),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_155),
.B(n_118),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_150),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_166),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_134),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_170),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_139),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_119),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_155),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_171),
.Y(n_185)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_172),
.B(n_174),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_121),
.C(n_119),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_135),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_121),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_175),
.A2(n_154),
.B(n_139),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_120),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_146),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_SL g203 ( 
.A1(n_178),
.A2(n_169),
.B(n_172),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_174),
.A2(n_135),
.B1(n_153),
.B2(n_141),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_188),
.B1(n_192),
.B2(n_158),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_182),
.A2(n_170),
.B(n_163),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_191),
.C(n_194),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_159),
.A2(n_147),
.B1(n_145),
.B2(n_148),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_175),
.B(n_153),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_159),
.A2(n_148),
.B1(n_146),
.B2(n_101),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_104),
.C(n_156),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_133),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_177),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_165),
.Y(n_196)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_196),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_SL g197 ( 
.A1(n_180),
.A2(n_161),
.B(n_162),
.C(n_158),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_197),
.A2(n_193),
.B1(n_184),
.B2(n_187),
.Y(n_211)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_177),
.C(n_167),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_198),
.A2(n_202),
.B(n_206),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_173),
.Y(n_199)
);

BUFx24_ASAP7_75t_SL g217 ( 
.A(n_199),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_204),
.C(n_208),
.Y(n_213)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_176),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_205),
.A2(n_207),
.B1(n_210),
.B2(n_178),
.Y(n_219)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_187),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_164),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_181),
.A2(n_160),
.B(n_171),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_209),
.A2(n_142),
.B1(n_88),
.B2(n_116),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_181),
.A2(n_161),
.B(n_169),
.Y(n_210)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_198),
.A2(n_193),
.B1(n_185),
.B2(n_203),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_214),
.A2(n_216),
.B(n_218),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_197),
.A2(n_184),
.B1(n_179),
.B2(n_191),
.Y(n_215)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_195),
.C(n_194),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_197),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_219),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_200),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_4),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_201),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_216),
.C(n_217),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_212),
.B(n_197),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_230),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_221),
.B(n_11),
.Y(n_230)
);

NAND3xp33_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_13),
.C(n_14),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_13),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_88),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_222),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_228),
.A2(n_218),
.B1(n_215),
.B2(n_211),
.Y(n_233)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_233),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_234),
.A2(n_238),
.B(n_237),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_235),
.B(n_236),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_214),
.C(n_109),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_239),
.A2(n_240),
.B(n_224),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_223),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_229),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_231),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_109),
.C(n_6),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_246),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_238),
.B(n_232),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_247),
.A2(n_9),
.B(n_14),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_234),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_249),
.A2(n_250),
.B(n_242),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_252),
.Y(n_255)
);

OAI21x1_ASAP7_75t_L g253 ( 
.A1(n_248),
.A2(n_109),
.B(n_9),
.Y(n_253)
);

AOI21x1_ASAP7_75t_L g254 ( 
.A1(n_253),
.A2(n_14),
.B(n_109),
.Y(n_254)
);

NOR5xp2_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_5),
.C(n_6),
.D(n_66),
.E(n_231),
.Y(n_256)
);

BUFx24_ASAP7_75t_SL g257 ( 
.A(n_256),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_255),
.Y(n_258)
);


endmodule