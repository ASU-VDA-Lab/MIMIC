module fake_aes_3903_n_31 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_31);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_31;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
INVx1_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
HB1xp67_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_7), .Y(n_14) );
INVx5_ASAP7_75t_L g15 ( .A(n_10), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_6), .Y(n_16) );
AND2x6_ASAP7_75t_L g17 ( .A(n_2), .B(n_0), .Y(n_17) );
INVx5_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_13), .B(n_0), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_18), .B(n_12), .Y(n_21) );
AND2x4_ASAP7_75t_L g22 ( .A(n_20), .B(n_16), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_23), .B(n_22), .Y(n_24) );
INVxp67_ASAP7_75t_SL g25 ( .A(n_24), .Y(n_25) );
OAI22xp5_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_21), .B1(n_14), .B2(n_15), .Y(n_26) );
NAND3xp33_ASAP7_75t_SL g27 ( .A(n_26), .B(n_21), .C(n_17), .Y(n_27) );
BUFx6f_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
OAI22xp5_ASAP7_75t_SL g29 ( .A1(n_28), .A2(n_1), .B1(n_3), .B2(n_5), .Y(n_29) );
INVx1_ASAP7_75t_SL g30 ( .A(n_29), .Y(n_30) );
AOI22xp33_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_27), .B1(n_9), .B2(n_11), .Y(n_31) );
endmodule