module fake_netlist_1_2320_n_32 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_32);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_32;
wire n_20;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_30;
wire n_16;
wire n_26;
wire n_13;
wire n_25;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_1), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_0), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_10), .Y(n_14) );
AND2x2_ASAP7_75t_L g15 ( .A(n_3), .B(n_2), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_2), .B(n_4), .Y(n_16) );
AND2x2_ASAP7_75t_SL g17 ( .A(n_14), .B(n_9), .Y(n_17) );
AND2x4_ASAP7_75t_L g18 ( .A(n_13), .B(n_14), .Y(n_18) );
NOR3xp33_ASAP7_75t_SL g19 ( .A(n_11), .B(n_0), .C(n_1), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_13), .B(n_3), .Y(n_20) );
AOI221xp5_ASAP7_75t_SL g21 ( .A1(n_20), .A2(n_12), .B1(n_15), .B2(n_16), .C(n_11), .Y(n_21) );
AOI21xp5_ASAP7_75t_L g22 ( .A1(n_18), .A2(n_15), .B(n_7), .Y(n_22) );
AOI22xp33_ASAP7_75t_L g23 ( .A1(n_17), .A2(n_5), .B1(n_6), .B2(n_8), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_18), .B(n_5), .Y(n_24) );
BUFx3_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_22), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_27), .B(n_21), .Y(n_28) );
CKINVDCx6p67_ASAP7_75t_R g29 ( .A(n_28), .Y(n_29) );
NAND4xp25_ASAP7_75t_SL g30 ( .A(n_29), .B(n_23), .C(n_19), .D(n_18), .Y(n_30) );
XNOR2x1_ASAP7_75t_L g31 ( .A(n_30), .B(n_19), .Y(n_31) );
XNOR2xp5_ASAP7_75t_L g32 ( .A(n_31), .B(n_25), .Y(n_32) );
endmodule