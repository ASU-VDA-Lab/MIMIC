module fake_jpeg_20046_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx6_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_21),
.B(n_24),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_23),
.B1(n_26),
.B2(n_14),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_10),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_20),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_1),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_25),
.B(n_3),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_11),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_23),
.A2(n_14),
.B1(n_16),
.B2(n_18),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_28),
.A2(n_35),
.B1(n_12),
.B2(n_15),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_21),
.A2(n_16),
.B(n_17),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_37),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_27),
.A2(n_12),
.B1(n_15),
.B2(n_17),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_41),
.B1(n_42),
.B2(n_28),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_24),
.B1(n_26),
.B2(n_25),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_35),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_43),
.B(n_34),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_25),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_30),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_13),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_13),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_48),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_50),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_34),
.B1(n_32),
.B2(n_18),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_47),
.A2(n_32),
.B1(n_13),
.B2(n_37),
.Y(n_53)
);

MAJx2_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_32),
.C(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_53),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_61),
.Y(n_63)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_59),
.B(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_64),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_56),
.A2(n_45),
.B(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_40),
.Y(n_65)
);

AOI322xp5_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_57),
.A3(n_61),
.B1(n_50),
.B2(n_60),
.C1(n_38),
.C2(n_29),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_39),
.B1(n_60),
.B2(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_66),
.B(n_57),
.Y(n_69)
);

NAND3xp33_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_29),
.C(n_9),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_70),
.C(n_67),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_66),
.C(n_29),
.Y(n_72)
);


endmodule