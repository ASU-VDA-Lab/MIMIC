module fake_jpeg_17925_n_301 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_301);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

BUFx12_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_24),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_29),
.Y(n_40)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_24),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_32),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_34),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_37),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_28),
.B(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_46),
.Y(n_58)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_28),
.B(n_14),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_28),
.B(n_19),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_34),
.Y(n_54)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_42),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_20),
.B(n_29),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_55),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_32),
.C(n_33),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_56),
.A2(n_74),
.B1(n_31),
.B2(n_38),
.Y(n_83)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_65),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_30),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_42),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_18),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_18),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_69),
.Y(n_88)
);

AOI22x1_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_31),
.B1(n_37),
.B2(n_32),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_67),
.A2(n_36),
.B1(n_50),
.B2(n_52),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_22),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_70),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_32),
.C(n_33),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_37),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_36),
.B1(n_27),
.B2(n_25),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_79),
.A2(n_82),
.B1(n_85),
.B2(n_86),
.Y(n_112)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_67),
.A2(n_25),
.B1(n_36),
.B2(n_30),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_74),
.Y(n_103)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_55),
.A2(n_36),
.B1(n_27),
.B2(n_25),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_89),
.B(n_98),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_97),
.Y(n_101)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_40),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_93),
.B(n_72),
.Y(n_120)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_57),
.A2(n_27),
.B1(n_19),
.B2(n_39),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_36),
.B1(n_73),
.B2(n_60),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_76),
.B1(n_60),
.B2(n_73),
.Y(n_125)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_108),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_120),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_58),
.Y(n_105)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_75),
.Y(n_106)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_93),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_20),
.B(n_37),
.Y(n_138)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_113),
.Y(n_124)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_94),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_115),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_71),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_72),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_117),
.B(n_121),
.Y(n_143)
);

BUFx24_ASAP7_75t_SL g118 ( 
.A(n_92),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_22),
.Y(n_139)
);

NOR2x1_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_31),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_122),
.B(n_139),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_129),
.B1(n_113),
.B2(n_102),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_121),
.A2(n_91),
.B1(n_85),
.B2(n_98),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_126),
.A2(n_130),
.B(n_134),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_127),
.Y(n_148)
);

AO21x2_ASAP7_75t_SL g129 ( 
.A1(n_112),
.A2(n_97),
.B(n_84),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_110),
.A2(n_89),
.B(n_30),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_99),
.A2(n_45),
.B(n_41),
.C(n_76),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_133),
.A2(n_135),
.B1(n_140),
.B2(n_104),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_78),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_110),
.A2(n_78),
.B1(n_96),
.B2(n_41),
.Y(n_135)
);

AO22x1_ASAP7_75t_L g136 ( 
.A1(n_119),
.A2(n_37),
.B1(n_68),
.B2(n_63),
.Y(n_136)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_138),
.A2(n_141),
.B(n_26),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_SL g140 ( 
.A1(n_116),
.A2(n_37),
.B(n_81),
.C(n_35),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_34),
.B(n_21),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_34),
.Y(n_142)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_20),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_64),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_87),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_146),
.B(n_17),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_147),
.A2(n_151),
.B1(n_171),
.B2(n_133),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_149),
.A2(n_157),
.B1(n_166),
.B2(n_136),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_116),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_150),
.A2(n_156),
.B(n_172),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_104),
.B1(n_100),
.B2(n_111),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_130),
.B(n_100),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_152),
.B(n_154),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_144),
.B(n_23),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_0),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_129),
.A2(n_21),
.B1(n_23),
.B2(n_19),
.Y(n_157)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_124),
.Y(n_159)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_70),
.Y(n_160)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_20),
.Y(n_161)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_61),
.Y(n_162)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_132),
.Y(n_163)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_163),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_168),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_129),
.A2(n_21),
.B1(n_26),
.B2(n_61),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_122),
.B(n_15),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_169),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_141),
.B(n_136),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_133),
.A2(n_64),
.B1(n_17),
.B2(n_33),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_0),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_17),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_128),
.C(n_138),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_186),
.C(n_190),
.Y(n_201)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_182),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_134),
.B(n_133),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_195),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_166),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_183),
.A2(n_189),
.B1(n_168),
.B2(n_172),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_128),
.C(n_134),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_149),
.A2(n_140),
.B1(n_1),
.B2(n_2),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_33),
.C(n_140),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_140),
.C(n_37),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_155),
.C(n_158),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_17),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_198),
.Y(n_202)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

MAJx2_ASAP7_75t_L g196 ( 
.A(n_156),
.B(n_15),
.C(n_13),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_196),
.B(n_172),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_150),
.B(n_0),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_208),
.C(n_212),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_154),
.Y(n_204)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_165),
.Y(n_205)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_206),
.A2(n_189),
.B1(n_194),
.B2(n_178),
.Y(n_226)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_152),
.C(n_170),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_148),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_209),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_214),
.Y(n_220)
);

AND2x6_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_156),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_211),
.A2(n_193),
.B(n_180),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_153),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_157),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_215),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_35),
.C(n_15),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_201),
.C(n_214),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_8),
.Y(n_217)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_217),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_13),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_218),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_221),
.A2(n_7),
.B1(n_12),
.B2(n_11),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_199),
.A2(n_176),
.B(n_188),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_176),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_200),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_192),
.Y(n_227)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_203),
.A2(n_188),
.B1(n_190),
.B2(n_198),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_231),
.A2(n_234),
.B1(n_1),
.B2(n_2),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_211),
.A2(n_184),
.B1(n_182),
.B2(n_196),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_201),
.Y(n_241)
);

XNOR2x2_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_184),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_236),
.A2(n_10),
.B1(n_12),
.B2(n_6),
.Y(n_251)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_228),
.B(n_208),
.Y(n_238)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_219),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_242),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_243),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_229),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_216),
.C(n_9),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_235),
.C(n_221),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_220),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_250),
.Y(n_262)
);

AO22x1_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_247)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_249),
.A2(n_232),
.B1(n_225),
.B2(n_224),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_251),
.A2(n_228),
.B1(n_222),
.B2(n_230),
.Y(n_257)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_239),
.A2(n_249),
.B1(n_248),
.B2(n_244),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_255),
.B(n_263),
.Y(n_273)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_257),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_245),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_259),
.B(n_1),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_248),
.A2(n_234),
.B1(n_226),
.B2(n_231),
.Y(n_261)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_261),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_220),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_6),
.C(n_5),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_265),
.B(n_266),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_258),
.C(n_255),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_6),
.C(n_5),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_269),
.Y(n_276)
);

AO21x1_ASAP7_75t_L g268 ( 
.A1(n_256),
.A2(n_260),
.B(n_262),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_268),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_5),
.C(n_13),
.Y(n_269)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_270),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_13),
.C(n_15),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_273),
.Y(n_278)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_275),
.B(n_257),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_280),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_272),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_13),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_3),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_283),
.C(n_15),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_271),
.A2(n_3),
.B(n_4),
.Y(n_283)
);

NAND3xp33_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_287),
.C(n_276),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_284),
.A2(n_3),
.B(n_4),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_286),
.A2(n_280),
.B(n_35),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_15),
.Y(n_287)
);

AOI21x1_ASAP7_75t_L g292 ( 
.A1(n_288),
.A2(n_282),
.B(n_279),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_292),
.C(n_293),
.Y(n_294)
);

OAI21xp33_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_290),
.B(n_289),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_295),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_289),
.C(n_35),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_297),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_35),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_299),
.B(n_35),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_35),
.C(n_148),
.Y(n_301)
);


endmodule