module fake_jpeg_10571_n_297 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_39),
.Y(n_47)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_19),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_42),
.B1(n_26),
.B2(n_21),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_32),
.Y(n_53)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_53),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_51),
.A2(n_33),
.B1(n_29),
.B2(n_66),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_56),
.Y(n_83)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_26),
.B1(n_21),
.B2(n_18),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_69),
.B1(n_26),
.B2(n_21),
.Y(n_70)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_60),
.Y(n_84)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_62),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_35),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_68),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_64),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_67),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_35),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_37),
.A2(n_26),
.B1(n_21),
.B2(n_18),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_70),
.A2(n_82),
.B1(n_99),
.B2(n_101),
.Y(n_132)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_71),
.B(n_76),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_18),
.B1(n_34),
.B2(n_23),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_73),
.A2(n_79),
.B1(n_97),
.B2(n_1),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_34),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_75),
.B(n_80),
.Y(n_120)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_55),
.A2(n_18),
.B1(n_34),
.B2(n_23),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_45),
.B(n_44),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_55),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_81),
.B(n_87),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_66),
.A2(n_32),
.B1(n_27),
.B2(n_23),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_64),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_64),
.A2(n_32),
.B(n_33),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_90),
.B(n_95),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_29),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_29),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_91),
.B(n_92),
.Y(n_123)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_96),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_33),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_22),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_50),
.A2(n_27),
.B1(n_30),
.B2(n_24),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_50),
.A2(n_30),
.B1(n_24),
.B2(n_17),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_56),
.A2(n_24),
.B1(n_30),
.B2(n_17),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_59),
.A2(n_19),
.B1(n_31),
.B2(n_20),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_102),
.A2(n_20),
.B1(n_28),
.B2(n_25),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_63),
.A2(n_44),
.B1(n_43),
.B2(n_25),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_105),
.A2(n_25),
.B1(n_22),
.B2(n_31),
.Y(n_114)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_106),
.B(n_121),
.Y(n_154)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_110),
.B(n_116),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_0),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_98),
.Y(n_135)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_70),
.A2(n_43),
.B(n_25),
.C(n_31),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_112),
.A2(n_128),
.B1(n_133),
.B2(n_103),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_114),
.A2(n_115),
.B1(n_117),
.B2(n_122),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_71),
.A2(n_20),
.B1(n_19),
.B2(n_31),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_73),
.A2(n_78),
.B1(n_94),
.B2(n_83),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_0),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_118),
.A2(n_76),
.B(n_101),
.Y(n_164)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_124),
.B(n_126),
.Y(n_156)
);

NOR3xp33_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_28),
.C(n_25),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_13),
.Y(n_163)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_80),
.A2(n_20),
.B1(n_25),
.B2(n_28),
.Y(n_128)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_129),
.Y(n_142)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

AO21x1_ASAP7_75t_L g137 ( 
.A1(n_130),
.A2(n_88),
.B(n_90),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_131),
.Y(n_140)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_134),
.B(n_137),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_135),
.B(n_136),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_110),
.B(n_86),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_138),
.B(n_141),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_96),
.C(n_104),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_139),
.B(n_87),
.C(n_77),
.Y(n_182)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_104),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_145),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_129),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_146),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_95),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_107),
.A2(n_85),
.B(n_95),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_164),
.B(n_151),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_97),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_151),
.Y(n_180)
);

MAJx2_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_105),
.C(n_79),
.Y(n_150)
);

XNOR2x1_ASAP7_75t_L g193 ( 
.A(n_150),
.B(n_74),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_105),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_155),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_153),
.A2(n_89),
.B1(n_74),
.B2(n_93),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_131),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_112),
.A2(n_81),
.B1(n_103),
.B2(n_105),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_158),
.A2(n_114),
.B1(n_128),
.B2(n_108),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_115),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_160),
.Y(n_189)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_111),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_161),
.B(n_1),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_105),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_162),
.A2(n_1),
.B(n_2),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_SL g170 ( 
.A1(n_163),
.A2(n_119),
.B(n_14),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_156),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_166),
.Y(n_207)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_167),
.A2(n_194),
.B(n_164),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_168),
.A2(n_184),
.B1(n_142),
.B2(n_144),
.Y(n_208)
);

AOI322xp5_ASAP7_75t_SL g169 ( 
.A1(n_138),
.A2(n_116),
.A3(n_118),
.B1(n_119),
.B2(n_108),
.C1(n_126),
.C2(n_124),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_170),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_132),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_172),
.B(n_176),
.C(n_182),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_156),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_174),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_149),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_160),
.A2(n_106),
.B1(n_121),
.B2(n_92),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_175),
.A2(n_158),
.B1(n_159),
.B2(n_153),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_72),
.Y(n_176)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_183),
.B(n_188),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_143),
.Y(n_185)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_89),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_186),
.B(n_164),
.Y(n_198)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_136),
.Y(n_188)
);

AO21x1_ASAP7_75t_L g190 ( 
.A1(n_135),
.A2(n_77),
.B(n_89),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_190),
.A2(n_191),
.B(n_193),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_140),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_161),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_193),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_195),
.B(n_197),
.Y(n_232)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_204),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_199),
.A2(n_178),
.B1(n_174),
.B2(n_183),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_212),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_181),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_201),
.B(n_202),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_185),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_157),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_189),
.A2(n_143),
.B1(n_157),
.B2(n_150),
.Y(n_205)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

OAI21xp33_ASAP7_75t_L g206 ( 
.A1(n_177),
.A2(n_152),
.B(n_137),
.Y(n_206)
);

AOI322xp5_ASAP7_75t_L g235 ( 
.A1(n_206),
.A2(n_190),
.A3(n_180),
.B1(n_142),
.B2(n_192),
.C1(n_140),
.C2(n_8),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_208),
.A2(n_210),
.B1(n_218),
.B2(n_194),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_168),
.A2(n_150),
.B1(n_137),
.B2(n_134),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_179),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_213),
.B(n_191),
.Y(n_228)
);

AO21x1_ASAP7_75t_L g220 ( 
.A1(n_214),
.A2(n_216),
.B(n_171),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_167),
.A2(n_162),
.B(n_141),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_171),
.A2(n_162),
.B(n_155),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_186),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_227),
.C(n_230),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_220),
.B(n_224),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_221),
.A2(n_223),
.B1(n_236),
.B2(n_210),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_201),
.A2(n_165),
.B1(n_188),
.B2(n_190),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_213),
.B(n_178),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_182),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_228),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_229),
.A2(n_209),
.B(n_205),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_176),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_203),
.B(n_207),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_234),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_212),
.B(n_166),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_211),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_199),
.A2(n_180),
.B1(n_140),
.B2(n_5),
.Y(n_236)
);

MAJx2_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_9),
.C(n_14),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_214),
.Y(n_240)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_215),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_240),
.B(n_221),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_230),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_244),
.A2(n_247),
.B(n_252),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_204),
.C(n_218),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_249),
.C(n_250),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_222),
.A2(n_202),
.B1(n_196),
.B2(n_197),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_246),
.A2(n_236),
.B1(n_226),
.B2(n_231),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_209),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_237),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_196),
.C(n_195),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_208),
.C(n_211),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_238),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_232),
.A2(n_200),
.B(n_4),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_222),
.A2(n_3),
.B(n_4),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_253),
.A2(n_3),
.B(n_4),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_259),
.Y(n_276)
);

OAI31xp33_ASAP7_75t_L g256 ( 
.A1(n_247),
.A2(n_220),
.A3(n_231),
.B(n_223),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_256),
.A2(n_266),
.B(n_5),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_258),
.B(n_249),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_263),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_254),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_252),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_246),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_248),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_241),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_265),
.A2(n_253),
.B1(n_244),
.B2(n_250),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_10),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_267),
.B(n_240),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_268),
.B(n_269),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_271),
.B(n_273),
.Y(n_282)
);

AND2x4_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_5),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_242),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_258),
.B(n_245),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_275),
.B(n_264),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_242),
.C(n_6),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_277),
.A2(n_6),
.B(n_7),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_272),
.A2(n_256),
.B1(n_257),
.B2(n_262),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_L g288 ( 
.A1(n_278),
.A2(n_284),
.B1(n_10),
.B2(n_11),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_279),
.B(n_281),
.Y(n_286)
);

OAI221xp5_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_265),
.B1(n_266),
.B2(n_257),
.C(n_8),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_283),
.A2(n_11),
.B(n_12),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_7),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_11),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_288),
.A2(n_289),
.B(n_282),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_276),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_284),
.B(n_278),
.Y(n_291)
);

OAI321xp33_ASAP7_75t_L g295 ( 
.A1(n_291),
.A2(n_292),
.A3(n_293),
.B1(n_12),
.B2(n_16),
.C(n_274),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_292),
.B(n_277),
.C(n_286),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_295),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_12),
.Y(n_297)
);


endmodule