module real_aes_9502_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_1380;
wire n_488;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1004;
wire n_580;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_720;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_1463;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_1172;
wire n_459;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_769;
wire n_434;
wire n_250;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1151;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1352;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
CKINVDCx5p33_ASAP7_75t_R g926 ( .A(n_0), .Y(n_926) );
AO221x1_ASAP7_75t_L g1203 ( .A1(n_1), .A2(n_149), .B1(n_1176), .B2(n_1204), .C(n_1206), .Y(n_1203) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_2), .A2(n_67), .B1(n_806), .B2(n_807), .Y(n_805) );
INVx1_ASAP7_75t_L g841 ( .A(n_2), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_3), .A2(n_234), .B1(n_892), .B2(n_893), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_3), .A2(n_234), .B1(n_901), .B2(n_902), .Y(n_900) );
AO22x2_ASAP7_75t_L g642 ( .A1(n_4), .A2(n_643), .B1(n_697), .B2(n_698), .Y(n_642) );
INVxp67_ASAP7_75t_L g697 ( .A(n_4), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_5), .A2(n_202), .B1(n_283), .B2(n_291), .Y(n_282) );
INVx1_ASAP7_75t_L g405 ( .A(n_5), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_6), .A2(n_213), .B1(n_687), .B2(n_723), .Y(n_1041) );
INVx1_ASAP7_75t_L g1049 ( .A(n_6), .Y(n_1049) );
CKINVDCx5p33_ASAP7_75t_R g943 ( .A(n_7), .Y(n_943) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_8), .Y(n_261) );
INVx1_ASAP7_75t_L g449 ( .A(n_8), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_8), .B(n_178), .Y(n_491) );
AND2x2_ASAP7_75t_L g495 ( .A(n_8), .B(n_287), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g1104 ( .A(n_9), .Y(n_1104) );
CKINVDCx5p33_ASAP7_75t_R g868 ( .A(n_10), .Y(n_868) );
AOI22xp5_ASAP7_75t_L g1185 ( .A1(n_11), .A2(n_117), .B1(n_1176), .B2(n_1180), .Y(n_1185) );
INVx1_ASAP7_75t_L g592 ( .A(n_12), .Y(n_592) );
OAI22xp33_ASAP7_75t_L g627 ( .A1(n_12), .A2(n_137), .B1(n_628), .B2(n_631), .Y(n_627) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_13), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g942 ( .A(n_14), .Y(n_942) );
INVx1_ASAP7_75t_L g1022 ( .A(n_15), .Y(n_1022) );
OAI22xp5_ASAP7_75t_L g1046 ( .A1(n_15), .A2(n_74), .B1(n_981), .B2(n_1047), .Y(n_1046) );
XNOR2x2_ASAP7_75t_L g452 ( .A(n_16), .B(n_453), .Y(n_452) );
AOI22xp33_ASAP7_75t_SL g1375 ( .A1(n_17), .A2(n_211), .B1(n_477), .B2(n_599), .Y(n_1375) );
AOI221xp5_ASAP7_75t_L g1411 ( .A1(n_17), .A2(n_72), .B1(n_359), .B2(n_513), .C(n_1412), .Y(n_1411) );
CKINVDCx5p33_ASAP7_75t_R g1069 ( .A(n_18), .Y(n_1069) );
AOI21xp33_ASAP7_75t_L g476 ( .A1(n_19), .A2(n_477), .B(n_478), .Y(n_476) );
INVx1_ASAP7_75t_L g556 ( .A(n_19), .Y(n_556) );
INVxp67_ASAP7_75t_SL g577 ( .A(n_20), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_20), .A2(n_219), .B1(n_612), .B2(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g984 ( .A(n_21), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_21), .A2(n_176), .B1(n_723), .B2(n_725), .Y(n_1012) );
AO221x2_ASAP7_75t_L g1324 ( .A1(n_22), .A2(n_158), .B1(n_1204), .B2(n_1325), .C(n_1327), .Y(n_1324) );
AOI22xp33_ASAP7_75t_L g1376 ( .A1(n_23), .A2(n_72), .B1(n_1377), .B2(n_1379), .Y(n_1376) );
AOI22xp33_ASAP7_75t_L g1414 ( .A1(n_23), .A2(n_211), .B1(n_618), .B2(n_1415), .Y(n_1414) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_24), .A2(n_44), .B1(n_336), .B2(n_344), .Y(n_335) );
INVx1_ASAP7_75t_L g437 ( .A(n_24), .Y(n_437) );
INVx2_ASAP7_75t_L g330 ( .A(n_25), .Y(n_330) );
OR2x2_ASAP7_75t_L g555 ( .A(n_25), .B(n_540), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_26), .A2(n_151), .B1(n_493), .B2(n_499), .Y(n_492) );
INVx1_ASAP7_75t_L g531 ( .A(n_26), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_27), .Y(n_480) );
AOI22xp33_ASAP7_75t_SL g604 ( .A1(n_28), .A2(n_77), .B1(n_601), .B2(n_605), .Y(n_604) );
INVxp33_ASAP7_75t_L g638 ( .A(n_28), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_29), .A2(n_195), .B1(n_723), .B2(n_725), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g849 ( .A1(n_29), .A2(n_195), .B1(n_499), .B2(n_781), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_30), .A2(n_99), .B1(n_993), .B2(n_994), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_30), .A2(n_99), .B1(n_1009), .B2(n_1036), .Y(n_1035) );
INVx1_ASAP7_75t_L g1369 ( .A(n_31), .Y(n_1369) );
OAI221xp5_ASAP7_75t_L g1398 ( .A1(n_31), .A2(n_54), .B1(n_1399), .B2(n_1401), .C(n_1403), .Y(n_1398) );
BUFx2_ASAP7_75t_L g278 ( .A(n_32), .Y(n_278) );
BUFx2_ASAP7_75t_L g376 ( .A(n_32), .Y(n_376) );
INVx1_ASAP7_75t_L g447 ( .A(n_32), .Y(n_447) );
OR2x2_ASAP7_75t_L g1078 ( .A(n_32), .B(n_491), .Y(n_1078) );
INVx1_ASAP7_75t_L g585 ( .A(n_33), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_33), .A2(n_61), .B1(n_618), .B2(n_619), .Y(n_617) );
OAI221xp5_ASAP7_75t_L g652 ( .A1(n_34), .A2(n_209), .B1(n_631), .B2(n_653), .C(n_654), .Y(n_652) );
INVx1_ASAP7_75t_L g664 ( .A(n_34), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_35), .A2(n_101), .B1(n_615), .B2(n_918), .Y(n_917) );
AOI221xp5_ASAP7_75t_L g936 ( .A1(n_35), .A2(n_101), .B1(n_415), .B2(n_481), .C(n_937), .Y(n_936) );
OAI22xp33_ASAP7_75t_L g503 ( .A1(n_36), .A2(n_42), .B1(n_504), .B2(n_506), .Y(n_503) );
AOI221xp5_ASAP7_75t_L g524 ( .A1(n_36), .A2(n_42), .B1(n_513), .B2(n_525), .C(n_527), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g1466 ( .A1(n_37), .A2(n_231), .B1(n_1464), .B2(n_1467), .Y(n_1466) );
INVxp67_ASAP7_75t_SL g1472 ( .A(n_37), .Y(n_1472) );
INVx1_ASAP7_75t_L g752 ( .A(n_38), .Y(n_752) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_38), .A2(n_56), .B1(n_788), .B2(n_790), .Y(n_787) );
CKINVDCx5p33_ASAP7_75t_R g927 ( .A(n_39), .Y(n_927) );
XNOR2xp5_ASAP7_75t_L g792 ( .A(n_40), .B(n_793), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g1381 ( .A1(n_41), .A2(n_53), .B1(n_607), .B2(n_831), .Y(n_1381) );
INVx1_ASAP7_75t_L g1419 ( .A(n_41), .Y(n_1419) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_43), .Y(n_459) );
INVx1_ASAP7_75t_L g315 ( .A(n_44), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_45), .A2(n_78), .B1(n_601), .B2(n_603), .Y(n_600) );
AOI22xp33_ASAP7_75t_SL g611 ( .A1(n_45), .A2(n_78), .B1(n_612), .B2(n_613), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_46), .A2(n_241), .B1(n_996), .B2(n_997), .Y(n_995) );
AOI22xp33_ASAP7_75t_SL g1007 ( .A1(n_46), .A2(n_241), .B1(n_736), .B2(n_804), .Y(n_1007) );
AOI22xp33_ASAP7_75t_SL g923 ( .A1(n_47), .A2(n_244), .B1(n_558), .B2(n_613), .Y(n_923) );
INVx1_ASAP7_75t_L g931 ( .A(n_47), .Y(n_931) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_48), .Y(n_384) );
INVx1_ASAP7_75t_L g1027 ( .A(n_49), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_49), .A2(n_220), .B1(n_847), .B2(n_1000), .Y(n_1032) );
INVx1_ASAP7_75t_L g965 ( .A(n_50), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_50), .A2(n_143), .B1(n_847), .B2(n_1000), .Y(n_999) );
INVx1_ASAP7_75t_L g1207 ( .A(n_51), .Y(n_1207) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_52), .Y(n_462) );
INVx1_ASAP7_75t_L g1410 ( .A(n_53), .Y(n_1410) );
INVx1_ASAP7_75t_L g1371 ( .A(n_54), .Y(n_1371) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_55), .A2(n_89), .B1(n_598), .B2(n_607), .Y(n_606) );
INVxp67_ASAP7_75t_SL g626 ( .A(n_55), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g756 ( .A1(n_56), .A2(n_65), .B1(n_598), .B2(n_607), .C(n_757), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_57), .A2(n_141), .B1(n_723), .B2(n_725), .Y(n_722) );
INVx1_ASAP7_75t_L g774 ( .A(n_57), .Y(n_774) );
INVx1_ASAP7_75t_L g970 ( .A(n_58), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_58), .A2(n_115), .B1(n_586), .B2(n_1004), .Y(n_1003) );
AOI22xp33_ASAP7_75t_SL g1452 ( .A1(n_59), .A2(n_111), .B1(n_588), .B2(n_1453), .Y(n_1452) );
AOI22xp33_ASAP7_75t_L g1463 ( .A1(n_59), .A2(n_111), .B1(n_1464), .B2(n_1465), .Y(n_1463) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_60), .Y(n_470) );
INVxp33_ASAP7_75t_L g580 ( .A(n_61), .Y(n_580) );
AO22x2_ASAP7_75t_L g1013 ( .A1(n_62), .A2(n_1014), .B1(n_1053), .B2(n_1054), .Y(n_1013) );
INVxp67_ASAP7_75t_SL g1053 ( .A(n_62), .Y(n_1053) );
AO221x1_ASAP7_75t_L g940 ( .A1(n_63), .A2(n_84), .B1(n_477), .B2(n_478), .C(n_608), .Y(n_940) );
INVx1_ASAP7_75t_L g951 ( .A(n_63), .Y(n_951) );
CKINVDCx5p33_ASAP7_75t_R g819 ( .A(n_64), .Y(n_819) );
OAI22xp5_ASAP7_75t_L g785 ( .A1(n_65), .A2(n_175), .B1(n_566), .B2(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g875 ( .A(n_66), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_66), .A2(n_131), .B1(n_612), .B2(n_902), .Y(n_905) );
INVx1_ASAP7_75t_L g838 ( .A(n_67), .Y(n_838) );
INVx1_ASAP7_75t_L g1062 ( .A(n_68), .Y(n_1062) );
AOI221xp5_ASAP7_75t_L g1121 ( .A1(n_68), .A2(n_130), .B1(n_1039), .B2(n_1122), .C(n_1124), .Y(n_1121) );
INVx1_ASAP7_75t_L g1208 ( .A(n_69), .Y(n_1208) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_70), .A2(n_215), .B1(n_551), .B2(n_810), .Y(n_809) );
OAI211xp5_ASAP7_75t_SL g823 ( .A1(n_70), .A2(n_506), .B(n_824), .C(n_834), .Y(n_823) );
INVx1_ASAP7_75t_L g662 ( .A(n_71), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_71), .A2(n_188), .B1(n_558), .B2(n_687), .Y(n_696) );
INVxp67_ASAP7_75t_SL g1439 ( .A(n_73), .Y(n_1439) );
AOI22xp33_ASAP7_75t_SL g1456 ( .A1(n_73), .A2(n_107), .B1(n_994), .B2(n_1453), .Y(n_1456) );
INVx1_ASAP7_75t_L g1024 ( .A(n_74), .Y(n_1024) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_75), .A2(n_198), .B1(n_601), .B2(n_675), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_75), .A2(n_198), .B1(n_612), .B2(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g877 ( .A(n_76), .Y(n_877) );
AOI22xp33_ASAP7_75t_SL g904 ( .A1(n_76), .A2(n_182), .B1(n_513), .B2(n_695), .Y(n_904) );
INVxp67_ASAP7_75t_SL g639 ( .A(n_77), .Y(n_639) );
INVx1_ASAP7_75t_L g871 ( .A(n_79), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_79), .A2(n_125), .B1(n_601), .B2(n_888), .Y(n_887) );
XNOR2x2_ASAP7_75t_L g960 ( .A(n_80), .B(n_961), .Y(n_960) );
AO221x1_ASAP7_75t_L g1187 ( .A1(n_80), .A2(n_121), .B1(n_1176), .B2(n_1180), .C(n_1188), .Y(n_1187) );
INVx1_ASAP7_75t_L g1329 ( .A(n_81), .Y(n_1329) );
AOI22xp33_ASAP7_75t_L g1469 ( .A1(n_82), .A2(n_118), .B1(n_723), .B2(n_725), .Y(n_1469) );
INVxp33_ASAP7_75t_SL g1475 ( .A(n_82), .Y(n_1475) );
INVx1_ASAP7_75t_L g816 ( .A(n_83), .Y(n_816) );
AOI221xp5_ASAP7_75t_L g830 ( .A1(n_83), .A2(n_161), .B1(n_608), .B2(n_757), .C(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g953 ( .A(n_84), .Y(n_953) );
INVx1_ASAP7_75t_L g1088 ( .A(n_85), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g1137 ( .A1(n_85), .A2(n_242), .B1(n_1138), .B2(n_1140), .Y(n_1137) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_86), .Y(n_396) );
AO22x2_ASAP7_75t_L g857 ( .A1(n_87), .A2(n_858), .B1(n_859), .B2(n_908), .Y(n_857) );
INVxp67_ASAP7_75t_SL g858 ( .A(n_87), .Y(n_858) );
AO221x1_ASAP7_75t_L g1192 ( .A1(n_87), .A2(n_154), .B1(n_1176), .B2(n_1180), .C(n_1193), .Y(n_1192) );
OAI222xp33_ASAP7_75t_L g862 ( .A1(n_88), .A2(n_162), .B1(n_196), .B2(n_628), .C1(n_631), .C2(n_863), .Y(n_862) );
INVx1_ASAP7_75t_L g878 ( .A(n_88), .Y(n_878) );
INVxp33_ASAP7_75t_L g633 ( .A(n_89), .Y(n_633) );
INVx1_ASAP7_75t_L g374 ( .A(n_90), .Y(n_374) );
INVx1_ASAP7_75t_L g540 ( .A(n_90), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_91), .A2(n_104), .B1(n_677), .B2(n_896), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_91), .A2(n_104), .B1(n_513), .B2(n_615), .Y(n_899) );
CKINVDCx5p33_ASAP7_75t_R g945 ( .A(n_92), .Y(n_945) );
INVx1_ASAP7_75t_L g1195 ( .A(n_93), .Y(n_1195) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_94), .A2(n_95), .B1(n_542), .B2(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g760 ( .A(n_94), .Y(n_760) );
INVx1_ASAP7_75t_L g763 ( .A(n_95), .Y(n_763) );
AOI22x1_ASAP7_75t_L g910 ( .A1(n_96), .A2(n_911), .B1(n_912), .B2(n_954), .Y(n_910) );
INVxp67_ASAP7_75t_SL g954 ( .A(n_96), .Y(n_954) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_97), .Y(n_393) );
INVx1_ASAP7_75t_L g867 ( .A(n_98), .Y(n_867) );
AOI22xp33_ASAP7_75t_SL g885 ( .A1(n_98), .A2(n_196), .B1(n_677), .B2(n_886), .Y(n_885) );
CKINVDCx5p33_ASAP7_75t_R g798 ( .A(n_100), .Y(n_798) );
CKINVDCx5p33_ASAP7_75t_R g797 ( .A(n_102), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_103), .A2(n_160), .B1(n_803), .B2(n_804), .Y(n_802) );
INVx1_ASAP7_75t_L g843 ( .A(n_103), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g1219 ( .A1(n_105), .A2(n_200), .B1(n_1176), .B2(n_1180), .Y(n_1219) );
INVx1_ASAP7_75t_L g730 ( .A(n_106), .Y(n_730) );
OAI221xp5_ASAP7_75t_L g766 ( .A1(n_106), .A2(n_504), .B1(n_767), .B2(n_770), .C(n_779), .Y(n_766) );
INVxp33_ASAP7_75t_SL g1433 ( .A(n_107), .Y(n_1433) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_108), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g435 ( .A(n_108), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_109), .A2(n_237), .B1(n_598), .B2(n_599), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_109), .A2(n_237), .B1(n_355), .B2(n_615), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_110), .A2(n_163), .B1(n_513), .B2(n_920), .Y(n_919) );
OAI221xp5_ASAP7_75t_L g939 ( .A1(n_110), .A2(n_506), .B1(n_940), .B2(n_941), .C(n_944), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_112), .A2(n_192), .B1(n_902), .B2(n_916), .Y(n_915) );
AOI22xp33_ASAP7_75t_SL g934 ( .A1(n_112), .A2(n_192), .B1(n_848), .B2(n_935), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_113), .A2(n_218), .B1(n_996), .B2(n_997), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_113), .A2(n_218), .B1(n_687), .B2(n_1039), .Y(n_1038) );
INVx1_ASAP7_75t_L g1190 ( .A(n_114), .Y(n_1190) );
INVx1_ASAP7_75t_L g964 ( .A(n_115), .Y(n_964) );
INVx1_ASAP7_75t_L g253 ( .A(n_116), .Y(n_253) );
OA22x2_ASAP7_75t_L g275 ( .A1(n_117), .A2(n_276), .B1(n_450), .B2(n_451), .Y(n_275) );
INVxp67_ASAP7_75t_SL g451 ( .A(n_117), .Y(n_451) );
INVxp67_ASAP7_75t_SL g1476 ( .A(n_118), .Y(n_1476) );
CKINVDCx5p33_ASAP7_75t_R g1017 ( .A(n_119), .Y(n_1017) );
AOI22xp5_ASAP7_75t_L g1168 ( .A1(n_120), .A2(n_179), .B1(n_1169), .B2(n_1172), .Y(n_1168) );
INVx1_ASAP7_75t_L g1189 ( .A(n_122), .Y(n_1189) );
INVx1_ASAP7_75t_L g655 ( .A(n_123), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_123), .A2(n_140), .B1(n_598), .B2(n_678), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g1380 ( .A1(n_124), .A2(n_171), .B1(n_601), .B2(n_893), .Y(n_1380) );
INVx1_ASAP7_75t_L g1420 ( .A(n_124), .Y(n_1420) );
INVx1_ASAP7_75t_L g870 ( .A(n_125), .Y(n_870) );
CKINVDCx5p33_ASAP7_75t_R g1110 ( .A(n_126), .Y(n_1110) );
CKINVDCx5p33_ASAP7_75t_R g1098 ( .A(n_127), .Y(n_1098) );
INVx1_ASAP7_75t_L g979 ( .A(n_128), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_128), .A2(n_181), .B1(n_806), .B2(n_807), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_129), .A2(n_223), .B1(n_806), .B2(n_1036), .Y(n_1040) );
INVx1_ASAP7_75t_L g1052 ( .A(n_129), .Y(n_1052) );
INVx1_ASAP7_75t_L g1071 ( .A(n_130), .Y(n_1071) );
INVx1_ASAP7_75t_L g874 ( .A(n_131), .Y(n_874) );
CKINVDCx5p33_ASAP7_75t_R g485 ( .A(n_132), .Y(n_485) );
OAI221xp5_ASAP7_75t_L g532 ( .A1(n_132), .A2(n_533), .B1(n_541), .B2(n_542), .C(n_545), .Y(n_532) );
CKINVDCx5p33_ASAP7_75t_R g1102 ( .A(n_133), .Y(n_1102) );
AOI22xp5_ASAP7_75t_L g1175 ( .A1(n_134), .A2(n_165), .B1(n_1176), .B2(n_1180), .Y(n_1175) );
AOI22xp5_ASAP7_75t_L g1220 ( .A1(n_135), .A2(n_246), .B1(n_1169), .B2(n_1172), .Y(n_1220) );
CKINVDCx5p33_ASAP7_75t_R g1385 ( .A(n_136), .Y(n_1385) );
INVxp67_ASAP7_75t_SL g589 ( .A(n_137), .Y(n_589) );
INVx1_ASAP7_75t_L g671 ( .A(n_138), .Y(n_671) );
AOI22xp33_ASAP7_75t_SL g694 ( .A1(n_138), .A2(n_142), .B1(n_513), .B2(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g1328 ( .A(n_139), .Y(n_1328) );
AOI222xp33_ASAP7_75t_L g1362 ( .A1(n_139), .A2(n_1363), .B1(n_1423), .B2(n_1427), .C1(n_1480), .C2(n_1482), .Y(n_1362) );
INVx1_ASAP7_75t_L g647 ( .A(n_140), .Y(n_647) );
INVx1_ASAP7_75t_L g778 ( .A(n_141), .Y(n_778) );
INVx1_ASAP7_75t_L g666 ( .A(n_142), .Y(n_666) );
INVx1_ASAP7_75t_L g968 ( .A(n_143), .Y(n_968) );
INVx1_ASAP7_75t_L g1383 ( .A(n_144), .Y(n_1383) );
AOI22xp33_ASAP7_75t_L g1405 ( .A1(n_144), .A2(n_208), .B1(n_331), .B2(n_360), .Y(n_1405) );
CKINVDCx5p33_ASAP7_75t_R g967 ( .A(n_145), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_146), .A2(n_167), .B1(n_677), .B2(n_678), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_146), .A2(n_167), .B1(n_513), .B2(n_615), .Y(n_689) );
CKINVDCx5p33_ASAP7_75t_R g472 ( .A(n_147), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_148), .A2(n_164), .B1(n_993), .B2(n_994), .Y(n_992) );
AOI22xp33_ASAP7_75t_SL g1008 ( .A1(n_148), .A2(n_164), .B1(n_807), .B2(n_1009), .Y(n_1008) );
INVxp33_ASAP7_75t_SL g1434 ( .A(n_150), .Y(n_1434) );
AOI22xp33_ASAP7_75t_SL g1454 ( .A1(n_150), .A2(n_177), .B1(n_1449), .B2(n_1455), .Y(n_1454) );
INVx1_ASAP7_75t_L g528 ( .A(n_151), .Y(n_528) );
INVx1_ASAP7_75t_L g821 ( .A(n_152), .Y(n_821) );
CKINVDCx5p33_ASAP7_75t_R g1066 ( .A(n_153), .Y(n_1066) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_155), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g1156 ( .A(n_155), .B(n_253), .Y(n_1156) );
AND3x2_ASAP7_75t_L g1179 ( .A(n_155), .B(n_253), .C(n_1159), .Y(n_1179) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_156), .Y(n_316) );
INVx2_ASAP7_75t_L g266 ( .A(n_157), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g650 ( .A(n_159), .Y(n_650) );
INVx1_ASAP7_75t_L g845 ( .A(n_160), .Y(n_845) );
INVx1_ASAP7_75t_L g818 ( .A(n_161), .Y(n_818) );
INVx1_ASAP7_75t_L g879 ( .A(n_162), .Y(n_879) );
INVx1_ASAP7_75t_L g938 ( .A(n_163), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g1448 ( .A1(n_166), .A2(n_184), .B1(n_1449), .B2(n_1450), .Y(n_1448) );
AOI22xp33_ASAP7_75t_L g1458 ( .A1(n_166), .A2(n_184), .B1(n_1459), .B2(n_1461), .Y(n_1458) );
INVx1_ASAP7_75t_L g1159 ( .A(n_168), .Y(n_1159) );
INVx1_ASAP7_75t_L g971 ( .A(n_169), .Y(n_971) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_169), .A2(n_193), .B1(n_981), .B2(n_982), .Y(n_980) );
CKINVDCx16_ASAP7_75t_R g569 ( .A(n_170), .Y(n_569) );
INVx1_ASAP7_75t_L g1397 ( .A(n_171), .Y(n_1397) );
CKINVDCx5p33_ASAP7_75t_R g1421 ( .A(n_172), .Y(n_1421) );
INVx1_ASAP7_75t_L g741 ( .A(n_173), .Y(n_741) );
INVx1_ASAP7_75t_L g1091 ( .A(n_174), .Y(n_1091) );
AOI221xp5_ASAP7_75t_L g1133 ( .A1(n_174), .A2(n_238), .B1(n_1039), .B2(n_1134), .C(n_1136), .Y(n_1133) );
INVx1_ASAP7_75t_L g755 ( .A(n_175), .Y(n_755) );
INVx1_ASAP7_75t_L g985 ( .A(n_176), .Y(n_985) );
INVxp33_ASAP7_75t_L g1437 ( .A(n_177), .Y(n_1437) );
INVx1_ASAP7_75t_L g268 ( .A(n_178), .Y(n_268) );
INVx2_ASAP7_75t_L g287 ( .A(n_178), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_180), .A2(n_207), .B1(n_736), .B2(n_738), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_180), .A2(n_207), .B1(n_781), .B2(n_782), .Y(n_780) );
INVx1_ASAP7_75t_L g987 ( .A(n_181), .Y(n_987) );
INVx1_ASAP7_75t_L g881 ( .A(n_182), .Y(n_881) );
AOI22xp5_ASAP7_75t_L g1184 ( .A1(n_183), .A2(n_199), .B1(n_1169), .B2(n_1172), .Y(n_1184) );
CKINVDCx5p33_ASAP7_75t_R g720 ( .A(n_185), .Y(n_720) );
INVx1_ASAP7_75t_L g464 ( .A(n_186), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g512 ( .A1(n_186), .A2(n_210), .B1(n_513), .B2(n_515), .C(n_518), .Y(n_512) );
INVx1_ASAP7_75t_L g1194 ( .A(n_187), .Y(n_1194) );
INVx1_ASAP7_75t_L g661 ( .A(n_188), .Y(n_661) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_189), .Y(n_281) );
INVx1_ASAP7_75t_L g1387 ( .A(n_190), .Y(n_1387) );
AOI21xp33_ASAP7_75t_L g1406 ( .A1(n_190), .A2(n_922), .B(n_1407), .Y(n_1406) );
XNOR2x1_ASAP7_75t_L g1057 ( .A(n_191), .B(n_1058), .Y(n_1057) );
INVx1_ASAP7_75t_L g975 ( .A(n_193), .Y(n_975) );
INVx1_ASAP7_75t_L g1026 ( .A(n_194), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_194), .A2(n_203), .B1(n_993), .B2(n_994), .Y(n_1033) );
INVx1_ASAP7_75t_L g734 ( .A(n_197), .Y(n_734) );
OAI211xp5_ASAP7_75t_SL g747 ( .A1(n_197), .A2(n_506), .B(n_748), .C(n_759), .Y(n_747) );
CKINVDCx5p33_ASAP7_75t_R g474 ( .A(n_201), .Y(n_474) );
INVx1_ASAP7_75t_L g407 ( .A(n_202), .Y(n_407) );
INVx1_ASAP7_75t_L g1020 ( .A(n_203), .Y(n_1020) );
INVx1_ASAP7_75t_L g484 ( .A(n_204), .Y(n_484) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_204), .Y(n_541) );
OAI211xp5_ASAP7_75t_L g352 ( .A1(n_205), .A2(n_353), .B(n_358), .C(n_369), .Y(n_352) );
INVx1_ASAP7_75t_L g442 ( .A(n_205), .Y(n_442) );
INVx1_ASAP7_75t_L g581 ( .A(n_206), .Y(n_581) );
INVx1_ASAP7_75t_L g1388 ( .A(n_208), .Y(n_1388) );
INVx1_ASAP7_75t_L g665 ( .A(n_209), .Y(n_665) );
AOI21xp33_ASAP7_75t_L g466 ( .A1(n_210), .A2(n_415), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g1160 ( .A(n_212), .Y(n_1160) );
NAND2xp5_ASAP7_75t_L g1174 ( .A(n_212), .B(n_1158), .Y(n_1174) );
INVx1_ASAP7_75t_L g1050 ( .A(n_213), .Y(n_1050) );
INVx1_ASAP7_75t_L g1440 ( .A(n_214), .Y(n_1440) );
OAI22xp5_ASAP7_75t_L g1473 ( .A1(n_214), .A2(n_230), .B1(n_591), .B2(n_1047), .Y(n_1473) );
OAI221xp5_ASAP7_75t_L g835 ( .A1(n_215), .A2(n_504), .B1(n_779), .B2(n_836), .C(n_842), .Y(n_835) );
INVx1_ASAP7_75t_L g1436 ( .A(n_216), .Y(n_1436) );
OAI211xp5_ASAP7_75t_L g297 ( .A1(n_217), .A2(n_298), .B(n_303), .C(n_310), .Y(n_297) );
INVx1_ASAP7_75t_L g403 ( .A(n_217), .Y(n_403) );
INVx1_ASAP7_75t_L g575 ( .A(n_219), .Y(n_575) );
INVx1_ASAP7_75t_L g1018 ( .A(n_220), .Y(n_1018) );
AO22x1_ASAP7_75t_L g1212 ( .A1(n_221), .A2(n_228), .B1(n_1180), .B2(n_1213), .Y(n_1212) );
CKINVDCx5p33_ASAP7_75t_R g721 ( .A(n_222), .Y(n_721) );
INVx1_ASAP7_75t_L g1044 ( .A(n_223), .Y(n_1044) );
INVx2_ASAP7_75t_L g265 ( .A(n_224), .Y(n_265) );
AO22x1_ASAP7_75t_L g1214 ( .A1(n_225), .A2(n_236), .B1(n_1169), .B2(n_1172), .Y(n_1214) );
CKINVDCx5p33_ASAP7_75t_R g1100 ( .A(n_226), .Y(n_1100) );
OAI221xp5_ASAP7_75t_L g1073 ( .A1(n_227), .A2(n_229), .B1(n_1074), .B2(n_1079), .C(n_1081), .Y(n_1073) );
OAI22xp5_ASAP7_75t_L g1115 ( .A1(n_227), .A2(n_229), .B1(n_1116), .B2(n_1119), .Y(n_1115) );
INVx1_ASAP7_75t_L g1441 ( .A(n_230), .Y(n_1441) );
INVxp33_ASAP7_75t_L g1478 ( .A(n_231), .Y(n_1478) );
INVx1_ASAP7_75t_L g651 ( .A(n_232), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_232), .A2(n_233), .B1(n_601), .B2(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g648 ( .A(n_233), .Y(n_648) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_235), .Y(n_388) );
INVx1_ASAP7_75t_L g1093 ( .A(n_238), .Y(n_1093) );
INVx1_ASAP7_75t_L g334 ( .A(n_239), .Y(n_334) );
BUFx3_ASAP7_75t_L g350 ( .A(n_239), .Y(n_350) );
BUFx3_ASAP7_75t_L g333 ( .A(n_240), .Y(n_333) );
INVx1_ASAP7_75t_L g343 ( .A(n_240), .Y(n_343) );
INVx1_ASAP7_75t_L g1095 ( .A(n_242), .Y(n_1095) );
OAI22xp5_ASAP7_75t_L g1427 ( .A1(n_243), .A2(n_1428), .B1(n_1429), .B2(n_1479), .Y(n_1427) );
INVx1_ASAP7_75t_L g1428 ( .A(n_243), .Y(n_1428) );
INVx1_ASAP7_75t_L g932 ( .A(n_244), .Y(n_932) );
CKINVDCx5p33_ASAP7_75t_R g815 ( .A(n_245), .Y(n_815) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_247), .Y(n_362) );
XNOR2xp5_ASAP7_75t_L g705 ( .A(n_248), .B(n_706), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_269), .B(n_1150), .Y(n_249) );
AND2x4_ASAP7_75t_L g250 ( .A(n_251), .B(n_256), .Y(n_250) );
AND2x4_ASAP7_75t_L g1426 ( .A(n_251), .B(n_257), .Y(n_1426) );
NOR2xp33_ASAP7_75t_SL g251 ( .A(n_252), .B(n_254), .Y(n_251) );
INVx1_ASAP7_75t_SL g1481 ( .A(n_252), .Y(n_1481) );
NAND2xp5_ASAP7_75t_L g1483 ( .A(n_252), .B(n_254), .Y(n_1483) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g1480 ( .A(n_254), .B(n_1481), .Y(n_1480) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_258), .B(n_262), .Y(n_257) );
INVxp67_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g277 ( .A(n_259), .B(n_278), .Y(n_277) );
OR2x6_ASAP7_75t_L g572 ( .A(n_259), .B(n_278), .Y(n_572) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g596 ( .A(n_260), .B(n_268), .Y(n_596) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g415 ( .A(n_261), .B(n_286), .Y(n_415) );
INVx8_ASAP7_75t_L g280 ( .A(n_262), .Y(n_280) );
OR2x6_ASAP7_75t_L g262 ( .A(n_263), .B(n_267), .Y(n_262) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_263), .Y(n_417) );
OR2x6_ASAP7_75t_L g583 ( .A(n_263), .B(n_285), .Y(n_583) );
INVx1_ASAP7_75t_L g840 ( .A(n_263), .Y(n_840) );
INVx2_ASAP7_75t_SL g1087 ( .A(n_263), .Y(n_1087) );
OR2x2_ASAP7_75t_L g1108 ( .A(n_263), .B(n_1078), .Y(n_1108) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g290 ( .A(n_265), .Y(n_290) );
AND2x4_ASAP7_75t_L g295 ( .A(n_265), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g302 ( .A(n_265), .Y(n_302) );
INVx1_ASAP7_75t_L g309 ( .A(n_265), .Y(n_309) );
AND2x2_ASAP7_75t_L g314 ( .A(n_265), .B(n_266), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_266), .B(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g296 ( .A(n_266), .Y(n_296) );
INVx1_ASAP7_75t_L g301 ( .A(n_266), .Y(n_301) );
INVx1_ASAP7_75t_L g318 ( .A(n_266), .Y(n_318) );
INVx1_ASAP7_75t_L g498 ( .A(n_266), .Y(n_498) );
AND2x4_ASAP7_75t_L g317 ( .A(n_267), .B(n_318), .Y(n_317) );
INVx2_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g982 ( .A(n_268), .B(n_321), .Y(n_982) );
OR2x2_ASAP7_75t_L g1047 ( .A(n_268), .B(n_321), .Y(n_1047) );
XNOR2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_700), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
XNOR2x1_ASAP7_75t_L g273 ( .A(n_274), .B(n_567), .Y(n_273) );
XNOR2x1_ASAP7_75t_L g274 ( .A(n_275), .B(n_452), .Y(n_274) );
INVx1_ASAP7_75t_L g450 ( .A(n_276), .Y(n_450) );
OAI211xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_279), .B(n_324), .C(n_377), .Y(n_276) );
AOI31xp33_ASAP7_75t_L g1042 ( .A1(n_277), .A2(n_1043), .A3(n_1048), .B(n_1051), .Y(n_1042) );
AOI31xp33_ASAP7_75t_L g1470 ( .A1(n_277), .A2(n_1471), .A3(n_1474), .B(n_1477), .Y(n_1470) );
AND2x4_ASAP7_75t_L g410 ( .A(n_278), .B(n_411), .Y(n_410) );
AND2x4_ASAP7_75t_L g559 ( .A(n_278), .B(n_560), .Y(n_559) );
AND2x4_ASAP7_75t_L g623 ( .A(n_278), .B(n_411), .Y(n_623) );
AOI211xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_281), .B(n_282), .C(n_297), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_280), .A2(n_580), .B1(n_581), .B2(n_582), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_280), .A2(n_582), .B1(n_650), .B2(n_671), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_280), .A2(n_868), .B1(n_881), .B2(n_882), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g986 ( .A1(n_280), .A2(n_582), .B1(n_967), .B2(n_987), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_280), .A2(n_882), .B1(n_1017), .B2(n_1052), .Y(n_1051) );
AOI22xp33_ASAP7_75t_SL g1477 ( .A1(n_280), .A2(n_882), .B1(n_1436), .B2(n_1478), .Y(n_1477) );
OAI22xp33_ASAP7_75t_L g400 ( .A1(n_281), .A2(n_394), .B1(n_401), .B2(n_403), .Y(n_400) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_288), .Y(n_283) );
AOI322xp5_ASAP7_75t_L g310 ( .A1(n_284), .A2(n_311), .A3(n_315), .B1(n_316), .B2(n_317), .C1(n_319), .C2(n_323), .Y(n_310) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x4_ASAP7_75t_L g292 ( .A(n_285), .B(n_293), .Y(n_292) );
AND2x4_ASAP7_75t_L g576 ( .A(n_285), .B(n_496), .Y(n_576) );
AND2x4_ASAP7_75t_L g578 ( .A(n_285), .B(n_293), .Y(n_578) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g307 ( .A(n_287), .Y(n_307) );
INVx2_ASAP7_75t_L g423 ( .A(n_288), .Y(n_423) );
BUFx2_ASAP7_75t_L g1094 ( .A(n_288), .Y(n_1094) );
BUFx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g430 ( .A(n_289), .Y(n_430) );
INVx1_ASAP7_75t_L g458 ( .A(n_289), .Y(n_458) );
INVx1_ASAP7_75t_L g487 ( .A(n_290), .Y(n_487) );
AND2x4_ASAP7_75t_L g496 ( .A(n_290), .B(n_497), .Y(n_496) );
INVx5_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g1048 ( .A1(n_292), .A2(n_576), .B1(n_1049), .B2(n_1050), .Y(n_1048) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g426 ( .A(n_295), .Y(n_426) );
INVx3_ASAP7_75t_L g434 ( .A(n_295), .Y(n_434) );
BUFx6f_ASAP7_75t_L g848 ( .A(n_295), .Y(n_848) );
AND2x4_ASAP7_75t_L g308 ( .A(n_296), .B(n_309), .Y(n_308) );
OAI221xp5_ASAP7_75t_L g767 ( .A1(n_298), .A2(n_720), .B1(n_721), .B2(n_768), .C(n_769), .Y(n_767) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g420 ( .A(n_300), .Y(n_420) );
INVx3_ASAP7_75t_L g465 ( .A(n_300), .Y(n_465) );
INVx2_ASAP7_75t_L g475 ( .A(n_300), .Y(n_475) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_301), .B(n_302), .Y(n_441) );
INVx1_ASAP7_75t_L g321 ( .A(n_302), .Y(n_321) );
NAND4xp25_ASAP7_75t_SL g573 ( .A(n_303), .B(n_574), .C(n_579), .D(n_584), .Y(n_573) );
NAND4xp25_ASAP7_75t_SL g659 ( .A(n_303), .B(n_660), .C(n_663), .D(n_670), .Y(n_659) );
NAND4xp25_ASAP7_75t_SL g872 ( .A(n_303), .B(n_873), .C(n_876), .D(n_880), .Y(n_872) );
CKINVDCx11_ASAP7_75t_R g303 ( .A(n_304), .Y(n_303) );
AOI211xp5_ASAP7_75t_L g978 ( .A1(n_304), .A2(n_678), .B(n_979), .C(n_980), .Y(n_978) );
AOI211xp5_ASAP7_75t_L g1043 ( .A1(n_304), .A2(n_1044), .B(n_1045), .C(n_1046), .Y(n_1043) );
AOI211xp5_ASAP7_75t_L g1471 ( .A1(n_304), .A2(n_1045), .B(n_1472), .C(n_1473), .Y(n_1471) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_308), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVxp67_ASAP7_75t_L g322 ( .A(n_306), .Y(n_322) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2x1p5_ASAP7_75t_L g448 ( .A(n_307), .B(n_449), .Y(n_448) );
BUFx3_ASAP7_75t_L g508 ( .A(n_308), .Y(n_508) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_308), .Y(n_588) );
BUFx6f_ASAP7_75t_L g608 ( .A(n_308), .Y(n_608) );
BUFx2_ASAP7_75t_L g669 ( .A(n_308), .Y(n_669) );
BUFx3_ASAP7_75t_L g937 ( .A(n_308), .Y(n_937) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g677 ( .A(n_312), .Y(n_677) );
INVx3_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
BUFx6f_ASAP7_75t_L g481 ( .A(n_313), .Y(n_481) );
AND2x4_ASAP7_75t_L g505 ( .A(n_313), .B(n_495), .Y(n_505) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx3_ASAP7_75t_L g468 ( .A(n_314), .Y(n_468) );
AOI322xp5_ASAP7_75t_L g358 ( .A1(n_316), .A2(n_323), .A3(n_359), .B1(n_361), .B2(n_362), .C1(n_363), .C2(n_367), .Y(n_358) );
INVx2_ASAP7_75t_L g591 ( .A(n_317), .Y(n_591) );
AOI222xp33_ASAP7_75t_L g663 ( .A1(n_317), .A2(n_319), .B1(n_664), .B2(n_665), .C1(n_666), .C2(n_667), .Y(n_663) );
INVx2_ASAP7_75t_L g981 ( .A(n_317), .Y(n_981) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_318), .A2(n_484), .B1(n_485), .B2(n_486), .Y(n_483) );
HB1xp67_ASAP7_75t_L g762 ( .A(n_318), .Y(n_762) );
INVx1_ASAP7_75t_L g949 ( .A(n_318), .Y(n_949) );
AOI222xp33_ASAP7_75t_L g584 ( .A1(n_319), .A2(n_585), .B1(n_586), .B2(n_589), .C1(n_590), .C2(n_592), .Y(n_584) );
AOI222xp33_ASAP7_75t_L g876 ( .A1(n_319), .A2(n_586), .B1(n_590), .B2(n_877), .C1(n_878), .C2(n_879), .Y(n_876) );
AND2x4_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g947 ( .A1(n_320), .A2(n_926), .B1(n_927), .B2(n_948), .Y(n_947) );
AND2x4_ASAP7_75t_L g1370 ( .A(n_320), .B(n_1077), .Y(n_1370) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OAI31xp33_ASAP7_75t_SL g324 ( .A1(n_325), .A2(n_335), .A3(n_352), .B(n_372), .Y(n_324) );
INVx4_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_327), .A2(n_637), .B1(n_638), .B2(n_639), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_327), .A2(n_646), .B1(n_647), .B2(n_648), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_327), .A2(n_637), .B1(n_870), .B2(n_871), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_327), .A2(n_345), .B1(n_967), .B2(n_968), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_327), .A2(n_345), .B1(n_1017), .B2(n_1018), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1435 ( .A1(n_327), .A2(n_345), .B1(n_1436), .B2(n_1437), .Y(n_1435) );
AND2x6_ASAP7_75t_L g327 ( .A(n_328), .B(n_331), .Y(n_327) );
AND2x4_ASAP7_75t_L g634 ( .A(n_328), .B(n_635), .Y(n_634) );
AND2x4_ASAP7_75t_L g646 ( .A(n_328), .B(n_635), .Y(n_646) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g629 ( .A(n_329), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g339 ( .A(n_330), .Y(n_339) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_330), .Y(n_347) );
AND2x2_ASAP7_75t_L g381 ( .A(n_330), .B(n_374), .Y(n_381) );
INVx2_ASAP7_75t_L g412 ( .A(n_330), .Y(n_412) );
INVx1_ASAP7_75t_L g408 ( .A(n_331), .Y(n_408) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_331), .Y(n_613) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_331), .Y(n_622) );
INVx2_ASAP7_75t_L g739 ( .A(n_331), .Y(n_739) );
INVx1_ASAP7_75t_L g1462 ( .A(n_331), .Y(n_1462) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g391 ( .A(n_332), .Y(n_391) );
INVx1_ASAP7_75t_L g521 ( .A(n_332), .Y(n_521) );
INVx1_ASAP7_75t_L g564 ( .A(n_332), .Y(n_564) );
BUFx6f_ASAP7_75t_L g688 ( .A(n_332), .Y(n_688) );
AND2x4_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx2_ASAP7_75t_L g351 ( .A(n_333), .Y(n_351) );
AND2x2_ASAP7_75t_L g357 ( .A(n_333), .B(n_350), .Y(n_357) );
INVx1_ASAP7_75t_L g341 ( .A(n_334), .Y(n_341) );
OR2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_340), .Y(n_336) );
INVx1_ASAP7_75t_L g361 ( .A(n_337), .Y(n_361) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g354 ( .A(n_338), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g371 ( .A(n_338), .Y(n_371) );
AND2x6_ASAP7_75t_L g637 ( .A(n_338), .B(n_360), .Y(n_637) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x6_ASAP7_75t_L g367 ( .A(n_339), .B(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g395 ( .A(n_340), .Y(n_395) );
INVx1_ASAP7_75t_L g719 ( .A(n_340), .Y(n_719) );
BUFx2_ASAP7_75t_L g1126 ( .A(n_340), .Y(n_1126) );
OR2x2_ASAP7_75t_L g1145 ( .A(n_340), .B(n_555), .Y(n_1145) );
OR2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
AND2x2_ASAP7_75t_L g399 ( .A(n_341), .B(n_342), .Y(n_399) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g360 ( .A(n_343), .B(n_350), .Y(n_360) );
INVx4_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_345), .A2(n_581), .B1(n_633), .B2(n_634), .Y(n_632) );
AOI221xp5_ASAP7_75t_L g649 ( .A1(n_345), .A2(n_637), .B1(n_650), .B2(n_651), .C(n_652), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_345), .A2(n_646), .B1(n_867), .B2(n_868), .Y(n_866) );
AND2x4_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
AND2x2_ASAP7_75t_SL g363 ( .A(n_346), .B(n_364), .Y(n_363) );
AND2x4_ASAP7_75t_L g974 ( .A(n_346), .B(n_364), .Y(n_974) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx6_ASAP7_75t_L g517 ( .A(n_348), .Y(n_517) );
INVx2_ASAP7_75t_L g552 ( .A(n_348), .Y(n_552) );
AND2x2_ASAP7_75t_L g560 ( .A(n_348), .B(n_538), .Y(n_560) );
BUFx2_ASAP7_75t_L g618 ( .A(n_348), .Y(n_618) );
AND2x4_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
INVx1_ASAP7_75t_L g368 ( .A(n_349), .Y(n_368) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g366 ( .A(n_351), .Y(n_366) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AOI211xp5_ASAP7_75t_L g625 ( .A1(n_354), .A2(n_370), .B(n_626), .C(n_627), .Y(n_625) );
HB1xp67_ASAP7_75t_L g1021 ( .A(n_355), .Y(n_1021) );
HB1xp67_ASAP7_75t_L g1465 ( .A(n_355), .Y(n_1465) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x4_ASAP7_75t_L g370 ( .A(n_356), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g514 ( .A(n_356), .Y(n_514) );
BUFx6f_ASAP7_75t_L g656 ( .A(n_356), .Y(n_656) );
INVx1_ASAP7_75t_L g711 ( .A(n_356), .Y(n_711) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_357), .Y(n_547) );
INVx2_ASAP7_75t_L g387 ( .A(n_359), .Y(n_387) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_SL g406 ( .A(n_360), .Y(n_406) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_360), .Y(n_520) );
BUFx2_ASAP7_75t_L g612 ( .A(n_360), .Y(n_612) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_360), .Y(n_724) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_360), .Y(n_737) );
BUFx2_ASAP7_75t_L g901 ( .A(n_360), .Y(n_901) );
BUFx3_ASAP7_75t_L g1460 ( .A(n_360), .Y(n_1460) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_362), .A2(n_428), .B1(n_431), .B2(n_435), .Y(n_427) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g630 ( .A(n_365), .Y(n_630) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g535 ( .A(n_366), .Y(n_535) );
INVx3_ASAP7_75t_L g631 ( .A(n_367), .Y(n_631) );
AOI222xp33_ASAP7_75t_L g969 ( .A1(n_367), .A2(n_918), .B1(n_970), .B2(n_971), .C1(n_972), .C2(n_975), .Y(n_969) );
AOI222xp33_ASAP7_75t_L g1019 ( .A1(n_367), .A2(n_1020), .B1(n_1021), .B2(n_1022), .C1(n_1023), .C2(n_1024), .Y(n_1019) );
AOI222xp33_ASAP7_75t_L g1438 ( .A1(n_367), .A2(n_810), .B1(n_974), .B2(n_1439), .C1(n_1440), .C2(n_1441), .Y(n_1438) );
BUFx3_ASAP7_75t_L g544 ( .A(n_368), .Y(n_544) );
CKINVDCx8_ASAP7_75t_R g369 ( .A(n_370), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g861 ( .A(n_370), .B(n_862), .Y(n_861) );
INVx5_ASAP7_75t_L g976 ( .A(n_370), .Y(n_976) );
OAI21xp33_ASAP7_75t_L g654 ( .A1(n_371), .A2(n_655), .B(n_656), .Y(n_654) );
INVx1_ASAP7_75t_SL g640 ( .A(n_372), .Y(n_640) );
AND2x4_ASAP7_75t_L g372 ( .A(n_373), .B(n_375), .Y(n_372) );
AND2x4_ASAP7_75t_L g658 ( .A(n_373), .B(n_375), .Y(n_658) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x4_ASAP7_75t_L g411 ( .A(n_374), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g851 ( .A(n_375), .Y(n_851) );
BUFx2_ASAP7_75t_L g1149 ( .A(n_375), .Y(n_1149) );
BUFx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g382 ( .A(n_376), .Y(n_382) );
OR2x6_ASAP7_75t_L g414 ( .A(n_376), .B(n_415), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_378), .B(n_413), .Y(n_377) );
OAI33xp33_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_383), .A3(n_392), .B1(n_400), .B2(n_404), .B3(n_409), .Y(n_378) );
INVx1_ASAP7_75t_SL g610 ( .A(n_379), .Y(n_610) );
OR2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
OR2x6_ASAP7_75t_L g523 ( .A(n_380), .B(n_382), .Y(n_523) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g692 ( .A(n_381), .Y(n_692) );
INVx2_ASAP7_75t_SL g1136 ( .A(n_381), .Y(n_1136) );
BUFx3_ASAP7_75t_L g1413 ( .A(n_381), .Y(n_1413) );
INVx2_ASAP7_75t_L g510 ( .A(n_382), .Y(n_510) );
AND2x4_ASAP7_75t_L g595 ( .A(n_382), .B(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g691 ( .A(n_382), .B(n_692), .Y(n_691) );
BUFx2_ASAP7_75t_L g783 ( .A(n_382), .Y(n_783) );
AND2x4_ASAP7_75t_L g991 ( .A(n_382), .B(n_596), .Y(n_991) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B1(n_388), .B2(n_389), .Y(n_383) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_384), .A2(n_388), .B1(n_422), .B2(n_424), .Y(n_421) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_387), .A2(n_528), .B1(n_529), .B2(n_531), .Y(n_527) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g530 ( .A(n_391), .Y(n_530) );
OR2x2_ASAP7_75t_L g1147 ( .A(n_391), .B(n_555), .Y(n_1147) );
OAI22xp33_ASAP7_75t_SL g392 ( .A1(n_393), .A2(n_394), .B1(n_396), .B2(n_397), .Y(n_392) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_393), .A2(n_396), .B1(n_417), .B2(n_418), .Y(n_416) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g729 ( .A(n_395), .Y(n_729) );
INVx1_ASAP7_75t_L g789 ( .A(n_395), .Y(n_789) );
BUFx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g402 ( .A(n_399), .Y(n_402) );
BUFx4f_ASAP7_75t_L g733 ( .A(n_399), .Y(n_733) );
INVx1_ASAP7_75t_L g865 ( .A(n_399), .Y(n_865) );
INVx1_ASAP7_75t_L g1404 ( .A(n_399), .Y(n_1404) );
BUFx3_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OR2x6_ASAP7_75t_L g566 ( .A(n_402), .B(n_554), .Y(n_566) );
OAI221xp5_ASAP7_75t_L g716 ( .A1(n_402), .A2(n_717), .B1(n_720), .B2(n_721), .C(n_722), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_406), .B1(n_407), .B2(n_408), .Y(n_404) );
INVx2_ASAP7_75t_L g558 ( .A(n_406), .Y(n_558) );
INVx1_ASAP7_75t_L g916 ( .A(n_406), .Y(n_916) );
INVx4_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AOI221xp5_ASAP7_75t_L g511 ( .A1(n_410), .A2(n_512), .B1(n_522), .B2(n_524), .C(n_532), .Y(n_511) );
BUFx4f_ASAP7_75t_L g727 ( .A(n_410), .Y(n_727) );
BUFx4f_ASAP7_75t_L g812 ( .A(n_410), .Y(n_812) );
AOI33xp33_ASAP7_75t_L g1034 ( .A1(n_410), .A2(n_801), .A3(n_1035), .B1(n_1038), .B2(n_1040), .B3(n_1041), .Y(n_1034) );
AOI33xp33_ASAP7_75t_L g1457 ( .A1(n_410), .A2(n_801), .A3(n_1458), .B1(n_1463), .B2(n_1466), .B3(n_1469), .Y(n_1457) );
INVx2_ASAP7_75t_L g1128 ( .A(n_411), .Y(n_1128) );
CKINVDCx5p33_ASAP7_75t_R g1407 ( .A(n_411), .Y(n_1407) );
AND2x4_ASAP7_75t_L g538 ( .A(n_412), .B(n_539), .Y(n_538) );
OAI33xp33_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_416), .A3(n_421), .B1(n_427), .B2(n_436), .B3(n_443), .Y(n_413) );
OAI33xp33_ASAP7_75t_L g1083 ( .A1(n_414), .A2(n_443), .A3(n_1084), .B1(n_1092), .B2(n_1097), .B3(n_1101), .Y(n_1083) );
OAI22xp33_ASAP7_75t_L g436 ( .A1(n_417), .A2(n_437), .B1(n_438), .B2(n_442), .Y(n_436) );
BUFx2_ASAP7_75t_L g768 ( .A(n_417), .Y(n_768) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_420), .B(n_483), .Y(n_482) );
OR2x2_ASAP7_75t_L g779 ( .A(n_420), .B(n_489), .Y(n_779) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g754 ( .A(n_424), .Y(n_754) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AND2x4_ASAP7_75t_L g500 ( .A(n_425), .B(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g829 ( .A(n_426), .Y(n_829) );
INVx2_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g844 ( .A(n_429), .Y(n_844) );
BUFx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g751 ( .A(n_430), .Y(n_751) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g682 ( .A(n_433), .Y(n_682) );
INVx2_ASAP7_75t_L g1451 ( .A(n_433), .Y(n_1451) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx3_ASAP7_75t_L g461 ( .A(n_434), .Y(n_461) );
INVx3_ASAP7_75t_L g777 ( .A(n_434), .Y(n_777) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_440), .B(n_947), .Y(n_946) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AOI33xp33_ASAP7_75t_L g594 ( .A1(n_444), .A2(n_595), .A3(n_597), .B1(n_600), .B2(n_604), .B3(n_606), .Y(n_594) );
AOI33xp33_ASAP7_75t_L g989 ( .A1(n_444), .A2(n_990), .A3(n_992), .B1(n_995), .B2(n_999), .B3(n_1003), .Y(n_989) );
AOI33xp33_ASAP7_75t_L g1029 ( .A1(n_444), .A2(n_990), .A3(n_1030), .B1(n_1031), .B2(n_1032), .B3(n_1033), .Y(n_1029) );
AOI33xp33_ASAP7_75t_L g1373 ( .A1(n_444), .A2(n_1374), .A3(n_1375), .B1(n_1376), .B2(n_1380), .B3(n_1381), .Y(n_1373) );
INVx6_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx5_ASAP7_75t_L g684 ( .A(n_445), .Y(n_684) );
OR2x6_ASAP7_75t_L g445 ( .A(n_446), .B(n_448), .Y(n_445) );
NAND2x1p5_ASAP7_75t_L g537 ( .A(n_446), .B(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g554 ( .A(n_447), .B(n_555), .Y(n_554) );
AND2x4_ASAP7_75t_L g1065 ( .A(n_447), .B(n_495), .Y(n_1065) );
BUFx2_ASAP7_75t_L g478 ( .A(n_448), .Y(n_478) );
INVx2_ASAP7_75t_L g758 ( .A(n_448), .Y(n_758) );
NAND4xp25_ASAP7_75t_L g453 ( .A(n_454), .B(n_511), .C(n_549), .D(n_561), .Y(n_453) );
OAI31xp33_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_492), .A3(n_503), .B(n_509), .Y(n_454) );
OAI221xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_463), .B1(n_469), .B2(n_473), .C(n_479), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_459), .B1(n_460), .B2(n_462), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_457), .A2(n_470), .B1(n_471), .B2(n_472), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g941 ( .A1(n_457), .A2(n_471), .B1(n_942), .B2(n_943), .Y(n_941) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g773 ( .A(n_458), .Y(n_773) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_459), .A2(n_462), .B1(n_519), .B2(n_521), .Y(n_518) );
INVx2_ASAP7_75t_L g605 ( .A(n_460), .Y(n_605) );
INVx2_ASAP7_75t_SL g675 ( .A(n_460), .Y(n_675) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g471 ( .A(n_461), .Y(n_471) );
INVx2_ASAP7_75t_L g889 ( .A(n_461), .Y(n_889) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B(n_466), .Y(n_463) );
BUFx2_ASAP7_75t_L g837 ( .A(n_465), .Y(n_837) );
INVx1_ASAP7_75t_L g1090 ( .A(n_465), .Y(n_1090) );
BUFx2_ASAP7_75t_L g598 ( .A(n_467), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_467), .B(n_745), .Y(n_744) );
INVx2_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g477 ( .A(n_468), .Y(n_477) );
INVx2_ASAP7_75t_SL g833 ( .A(n_468), .Y(n_833) );
AOI222xp33_ASAP7_75t_L g549 ( .A1(n_470), .A2(n_480), .B1(n_550), .B2(n_556), .C1(n_557), .C2(n_559), .Y(n_549) );
INVx1_ASAP7_75t_L g603 ( .A(n_471), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_472), .A2(n_474), .B1(n_562), .B2(n_565), .Y(n_561) );
OAI21xp33_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B(n_476), .Y(n_473) );
BUFx3_ASAP7_75t_L g993 ( .A(n_477), .Y(n_993) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B(n_482), .C(n_488), .Y(n_479) );
INVx1_ASAP7_75t_L g1005 ( .A(n_481), .Y(n_1005) );
NAND2x1p5_ASAP7_75t_L g1080 ( .A(n_486), .B(n_1077), .Y(n_1080) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OR2x6_ASAP7_75t_L g765 ( .A(n_487), .B(n_489), .Y(n_765) );
A2O1A1Ixp33_ASAP7_75t_L g944 ( .A1(n_488), .A2(n_677), .B(n_945), .C(n_946), .Y(n_944) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g745 ( .A(n_489), .Y(n_745) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx3_ASAP7_75t_L g781 ( .A(n_494), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_494), .A2(n_500), .B1(n_931), .B2(n_932), .Y(n_930) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
INVx2_ASAP7_75t_L g502 ( .A(n_495), .Y(n_502) );
INVx1_ASAP7_75t_L g602 ( .A(n_496), .Y(n_602) );
BUFx2_ASAP7_75t_L g892 ( .A(n_496), .Y(n_892) );
BUFx6f_ASAP7_75t_L g935 ( .A(n_496), .Y(n_935) );
BUFx2_ASAP7_75t_L g996 ( .A(n_496), .Y(n_996) );
BUFx6f_ASAP7_75t_L g1002 ( .A(n_496), .Y(n_1002) );
INVx1_ASAP7_75t_L g1378 ( .A(n_496), .Y(n_1378) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx3_ASAP7_75t_L g782 ( .A(n_500), .Y(n_782) );
AND2x4_ASAP7_75t_L g507 ( .A(n_501), .B(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
CKINVDCx6p67_ASAP7_75t_R g504 ( .A(n_505), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g933 ( .A1(n_505), .A2(n_934), .B1(n_936), .B2(n_938), .Y(n_933) );
INVx8_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g897 ( .A(n_508), .Y(n_897) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NOR2xp67_ASAP7_75t_L g743 ( .A(n_510), .B(n_744), .Y(n_743) );
INVx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_517), .Y(n_526) );
INVx2_ASAP7_75t_L g616 ( .A(n_517), .Y(n_616) );
INVx2_ASAP7_75t_L g635 ( .A(n_517), .Y(n_635) );
INVx1_ASAP7_75t_L g695 ( .A(n_517), .Y(n_695) );
INVx2_ASAP7_75t_SL g922 ( .A(n_517), .Y(n_922) );
INVx2_ASAP7_75t_L g1010 ( .A(n_517), .Y(n_1010) );
INVx1_ASAP7_75t_L g803 ( .A(n_519), .Y(n_803) );
INVx2_ASAP7_75t_SL g519 ( .A(n_520), .Y(n_519) );
BUFx3_ASAP7_75t_L g1039 ( .A(n_520), .Y(n_1039) );
AND2x4_ASAP7_75t_L g1113 ( .A(n_520), .B(n_1114), .Y(n_1113) );
INVx1_ASAP7_75t_L g725 ( .A(n_521), .Y(n_725) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
OAI22xp5_ASAP7_75t_SL g715 ( .A1(n_523), .A2(n_716), .B1(n_726), .B2(n_728), .Y(n_715) );
CKINVDCx5p33_ASAP7_75t_R g801 ( .A(n_523), .Y(n_801) );
INVx4_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g902 ( .A(n_529), .Y(n_902) );
INVx1_ASAP7_75t_L g1415 ( .A(n_529), .Y(n_1415) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g714 ( .A(n_533), .Y(n_714) );
INVx2_ASAP7_75t_L g925 ( .A(n_533), .Y(n_925) );
NAND2x1p5_ASAP7_75t_L g533 ( .A(n_534), .B(n_536), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g1118 ( .A(n_535), .Y(n_1118) );
INVx2_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
OR2x6_ASAP7_75t_L g542 ( .A(n_537), .B(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g548 ( .A(n_537), .Y(n_548) );
AND2x4_ASAP7_75t_L g1117 ( .A(n_538), .B(n_1118), .Y(n_1117) );
INVx1_ASAP7_75t_L g1120 ( .A(n_538), .Y(n_1120) );
AND2x4_ASAP7_75t_L g1400 ( .A(n_538), .B(n_1118), .Y(n_1400) );
AND2x4_ASAP7_75t_L g1402 ( .A(n_538), .B(n_544), .Y(n_1402) );
BUFx2_ASAP7_75t_L g1417 ( .A(n_538), .Y(n_1417) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g799 ( .A(n_542), .Y(n_799) );
OR2x2_ASAP7_75t_L g1119 ( .A(n_543), .B(n_1120), .Y(n_1119) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NAND3xp33_ASAP7_75t_SL g795 ( .A(n_545), .B(n_796), .C(n_800), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_548), .Y(n_545) );
INVx1_ASAP7_75t_L g1468 ( .A(n_546), .Y(n_1468) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g620 ( .A(n_547), .Y(n_620) );
INVx2_ASAP7_75t_SL g808 ( .A(n_547), .Y(n_808) );
BUFx3_ASAP7_75t_L g810 ( .A(n_547), .Y(n_810) );
BUFx4f_ASAP7_75t_L g918 ( .A(n_547), .Y(n_918) );
AND2x4_ASAP7_75t_L g1132 ( .A(n_547), .B(n_1114), .Y(n_1132) );
INVx1_ASAP7_75t_L g1135 ( .A(n_547), .Y(n_1135) );
AND2x4_ASAP7_75t_L g1416 ( .A(n_547), .B(n_1417), .Y(n_1416) );
AND2x2_ASAP7_75t_L g709 ( .A(n_548), .B(n_710), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_550), .A2(n_557), .B1(n_818), .B2(n_819), .Y(n_817) );
AOI222xp33_ASAP7_75t_L g950 ( .A1(n_550), .A2(n_559), .B1(n_562), .B2(n_942), .C1(n_945), .C2(n_951), .Y(n_950) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_553), .Y(n_550) );
BUFx2_ASAP7_75t_L g1464 ( .A(n_551), .Y(n_1464) );
INVx2_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g806 ( .A(n_552), .Y(n_806) );
AND2x2_ASAP7_75t_L g557 ( .A(n_553), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
OR2x6_ASAP7_75t_L g563 ( .A(n_554), .B(n_564), .Y(n_563) );
OR2x2_ASAP7_75t_L g786 ( .A(n_554), .B(n_564), .Y(n_786) );
OR2x2_ASAP7_75t_L g788 ( .A(n_554), .B(n_789), .Y(n_788) );
OR2x2_ASAP7_75t_L g790 ( .A(n_554), .B(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g1114 ( .A(n_555), .Y(n_1114) );
AOI22xp5_ASAP7_75t_L g952 ( .A1(n_557), .A2(n_565), .B1(n_943), .B2(n_953), .Y(n_952) );
OR2x6_ASAP7_75t_L g742 ( .A(n_559), .B(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g1109 ( .A(n_559), .Y(n_1109) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_562), .A2(n_565), .B1(n_815), .B2(n_816), .Y(n_814) );
CKINVDCx6p67_ASAP7_75t_R g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g1140 ( .A(n_564), .Y(n_1140) );
CKINVDCx6p67_ASAP7_75t_R g565 ( .A(n_566), .Y(n_565) );
OA22x2_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_641), .B1(n_642), .B2(n_699), .Y(n_567) );
INVx1_ASAP7_75t_L g699 ( .A(n_568), .Y(n_699) );
XNOR2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
AOI211xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_573), .B(n_593), .C(n_624), .Y(n_570) );
AOI221x1_ASAP7_75t_L g643 ( .A1(n_571), .A2(n_644), .B1(n_657), .B2(n_659), .C(n_672), .Y(n_643) );
AOI221x1_ASAP7_75t_L g859 ( .A1(n_571), .A2(n_657), .B1(n_860), .B2(n_872), .C(n_883), .Y(n_859) );
CKINVDCx16_ASAP7_75t_R g571 ( .A(n_572), .Y(n_571) );
AOI31xp33_ASAP7_75t_L g977 ( .A1(n_572), .A2(n_978), .A3(n_983), .B(n_986), .Y(n_977) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .B1(n_577), .B2(n_578), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_576), .A2(n_578), .B1(n_661), .B2(n_662), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_576), .A2(n_578), .B1(n_874), .B2(n_875), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_576), .A2(n_578), .B1(n_984), .B2(n_985), .Y(n_983) );
AOI22xp33_ASAP7_75t_SL g1474 ( .A1(n_576), .A2(n_578), .B1(n_1475), .B2(n_1476), .Y(n_1474) );
INVx4_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx5_ASAP7_75t_L g882 ( .A(n_583), .Y(n_882) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_SL g994 ( .A(n_587), .Y(n_994) );
INVx2_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_588), .Y(n_599) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_594), .B(n_609), .Y(n_593) );
NAND3xp33_ASAP7_75t_L g673 ( .A(n_595), .B(n_674), .C(n_676), .Y(n_673) );
NAND3xp33_ASAP7_75t_L g890 ( .A(n_595), .B(n_891), .C(n_895), .Y(n_890) );
BUFx2_ASAP7_75t_L g1374 ( .A(n_595), .Y(n_1374) );
BUFx2_ASAP7_75t_SL g769 ( .A(n_596), .Y(n_769) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
BUFx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_SL g679 ( .A(n_608), .Y(n_679) );
HB1xp67_ASAP7_75t_L g886 ( .A(n_608), .Y(n_886) );
AOI33xp33_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .A3(n_614), .B1(n_617), .B2(n_621), .B3(n_623), .Y(n_609) );
AOI33xp33_ASAP7_75t_L g914 ( .A1(n_610), .A2(n_623), .A3(n_915), .B1(n_917), .B2(n_919), .B3(n_923), .Y(n_914) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g1139 ( .A(n_616), .Y(n_1139) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND3xp33_ASAP7_75t_L g693 ( .A(n_623), .B(n_694), .C(n_696), .Y(n_693) );
INVx1_ASAP7_75t_L g907 ( .A(n_623), .Y(n_907) );
AOI31xp33_ASAP7_75t_SL g624 ( .A1(n_625), .A2(n_632), .A3(n_636), .B(n_640), .Y(n_624) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g653 ( .A(n_629), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g1432 ( .A1(n_634), .A2(n_637), .B1(n_1433), .B2(n_1434), .Y(n_1432) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_637), .A2(n_646), .B1(n_964), .B2(n_965), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_637), .A2(n_646), .B1(n_1026), .B2(n_1027), .Y(n_1025) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g698 ( .A(n_643), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_649), .Y(n_644) );
INVx1_ASAP7_75t_L g1037 ( .A(n_656), .Y(n_1037) );
AND2x4_ASAP7_75t_L g1141 ( .A(n_656), .B(n_1142), .Y(n_1141) );
AOI211x1_ASAP7_75t_L g961 ( .A1(n_657), .A2(n_962), .B(n_977), .C(n_988), .Y(n_961) );
BUFx6f_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AOI211x1_ASAP7_75t_SL g1014 ( .A1(n_658), .A2(n_1015), .B(n_1028), .C(n_1042), .Y(n_1014) );
INVx1_ASAP7_75t_L g1443 ( .A(n_658), .Y(n_1443) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AND2x4_ASAP7_75t_L g1372 ( .A(n_669), .B(n_1077), .Y(n_1372) );
NAND4xp25_ASAP7_75t_L g672 ( .A(n_673), .B(n_680), .C(n_685), .D(n_693), .Y(n_672) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NAND3xp33_ASAP7_75t_L g680 ( .A(n_681), .B(n_683), .C(n_684), .Y(n_680) );
NAND3xp33_ASAP7_75t_L g884 ( .A(n_684), .B(n_885), .C(n_887), .Y(n_884) );
AOI33xp33_ASAP7_75t_L g1445 ( .A1(n_684), .A2(n_1446), .A3(n_1448), .B1(n_1452), .B2(n_1454), .B3(n_1456), .Y(n_1445) );
NAND3xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_689), .C(n_690), .Y(n_685) );
BUFx6f_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g1123 ( .A(n_688), .Y(n_1123) );
NAND3xp33_ASAP7_75t_L g898 ( .A(n_690), .B(n_899), .C(n_900), .Y(n_898) );
INVx3_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_702), .B1(n_955), .B2(n_956), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AO22x2_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_704), .B1(n_854), .B2(n_855), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AO22x1_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_792), .B1(n_852), .B2(n_853), .Y(n_704) );
INVx1_ASAP7_75t_L g853 ( .A(n_705), .Y(n_853) );
AND4x1_ASAP7_75t_L g706 ( .A(n_707), .B(n_740), .C(n_746), .D(n_784), .Y(n_706) );
NOR3xp33_ASAP7_75t_SL g707 ( .A(n_708), .B(n_712), .C(n_715), .Y(n_707) );
BUFx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AOI221xp5_ASAP7_75t_L g924 ( .A1(n_709), .A2(n_799), .B1(n_925), .B2(n_926), .C(n_927), .Y(n_924) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_714), .A2(n_797), .B1(n_798), .B2(n_799), .Y(n_796) );
BUFx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
BUFx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g791 ( .A(n_724), .Y(n_791) );
AND2x2_ASAP7_75t_L g1396 ( .A(n_724), .B(n_1114), .Y(n_1396) );
CKINVDCx5p33_ASAP7_75t_R g726 ( .A(n_727), .Y(n_726) );
OAI221xp5_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_730), .B1(n_731), .B2(n_734), .C(n_735), .Y(n_728) );
BUFx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g1125 ( .A(n_733), .Y(n_1125) );
BUFx3_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g804 ( .A(n_739), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_742), .B(n_821), .Y(n_820) );
AND2x2_ASAP7_75t_L g761 ( .A(n_745), .B(n_762), .Y(n_761) );
OAI31xp33_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_766), .A3(n_780), .B(n_783), .Y(n_746) );
OAI221xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_752), .B1(n_753), .B2(n_755), .C(n_756), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
BUFx2_ASAP7_75t_L g825 ( .A(n_751), .Y(n_825) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_761), .B1(n_763), .B2(n_764), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_761), .A2(n_764), .B1(n_797), .B2(n_798), .Y(n_834) );
AND2x4_ASAP7_75t_L g1368 ( .A(n_762), .B(n_1077), .Y(n_1368) );
CKINVDCx11_ASAP7_75t_R g764 ( .A(n_765), .Y(n_764) );
OAI221xp5_ASAP7_75t_L g836 ( .A1(n_769), .A2(n_837), .B1(n_838), .B2(n_839), .C(n_841), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_774), .B1(n_775), .B2(n_778), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
CKINVDCx5p33_ASAP7_75t_R g775 ( .A(n_776), .Y(n_775) );
BUFx3_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx2_ASAP7_75t_L g894 ( .A(n_777), .Y(n_894) );
AND2x4_ASAP7_75t_L g1064 ( .A(n_777), .B(n_1065), .Y(n_1064) );
NOR2xp33_ASAP7_75t_L g784 ( .A(n_785), .B(n_787), .Y(n_784) );
INVx1_ASAP7_75t_L g852 ( .A(n_792), .Y(n_852) );
AND3x1_ASAP7_75t_L g793 ( .A(n_794), .B(n_820), .C(n_822), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g794 ( .A(n_795), .B(n_813), .Y(n_794) );
AOI33xp33_ASAP7_75t_L g800 ( .A1(n_801), .A2(n_802), .A3(n_805), .B1(n_809), .B2(n_811), .B3(n_812), .Y(n_800) );
AOI33xp33_ASAP7_75t_L g1006 ( .A1(n_801), .A2(n_812), .A3(n_1007), .B1(n_1008), .B2(n_1011), .B3(n_1012), .Y(n_1006) );
INVx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_814), .B(n_817), .Y(n_813) );
OAI221xp5_ASAP7_75t_L g824 ( .A1(n_815), .A2(n_819), .B1(n_825), .B2(n_826), .C(n_830), .Y(n_824) );
OAI31xp33_ASAP7_75t_L g822 ( .A1(n_823), .A2(n_835), .A3(n_849), .B(n_850), .Y(n_822) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
HB1xp67_ASAP7_75t_L g1379 ( .A(n_829), .Y(n_1379) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
AND2x4_ASAP7_75t_L g1070 ( .A(n_833), .B(n_1065), .Y(n_1070) );
BUFx3_ASAP7_75t_L g1453 ( .A(n_833), .Y(n_1453) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g842 ( .A1(n_843), .A2(n_844), .B1(n_845), .B2(n_846), .Y(n_842) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
BUFx3_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx4_ASAP7_75t_L g998 ( .A(n_848), .Y(n_998) );
INVx2_ASAP7_75t_SL g1096 ( .A(n_848), .Y(n_1096) );
INVx2_ASAP7_75t_SL g1099 ( .A(n_848), .Y(n_1099) );
OAI21xp5_ASAP7_75t_L g928 ( .A1(n_850), .A2(n_929), .B(n_939), .Y(n_928) );
BUFx8_ASAP7_75t_SL g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
OAI22x1_ASAP7_75t_L g855 ( .A1(n_856), .A2(n_857), .B1(n_909), .B2(n_910), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g908 ( .A(n_859), .Y(n_908) );
NAND3xp33_ASAP7_75t_L g860 ( .A(n_861), .B(n_866), .C(n_869), .Y(n_860) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
NAND4xp25_ASAP7_75t_L g883 ( .A(n_884), .B(n_890), .C(n_898), .D(n_903), .Y(n_883) );
INVx2_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
INVx1_ASAP7_75t_L g1045 ( .A(n_897), .Y(n_1045) );
NAND3xp33_ASAP7_75t_L g903 ( .A(n_904), .B(n_905), .C(n_906), .Y(n_903) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
INVx2_ASAP7_75t_SL g909 ( .A(n_910), .Y(n_909) );
INVx2_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
NAND4xp75_ASAP7_75t_L g912 ( .A(n_913), .B(n_928), .C(n_950), .D(n_952), .Y(n_912) );
AND2x2_ASAP7_75t_L g913 ( .A(n_914), .B(n_924), .Y(n_913) );
INVx2_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_930), .B(n_933), .Y(n_929) );
BUFx3_ASAP7_75t_L g1449 ( .A(n_935), .Y(n_1449) );
AND2x6_ASAP7_75t_L g1067 ( .A(n_937), .B(n_1065), .Y(n_1067) );
NAND2x1p5_ASAP7_75t_L g1082 ( .A(n_937), .B(n_1077), .Y(n_1082) );
NAND2x1_ASAP7_75t_SL g1076 ( .A(n_948), .B(n_1077), .Y(n_1076) );
INVx2_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
INVx1_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
AOI22xp33_ASAP7_75t_SL g956 ( .A1(n_957), .A2(n_958), .B1(n_1056), .B2(n_1057), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
OAI22xp5_ASAP7_75t_L g958 ( .A1(n_959), .A2(n_960), .B1(n_1013), .B2(n_1055), .Y(n_958) );
INVx2_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
NAND4xp25_ASAP7_75t_SL g962 ( .A(n_963), .B(n_966), .C(n_969), .D(n_976), .Y(n_962) );
INVx1_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
BUFx4f_ASAP7_75t_L g1023 ( .A(n_974), .Y(n_1023) );
NAND4xp25_ASAP7_75t_L g1015 ( .A(n_976), .B(n_1016), .C(n_1019), .D(n_1025), .Y(n_1015) );
NAND4xp25_ASAP7_75t_L g1431 ( .A(n_976), .B(n_1432), .C(n_1435), .D(n_1438), .Y(n_1431) );
NAND2xp5_ASAP7_75t_L g988 ( .A(n_989), .B(n_1006), .Y(n_988) );
BUFx3_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
INVx2_ASAP7_75t_L g1447 ( .A(n_991), .Y(n_1447) );
INVx2_ASAP7_75t_SL g997 ( .A(n_998), .Y(n_997) );
INVx3_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
INVx2_ASAP7_75t_SL g1001 ( .A(n_1002), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_1002), .B(n_1065), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1389 ( .A(n_1002), .B(n_1065), .Y(n_1389) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
BUFx3_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
INVx2_ASAP7_75t_L g1055 ( .A(n_1013), .Y(n_1055) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1014), .Y(n_1054) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1034), .Y(n_1028) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
INVx3_ASAP7_75t_SL g1056 ( .A(n_1057), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1105), .Y(n_1058) );
NOR3xp33_ASAP7_75t_L g1059 ( .A(n_1060), .B(n_1073), .C(n_1083), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1068), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g1061 ( .A1(n_1062), .A2(n_1063), .B1(n_1066), .B2(n_1067), .Y(n_1061) );
BUFx2_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
BUFx2_ASAP7_75t_L g1384 ( .A(n_1064), .Y(n_1384) );
OAI221xp5_ASAP7_75t_L g1124 ( .A1(n_1066), .A2(n_1069), .B1(n_1125), .B2(n_1126), .C(n_1127), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g1382 ( .A1(n_1067), .A2(n_1383), .B1(n_1384), .B2(n_1385), .Y(n_1382) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_1069), .A2(n_1070), .B1(n_1071), .B2(n_1072), .Y(n_1068) );
AOI22xp33_ASAP7_75t_L g1386 ( .A1(n_1070), .A2(n_1387), .B1(n_1388), .B2(n_1389), .Y(n_1386) );
INVx2_ASAP7_75t_L g1074 ( .A(n_1075), .Y(n_1074) );
INVx2_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
INVx3_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
BUFx4f_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
BUFx2_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
OAI22xp33_ASAP7_75t_L g1084 ( .A1(n_1085), .A2(n_1088), .B1(n_1089), .B2(n_1091), .Y(n_1084) );
OAI22xp33_ASAP7_75t_L g1101 ( .A1(n_1085), .A2(n_1102), .B1(n_1103), .B2(n_1104), .Y(n_1101) );
BUFx2_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
INVx2_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1090), .Y(n_1103) );
OAI22xp5_ASAP7_75t_L g1092 ( .A1(n_1093), .A2(n_1094), .B1(n_1095), .B2(n_1096), .Y(n_1092) );
OAI22xp5_ASAP7_75t_L g1097 ( .A1(n_1094), .A2(n_1098), .B1(n_1099), .B2(n_1100), .Y(n_1097) );
AOI211xp5_ASAP7_75t_L g1112 ( .A1(n_1098), .A2(n_1113), .B(n_1115), .C(n_1121), .Y(n_1112) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1099), .Y(n_1455) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_1100), .A2(n_1102), .B1(n_1144), .B2(n_1146), .Y(n_1143) );
AOI221xp5_ASAP7_75t_L g1129 ( .A1(n_1104), .A2(n_1130), .B1(n_1133), .B2(n_1137), .C(n_1141), .Y(n_1129) );
AOI21xp5_ASAP7_75t_L g1105 ( .A1(n_1106), .A2(n_1110), .B(n_1111), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
INVx2_ASAP7_75t_L g1422 ( .A(n_1107), .Y(n_1422) );
AND2x4_ASAP7_75t_L g1107 ( .A(n_1108), .B(n_1109), .Y(n_1107) );
AOI31xp33_ASAP7_75t_L g1111 ( .A1(n_1112), .A2(n_1129), .A3(n_1143), .B(n_1148), .Y(n_1111) );
INVx2_ASAP7_75t_SL g1116 ( .A(n_1117), .Y(n_1116) );
INVx1_ASAP7_75t_SL g1142 ( .A(n_1120), .Y(n_1142) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1131), .Y(n_1130) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
HB1xp67_ASAP7_75t_L g1409 ( .A(n_1132), .Y(n_1409) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
INVx2_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
AOI22xp33_ASAP7_75t_L g1418 ( .A1(n_1144), .A2(n_1146), .B1(n_1419), .B2(n_1420), .Y(n_1418) );
INVx6_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
INVx4_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1148), .Y(n_1391) );
INVx2_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
OAI21xp5_ASAP7_75t_L g1150 ( .A1(n_1151), .A2(n_1161), .B(n_1362), .Y(n_1150) );
CKINVDCx16_ASAP7_75t_R g1151 ( .A(n_1152), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
OAI22xp33_ASAP7_75t_L g1327 ( .A1(n_1153), .A2(n_1328), .B1(n_1329), .B2(n_1330), .Y(n_1327) );
BUFx3_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
OAI22xp5_ASAP7_75t_L g1188 ( .A1(n_1154), .A2(n_1189), .B1(n_1190), .B2(n_1191), .Y(n_1188) );
OAI22xp33_ASAP7_75t_L g1193 ( .A1(n_1154), .A2(n_1191), .B1(n_1194), .B2(n_1195), .Y(n_1193) );
OAI22xp33_ASAP7_75t_L g1206 ( .A1(n_1154), .A2(n_1207), .B1(n_1208), .B2(n_1209), .Y(n_1206) );
BUFx6f_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
OR2x2_ASAP7_75t_L g1155 ( .A(n_1156), .B(n_1157), .Y(n_1155) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1156), .Y(n_1171) );
OR2x2_ASAP7_75t_L g1191 ( .A(n_1156), .B(n_1174), .Y(n_1191) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1157), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1158), .B(n_1160), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1160), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1162), .B(n_1290), .Y(n_1161) );
NOR2xp33_ASAP7_75t_L g1162 ( .A(n_1163), .B(n_1272), .Y(n_1162) );
NAND3xp33_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1229), .C(n_1258), .Y(n_1163) );
O2A1O1Ixp33_ASAP7_75t_L g1164 ( .A1(n_1165), .A2(n_1196), .B(n_1201), .C(n_1215), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1166), .B(n_1181), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1217 ( .A(n_1166), .B(n_1218), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1166), .B(n_1239), .Y(n_1238) );
NOR2xp33_ASAP7_75t_L g1256 ( .A(n_1166), .B(n_1202), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1166), .B(n_1182), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_1166), .B(n_1257), .Y(n_1271) );
OAI332xp33_ASAP7_75t_L g1294 ( .A1(n_1166), .A2(n_1226), .A3(n_1245), .B1(n_1246), .B2(n_1295), .B3(n_1298), .C1(n_1299), .C2(n_1301), .Y(n_1294) );
OAI32xp33_ASAP7_75t_L g1355 ( .A1(n_1166), .A2(n_1287), .A3(n_1312), .B1(n_1341), .B2(n_1356), .Y(n_1355) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1166), .Y(n_1357) );
INVx4_ASAP7_75t_L g1166 ( .A(n_1167), .Y(n_1166) );
NAND2xp5_ASAP7_75t_L g1198 ( .A(n_1167), .B(n_1199), .Y(n_1198) );
NAND2xp5_ASAP7_75t_L g1226 ( .A(n_1167), .B(n_1218), .Y(n_1226) );
INVx3_ASAP7_75t_L g1244 ( .A(n_1167), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1167), .B(n_1246), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1167), .B(n_1266), .Y(n_1281) );
OR2x2_ASAP7_75t_L g1310 ( .A(n_1167), .B(n_1218), .Y(n_1310) );
NOR2xp33_ASAP7_75t_L g1352 ( .A(n_1167), .B(n_1297), .Y(n_1352) );
NAND3xp33_ASAP7_75t_L g1359 ( .A(n_1167), .B(n_1342), .C(n_1353), .Y(n_1359) );
NOR3xp33_ASAP7_75t_L g1360 ( .A(n_1167), .B(n_1240), .C(n_1361), .Y(n_1360) );
AND2x4_ASAP7_75t_L g1167 ( .A(n_1168), .B(n_1175), .Y(n_1167) );
AND2x4_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1171), .Y(n_1169) );
OAI21xp33_ASAP7_75t_SL g1482 ( .A1(n_1170), .A2(n_1481), .B(n_1483), .Y(n_1482) );
AND2x4_ASAP7_75t_L g1172 ( .A(n_1171), .B(n_1173), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1176), .Y(n_1326) );
AND2x4_ASAP7_75t_L g1176 ( .A(n_1177), .B(n_1179), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1177), .B(n_1179), .Y(n_1213) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
AND2x4_ASAP7_75t_L g1180 ( .A(n_1178), .B(n_1179), .Y(n_1180) );
INVx2_ASAP7_75t_L g1205 ( .A(n_1180), .Y(n_1205) );
OAI21xp5_ASAP7_75t_L g1223 ( .A1(n_1181), .A2(n_1224), .B(n_1225), .Y(n_1223) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1181), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1181), .B(n_1243), .Y(n_1315) );
AOI221xp5_ASAP7_75t_L g1350 ( .A1(n_1181), .A2(n_1249), .B1(n_1344), .B2(n_1351), .C(n_1352), .Y(n_1350) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1182), .B(n_1186), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1182), .B(n_1197), .Y(n_1196) );
NOR2x1_ASAP7_75t_L g1239 ( .A(n_1182), .B(n_1240), .Y(n_1239) );
NAND2xp5_ASAP7_75t_L g1254 ( .A(n_1182), .B(n_1240), .Y(n_1254) );
NAND2xp5_ASAP7_75t_L g1275 ( .A(n_1182), .B(n_1265), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1182), .B(n_1235), .Y(n_1300) );
OR2x2_ASAP7_75t_L g1303 ( .A(n_1182), .B(n_1304), .Y(n_1303) );
INVx2_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1183), .B(n_1186), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1224 ( .A(n_1183), .B(n_1199), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1183), .B(n_1234), .Y(n_1233) );
BUFx3_ASAP7_75t_L g1246 ( .A(n_1183), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1183), .B(n_1240), .Y(n_1270) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1183), .B(n_1265), .Y(n_1279) );
OR2x2_ASAP7_75t_L g1339 ( .A(n_1183), .B(n_1340), .Y(n_1339) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1184), .B(n_1185), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1186), .B(n_1252), .Y(n_1251) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1186), .Y(n_1297) );
OAI21xp5_ASAP7_75t_L g1343 ( .A1(n_1186), .A2(n_1300), .B(n_1344), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1192), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1199 ( .A(n_1187), .B(n_1200), .Y(n_1199) );
INVx2_ASAP7_75t_L g1235 ( .A(n_1187), .Y(n_1235) );
HB1xp67_ASAP7_75t_L g1209 ( .A(n_1191), .Y(n_1209) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1191), .Y(n_1331) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1192), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1192), .B(n_1235), .Y(n_1234) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1192), .Y(n_1240) );
AOI221xp5_ASAP7_75t_L g1276 ( .A1(n_1196), .A2(n_1257), .B1(n_1277), .B2(n_1281), .C(n_1282), .Y(n_1276) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1198), .Y(n_1197) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1199), .Y(n_1340) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1200), .B(n_1235), .Y(n_1265) );
NAND3xp33_ASAP7_75t_L g1250 ( .A(n_1201), .B(n_1248), .C(n_1251), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g1319 ( .A(n_1201), .B(n_1249), .Y(n_1319) );
AND2x4_ASAP7_75t_SL g1201 ( .A(n_1202), .B(n_1210), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1202), .B(n_1211), .Y(n_1231) );
OR2x2_ASAP7_75t_L g1287 ( .A(n_1202), .B(n_1210), .Y(n_1287) );
INVx2_ASAP7_75t_SL g1202 ( .A(n_1203), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1203), .B(n_1210), .Y(n_1228) );
OR2x2_ASAP7_75t_L g1247 ( .A(n_1203), .B(n_1248), .Y(n_1247) );
INVx2_ASAP7_75t_L g1284 ( .A(n_1203), .Y(n_1284) );
INVx2_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1210), .B(n_1249), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1342 ( .A(n_1210), .B(n_1218), .Y(n_1342) );
CKINVDCx6p67_ASAP7_75t_R g1210 ( .A(n_1211), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1211), .B(n_1218), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1211), .B(n_1267), .Y(n_1266) );
CKINVDCx5p33_ASAP7_75t_R g1301 ( .A(n_1211), .Y(n_1301) );
OR2x6_ASAP7_75t_L g1211 ( .A(n_1212), .B(n_1214), .Y(n_1211) );
O2A1O1Ixp33_ASAP7_75t_L g1215 ( .A1(n_1216), .A2(n_1221), .B(n_1223), .C(n_1227), .Y(n_1215) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1217), .B(n_1265), .Y(n_1306) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1218), .Y(n_1232) );
CKINVDCx5p33_ASAP7_75t_R g1249 ( .A(n_1218), .Y(n_1249) );
INVx1_ASAP7_75t_SL g1267 ( .A(n_1218), .Y(n_1267) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1219), .B(n_1220), .Y(n_1218) );
AOI21xp33_ASAP7_75t_SL g1253 ( .A1(n_1221), .A2(n_1254), .B(n_1255), .Y(n_1253) );
NOR2xp33_ASAP7_75t_L g1337 ( .A(n_1221), .B(n_1249), .Y(n_1337) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1222), .Y(n_1221) );
AOI21xp5_ASAP7_75t_L g1316 ( .A1(n_1222), .A2(n_1317), .B(n_1318), .Y(n_1316) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_1222), .B(n_1293), .Y(n_1336) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1224), .B(n_1283), .Y(n_1282) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1226), .Y(n_1225) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1228), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1273 ( .A(n_1228), .B(n_1267), .Y(n_1273) );
NAND2xp5_ASAP7_75t_L g1305 ( .A(n_1228), .B(n_1306), .Y(n_1305) );
NAND2xp5_ASAP7_75t_L g1335 ( .A(n_1228), .B(n_1244), .Y(n_1335) );
AOI211xp5_ASAP7_75t_SL g1229 ( .A1(n_1230), .A2(n_1233), .B(n_1236), .C(n_1253), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1231), .B(n_1232), .Y(n_1230) );
INVx2_ASAP7_75t_L g1241 ( .A(n_1231), .Y(n_1241) );
NAND3xp33_ASAP7_75t_L g1356 ( .A(n_1232), .B(n_1351), .C(n_1357), .Y(n_1356) );
NAND2xp5_ASAP7_75t_L g1260 ( .A(n_1234), .B(n_1261), .Y(n_1260) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_1234), .B(n_1244), .Y(n_1304) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1234), .Y(n_1321) );
INVx2_ASAP7_75t_L g1351 ( .A(n_1235), .Y(n_1351) );
OAI221xp5_ASAP7_75t_L g1236 ( .A1(n_1237), .A2(n_1241), .B1(n_1242), .B2(n_1247), .C(n_1250), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
OR2x2_ASAP7_75t_L g1245 ( .A(n_1240), .B(n_1246), .Y(n_1245) );
AOI222xp33_ASAP7_75t_L g1354 ( .A1(n_1240), .A2(n_1262), .B1(n_1324), .B2(n_1355), .C1(n_1358), .C2(n_1360), .Y(n_1354) );
OR2x2_ASAP7_75t_L g1242 ( .A(n_1243), .B(n_1245), .Y(n_1242) );
NAND2xp5_ASAP7_75t_L g1311 ( .A(n_1243), .B(n_1262), .Y(n_1311) );
INVx2_ASAP7_75t_L g1243 ( .A(n_1244), .Y(n_1243) );
OR2x2_ASAP7_75t_L g1274 ( .A(n_1244), .B(n_1275), .Y(n_1274) );
NAND2xp5_ASAP7_75t_L g1289 ( .A(n_1244), .B(n_1279), .Y(n_1289) );
NAND2xp5_ASAP7_75t_L g1348 ( .A(n_1244), .B(n_1300), .Y(n_1348) );
OR2x2_ASAP7_75t_L g1320 ( .A(n_1246), .B(n_1321), .Y(n_1320) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1247), .Y(n_1317) );
INVx3_ASAP7_75t_L g1248 ( .A(n_1249), .Y(n_1248) );
NOR2xp33_ASAP7_75t_L g1346 ( .A(n_1249), .B(n_1289), .Y(n_1346) );
NAND2xp5_ASAP7_75t_L g1255 ( .A(n_1256), .B(n_1257), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1257), .B(n_1284), .Y(n_1283) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1257), .Y(n_1298) );
AOI221xp5_ASAP7_75t_L g1258 ( .A1(n_1259), .A2(n_1262), .B1(n_1263), .B2(n_1266), .C(n_1268), .Y(n_1258) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
NAND2xp5_ASAP7_75t_L g1264 ( .A(n_1261), .B(n_1265), .Y(n_1264) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1265), .Y(n_1296) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1266), .Y(n_1349) );
INVxp67_ASAP7_75t_SL g1268 ( .A(n_1269), .Y(n_1268) );
NAND2xp5_ASAP7_75t_L g1269 ( .A(n_1270), .B(n_1271), .Y(n_1269) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1270), .Y(n_1312) );
OAI211xp5_ASAP7_75t_L g1272 ( .A1(n_1273), .A2(n_1274), .B(n_1276), .C(n_1285), .Y(n_1272) );
OAI221xp5_ASAP7_75t_L g1334 ( .A1(n_1273), .A2(n_1299), .B1(n_1320), .B2(n_1335), .C(n_1336), .Y(n_1334) );
NAND2xp5_ASAP7_75t_L g1277 ( .A(n_1278), .B(n_1280), .Y(n_1277) );
OAI221xp5_ASAP7_75t_L g1302 ( .A1(n_1278), .A2(n_1287), .B1(n_1301), .B2(n_1303), .C(n_1305), .Y(n_1302) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
INVx2_ASAP7_75t_L g1293 ( .A(n_1284), .Y(n_1293) );
NOR2xp33_ASAP7_75t_L g1309 ( .A(n_1284), .B(n_1310), .Y(n_1309) );
INVx2_ASAP7_75t_L g1314 ( .A(n_1284), .Y(n_1314) );
OAI31xp33_ASAP7_75t_L g1338 ( .A1(n_1284), .A2(n_1339), .A3(n_1341), .B(n_1343), .Y(n_1338) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1284), .B(n_1324), .Y(n_1353) );
NAND2xp5_ASAP7_75t_L g1285 ( .A(n_1286), .B(n_1288), .Y(n_1285) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
AOI21xp5_ASAP7_75t_L g1290 ( .A1(n_1291), .A2(n_1322), .B(n_1332), .Y(n_1290) );
NAND3xp33_ASAP7_75t_L g1291 ( .A(n_1292), .B(n_1313), .C(n_1316), .Y(n_1291) );
AOI211xp5_ASAP7_75t_L g1292 ( .A1(n_1293), .A2(n_1294), .B(n_1302), .C(n_1307), .Y(n_1292) );
NAND2xp5_ASAP7_75t_L g1295 ( .A(n_1296), .B(n_1297), .Y(n_1295) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1300), .Y(n_1299) );
OAI221xp5_ASAP7_75t_SL g1347 ( .A1(n_1301), .A2(n_1321), .B1(n_1348), .B2(n_1349), .C(n_1350), .Y(n_1347) );
AOI21xp33_ASAP7_75t_SL g1307 ( .A1(n_1308), .A2(n_1311), .B(n_1312), .Y(n_1307) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1309), .Y(n_1308) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1310), .Y(n_1344) );
NAND2xp5_ASAP7_75t_L g1313 ( .A(n_1314), .B(n_1315), .Y(n_1313) );
NOR2xp33_ASAP7_75t_L g1318 ( .A(n_1319), .B(n_1320), .Y(n_1318) );
INVx2_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
OAI31xp33_ASAP7_75t_L g1333 ( .A1(n_1323), .A2(n_1334), .A3(n_1337), .B(n_1338), .Y(n_1333) );
BUFx3_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1324), .Y(n_1361) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
XNOR2x1_ASAP7_75t_L g1364 ( .A(n_1328), .B(n_1365), .Y(n_1364) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
NAND3xp33_ASAP7_75t_L g1332 ( .A(n_1333), .B(n_1345), .C(n_1354), .Y(n_1332) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
OAI21xp33_ASAP7_75t_L g1345 ( .A1(n_1346), .A2(n_1347), .B(n_1353), .Y(n_1345) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1364), .Y(n_1363) );
NAND2x1_ASAP7_75t_L g1365 ( .A(n_1366), .B(n_1390), .Y(n_1365) );
AND4x1_ASAP7_75t_L g1366 ( .A(n_1367), .B(n_1373), .C(n_1382), .D(n_1386), .Y(n_1366) );
AOI221xp5_ASAP7_75t_L g1367 ( .A1(n_1368), .A2(n_1369), .B1(n_1370), .B2(n_1371), .C(n_1372), .Y(n_1367) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
OAI211xp5_ASAP7_75t_L g1403 ( .A1(n_1385), .A2(n_1404), .B(n_1405), .C(n_1406), .Y(n_1403) );
AOI22xp5_ASAP7_75t_L g1390 ( .A1(n_1391), .A2(n_1392), .B1(n_1421), .B2(n_1422), .Y(n_1390) );
NAND3xp33_ASAP7_75t_L g1392 ( .A(n_1393), .B(n_1408), .C(n_1418), .Y(n_1392) );
AOI21xp5_ASAP7_75t_SL g1393 ( .A1(n_1394), .A2(n_1397), .B(n_1398), .Y(n_1393) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1395), .Y(n_1394) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1396), .Y(n_1395) );
INVx4_ASAP7_75t_L g1399 ( .A(n_1400), .Y(n_1399) );
INVx2_ASAP7_75t_SL g1401 ( .A(n_1402), .Y(n_1401) );
AOI221xp5_ASAP7_75t_L g1408 ( .A1(n_1409), .A2(n_1410), .B1(n_1411), .B2(n_1414), .C(n_1416), .Y(n_1408) );
INVxp67_ASAP7_75t_L g1412 ( .A(n_1413), .Y(n_1412) );
BUFx2_ASAP7_75t_L g1423 ( .A(n_1424), .Y(n_1423) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1425), .Y(n_1424) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1426), .Y(n_1425) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1429), .Y(n_1479) );
HB1xp67_ASAP7_75t_L g1429 ( .A(n_1430), .Y(n_1429) );
AOI211x1_ASAP7_75t_L g1430 ( .A1(n_1431), .A2(n_1442), .B(n_1444), .C(n_1470), .Y(n_1430) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1443), .Y(n_1442) );
NAND2xp5_ASAP7_75t_L g1444 ( .A(n_1445), .B(n_1457), .Y(n_1444) );
INVx2_ASAP7_75t_L g1446 ( .A(n_1447), .Y(n_1446) );
HB1xp67_ASAP7_75t_L g1450 ( .A(n_1451), .Y(n_1450) );
BUFx3_ASAP7_75t_L g1459 ( .A(n_1460), .Y(n_1459) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1462), .Y(n_1461) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
endmodule