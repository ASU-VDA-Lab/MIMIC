module fake_jpeg_12067_n_632 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_632);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_632;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_0),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_10),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_62),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_63),
.B(n_75),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_64),
.Y(n_175)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_65),
.Y(n_157)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

BUFx8_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_67),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_68),
.Y(n_188)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_69),
.Y(n_189)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_70),
.Y(n_134)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_73),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_74),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_9),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_76),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_77),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_78),
.Y(n_199)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_23),
.B(n_9),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_80),
.B(n_92),
.Y(n_174)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_82),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_83),
.Y(n_187)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_87),
.Y(n_159)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_88),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_59),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_89),
.A2(n_35),
.B1(n_55),
.B2(n_33),
.Y(n_164)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_90),
.Y(n_168)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_91),
.Y(n_150)
);

BUFx4f_ASAP7_75t_SL g92 ( 
.A(n_48),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_93),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_23),
.B(n_36),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_94),
.B(n_97),
.Y(n_178)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_96),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_34),
.B(n_8),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_98),
.Y(n_180)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_99),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_34),
.B(n_8),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_100),
.B(n_12),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_101),
.Y(n_195)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_25),
.Y(n_105)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

INVx6_ASAP7_75t_SL g106 ( 
.A(n_37),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_106),
.Y(n_165)
);

AOI21xp33_ASAP7_75t_SL g107 ( 
.A1(n_37),
.A2(n_7),
.B(n_16),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g145 ( 
.A(n_107),
.B(n_10),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_42),
.Y(n_108)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_108),
.Y(n_205)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_22),
.Y(n_109)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_109),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_22),
.Y(n_110)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_111),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_45),
.Y(n_112)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_112),
.Y(n_202)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_45),
.Y(n_113)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_45),
.Y(n_114)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_114),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_45),
.Y(n_115)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_115),
.Y(n_192)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_25),
.Y(n_116)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_21),
.Y(n_117)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_22),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_118),
.B(n_25),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_21),
.Y(n_119)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_49),
.Y(n_120)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_21),
.Y(n_121)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_121),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_122),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_19),
.Y(n_123)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_123),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_124),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_75),
.B(n_36),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_131),
.B(n_138),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_65),
.A2(n_59),
.B1(n_35),
.B2(n_50),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_136),
.A2(n_179),
.B1(n_184),
.B2(n_190),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_46),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_119),
.A2(n_58),
.B1(n_46),
.B2(n_57),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_139),
.A2(n_164),
.B1(n_170),
.B2(n_198),
.Y(n_261)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_141),
.Y(n_207)
);

HAxp5_ASAP7_75t_SL g144 ( 
.A(n_89),
.B(n_59),
.CON(n_144),
.SN(n_144)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_144),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_145),
.B(n_7),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_69),
.A2(n_35),
.B1(n_30),
.B2(n_18),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_166),
.A2(n_38),
.B1(n_33),
.B2(n_55),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_L g170 ( 
.A1(n_62),
.A2(n_50),
.B1(n_35),
.B2(n_57),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_88),
.B(n_18),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_173),
.B(n_25),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_76),
.A2(n_50),
.B1(n_57),
.B2(n_28),
.Y(n_179)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_121),
.Y(n_183)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_60),
.A2(n_28),
.B1(n_25),
.B2(n_31),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_122),
.Y(n_185)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_185),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_78),
.A2(n_28),
.B1(n_25),
.B2(n_31),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_124),
.Y(n_191)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_191),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_194),
.Y(n_240)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_117),
.Y(n_197)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_197),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_64),
.A2(n_38),
.B1(n_30),
.B2(n_56),
.Y(n_198)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_68),
.Y(n_200)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_200),
.Y(n_242)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_73),
.Y(n_201)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_203),
.B(n_11),
.Y(n_247)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_146),
.Y(n_206)
);

INVx6_ASAP7_75t_L g306 ( 
.A(n_206),
.Y(n_306)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_156),
.Y(n_208)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_208),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_209),
.A2(n_221),
.B1(n_228),
.B2(n_244),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_118),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_211),
.B(n_218),
.Y(n_287)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_213),
.Y(n_293)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_129),
.Y(n_214)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_214),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_216),
.B(n_247),
.Y(n_316)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_125),
.Y(n_217)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_217),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_178),
.B(n_56),
.Y(n_218)
);

AOI21xp33_ASAP7_75t_L g312 ( 
.A1(n_219),
.A2(n_273),
.B(n_280),
.Y(n_312)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_132),
.Y(n_220)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_220),
.Y(n_324)
);

OAI22xp33_ASAP7_75t_L g221 ( 
.A1(n_166),
.A2(n_83),
.B1(n_115),
.B2(n_114),
.Y(n_221)
);

INVx11_ASAP7_75t_L g222 ( 
.A(n_157),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_222),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_145),
.B(n_51),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_223),
.B(n_248),
.C(n_111),
.Y(n_326)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_151),
.Y(n_224)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_224),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_143),
.B(n_67),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_225),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_169),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_226),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_143),
.A2(n_77),
.B1(n_93),
.B2(n_112),
.Y(n_228)
);

INVx11_ASAP7_75t_L g229 ( 
.A(n_157),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_229),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_174),
.B(n_118),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_230),
.B(n_245),
.Y(n_289)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_159),
.Y(n_231)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_231),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_169),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_232),
.B(n_237),
.Y(n_285)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_130),
.Y(n_233)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_233),
.Y(n_291)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_204),
.Y(n_235)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_235),
.Y(n_317)
);

OAI32xp33_ASAP7_75t_L g237 ( 
.A1(n_174),
.A2(n_113),
.A3(n_96),
.B1(n_108),
.B2(n_101),
.Y(n_237)
);

INVx13_ASAP7_75t_L g238 ( 
.A(n_181),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_238),
.Y(n_295)
);

BUFx4f_ASAP7_75t_L g239 ( 
.A(n_172),
.Y(n_239)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_239),
.Y(n_299)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_154),
.Y(n_241)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_241),
.Y(n_300)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_179),
.A2(n_98),
.B1(n_110),
.B2(n_19),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_128),
.B(n_40),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_150),
.Y(n_246)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_246),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_133),
.B(n_26),
.C(n_40),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_155),
.Y(n_249)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_249),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_165),
.B(n_92),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_251),
.Y(n_305)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_153),
.Y(n_252)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_252),
.Y(n_335)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_181),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_253),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_142),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_254),
.Y(n_340)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_177),
.Y(n_255)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_255),
.Y(n_325)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_158),
.Y(n_256)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_256),
.Y(n_339)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_186),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_257),
.B(n_264),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_144),
.A2(n_47),
.B1(n_31),
.B2(n_29),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_258),
.A2(n_55),
.B1(n_33),
.B2(n_127),
.Y(n_290)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_146),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_259),
.Y(n_309)
);

BUFx10_ASAP7_75t_L g260 ( 
.A(n_148),
.Y(n_260)
);

INVx8_ASAP7_75t_L g308 ( 
.A(n_260),
.Y(n_308)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_163),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_262),
.B(n_272),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_135),
.A2(n_52),
.B1(n_47),
.B2(n_29),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_263),
.A2(n_278),
.B(n_82),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_175),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_134),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_265),
.B(n_266),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_194),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_137),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_267),
.B(n_269),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_170),
.A2(n_176),
.B1(n_161),
.B2(n_171),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_268),
.A2(n_189),
.B1(n_188),
.B2(n_175),
.Y(n_319)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_140),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_180),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_270),
.B(n_271),
.Y(n_337)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_147),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_162),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_136),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_195),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_274),
.Y(n_286)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_182),
.Y(n_275)
);

NAND2xp33_ASAP7_75t_R g323 ( 
.A(n_275),
.B(n_276),
.Y(n_323)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_202),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_199),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_277),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_184),
.A2(n_52),
.B1(n_47),
.B2(n_29),
.Y(n_278)
);

O2A1O1Ixp33_ASAP7_75t_L g279 ( 
.A1(n_190),
.A2(n_67),
.B(n_52),
.C(n_26),
.Y(n_279)
);

O2A1O1Ixp33_ASAP7_75t_L g294 ( 
.A1(n_279),
.A2(n_273),
.B(n_222),
.C(n_229),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_126),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_210),
.B(n_167),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_282),
.B(n_296),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_290),
.A2(n_297),
.B1(n_311),
.B2(n_322),
.Y(n_358)
);

O2A1O1Ixp33_ASAP7_75t_L g385 ( 
.A1(n_294),
.A2(n_281),
.B(n_295),
.C(n_323),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_223),
.B(n_192),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_250),
.A2(n_149),
.B1(n_196),
.B2(n_160),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_248),
.B(n_187),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_301),
.B(n_307),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_219),
.B(n_187),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_221),
.A2(n_196),
.B1(n_160),
.B2(n_149),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_225),
.B(n_152),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_313),
.B(n_224),
.C(n_214),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_238),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_314),
.B(n_333),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_240),
.B(n_189),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_318),
.B(n_320),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_319),
.A2(n_259),
.B1(n_206),
.B2(n_264),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_240),
.B(n_207),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_244),
.A2(n_188),
.B1(n_205),
.B2(n_168),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_326),
.B(n_213),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_261),
.B(n_0),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_327),
.B(n_311),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_212),
.A2(n_82),
.B1(n_6),
.B2(n_12),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_331),
.A2(n_334),
.B(n_268),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_260),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_261),
.A2(n_14),
.B1(n_17),
.B2(n_2),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_336),
.A2(n_243),
.B1(n_242),
.B2(n_215),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_334),
.A2(n_212),
.B(n_279),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_344),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g345 ( 
.A(n_320),
.B(n_278),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_345),
.B(n_364),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_327),
.A2(n_285),
.B1(n_288),
.B2(n_301),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_346),
.A2(n_352),
.B1(n_365),
.B2(n_315),
.Y(n_400)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_332),
.Y(n_347)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_347),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_348),
.B(n_359),
.Y(n_391)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_321),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_349),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g412 ( 
.A(n_350),
.B(n_341),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_351),
.B(n_388),
.C(n_313),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_288),
.A2(n_263),
.B1(n_227),
.B2(n_234),
.Y(n_352)
);

BUFx5_ASAP7_75t_L g354 ( 
.A(n_306),
.Y(n_354)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_354),
.Y(n_398)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_332),
.Y(n_355)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_355),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_356),
.A2(n_360),
.B1(n_387),
.B2(n_315),
.Y(n_401)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_335),
.Y(n_357)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_357),
.Y(n_423)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_335),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_294),
.A2(n_254),
.B1(n_270),
.B2(n_274),
.Y(n_360)
);

BUFx24_ASAP7_75t_L g361 ( 
.A(n_295),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_361),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_362),
.A2(n_299),
.B1(n_302),
.B2(n_300),
.Y(n_430)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_317),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_282),
.A2(n_236),
.B1(n_231),
.B2(n_220),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_287),
.B(n_241),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_366),
.B(n_376),
.Y(n_406)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_317),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_367),
.B(n_369),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_328),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_368),
.B(n_370),
.Y(n_417)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_325),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_312),
.A2(n_305),
.B(n_289),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_371),
.B(n_374),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_292),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_372),
.B(n_373),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_337),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_321),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_325),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_375),
.B(n_378),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_305),
.B(n_280),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_284),
.B(n_277),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_377),
.B(n_379),
.Y(n_429)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_304),
.Y(n_378)
);

AOI32xp33_ASAP7_75t_L g379 ( 
.A1(n_316),
.A2(n_260),
.A3(n_208),
.B1(n_262),
.B2(n_239),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g380 ( 
.A(n_297),
.B(n_303),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_380),
.B(n_382),
.Y(n_411)
);

AO21x2_ASAP7_75t_L g381 ( 
.A1(n_322),
.A2(n_239),
.B(n_1),
.Y(n_381)
);

OA22x2_ASAP7_75t_L g405 ( 
.A1(n_381),
.A2(n_385),
.B1(n_386),
.B2(n_308),
.Y(n_405)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_304),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_296),
.B(n_307),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_383),
.B(n_384),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_310),
.B(n_14),
.Y(n_384)
);

OA22x2_ASAP7_75t_L g386 ( 
.A1(n_290),
.A2(n_14),
.B1(n_17),
.B2(n_3),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_318),
.A2(n_14),
.B1(n_17),
.B2(n_3),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_326),
.B(n_0),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_298),
.B(n_0),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_389),
.B(n_0),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_343),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_395),
.B(n_427),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_397),
.B(n_413),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_351),
.B(n_291),
.C(n_329),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_399),
.B(n_404),
.C(n_409),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_400),
.B(n_422),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_401),
.A2(n_407),
.B1(n_408),
.B2(n_428),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_346),
.A2(n_331),
.B1(n_286),
.B2(n_306),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_402),
.A2(n_421),
.B1(n_381),
.B2(n_387),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_353),
.B(n_342),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g435 ( 
.A(n_405),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_371),
.A2(n_309),
.B1(n_281),
.B2(n_315),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_345),
.A2(n_309),
.B1(n_338),
.B2(n_341),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_353),
.B(n_304),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_412),
.B(n_419),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_388),
.B(n_342),
.C(n_383),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_344),
.A2(n_340),
.B(n_338),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_418),
.A2(n_390),
.B(n_392),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_350),
.B(n_363),
.C(n_370),
.Y(n_419)
);

OAI22x1_ASAP7_75t_L g420 ( 
.A1(n_380),
.A2(n_308),
.B1(n_324),
.B2(n_293),
.Y(n_420)
);

OA21x2_ASAP7_75t_L g438 ( 
.A1(n_420),
.A2(n_356),
.B(n_382),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_352),
.A2(n_293),
.B1(n_324),
.B2(n_283),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_363),
.B(n_339),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_425),
.B(n_389),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_378),
.B(n_340),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_426),
.B(n_361),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_361),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_381),
.A2(n_283),
.B1(n_339),
.B2(n_302),
.Y(n_428)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_430),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_406),
.B(n_372),
.Y(n_431)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_431),
.Y(n_472)
);

XNOR2x1_ASAP7_75t_SL g432 ( 
.A(n_419),
.B(n_385),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_432),
.B(n_412),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_434),
.B(n_452),
.Y(n_490)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_436),
.Y(n_498)
);

INVx8_ASAP7_75t_L g437 ( 
.A(n_398),
.Y(n_437)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_437),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_438),
.Y(n_492)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_414),
.Y(n_439)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_439),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_391),
.A2(n_358),
.B1(n_348),
.B2(n_373),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_442),
.A2(n_456),
.B1(n_418),
.B2(n_421),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_393),
.Y(n_443)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_443),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_390),
.A2(n_391),
.B(n_411),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_444),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_424),
.B(n_368),
.Y(n_446)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_446),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_447),
.A2(n_459),
.B1(n_462),
.B2(n_428),
.Y(n_468)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_403),
.Y(n_448)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_448),
.Y(n_496)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_403),
.Y(n_449)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_449),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_417),
.B(n_330),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_450),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_404),
.B(n_425),
.Y(n_451)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_451),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_410),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_415),
.Y(n_453)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_453),
.Y(n_483)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_415),
.Y(n_455)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_455),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_391),
.A2(n_381),
.B1(n_357),
.B2(n_367),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_416),
.B(n_330),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_457),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_400),
.A2(n_381),
.B1(n_355),
.B2(n_364),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_396),
.B(n_359),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_460),
.B(n_461),
.Y(n_497)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_423),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_402),
.A2(n_347),
.B1(n_386),
.B2(n_369),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_396),
.B(n_375),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_463),
.Y(n_479)
);

XNOR2x1_ASAP7_75t_L g499 ( 
.A(n_464),
.B(n_374),
.Y(n_499)
);

NOR2x1_ASAP7_75t_L g465 ( 
.A(n_411),
.B(n_361),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g482 ( 
.A(n_465),
.B(n_466),
.Y(n_482)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_423),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_468),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_459),
.A2(n_408),
.B1(n_409),
.B2(n_426),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_469),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_470),
.A2(n_473),
.B1(n_495),
.B2(n_462),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_440),
.A2(n_429),
.B1(n_416),
.B2(n_410),
.Y(n_471)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_471),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_442),
.A2(n_405),
.B1(n_399),
.B2(n_413),
.Y(n_473)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_437),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_481),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_SL g512 ( 
.A(n_484),
.B(n_499),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_441),
.B(n_397),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_486),
.B(n_487),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_441),
.B(n_420),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_458),
.B(n_394),
.C(n_405),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_488),
.B(n_432),
.C(n_464),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_458),
.B(n_454),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_493),
.B(n_465),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_435),
.A2(n_405),
.B1(n_422),
.B2(n_398),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_494),
.B(n_438),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_467),
.A2(n_430),
.B1(n_394),
.B2(n_386),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g502 ( 
.A(n_497),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_502),
.B(n_514),
.Y(n_533)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_497),
.Y(n_503)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_503),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_504),
.B(n_518),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_475),
.B(n_445),
.Y(n_505)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_505),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_506),
.B(n_524),
.Y(n_540)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_477),
.Y(n_507)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_507),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_508),
.B(n_468),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_473),
.A2(n_435),
.B1(n_467),
.B2(n_452),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_509),
.B(n_521),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_493),
.B(n_454),
.C(n_436),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_510),
.B(n_511),
.C(n_517),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_486),
.B(n_444),
.C(n_451),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_482),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_474),
.Y(n_515)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_515),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_499),
.B(n_439),
.C(n_434),
.Y(n_517)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_474),
.Y(n_519)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_519),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_492),
.A2(n_435),
.B1(n_447),
.B2(n_438),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_484),
.B(n_460),
.C(n_463),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_522),
.B(n_529),
.C(n_530),
.Y(n_535)
);

CKINVDCx16_ASAP7_75t_R g523 ( 
.A(n_500),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_523),
.B(n_525),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_SL g524 ( 
.A(n_487),
.B(n_456),
.Y(n_524)
);

CKINVDCx14_ASAP7_75t_R g525 ( 
.A(n_490),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_488),
.B(n_440),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_526),
.B(n_494),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_492),
.A2(n_433),
.B1(n_466),
.B2(n_453),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_528),
.B(n_495),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_469),
.B(n_461),
.C(n_449),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_498),
.B(n_448),
.C(n_455),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_510),
.B(n_480),
.C(n_491),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_537),
.B(n_549),
.Y(n_571)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_538),
.Y(n_557)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_539),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_501),
.Y(n_541)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_541),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_528),
.B(n_479),
.Y(n_543)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_543),
.B(n_552),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_527),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g565 ( 
.A(n_544),
.B(n_550),
.Y(n_565)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_530),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_509),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_551),
.B(n_526),
.Y(n_556)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_529),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_513),
.B(n_480),
.C(n_490),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_553),
.B(n_555),
.C(n_522),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_516),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_554),
.A2(n_472),
.B1(n_481),
.B2(n_476),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_513),
.B(n_485),
.C(n_482),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_556),
.B(n_559),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_558),
.B(n_553),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_540),
.B(n_535),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_534),
.A2(n_504),
.B1(n_521),
.B2(n_520),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_560),
.A2(n_539),
.B1(n_543),
.B2(n_531),
.Y(n_580)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_562),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_539),
.A2(n_506),
.B1(n_511),
.B2(n_517),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_563),
.B(n_567),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_L g564 ( 
.A1(n_534),
.A2(n_524),
.B(n_518),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_L g579 ( 
.A1(n_564),
.A2(n_555),
.B(n_538),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_535),
.B(n_512),
.C(n_485),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_566),
.B(n_572),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_540),
.B(n_512),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_548),
.B(n_489),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_569),
.B(n_570),
.Y(n_591)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_548),
.B(n_483),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_532),
.B(n_483),
.C(n_496),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_551),
.B(n_433),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_573),
.B(n_537),
.C(n_542),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_532),
.B(n_478),
.C(n_349),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_574),
.B(n_478),
.Y(n_585)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_565),
.Y(n_577)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_577),
.Y(n_594)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_561),
.Y(n_578)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_578),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g597 ( 
.A(n_579),
.B(n_583),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_580),
.A2(n_587),
.B1(n_568),
.B2(n_557),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_581),
.B(n_586),
.Y(n_605)
);

OAI21x1_ASAP7_75t_L g599 ( 
.A1(n_585),
.A2(n_573),
.B(n_569),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_558),
.B(n_536),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_560),
.A2(n_554),
.B1(n_541),
.B2(n_533),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_SL g589 ( 
.A1(n_561),
.A2(n_547),
.B(n_546),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_L g602 ( 
.A1(n_589),
.A2(n_564),
.B(n_563),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_559),
.B(n_545),
.C(n_300),
.Y(n_590)
);

NOR2xp67_ASAP7_75t_SL g598 ( 
.A(n_590),
.B(n_556),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_574),
.B(n_572),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_592),
.B(n_567),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_583),
.B(n_571),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_593),
.B(n_595),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_590),
.B(n_575),
.Y(n_595)
);

NAND2xp33_ASAP7_75t_SL g607 ( 
.A(n_596),
.B(n_602),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g613 ( 
.A(n_598),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_599),
.B(n_601),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_584),
.B(n_566),
.C(n_570),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_603),
.B(n_604),
.Y(n_614)
);

OAI21xp5_ASAP7_75t_SL g604 ( 
.A1(n_582),
.A2(n_354),
.B(n_299),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_576),
.B(n_386),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_SL g610 ( 
.A(n_606),
.B(n_587),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g618 ( 
.A(n_610),
.Y(n_618)
);

XOR2xp5_ASAP7_75t_L g611 ( 
.A(n_597),
.B(n_579),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_611),
.B(n_616),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_597),
.B(n_589),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_612),
.A2(n_615),
.B(n_602),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_605),
.B(n_584),
.Y(n_615)
);

XOR2xp5_ASAP7_75t_L g616 ( 
.A(n_601),
.B(n_591),
.Y(n_616)
);

OAI221xp5_ASAP7_75t_L g623 ( 
.A1(n_617),
.A2(n_619),
.B1(n_621),
.B2(n_613),
.C(n_614),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_609),
.Y(n_619)
);

OAI21xp33_ASAP7_75t_L g621 ( 
.A1(n_608),
.A2(n_593),
.B(n_600),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_L g622 ( 
.A1(n_613),
.A2(n_596),
.B(n_594),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_SL g624 ( 
.A1(n_622),
.A2(n_607),
.B(n_611),
.Y(n_624)
);

AOI21x1_ASAP7_75t_L g628 ( 
.A1(n_623),
.A2(n_625),
.B(n_626),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_624),
.B(n_588),
.C(n_580),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_618),
.A2(n_616),
.B(n_588),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_620),
.B(n_591),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_627),
.B(n_1),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_629),
.B(n_3),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_630),
.A2(n_628),
.B(n_4),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_631),
.B(n_4),
.C(n_295),
.Y(n_632)
);


endmodule