module fake_ibex_222_n_2341 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_446, n_108, n_350, n_165, n_452, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_457, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_176, n_58, n_43, n_216, n_33, n_421, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_453, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_465, n_48, n_325, n_57, n_301, n_434, n_296, n_120, n_168, n_155, n_315, n_441, n_13, n_122, n_116, n_370, n_431, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_22, n_136, n_261, n_459, n_30, n_367, n_221, n_437, n_355, n_407, n_102, n_52, n_448, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_420, n_141, n_222, n_186, n_349, n_454, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_429, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_445, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_416, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_447, n_26, n_188, n_200, n_444, n_199, n_410, n_308, n_463, n_411, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_381, n_382, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_460, n_461, n_313, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_462, n_302, n_450, n_443, n_344, n_393, n_436, n_428, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_399, n_254, n_213, n_424, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_425, n_2341);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_446;
input n_108;
input n_350;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_457;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_453;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_434;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_116;
input n_370;
input n_431;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_22;
input n_136;
input n_261;
input n_459;
input n_30;
input n_367;
input n_221;
input n_437;
input n_355;
input n_407;
input n_102;
input n_52;
input n_448;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_141;
input n_222;
input n_186;
input n_349;
input n_454;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_429;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_416;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_199;
input n_410;
input n_308;
input n_463;
input n_411;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_381;
input n_382;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_460;
input n_461;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_462;
input n_302;
input n_450;
input n_443;
input n_344;
input n_393;
input n_436;
input n_428;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_399;
input n_254;
input n_213;
input n_424;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;
input n_425;

output n_2341;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_2201;
wire n_766;
wire n_2175;
wire n_2071;
wire n_1110;
wire n_1382;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_773;
wire n_2038;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_2183;
wire n_1954;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_2276;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2139;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_2151;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_1971;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_557;
wire n_641;
wire n_1937;
wire n_2311;
wire n_527;
wire n_893;
wire n_1654;
wire n_496;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_2015;
wire n_1130;
wire n_1228;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_538;
wire n_1155;
wire n_1292;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_1926;
wire n_904;
wire n_2003;
wire n_1970;
wire n_1778;
wire n_646;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_1955;
wire n_917;
wire n_2249;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_2090;
wire n_666;
wire n_2260;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1960;
wire n_1723;
wire n_793;
wire n_937;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_2283;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_554;
wire n_553;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_2275;
wire n_2189;
wire n_745;
wire n_2112;
wire n_1753;
wire n_562;
wire n_564;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2171;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_499;
wire n_971;
wire n_702;
wire n_1326;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_579;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_2203;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_1121;
wire n_693;
wire n_2256;
wire n_737;
wire n_606;
wire n_1571;
wire n_1980;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_1543;
wire n_823;
wire n_2233;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_1591;
wire n_583;
wire n_2289;
wire n_2288;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2101;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_1831;
wire n_864;
wire n_608;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_846;
wire n_471;
wire n_1793;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_1498;
wire n_2312;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_469;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_1589;
wire n_2204;
wire n_1210;
wire n_2319;
wire n_591;
wire n_1933;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2006;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2146;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1566;
wire n_1464;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_585;
wire n_2252;
wire n_1982;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_2294;
wire n_1977;
wire n_1200;
wire n_2295;
wire n_1120;
wire n_2300;
wire n_576;
wire n_1602;
wire n_1776;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_827;
wire n_607;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_2287;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_488;
wire n_705;
wire n_2142;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_472;
wire n_1704;
wire n_2160;
wire n_2234;
wire n_847;
wire n_1436;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_801;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1599;
wire n_1539;
wire n_1806;
wire n_650;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_517;
wire n_817;
wire n_2193;
wire n_2095;
wire n_555;
wire n_951;
wire n_2053;
wire n_468;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_502;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_532;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_863;
wire n_597;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_2170;
wire n_1785;
wire n_486;
wire n_1870;
wire n_1405;
wire n_997;
wire n_2308;
wire n_1428;
wire n_2243;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_1925;
wire n_2106;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_890;
wire n_628;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_2298;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2064;
wire n_1679;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1997;
wire n_1894;
wire n_2110;
wire n_961;
wire n_991;
wire n_634;
wire n_1331;
wire n_1223;
wire n_1349;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1694;
wire n_1458;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_1830;
wire n_2261;
wire n_1629;
wire n_2011;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_2317;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_1099;
wire n_598;
wire n_2141;
wire n_1422;
wire n_508;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2210;
wire n_1517;
wire n_690;
wire n_1225;
wire n_1962;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_2087;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_1348;
wire n_838;
wire n_1289;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_2309;
wire n_842;
wire n_2274;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_636;
wire n_1259;
wire n_490;
wire n_2108;
wire n_595;
wire n_1001;
wire n_570;
wire n_2143;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_1538;
wire n_487;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_993;
wire n_851;
wire n_2085;
wire n_1725;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_571;
wire n_648;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_473;
wire n_1241;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_826;
wire n_2154;
wire n_1976;
wire n_2035;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_1270;
wire n_834;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2012;
wire n_722;
wire n_2251;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_480;
wire n_2182;
wire n_1057;
wire n_1473;
wire n_516;
wire n_2125;
wire n_1403;
wire n_2181;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_2315;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_2272;
wire n_535;
wire n_1956;
wire n_681;
wire n_1718;
wire n_2225;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_786;
wire n_505;
wire n_2043;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_1085;
wire n_2222;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_2135;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2232;
wire n_2121;
wire n_1893;
wire n_1570;
wire n_2231;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1961;
wire n_1050;
wire n_2218;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_1632;
wire n_688;
wire n_1547;
wire n_946;
wire n_1542;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_1909;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_1940;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_1767;
wire n_1939;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_478;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2156;
wire n_753;
wire n_2126;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_682;
wire n_2061;
wire n_1373;
wire n_1686;
wire n_2131;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_755;
wire n_2091;
wire n_1029;
wire n_470;
wire n_770;
wire n_1635;
wire n_1572;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_2337;
wire n_854;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_2323;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_569;
wire n_2305;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_2048;
wire n_987;
wire n_750;
wire n_1299;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_2227;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_1692;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_689;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_2291;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2303;
wire n_924;
wire n_2331;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2092;
wire n_566;
wire n_581;
wire n_1365;
wire n_1472;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_548;
wire n_1158;
wire n_1974;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_888;
wire n_1325;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_1468;
wire n_2327;
wire n_913;
wire n_509;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_2321;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_519;
wire n_1843;
wire n_2186;
wire n_2030;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_2100;
wire n_1902;
wire n_683;
wire n_1194;
wire n_1150;
wire n_620;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_2282;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_438),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_92),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_19),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_397),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_338),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_185),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_361),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_374),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_396),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_347),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_157),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_99),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_255),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_181),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_277),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_161),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_401),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_24),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_244),
.Y(n_484)
);

BUFx5_ASAP7_75t_L g485 ( 
.A(n_280),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_461),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_390),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_429),
.Y(n_488)
);

CKINVDCx16_ASAP7_75t_R g489 ( 
.A(n_344),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_307),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_33),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_242),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_161),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_171),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_135),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_416),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_148),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_101),
.B(n_187),
.Y(n_498)
);

CKINVDCx14_ASAP7_75t_R g499 ( 
.A(n_313),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_71),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_103),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_457),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_424),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_54),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_195),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_373),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_311),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_383),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_16),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_325),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_434),
.Y(n_511)
);

CKINVDCx16_ASAP7_75t_R g512 ( 
.A(n_357),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_256),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_448),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_399),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_33),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_439),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_370),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_332),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_352),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_381),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_168),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_393),
.Y(n_523)
);

CKINVDCx16_ASAP7_75t_R g524 ( 
.A(n_58),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_377),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_388),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_85),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_95),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_261),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_142),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_353),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_432),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_456),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_179),
.Y(n_534)
);

BUFx10_ASAP7_75t_L g535 ( 
.A(n_403),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_335),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g537 ( 
.A(n_145),
.Y(n_537)
);

BUFx2_ASAP7_75t_SL g538 ( 
.A(n_200),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_105),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_421),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_459),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_464),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_452),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_108),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_280),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_303),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_413),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_224),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_418),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_228),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_450),
.Y(n_551)
);

BUFx8_ASAP7_75t_SL g552 ( 
.A(n_30),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_193),
.Y(n_553)
);

CKINVDCx16_ASAP7_75t_R g554 ( 
.A(n_398),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_465),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_18),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_230),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_274),
.Y(n_558)
);

INVx1_ASAP7_75t_SL g559 ( 
.A(n_78),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_147),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_440),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_385),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_46),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_164),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_150),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_378),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_38),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_276),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_2),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_247),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_375),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_4),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_50),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_47),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_256),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_408),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_132),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_376),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_71),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_35),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_177),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_326),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_255),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_241),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_216),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_437),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_345),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_94),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_322),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_153),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_400),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_230),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_73),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_305),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_216),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_143),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_8),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_444),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_341),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_212),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_157),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_317),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_386),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_292),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_333),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_50),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_46),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_250),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_205),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_304),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_36),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_190),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_443),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_266),
.Y(n_614)
);

INVxp67_ASAP7_75t_L g615 ( 
.A(n_58),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_61),
.Y(n_616)
);

NOR2xp67_ASAP7_75t_L g617 ( 
.A(n_241),
.B(n_91),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_364),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_312),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_171),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_337),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_262),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_44),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_134),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_236),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_284),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_28),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_233),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_442),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_422),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_53),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_179),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_215),
.B(n_38),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_145),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_296),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_405),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_279),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_342),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_458),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_252),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_371),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_225),
.Y(n_642)
);

INVxp33_ASAP7_75t_SL g643 ( 
.A(n_111),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_17),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_180),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_61),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_244),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_210),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_72),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_360),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_384),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_409),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_346),
.Y(n_653)
);

CKINVDCx16_ASAP7_75t_R g654 ( 
.A(n_414),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_151),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_162),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_175),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_94),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_301),
.Y(n_659)
);

INVx1_ASAP7_75t_SL g660 ( 
.A(n_57),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_290),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_97),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_72),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_234),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_288),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_273),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_324),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_366),
.B(n_42),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_410),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_379),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_53),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_30),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_198),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_404),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_261),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_319),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_133),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_211),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_36),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_126),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_7),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_198),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_169),
.Y(n_683)
);

CKINVDCx20_ASAP7_75t_R g684 ( 
.A(n_372),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_426),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_271),
.Y(n_686)
);

INVxp67_ASAP7_75t_L g687 ( 
.A(n_387),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_78),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_95),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_427),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_251),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_223),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_195),
.Y(n_693)
);

CKINVDCx20_ASAP7_75t_R g694 ( 
.A(n_220),
.Y(n_694)
);

INVxp67_ASAP7_75t_SL g695 ( 
.A(n_327),
.Y(n_695)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_57),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_237),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_389),
.Y(n_698)
);

HB1xp67_ASAP7_75t_L g699 ( 
.A(n_154),
.Y(n_699)
);

BUFx2_ASAP7_75t_L g700 ( 
.A(n_314),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_402),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_447),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_296),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_462),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_79),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_441),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_184),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_228),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_392),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_407),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_218),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_121),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_310),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_235),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_167),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_63),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_11),
.Y(n_717)
);

INVx1_ASAP7_75t_SL g718 ( 
.A(n_330),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_125),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_232),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_246),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_5),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_136),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_436),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_406),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_65),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_207),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_177),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_417),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_391),
.Y(n_730)
);

CKINVDCx16_ASAP7_75t_R g731 ( 
.A(n_158),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_395),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_363),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_15),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_221),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_90),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_215),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_349),
.Y(n_738)
);

BUFx10_ASAP7_75t_L g739 ( 
.A(n_85),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_62),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_11),
.Y(n_741)
);

CKINVDCx20_ASAP7_75t_R g742 ( 
.A(n_253),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_445),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_290),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_170),
.Y(n_745)
);

INVxp67_ASAP7_75t_SL g746 ( 
.A(n_303),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_86),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_144),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_0),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_268),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_321),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_394),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_118),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_187),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_605),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_470),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_485),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_552),
.Y(n_758)
);

BUFx8_ASAP7_75t_L g759 ( 
.A(n_514),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_691),
.B(n_1),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_SL g761 ( 
.A1(n_569),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_525),
.Y(n_762)
);

BUFx8_ASAP7_75t_L g763 ( 
.A(n_700),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_691),
.B(n_3),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_485),
.Y(n_765)
);

AND2x6_ASAP7_75t_L g766 ( 
.A(n_525),
.B(n_306),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_552),
.Y(n_767)
);

BUFx2_ASAP7_75t_L g768 ( 
.A(n_493),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_470),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_640),
.B(n_4),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_643),
.A2(n_489),
.B1(n_512),
.B2(n_496),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_470),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_485),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_485),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_738),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_485),
.Y(n_776)
);

OAI21x1_ASAP7_75t_L g777 ( 
.A1(n_474),
.A2(n_309),
.B(n_308),
.Y(n_777)
);

BUFx8_ASAP7_75t_L g778 ( 
.A(n_542),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_485),
.Y(n_779)
);

OA21x2_ASAP7_75t_L g780 ( 
.A1(n_474),
.A2(n_316),
.B(n_315),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_680),
.B(n_5),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_485),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_515),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_524),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_515),
.Y(n_785)
);

OAI21x1_ASAP7_75t_L g786 ( 
.A1(n_517),
.A2(n_320),
.B(n_318),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_696),
.B(n_6),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_534),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_517),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_629),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_731),
.B(n_9),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_699),
.B(n_735),
.Y(n_792)
);

AND2x6_ASAP7_75t_L g793 ( 
.A(n_533),
.B(n_323),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_470),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_579),
.Y(n_795)
);

AND2x6_ASAP7_75t_L g796 ( 
.A(n_676),
.B(n_328),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_708),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_468),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_739),
.Y(n_799)
);

BUFx2_ASAP7_75t_L g800 ( 
.A(n_708),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_560),
.B(n_10),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_560),
.Y(n_802)
);

OR2x6_ASAP7_75t_L g803 ( 
.A(n_538),
.B(n_10),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_554),
.B(n_12),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_629),
.Y(n_805)
);

OAI22xp33_ASAP7_75t_R g806 ( 
.A1(n_746),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_698),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_654),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_508),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_643),
.A2(n_17),
.B1(n_13),
.B2(n_14),
.Y(n_810)
);

BUFx12f_ASAP7_75t_L g811 ( 
.A(n_535),
.Y(n_811)
);

BUFx8_ASAP7_75t_L g812 ( 
.A(n_562),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_508),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_563),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_698),
.Y(n_815)
);

OA21x2_ASAP7_75t_L g816 ( 
.A1(n_469),
.A2(n_331),
.B(n_329),
.Y(n_816)
);

OAI22x1_ASAP7_75t_SL g817 ( 
.A1(n_569),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_676),
.Y(n_818)
);

BUFx3_ASAP7_75t_L g819 ( 
.A(n_472),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_567),
.B(n_20),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_597),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_473),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_570),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_615),
.B(n_21),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_597),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_468),
.B(n_22),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_491),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_475),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_482),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_508),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_486),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_508),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_490),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_502),
.Y(n_834)
);

BUFx2_ASAP7_75t_L g835 ( 
.A(n_491),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_623),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_566),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_499),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_492),
.B(n_23),
.Y(n_839)
);

CKINVDCx16_ASAP7_75t_R g840 ( 
.A(n_739),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_627),
.Y(n_841)
);

INVx5_ASAP7_75t_L g842 ( 
.A(n_566),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_627),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_692),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_492),
.B(n_25),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_692),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_703),
.B(n_25),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_703),
.B(n_26),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_757),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_760),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_757),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_765),
.Y(n_852)
);

INVxp33_ASAP7_75t_L g853 ( 
.A(n_835),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_760),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_760),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_765),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_764),
.Y(n_857)
);

NAND2xp33_ASAP7_75t_L g858 ( 
.A(n_766),
.B(n_566),
.Y(n_858)
);

BUFx2_ASAP7_75t_L g859 ( 
.A(n_808),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_798),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_764),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_773),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_811),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_840),
.B(n_739),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_792),
.Y(n_865)
);

INVx4_ASAP7_75t_L g866 ( 
.A(n_766),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_764),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_801),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_768),
.B(n_494),
.Y(n_869)
);

INVxp67_ASAP7_75t_SL g870 ( 
.A(n_768),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_811),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_801),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_801),
.Y(n_873)
);

OAI22xp33_ASAP7_75t_L g874 ( 
.A1(n_810),
.A2(n_803),
.B1(n_771),
.B2(n_784),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_808),
.Y(n_875)
);

NAND2xp33_ASAP7_75t_L g876 ( 
.A(n_766),
.B(n_566),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_767),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_773),
.Y(n_878)
);

INVx6_ASAP7_75t_L g879 ( 
.A(n_778),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_774),
.Y(n_880)
);

CKINVDCx14_ASAP7_75t_R g881 ( 
.A(n_838),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_800),
.B(n_494),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_820),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_776),
.B(n_518),
.Y(n_884)
);

BUFx4f_ASAP7_75t_L g885 ( 
.A(n_803),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_820),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_776),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_779),
.Y(n_888)
);

BUFx4f_ASAP7_75t_L g889 ( 
.A(n_803),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_779),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_782),
.B(n_520),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_755),
.B(n_754),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_782),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_822),
.B(n_523),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_756),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_756),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_838),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_847),
.Y(n_898)
);

NAND2xp33_ASAP7_75t_L g899 ( 
.A(n_766),
.B(n_793),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_756),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_800),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_759),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_775),
.B(n_687),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_847),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_848),
.B(n_716),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_822),
.B(n_828),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_759),
.Y(n_907)
);

BUFx10_ASAP7_75t_L g908 ( 
.A(n_848),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_756),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_848),
.Y(n_910)
);

BUFx10_ASAP7_75t_L g911 ( 
.A(n_766),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_772),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_788),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_788),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_828),
.B(n_526),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_788),
.Y(n_916)
);

BUFx10_ASAP7_75t_L g917 ( 
.A(n_766),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_799),
.A2(n_505),
.B1(n_509),
.B2(n_501),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_772),
.Y(n_919)
);

OR2x6_ASAP7_75t_L g920 ( 
.A(n_803),
.B(n_617),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_804),
.Y(n_921)
);

INVx5_ASAP7_75t_L g922 ( 
.A(n_793),
.Y(n_922)
);

BUFx3_ASAP7_75t_L g923 ( 
.A(n_778),
.Y(n_923)
);

BUFx2_ASAP7_75t_L g924 ( 
.A(n_759),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_819),
.B(n_762),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_821),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_829),
.B(n_532),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_772),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_791),
.B(n_535),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_795),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_772),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_797),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_770),
.A2(n_521),
.B1(n_639),
.B2(n_531),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_783),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_829),
.B(n_536),
.Y(n_935)
);

NAND2xp33_ASAP7_75t_SL g936 ( 
.A(n_791),
.B(n_521),
.Y(n_936)
);

OAI22xp33_ASAP7_75t_L g937 ( 
.A1(n_827),
.A2(n_574),
.B1(n_584),
.B2(n_570),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_794),
.Y(n_938)
);

AND2x6_ASAP7_75t_L g939 ( 
.A(n_793),
.B(n_540),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_831),
.B(n_541),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_831),
.B(n_535),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_812),
.Y(n_942)
);

INVx5_ASAP7_75t_L g943 ( 
.A(n_793),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_794),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_821),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_783),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_794),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_794),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_812),
.B(n_833),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_785),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_785),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_821),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_809),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_789),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_790),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_833),
.B(n_522),
.Y(n_956)
);

INVxp33_ASAP7_75t_L g957 ( 
.A(n_826),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_790),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_805),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_812),
.B(n_834),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_763),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_805),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_807),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_763),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_802),
.B(n_543),
.Y(n_965)
);

INVx1_ASAP7_75t_SL g966 ( 
.A(n_823),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_807),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_R g968 ( 
.A(n_763),
.B(n_531),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_813),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_815),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_814),
.B(n_547),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_830),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_781),
.A2(n_684),
.B1(n_690),
.B2(n_639),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_830),
.Y(n_974)
);

OR2x2_ASAP7_75t_L g975 ( 
.A(n_787),
.B(n_754),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_815),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_841),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_818),
.B(n_522),
.Y(n_978)
);

BUFx10_ASAP7_75t_L g979 ( 
.A(n_796),
.Y(n_979)
);

INVxp33_ASAP7_75t_L g980 ( 
.A(n_839),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_818),
.B(n_549),
.Y(n_981)
);

INVx4_ASAP7_75t_L g982 ( 
.A(n_796),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_825),
.Y(n_983)
);

INVx11_ASAP7_75t_L g984 ( 
.A(n_796),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_836),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_SL g986 ( 
.A1(n_761),
.A2(n_742),
.B1(n_584),
.B2(n_622),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_844),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_846),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_841),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_843),
.Y(n_990)
);

AOI22xp33_ASAP7_75t_L g991 ( 
.A1(n_796),
.A2(n_467),
.B1(n_478),
.B2(n_471),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_SL g992 ( 
.A1(n_845),
.A2(n_622),
.B1(n_637),
.B2(n_574),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_843),
.B(n_590),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_843),
.B(n_551),
.Y(n_994)
);

BUFx3_ASAP7_75t_L g995 ( 
.A(n_796),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_823),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_824),
.Y(n_997)
);

INVx2_ASAP7_75t_SL g998 ( 
.A(n_842),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_832),
.Y(n_999)
);

AOI21x1_ASAP7_75t_L g1000 ( 
.A1(n_777),
.A2(n_561),
.B(n_555),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_842),
.B(n_590),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_842),
.B(n_571),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_842),
.B(n_596),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_786),
.Y(n_1004)
);

INVx4_ASAP7_75t_L g1005 ( 
.A(n_796),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_832),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_780),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_842),
.B(n_578),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_780),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_837),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_837),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_837),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_780),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_SL g1014 ( 
.A1(n_885),
.A2(n_681),
.B1(n_683),
.B2(n_637),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_968),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_914),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_913),
.Y(n_1017)
);

OR2x2_ASAP7_75t_L g1018 ( 
.A(n_865),
.B(n_596),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_SL g1019 ( 
.A(n_879),
.B(n_690),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_885),
.A2(n_480),
.B1(n_481),
.B2(n_479),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_997),
.B(n_466),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_SL g1022 ( 
.A(n_879),
.B(n_729),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_956),
.B(n_488),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_941),
.B(n_503),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_860),
.Y(n_1025)
);

AOI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_889),
.A2(n_483),
.B1(n_500),
.B2(n_497),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_908),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_850),
.B(n_503),
.Y(n_1028)
);

AND2x6_ASAP7_75t_SL g1029 ( 
.A(n_920),
.B(n_758),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_854),
.B(n_507),
.Y(n_1030)
);

NAND3xp33_ASAP7_75t_L g1031 ( 
.A(n_991),
.B(n_607),
.C(n_601),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_855),
.B(n_510),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_861),
.B(n_510),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_916),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_867),
.B(n_511),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_873),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_857),
.B(n_511),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_923),
.B(n_519),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_926),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_853),
.B(n_607),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_SL g1041 ( 
.A(n_866),
.B(n_729),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_923),
.B(n_519),
.Y(n_1042)
);

NAND2xp33_ASAP7_75t_SL g1043 ( 
.A(n_964),
.B(n_498),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_857),
.A2(n_513),
.B(n_516),
.C(n_504),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_957),
.B(n_598),
.Y(n_1045)
);

AND2x6_ASAP7_75t_L g1046 ( 
.A(n_995),
.B(n_942),
.Y(n_1046)
);

INVxp67_ASAP7_75t_L g1047 ( 
.A(n_921),
.Y(n_1047)
);

AND2x2_ASAP7_75t_SL g1048 ( 
.A(n_889),
.B(n_758),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_942),
.B(n_610),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_911),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_980),
.B(n_709),
.Y(n_1051)
);

INVx2_ASAP7_75t_SL g1052 ( 
.A(n_863),
.Y(n_1052)
);

INVx2_ASAP7_75t_SL g1053 ( 
.A(n_871),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_873),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_898),
.Y(n_1055)
);

OR2x2_ASAP7_75t_L g1056 ( 
.A(n_892),
.B(n_601),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_945),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_945),
.Y(n_1058)
);

INVx5_ASAP7_75t_L g1059 ( 
.A(n_908),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_949),
.B(n_960),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_870),
.B(n_724),
.Y(n_1061)
);

INVx2_ASAP7_75t_SL g1062 ( 
.A(n_864),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_853),
.B(n_725),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_920),
.A2(n_711),
.B1(n_722),
.B2(n_707),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_869),
.B(n_730),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_911),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_898),
.Y(n_1067)
);

NOR3xp33_ASAP7_75t_L g1068 ( 
.A(n_933),
.B(n_559),
.C(n_537),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_882),
.B(n_743),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_952),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_952),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_901),
.B(n_743),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_905),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_903),
.B(n_752),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_874),
.A2(n_806),
.B1(n_736),
.B2(n_737),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_920),
.A2(n_736),
.B1(n_737),
.B2(n_734),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_977),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_929),
.B(n_487),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_975),
.B(n_506),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_868),
.A2(n_539),
.B(n_545),
.C(n_528),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1007),
.A2(n_816),
.B(n_695),
.Y(n_1081)
);

INVx8_ASAP7_75t_L g1082 ( 
.A(n_939),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_977),
.Y(n_1083)
);

INVx2_ASAP7_75t_SL g1084 ( 
.A(n_993),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_905),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_SL g1086 ( 
.A(n_905),
.Y(n_1086)
);

NOR2x1p5_ASAP7_75t_L g1087 ( 
.A(n_902),
.B(n_745),
.Y(n_1087)
);

INVx2_ASAP7_75t_SL g1088 ( 
.A(n_908),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_978),
.B(n_576),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_872),
.B(n_582),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_907),
.B(n_476),
.Y(n_1091)
);

BUFx8_ASAP7_75t_L g1092 ( 
.A(n_924),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_883),
.B(n_586),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_989),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_961),
.Y(n_1095)
);

INVxp33_ASAP7_75t_L g1096 ( 
.A(n_973),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_859),
.B(n_477),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_886),
.B(n_613),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_990),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_904),
.A2(n_548),
.B1(n_550),
.B2(n_546),
.Y(n_1100)
);

INVxp67_ASAP7_75t_L g1101 ( 
.A(n_875),
.Y(n_1101)
);

AND2x6_ASAP7_75t_L g1102 ( 
.A(n_984),
.B(n_587),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_910),
.A2(n_564),
.B1(n_568),
.B2(n_553),
.Y(n_1103)
);

BUFx5_ASAP7_75t_L g1104 ( 
.A(n_917),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_881),
.B(n_918),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_925),
.B(n_621),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_917),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_881),
.B(n_897),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_983),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_982),
.B(n_630),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_930),
.B(n_589),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_874),
.A2(n_484),
.B1(n_529),
.B2(n_527),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_985),
.Y(n_1113)
);

AOI221xp5_ASAP7_75t_L g1114 ( 
.A1(n_937),
.A2(n_817),
.B1(n_575),
.B2(n_577),
.C(n_573),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_987),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_1005),
.B(n_651),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_988),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_932),
.B(n_927),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_897),
.B(n_718),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_934),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_965),
.A2(n_581),
.B(n_592),
.C(n_572),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_922),
.B(n_667),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_992),
.B(n_530),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_877),
.B(n_994),
.Y(n_1124)
);

INVx2_ASAP7_75t_SL g1125 ( 
.A(n_1001),
.Y(n_1125)
);

AO221x1_ASAP7_75t_L g1126 ( 
.A1(n_937),
.A2(n_694),
.B1(n_719),
.B2(n_686),
.C(n_683),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1003),
.B(n_670),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_946),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1009),
.A2(n_594),
.B(n_591),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_950),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_922),
.B(n_593),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_877),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_971),
.A2(n_600),
.B(n_604),
.C(n_595),
.Y(n_1133)
);

AOI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_936),
.A2(n_556),
.B1(n_557),
.B2(n_544),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_951),
.Y(n_1135)
);

INVxp67_ASAP7_75t_L g1136 ( 
.A(n_936),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_954),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_955),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_894),
.B(n_701),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_915),
.B(n_706),
.Y(n_1140)
);

INVxp67_ASAP7_75t_SL g1141 ( 
.A(n_849),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_996),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_915),
.B(n_558),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_935),
.B(n_565),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_958),
.Y(n_1145)
);

INVx4_ASAP7_75t_L g1146 ( 
.A(n_922),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_940),
.B(n_580),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_966),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_959),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_962),
.B(n_583),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_963),
.B(n_585),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_943),
.B(n_599),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_967),
.B(n_588),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_939),
.B(n_602),
.Y(n_1154)
);

AOI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_991),
.A2(n_611),
.B1(n_624),
.B2(n_614),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_851),
.B(n_603),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_852),
.B(n_618),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_852),
.B(n_619),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_970),
.Y(n_1159)
);

AOI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_858),
.A2(n_625),
.B1(n_632),
.B2(n_631),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_856),
.B(n_636),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_976),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_856),
.B(n_638),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_943),
.B(n_641),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_906),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1004),
.A2(n_606),
.B(n_609),
.C(n_608),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_943),
.A2(n_646),
.B1(n_648),
.B2(n_642),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_986),
.B(n_649),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_862),
.B(n_650),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_878),
.B(n_652),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_878),
.Y(n_1171)
);

INVx2_ASAP7_75t_SL g1172 ( 
.A(n_981),
.Y(n_1172)
);

BUFx3_ASAP7_75t_L g1173 ( 
.A(n_880),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_943),
.B(n_669),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_880),
.B(n_674),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_906),
.B(n_655),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_887),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_888),
.B(n_685),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_979),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_884),
.B(n_702),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_888),
.B(n_710),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_890),
.B(n_713),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_890),
.B(n_656),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_891),
.A2(n_612),
.B(n_620),
.C(n_616),
.Y(n_1184)
);

AOI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_858),
.A2(n_662),
.B1(n_663),
.B2(n_657),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_893),
.B(n_732),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_893),
.B(n_733),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1002),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_876),
.B(n_666),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1002),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_SL g1191 ( 
.A(n_1008),
.B(n_686),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1013),
.B(n_751),
.Y(n_1192)
);

AND2x2_ASAP7_75t_SL g1193 ( 
.A(n_876),
.B(n_716),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1008),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1000),
.B(n_717),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_998),
.B(n_717),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_896),
.B(n_744),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_900),
.B(n_744),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_895),
.B(n_675),
.Y(n_1199)
);

OAI21xp33_ASAP7_75t_L g1200 ( 
.A1(n_909),
.A2(n_628),
.B(n_626),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_912),
.B(n_634),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_895),
.B(n_679),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_912),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_919),
.B(n_635),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_972),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_919),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_928),
.B(n_644),
.Y(n_1207)
);

OAI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_928),
.A2(n_719),
.B1(n_723),
.B2(n_694),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_931),
.A2(n_668),
.B(n_769),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_931),
.B(n_645),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_938),
.B(n_689),
.Y(n_1211)
);

BUFx5_ASAP7_75t_L g1212 ( 
.A(n_1006),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_938),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_944),
.B(n_647),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_944),
.A2(n_661),
.B1(n_664),
.B2(n_659),
.Y(n_1215)
);

INVx4_ASAP7_75t_L g1216 ( 
.A(n_1010),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_947),
.B(n_665),
.Y(n_1217)
);

NOR3xp33_ASAP7_75t_L g1218 ( 
.A(n_1025),
.B(n_1114),
.C(n_1208),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1040),
.B(n_723),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1192),
.A2(n_953),
.B(n_948),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1021),
.B(n_671),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1173),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1101),
.Y(n_1223)
);

INVx8_ASAP7_75t_L g1224 ( 
.A(n_1059),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1021),
.B(n_672),
.Y(n_1225)
);

O2A1O1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1121),
.A2(n_1133),
.B(n_1166),
.C(n_1080),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1129),
.A2(n_677),
.B(n_678),
.C(n_673),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1162),
.B(n_682),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_1148),
.Y(n_1229)
);

O2A1O1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1044),
.A2(n_693),
.B(n_697),
.C(n_688),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1092),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1018),
.B(n_742),
.Y(n_1232)
);

NAND2x1p5_ASAP7_75t_L g1233 ( 
.A(n_1059),
.B(n_705),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1183),
.B(n_712),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_1092),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1084),
.B(n_720),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1096),
.A2(n_721),
.B1(n_727),
.B2(n_726),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1036),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1054),
.Y(n_1239)
);

O2A1O1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1047),
.A2(n_740),
.B(n_741),
.C(n_728),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1055),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1067),
.Y(n_1242)
);

NAND3xp33_ASAP7_75t_L g1243 ( 
.A(n_1068),
.B(n_1063),
.C(n_1072),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1062),
.B(n_660),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1045),
.B(n_747),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1195),
.A2(n_974),
.B(n_969),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1051),
.B(n_748),
.Y(n_1247)
);

BUFx4f_ASAP7_75t_L g1248 ( 
.A(n_1048),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1060),
.A2(n_974),
.B(n_969),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1023),
.B(n_749),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1023),
.B(n_1024),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1136),
.B(n_750),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1097),
.B(n_753),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1024),
.B(n_633),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1056),
.B(n_495),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1029),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1031),
.A2(n_714),
.B1(n_715),
.B2(n_658),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1041),
.A2(n_714),
.B1(n_715),
.B2(n_658),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1120),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1149),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1028),
.A2(n_1011),
.B(n_999),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1028),
.A2(n_1032),
.B(n_1030),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1108),
.B(n_715),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1124),
.B(n_27),
.Y(n_1264)
);

AO21x1_ASAP7_75t_L g1265 ( 
.A1(n_1209),
.A2(n_1012),
.B(n_769),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1073),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1030),
.A2(n_1010),
.B(n_769),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1032),
.A2(n_1035),
.B(n_1033),
.Y(n_1268)
);

BUFx12f_ASAP7_75t_L g1269 ( 
.A(n_1142),
.Y(n_1269)
);

INVx3_ASAP7_75t_SL g1270 ( 
.A(n_1132),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1033),
.A2(n_1010),
.B(n_769),
.Y(n_1271)
);

OR2x6_ASAP7_75t_SL g1272 ( 
.A(n_1064),
.B(n_29),
.Y(n_1272)
);

A2O1A1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1184),
.A2(n_704),
.B(n_653),
.C(n_32),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1035),
.A2(n_704),
.B(n_653),
.Y(n_1274)
);

INVx3_ASAP7_75t_SL g1275 ( 
.A(n_1015),
.Y(n_1275)
);

INVx3_ASAP7_75t_L g1276 ( 
.A(n_1027),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1141),
.A2(n_35),
.B1(n_31),
.B2(n_34),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_1027),
.B(n_1088),
.Y(n_1278)
);

O2A1O1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1085),
.A2(n_40),
.B(n_37),
.C(n_39),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1037),
.A2(n_336),
.B(n_334),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1037),
.A2(n_340),
.B(n_339),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1154),
.A2(n_348),
.B(n_343),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1079),
.B(n_37),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1118),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1196),
.Y(n_1285)
);

O2A1O1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1076),
.A2(n_47),
.B(n_43),
.C(n_45),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1109),
.B(n_45),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1113),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1115),
.B(n_48),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_1095),
.Y(n_1290)
);

A2O1A1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_1188),
.A2(n_52),
.B(n_49),
.C(n_51),
.Y(n_1291)
);

INVx3_ASAP7_75t_L g1292 ( 
.A(n_1046),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1117),
.B(n_55),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1061),
.B(n_56),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1065),
.B(n_59),
.Y(n_1295)
);

OA22x2_ASAP7_75t_L g1296 ( 
.A1(n_1126),
.A2(n_62),
.B1(n_59),
.B2(n_60),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1091),
.B(n_60),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1043),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1069),
.B(n_64),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1052),
.B(n_64),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1100),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1017),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1190),
.A2(n_1194),
.B(n_1165),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_1019),
.Y(n_1304)
);

AO21x2_ASAP7_75t_L g1305 ( 
.A1(n_1156),
.A2(n_351),
.B(n_350),
.Y(n_1305)
);

A2O1A1Ixp33_ASAP7_75t_L g1306 ( 
.A1(n_1130),
.A2(n_69),
.B(n_67),
.C(n_68),
.Y(n_1306)
);

CKINVDCx20_ASAP7_75t_R g1307 ( 
.A(n_1053),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1123),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1105),
.B(n_69),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1034),
.Y(n_1310)
);

CKINVDCx10_ASAP7_75t_R g1311 ( 
.A(n_1086),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1103),
.A2(n_74),
.B1(n_70),
.B2(n_73),
.Y(n_1312)
);

OA22x2_ASAP7_75t_L g1313 ( 
.A1(n_1075),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1074),
.B(n_75),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1128),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1086),
.A2(n_1191),
.B1(n_1112),
.B2(n_1026),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1020),
.A2(n_79),
.B1(n_76),
.B2(n_77),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1094),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1150),
.A2(n_463),
.B(n_355),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1137),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1138),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_SL g1322 ( 
.A(n_1125),
.B(n_80),
.Y(n_1322)
);

AOI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1134),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1145),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1168),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_1325)
);

O2A1O1Ixp33_ASAP7_75t_L g1326 ( 
.A1(n_1111),
.A2(n_86),
.B(n_83),
.C(n_84),
.Y(n_1326)
);

NOR2x1_ASAP7_75t_R g1327 ( 
.A(n_1014),
.B(n_84),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1151),
.A2(n_356),
.B(n_354),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1153),
.B(n_87),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1119),
.B(n_1087),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_1046),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1078),
.B(n_88),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1135),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1099),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1090),
.A2(n_460),
.B(n_358),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1211),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1093),
.A2(n_362),
.B(n_359),
.Y(n_1337)
);

INVx4_ASAP7_75t_L g1338 ( 
.A(n_1046),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1155),
.B(n_89),
.Y(n_1339)
);

INVx2_ASAP7_75t_SL g1340 ( 
.A(n_1038),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_SL g1341 ( 
.A(n_1160),
.B(n_90),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1159),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_R g1343 ( 
.A(n_1193),
.B(n_93),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_1185),
.B(n_96),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1098),
.A2(n_367),
.B(n_365),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1172),
.A2(n_100),
.B1(n_97),
.B2(n_98),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1042),
.B(n_100),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1049),
.B(n_101),
.Y(n_1348)
);

A2O1A1Ixp33_ASAP7_75t_L g1349 ( 
.A1(n_1156),
.A2(n_105),
.B(n_102),
.C(n_104),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1176),
.A2(n_107),
.B1(n_104),
.B2(n_106),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1171),
.A2(n_369),
.B(n_368),
.Y(n_1351)
);

NAND2x1p5_ASAP7_75t_L g1352 ( 
.A(n_1131),
.B(n_107),
.Y(n_1352)
);

NAND2x1p5_ASAP7_75t_L g1353 ( 
.A(n_1131),
.B(n_108),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1143),
.B(n_1144),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1177),
.A2(n_382),
.B(n_380),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1111),
.B(n_109),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1046),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1039),
.B(n_110),
.Y(n_1358)
);

OAI22x1_ASAP7_75t_L g1359 ( 
.A1(n_1189),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1157),
.A2(n_1161),
.B(n_1158),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1147),
.B(n_114),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1089),
.B(n_115),
.Y(n_1362)
);

INVx2_ASAP7_75t_SL g1363 ( 
.A(n_1057),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_R g1364 ( 
.A(n_1102),
.B(n_116),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1158),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1161),
.A2(n_120),
.B1(n_117),
.B2(n_119),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1167),
.B(n_122),
.Y(n_1367)
);

CKINVDCx10_ASAP7_75t_R g1368 ( 
.A(n_1215),
.Y(n_1368)
);

AOI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1102),
.A2(n_1016),
.B1(n_1180),
.B2(n_1187),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1102),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1102),
.A2(n_126),
.B1(n_123),
.B2(n_124),
.Y(n_1371)
);

INVx3_ASAP7_75t_L g1372 ( 
.A(n_1146),
.Y(n_1372)
);

BUFx4f_ASAP7_75t_L g1373 ( 
.A(n_1102),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1163),
.B(n_127),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1200),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_1375)
);

A2O1A1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1163),
.A2(n_130),
.B(n_128),
.C(n_129),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1201),
.Y(n_1377)
);

OAI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1169),
.A2(n_1175),
.B(n_1170),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_SL g1379 ( 
.A1(n_1058),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1169),
.B(n_1170),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_1082),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1070),
.A2(n_134),
.B1(n_131),
.B2(n_133),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1175),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_SL g1384 ( 
.A(n_1082),
.B(n_137),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1204),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1178),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1071),
.B(n_139),
.Y(n_1387)
);

INVx3_ASAP7_75t_L g1388 ( 
.A(n_1146),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1077),
.B(n_140),
.Y(n_1389)
);

A2O1A1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1178),
.A2(n_141),
.B(n_142),
.C(n_143),
.Y(n_1390)
);

OAI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1181),
.A2(n_412),
.B(n_411),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1181),
.A2(n_141),
.B1(n_144),
.B2(n_146),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1083),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1182),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1182),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1186),
.B(n_149),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1110),
.A2(n_419),
.B(n_415),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1106),
.Y(n_1398)
);

AOI21xp33_ASAP7_75t_L g1399 ( 
.A1(n_1139),
.A2(n_151),
.B(n_152),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1116),
.A2(n_455),
.B(n_423),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1152),
.A2(n_454),
.B(n_425),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1207),
.B(n_154),
.Y(n_1402)
);

O2A1O1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1210),
.A2(n_155),
.B(n_156),
.C(n_158),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1140),
.B(n_155),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1197),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1164),
.A2(n_428),
.B(n_420),
.Y(n_1406)
);

NAND3xp33_ASAP7_75t_SL g1407 ( 
.A(n_1127),
.B(n_156),
.C(n_159),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1199),
.B(n_159),
.Y(n_1408)
);

INVxp67_ASAP7_75t_L g1409 ( 
.A(n_1202),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1174),
.A2(n_431),
.B(n_430),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1122),
.B(n_160),
.Y(n_1411)
);

OAI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1210),
.A2(n_435),
.B(n_433),
.Y(n_1412)
);

INVx1_ASAP7_75t_SL g1413 ( 
.A(n_1214),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_SL g1414 ( 
.A(n_1082),
.B(n_163),
.Y(n_1414)
);

O2A1O1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1214),
.A2(n_164),
.B(n_165),
.C(n_166),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_1050),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1217),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_1417)
);

NOR2xp67_ASAP7_75t_L g1418 ( 
.A(n_1197),
.B(n_168),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_SL g1419 ( 
.A1(n_1104),
.A2(n_169),
.B1(n_170),
.B2(n_172),
.Y(n_1419)
);

INVx1_ASAP7_75t_SL g1420 ( 
.A(n_1198),
.Y(n_1420)
);

AOI21xp33_ASAP7_75t_L g1421 ( 
.A1(n_1205),
.A2(n_173),
.B(n_174),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1198),
.Y(n_1422)
);

OAI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1203),
.A2(n_453),
.B(n_451),
.Y(n_1423)
);

AOI221xp5_ASAP7_75t_L g1424 ( 
.A1(n_1206),
.A2(n_175),
.B1(n_176),
.B2(n_178),
.C(n_180),
.Y(n_1424)
);

AOI21xp33_ASAP7_75t_L g1425 ( 
.A1(n_1066),
.A2(n_181),
.B(n_182),
.Y(n_1425)
);

INVx4_ASAP7_75t_L g1426 ( 
.A(n_1107),
.Y(n_1426)
);

OAI21xp33_ASAP7_75t_L g1427 ( 
.A1(n_1213),
.A2(n_182),
.B(n_183),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1216),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1107),
.A2(n_185),
.B1(n_186),
.B2(n_188),
.Y(n_1429)
);

A2O1A1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1107),
.A2(n_186),
.B(n_188),
.C(n_189),
.Y(n_1430)
);

CKINVDCx20_ASAP7_75t_R g1431 ( 
.A(n_1179),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_1179),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1179),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1104),
.B(n_191),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1104),
.A2(n_1212),
.B(n_449),
.Y(n_1435)
);

INVx4_ASAP7_75t_L g1436 ( 
.A(n_1212),
.Y(n_1436)
);

AOI33xp33_ASAP7_75t_L g1437 ( 
.A1(n_1212),
.A2(n_192),
.A3(n_193),
.B1(n_194),
.B2(n_196),
.B3(n_197),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1096),
.A2(n_192),
.B1(n_194),
.B2(n_196),
.Y(n_1438)
);

NOR2x1p5_ASAP7_75t_SL g1439 ( 
.A(n_1212),
.B(n_446),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1162),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1025),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_SL g1442 ( 
.A(n_1059),
.B(n_199),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_SL g1443 ( 
.A(n_1290),
.B(n_199),
.Y(n_1443)
);

NAND2xp33_ASAP7_75t_L g1444 ( 
.A(n_1331),
.B(n_201),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1394),
.B(n_202),
.Y(n_1445)
);

OA21x2_ASAP7_75t_L g1446 ( 
.A1(n_1246),
.A2(n_203),
.B(n_204),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1302),
.Y(n_1447)
);

NOR2xp67_ASAP7_75t_L g1448 ( 
.A(n_1441),
.B(n_203),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1219),
.B(n_206),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1380),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1262),
.B(n_1268),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1360),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_1452)
);

NAND3xp33_ASAP7_75t_SL g1453 ( 
.A(n_1304),
.B(n_212),
.C(n_213),
.Y(n_1453)
);

AO31x2_ASAP7_75t_L g1454 ( 
.A1(n_1265),
.A2(n_214),
.A3(n_217),
.B(n_218),
.Y(n_1454)
);

INVx4_ASAP7_75t_L g1455 ( 
.A(n_1224),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1310),
.Y(n_1456)
);

BUFx10_ASAP7_75t_L g1457 ( 
.A(n_1358),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1285),
.B(n_219),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1223),
.B(n_220),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_SL g1460 ( 
.A(n_1229),
.B(n_221),
.Y(n_1460)
);

INVxp67_ASAP7_75t_L g1461 ( 
.A(n_1327),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1318),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_SL g1463 ( 
.A1(n_1338),
.A2(n_222),
.B(n_225),
.Y(n_1463)
);

AOI221xp5_ASAP7_75t_L g1464 ( 
.A1(n_1237),
.A2(n_226),
.B1(n_227),
.B2(n_229),
.C(n_231),
.Y(n_1464)
);

BUFx12f_ASAP7_75t_L g1465 ( 
.A(n_1235),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1320),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1218),
.B(n_227),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1232),
.B(n_229),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1378),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_1469)
);

OAI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1248),
.A2(n_1384),
.B1(n_1414),
.B2(n_1316),
.Y(n_1470)
);

INVx2_ASAP7_75t_SL g1471 ( 
.A(n_1231),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1251),
.B(n_238),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_L g1473 ( 
.A(n_1224),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1413),
.B(n_239),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1321),
.Y(n_1475)
);

AO32x2_ASAP7_75t_L g1476 ( 
.A1(n_1277),
.A2(n_240),
.A3(n_242),
.B1(n_243),
.B2(n_245),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1440),
.B(n_246),
.Y(n_1477)
);

AOI221xp5_ASAP7_75t_SL g1478 ( 
.A1(n_1227),
.A2(n_248),
.B1(n_249),
.B2(n_251),
.C(n_252),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1336),
.B(n_248),
.Y(n_1479)
);

NAND3xp33_ASAP7_75t_L g1480 ( 
.A(n_1243),
.B(n_253),
.C(n_254),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1324),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1398),
.B(n_254),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1261),
.A2(n_257),
.B(n_258),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1377),
.B(n_257),
.Y(n_1484)
);

OAI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1267),
.A2(n_258),
.B(n_259),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1308),
.B(n_259),
.Y(n_1486)
);

AO31x2_ASAP7_75t_L g1487 ( 
.A1(n_1273),
.A2(n_260),
.A3(n_263),
.B(n_264),
.Y(n_1487)
);

A2O1A1Ixp33_ASAP7_75t_L g1488 ( 
.A1(n_1362),
.A2(n_265),
.B(n_267),
.C(n_269),
.Y(n_1488)
);

AO31x2_ASAP7_75t_L g1489 ( 
.A1(n_1280),
.A2(n_270),
.A3(n_271),
.B(n_272),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1311),
.Y(n_1490)
);

INVxp67_ASAP7_75t_SL g1491 ( 
.A(n_1431),
.Y(n_1491)
);

AOI22x1_ASAP7_75t_L g1492 ( 
.A1(n_1271),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1253),
.B(n_275),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1385),
.B(n_277),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1270),
.B(n_278),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1330),
.B(n_278),
.Y(n_1496)
);

INVx5_ASAP7_75t_L g1497 ( 
.A(n_1331),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1288),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1334),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_SL g1500 ( 
.A(n_1233),
.B(n_1248),
.Y(n_1500)
);

A2O1A1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1264),
.A2(n_281),
.B(n_282),
.C(n_283),
.Y(n_1501)
);

CKINVDCx11_ASAP7_75t_R g1502 ( 
.A(n_1275),
.Y(n_1502)
);

OAI22x1_ASAP7_75t_L g1503 ( 
.A1(n_1352),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1342),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_R g1505 ( 
.A(n_1307),
.B(n_289),
.Y(n_1505)
);

OA21x2_ASAP7_75t_L g1506 ( 
.A1(n_1391),
.A2(n_1412),
.B(n_1423),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_1269),
.Y(n_1507)
);

INVx4_ASAP7_75t_L g1508 ( 
.A(n_1381),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1228),
.B(n_291),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1315),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1420),
.B(n_293),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1272),
.B(n_294),
.Y(n_1512)
);

AO32x2_ASAP7_75t_L g1513 ( 
.A1(n_1365),
.A2(n_295),
.A3(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1220),
.A2(n_300),
.B(n_302),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1220),
.A2(n_302),
.B(n_1249),
.Y(n_1515)
);

AO32x2_ASAP7_75t_L g1516 ( 
.A1(n_1366),
.A2(n_1392),
.A3(n_1386),
.B1(n_1383),
.B2(n_1395),
.Y(n_1516)
);

BUFx2_ASAP7_75t_L g1517 ( 
.A(n_1364),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1221),
.B(n_1225),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1298),
.B(n_1244),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_SL g1520 ( 
.A(n_1373),
.B(n_1357),
.Y(n_1520)
);

CKINVDCx8_ASAP7_75t_R g1521 ( 
.A(n_1368),
.Y(n_1521)
);

OAI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1405),
.A2(n_1337),
.B(n_1335),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1333),
.Y(n_1523)
);

INVx1_ASAP7_75t_SL g1524 ( 
.A(n_1422),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1352),
.Y(n_1525)
);

CKINVDCx16_ASAP7_75t_R g1526 ( 
.A(n_1343),
.Y(n_1526)
);

INVx5_ASAP7_75t_L g1527 ( 
.A(n_1416),
.Y(n_1527)
);

BUFx4_ASAP7_75t_R g1528 ( 
.A(n_1222),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_1256),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1340),
.B(n_1236),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1287),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1358),
.A2(n_1389),
.B1(n_1353),
.B2(n_1402),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1389),
.Y(n_1533)
);

NAND3x1_ASAP7_75t_L g1534 ( 
.A(n_1309),
.B(n_1323),
.C(n_1437),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1339),
.B(n_1297),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1245),
.A2(n_1247),
.B(n_1250),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1266),
.B(n_1254),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1367),
.A2(n_1344),
.B1(n_1341),
.B2(n_1347),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1238),
.B(n_1239),
.Y(n_1539)
);

INVx2_ASAP7_75t_SL g1540 ( 
.A(n_1353),
.Y(n_1540)
);

INVxp67_ASAP7_75t_SL g1541 ( 
.A(n_1381),
.Y(n_1541)
);

AOI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1348),
.A2(n_1300),
.B1(n_1404),
.B2(n_1411),
.Y(n_1542)
);

A2O1A1Ixp33_ASAP7_75t_L g1543 ( 
.A1(n_1356),
.A2(n_1230),
.B(n_1295),
.C(n_1299),
.Y(n_1543)
);

AND2x2_ASAP7_75t_SL g1544 ( 
.A(n_1411),
.B(n_1370),
.Y(n_1544)
);

NAND3xp33_ASAP7_75t_L g1545 ( 
.A(n_1258),
.B(n_1257),
.C(n_1255),
.Y(n_1545)
);

OAI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1345),
.A2(n_1328),
.B(n_1319),
.Y(n_1546)
);

CKINVDCx14_ASAP7_75t_R g1547 ( 
.A(n_1379),
.Y(n_1547)
);

NOR2x1_ASAP7_75t_SL g1548 ( 
.A(n_1416),
.B(n_1432),
.Y(n_1548)
);

AO21x2_ASAP7_75t_L g1549 ( 
.A1(n_1351),
.A2(n_1355),
.B(n_1305),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1241),
.B(n_1242),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1289),
.Y(n_1551)
);

INVx3_ASAP7_75t_SL g1552 ( 
.A(n_1263),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1374),
.A2(n_1396),
.B1(n_1293),
.B2(n_1350),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1234),
.B(n_1252),
.Y(n_1554)
);

AO32x2_ASAP7_75t_L g1555 ( 
.A1(n_1284),
.A2(n_1317),
.A3(n_1417),
.B1(n_1312),
.B2(n_1301),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1276),
.B(n_1278),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1363),
.B(n_1292),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1332),
.B(n_1314),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1240),
.B(n_1409),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1294),
.B(n_1259),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1260),
.B(n_1361),
.Y(n_1561)
);

OAI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1282),
.A2(n_1397),
.B(n_1400),
.Y(n_1562)
);

AO31x2_ASAP7_75t_L g1563 ( 
.A1(n_1282),
.A2(n_1291),
.A3(n_1349),
.B(n_1390),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1322),
.B(n_1329),
.Y(n_1564)
);

NOR3xp33_ASAP7_75t_L g1565 ( 
.A(n_1407),
.B(n_1286),
.C(n_1279),
.Y(n_1565)
);

NAND2x1p5_ASAP7_75t_L g1566 ( 
.A(n_1426),
.B(n_1432),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1387),
.B(n_1393),
.Y(n_1567)
);

INVx5_ASAP7_75t_L g1568 ( 
.A(n_1432),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_SL g1569 ( 
.A(n_1436),
.B(n_1434),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_1433),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1313),
.Y(n_1571)
);

AO31x2_ASAP7_75t_L g1572 ( 
.A1(n_1376),
.A2(n_1401),
.A3(n_1410),
.B(n_1406),
.Y(n_1572)
);

AOI221x1_ASAP7_75t_L g1573 ( 
.A1(n_1427),
.A2(n_1359),
.B1(n_1421),
.B2(n_1430),
.C(n_1399),
.Y(n_1573)
);

CKINVDCx6p67_ASAP7_75t_R g1574 ( 
.A(n_1442),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1369),
.B(n_1428),
.Y(n_1575)
);

CKINVDCx16_ASAP7_75t_R g1576 ( 
.A(n_1346),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1372),
.Y(n_1577)
);

OAI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1438),
.A2(n_1325),
.B1(n_1371),
.B2(n_1313),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1296),
.Y(n_1579)
);

CKINVDCx11_ASAP7_75t_R g1580 ( 
.A(n_1429),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1296),
.Y(n_1581)
);

BUFx10_ASAP7_75t_L g1582 ( 
.A(n_1419),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1408),
.B(n_1424),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1388),
.B(n_1418),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1306),
.B(n_1382),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1305),
.A2(n_1403),
.B(n_1415),
.Y(n_1586)
);

AO31x2_ASAP7_75t_L g1587 ( 
.A1(n_1439),
.A2(n_1326),
.A3(n_1375),
.B(n_1425),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1290),
.B(n_1336),
.Y(n_1588)
);

NOR2xp67_ASAP7_75t_L g1589 ( 
.A(n_1441),
.B(n_964),
.Y(n_1589)
);

INVx2_ASAP7_75t_SL g1590 ( 
.A(n_1231),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1394),
.B(n_1262),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_1441),
.Y(n_1592)
);

AOI21x1_ASAP7_75t_L g1593 ( 
.A1(n_1435),
.A2(n_1081),
.B(n_1000),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1288),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1290),
.B(n_1025),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1441),
.Y(n_1596)
);

A2O1A1Ixp33_ASAP7_75t_L g1597 ( 
.A1(n_1262),
.A2(n_1268),
.B(n_1354),
.C(n_1226),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1441),
.B(n_865),
.Y(n_1598)
);

AOI21x1_ASAP7_75t_L g1599 ( 
.A1(n_1435),
.A2(n_1081),
.B(n_1000),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1441),
.B(n_865),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1441),
.Y(n_1601)
);

AO31x2_ASAP7_75t_L g1602 ( 
.A1(n_1265),
.A2(n_1274),
.A3(n_1081),
.B(n_1195),
.Y(n_1602)
);

INVx2_ASAP7_75t_SL g1603 ( 
.A(n_1231),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1394),
.B(n_1262),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1302),
.Y(n_1605)
);

AND3x4_ASAP7_75t_L g1606 ( 
.A(n_1231),
.B(n_1218),
.C(n_1068),
.Y(n_1606)
);

OAI21x1_ASAP7_75t_SL g1607 ( 
.A1(n_1262),
.A2(n_1268),
.B(n_1338),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1262),
.A2(n_1268),
.B(n_1303),
.Y(n_1608)
);

AOI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1262),
.A2(n_899),
.B(n_1268),
.Y(n_1609)
);

AOI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1262),
.A2(n_899),
.B(n_1268),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1288),
.Y(n_1611)
);

BUFx2_ASAP7_75t_R g1612 ( 
.A(n_1231),
.Y(n_1612)
);

AOI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1262),
.A2(n_1268),
.B(n_899),
.Y(n_1613)
);

INVx4_ASAP7_75t_L g1614 ( 
.A(n_1224),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1232),
.B(n_1025),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1441),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1394),
.B(n_1262),
.Y(n_1617)
);

BUFx2_ASAP7_75t_L g1618 ( 
.A(n_1441),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1394),
.B(n_1262),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1394),
.B(n_1262),
.Y(n_1620)
);

OAI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1262),
.A2(n_1268),
.B(n_1303),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1302),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_1311),
.Y(n_1623)
);

AOI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1262),
.A2(n_899),
.B(n_1268),
.Y(n_1624)
);

AO21x2_ASAP7_75t_L g1625 ( 
.A1(n_1274),
.A2(n_1081),
.B(n_1265),
.Y(n_1625)
);

AOI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1232),
.A2(n_1025),
.B1(n_973),
.B2(n_933),
.Y(n_1626)
);

A2O1A1Ixp33_ASAP7_75t_L g1627 ( 
.A1(n_1262),
.A2(n_1268),
.B(n_1354),
.C(n_1226),
.Y(n_1627)
);

INVx1_ASAP7_75t_SL g1628 ( 
.A(n_1441),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1288),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1394),
.B(n_1262),
.Y(n_1630)
);

BUFx6f_ASAP7_75t_L g1631 ( 
.A(n_1224),
.Y(n_1631)
);

NOR2x1_ASAP7_75t_L g1632 ( 
.A(n_1231),
.B(n_1025),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_SL g1633 ( 
.A(n_1290),
.B(n_1025),
.Y(n_1633)
);

AOI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1262),
.A2(n_1268),
.B(n_899),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1394),
.B(n_1262),
.Y(n_1635)
);

INVxp67_ASAP7_75t_SL g1636 ( 
.A(n_1441),
.Y(n_1636)
);

BUFx2_ASAP7_75t_SL g1637 ( 
.A(n_1231),
.Y(n_1637)
);

INVxp67_ASAP7_75t_SL g1638 ( 
.A(n_1441),
.Y(n_1638)
);

AO21x1_ASAP7_75t_L g1639 ( 
.A1(n_1280),
.A2(n_1281),
.B(n_1274),
.Y(n_1639)
);

INVx3_ASAP7_75t_SL g1640 ( 
.A(n_1231),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1441),
.B(n_865),
.Y(n_1641)
);

AOI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1262),
.A2(n_899),
.B(n_1268),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1311),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1394),
.B(n_1262),
.Y(n_1644)
);

O2A1O1Ixp5_ASAP7_75t_L g1645 ( 
.A1(n_1274),
.A2(n_1265),
.B(n_1283),
.C(n_1268),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1288),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1288),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1302),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1302),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1288),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1262),
.A2(n_899),
.B(n_1268),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1262),
.A2(n_899),
.B(n_1268),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1302),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1302),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_SL g1655 ( 
.A(n_1290),
.B(n_1025),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1441),
.B(n_865),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_SL g1657 ( 
.A(n_1290),
.B(n_1025),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1394),
.B(n_1262),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1302),
.Y(n_1659)
);

AO21x2_ASAP7_75t_L g1660 ( 
.A1(n_1274),
.A2(n_1081),
.B(n_1265),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1288),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1394),
.B(n_1262),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1394),
.B(n_1262),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1394),
.B(n_1262),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1302),
.Y(n_1665)
);

NOR2xp67_ASAP7_75t_L g1666 ( 
.A(n_1441),
.B(n_964),
.Y(n_1666)
);

NOR3xp33_ASAP7_75t_L g1667 ( 
.A(n_1327),
.B(n_1025),
.C(n_1232),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1262),
.A2(n_899),
.B(n_1268),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1302),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1394),
.B(n_1262),
.Y(n_1670)
);

OAI22x1_ASAP7_75t_L g1671 ( 
.A1(n_1304),
.A2(n_1025),
.B1(n_966),
.B2(n_996),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1262),
.A2(n_899),
.B(n_1268),
.Y(n_1672)
);

A2O1A1Ixp33_ASAP7_75t_L g1673 ( 
.A1(n_1262),
.A2(n_1268),
.B(n_1354),
.C(n_1226),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1394),
.B(n_1262),
.Y(n_1674)
);

AO31x2_ASAP7_75t_L g1675 ( 
.A1(n_1265),
.A2(n_1274),
.A3(n_1081),
.B(n_1195),
.Y(n_1675)
);

AO31x2_ASAP7_75t_L g1676 ( 
.A1(n_1265),
.A2(n_1274),
.A3(n_1081),
.B(n_1195),
.Y(n_1676)
);

NOR2xp67_ASAP7_75t_L g1677 ( 
.A(n_1441),
.B(n_964),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1262),
.A2(n_899),
.B(n_1268),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1380),
.A2(n_1360),
.B1(n_1378),
.B2(n_1358),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1262),
.A2(n_899),
.B(n_1268),
.Y(n_1680)
);

BUFx2_ASAP7_75t_L g1681 ( 
.A(n_1441),
.Y(n_1681)
);

AOI21x1_ASAP7_75t_L g1682 ( 
.A1(n_1435),
.A2(n_1081),
.B(n_1000),
.Y(n_1682)
);

AOI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1262),
.A2(n_899),
.B(n_1268),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1394),
.B(n_1262),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1441),
.B(n_865),
.Y(n_1685)
);

BUFx6f_ASAP7_75t_L g1686 ( 
.A(n_1224),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1394),
.B(n_1262),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1262),
.A2(n_899),
.B(n_1268),
.Y(n_1688)
);

BUFx2_ASAP7_75t_L g1689 ( 
.A(n_1441),
.Y(n_1689)
);

OAI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1262),
.A2(n_1268),
.B(n_1303),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_SL g1691 ( 
.A1(n_1338),
.A2(n_1357),
.B(n_1331),
.Y(n_1691)
);

OAI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1441),
.A2(n_1022),
.B1(n_1019),
.B2(n_973),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1290),
.B(n_1336),
.Y(n_1693)
);

AOI21x1_ASAP7_75t_L g1694 ( 
.A1(n_1435),
.A2(n_1081),
.B(n_1000),
.Y(n_1694)
);

NOR2xp67_ASAP7_75t_SL g1695 ( 
.A(n_1231),
.B(n_1025),
.Y(n_1695)
);

AO31x2_ASAP7_75t_L g1696 ( 
.A1(n_1265),
.A2(n_1274),
.A3(n_1081),
.B(n_1195),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1394),
.B(n_1262),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1302),
.Y(n_1698)
);

NAND3xp33_ASAP7_75t_SL g1699 ( 
.A(n_1304),
.B(n_968),
.C(n_1019),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1441),
.B(n_865),
.Y(n_1700)
);

OAI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1262),
.A2(n_1268),
.B(n_1303),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1447),
.Y(n_1702)
);

HB1xp67_ASAP7_75t_L g1703 ( 
.A(n_1524),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1456),
.Y(n_1704)
);

AOI22xp33_ASAP7_75t_L g1705 ( 
.A1(n_1544),
.A2(n_1565),
.B1(n_1606),
.B2(n_1467),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1462),
.Y(n_1706)
);

OAI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1534),
.A2(n_1536),
.B(n_1543),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1559),
.B(n_1535),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1598),
.B(n_1600),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_SL g1710 ( 
.A(n_1521),
.B(n_1490),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1641),
.B(n_1656),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1466),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1475),
.Y(n_1713)
);

AOI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1615),
.A2(n_1667),
.B1(n_1700),
.B2(n_1685),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1481),
.Y(n_1715)
);

HB1xp67_ASAP7_75t_L g1716 ( 
.A(n_1532),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1605),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1622),
.Y(n_1718)
);

AOI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1547),
.A2(n_1571),
.B1(n_1583),
.B2(n_1582),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1607),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1648),
.Y(n_1721)
);

AO21x1_ASAP7_75t_L g1722 ( 
.A1(n_1452),
.A2(n_1469),
.B(n_1532),
.Y(n_1722)
);

BUFx2_ASAP7_75t_L g1723 ( 
.A(n_1491),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1455),
.B(n_1614),
.Y(n_1724)
);

CKINVDCx20_ASAP7_75t_R g1725 ( 
.A(n_1623),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1649),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1597),
.A2(n_1673),
.B(n_1627),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1628),
.B(n_1482),
.Y(n_1728)
);

AO31x2_ASAP7_75t_L g1729 ( 
.A1(n_1639),
.A2(n_1451),
.A3(n_1634),
.B(n_1613),
.Y(n_1729)
);

BUFx3_ASAP7_75t_L g1730 ( 
.A(n_1473),
.Y(n_1730)
);

INVx1_ASAP7_75t_SL g1731 ( 
.A(n_1628),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1653),
.Y(n_1732)
);

INVx1_ASAP7_75t_SL g1733 ( 
.A(n_1528),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1592),
.B(n_1601),
.Y(n_1734)
);

OAI21x1_ASAP7_75t_L g1735 ( 
.A1(n_1621),
.A2(n_1701),
.B(n_1690),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1654),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1602),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1659),
.Y(n_1738)
);

NAND2x1p5_ASAP7_75t_L g1739 ( 
.A(n_1455),
.B(n_1614),
.Y(n_1739)
);

BUFx2_ASAP7_75t_L g1740 ( 
.A(n_1618),
.Y(n_1740)
);

CKINVDCx20_ASAP7_75t_R g1741 ( 
.A(n_1643),
.Y(n_1741)
);

AOI21x1_ASAP7_75t_L g1742 ( 
.A1(n_1593),
.A2(n_1682),
.B(n_1599),
.Y(n_1742)
);

NAND3xp33_ASAP7_75t_L g1743 ( 
.A(n_1573),
.B(n_1480),
.C(n_1478),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_SL g1744 ( 
.A(n_1569),
.B(n_1679),
.Y(n_1744)
);

INVx2_ASAP7_75t_SL g1745 ( 
.A(n_1473),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1665),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1554),
.B(n_1518),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1681),
.B(n_1689),
.Y(n_1748)
);

AO21x2_ASAP7_75t_L g1749 ( 
.A1(n_1546),
.A2(n_1549),
.B(n_1562),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1626),
.B(n_1554),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1669),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1482),
.B(n_1588),
.Y(n_1752)
);

OAI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1645),
.A2(n_1610),
.B(n_1609),
.Y(n_1753)
);

OAI21x1_ASAP7_75t_L g1754 ( 
.A1(n_1694),
.A2(n_1522),
.B(n_1624),
.Y(n_1754)
);

INVx3_ASAP7_75t_L g1755 ( 
.A(n_1631),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1576),
.B(n_1588),
.Y(n_1756)
);

OAI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1642),
.A2(n_1652),
.B(n_1651),
.Y(n_1757)
);

BUFx6f_ASAP7_75t_L g1758 ( 
.A(n_1631),
.Y(n_1758)
);

BUFx4f_ASAP7_75t_L g1759 ( 
.A(n_1640),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1698),
.Y(n_1760)
);

AOI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1668),
.A2(n_1678),
.B(n_1672),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1636),
.B(n_1638),
.Y(n_1762)
);

INVx3_ASAP7_75t_L g1763 ( 
.A(n_1631),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1537),
.B(n_1530),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1499),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1537),
.B(n_1493),
.Y(n_1766)
);

BUFx4f_ASAP7_75t_SL g1767 ( 
.A(n_1465),
.Y(n_1767)
);

INVx3_ASAP7_75t_L g1768 ( 
.A(n_1686),
.Y(n_1768)
);

OAI21xp5_ASAP7_75t_L g1769 ( 
.A1(n_1680),
.A2(n_1688),
.B(n_1683),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1504),
.Y(n_1770)
);

CKINVDCx20_ASAP7_75t_R g1771 ( 
.A(n_1502),
.Y(n_1771)
);

BUFx12f_ASAP7_75t_L g1772 ( 
.A(n_1507),
.Y(n_1772)
);

AO21x2_ASAP7_75t_L g1773 ( 
.A1(n_1625),
.A2(n_1660),
.B(n_1515),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1539),
.Y(n_1774)
);

AOI22xp33_ASAP7_75t_L g1775 ( 
.A1(n_1583),
.A2(n_1582),
.B1(n_1581),
.B2(n_1579),
.Y(n_1775)
);

BUFx3_ASAP7_75t_L g1776 ( 
.A(n_1527),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1550),
.B(n_1449),
.Y(n_1777)
);

OAI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1553),
.A2(n_1558),
.B(n_1585),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1550),
.Y(n_1779)
);

OAI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1553),
.A2(n_1558),
.B(n_1585),
.Y(n_1780)
);

AO31x2_ASAP7_75t_L g1781 ( 
.A1(n_1591),
.A2(n_1604),
.A3(n_1619),
.B(n_1617),
.Y(n_1781)
);

OR3x4_ASAP7_75t_SL g1782 ( 
.A(n_1612),
.B(n_1505),
.C(n_1526),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1458),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1458),
.Y(n_1784)
);

BUFx2_ASAP7_75t_R g1785 ( 
.A(n_1637),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1484),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1596),
.B(n_1616),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1675),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1676),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1484),
.Y(n_1790)
);

AOI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1506),
.A2(n_1630),
.B(n_1620),
.Y(n_1791)
);

AO31x2_ASAP7_75t_L g1792 ( 
.A1(n_1630),
.A2(n_1658),
.A3(n_1664),
.B(n_1663),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1494),
.Y(n_1793)
);

INVx2_ASAP7_75t_SL g1794 ( 
.A(n_1471),
.Y(n_1794)
);

HB1xp67_ASAP7_75t_L g1795 ( 
.A(n_1527),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1494),
.Y(n_1796)
);

AO21x2_ASAP7_75t_L g1797 ( 
.A1(n_1625),
.A2(n_1660),
.B(n_1485),
.Y(n_1797)
);

CKINVDCx20_ASAP7_75t_R g1798 ( 
.A(n_1529),
.Y(n_1798)
);

A2O1A1Ixp33_ASAP7_75t_L g1799 ( 
.A1(n_1635),
.A2(n_1662),
.B(n_1697),
.C(n_1644),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1498),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1445),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1595),
.B(n_1633),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1676),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1445),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1693),
.B(n_1459),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1474),
.Y(n_1806)
);

OR2x6_ASAP7_75t_L g1807 ( 
.A(n_1525),
.B(n_1500),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1693),
.B(n_1519),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1479),
.B(n_1512),
.Y(n_1809)
);

AO21x2_ASAP7_75t_L g1810 ( 
.A1(n_1670),
.A2(n_1684),
.B(n_1674),
.Y(n_1810)
);

OR2x6_ASAP7_75t_L g1811 ( 
.A(n_1479),
.B(n_1540),
.Y(n_1811)
);

OAI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1674),
.A2(n_1687),
.B(n_1684),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1696),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1696),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1474),
.Y(n_1815)
);

NAND2x1p5_ASAP7_75t_L g1816 ( 
.A(n_1568),
.B(n_1508),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1542),
.B(n_1692),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_1612),
.Y(n_1818)
);

OAI21x1_ASAP7_75t_SL g1819 ( 
.A1(n_1548),
.A2(n_1463),
.B(n_1469),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1696),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1509),
.B(n_1531),
.Y(n_1821)
);

INVx2_ASAP7_75t_SL g1822 ( 
.A(n_1590),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1511),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1511),
.Y(n_1824)
);

OAI21x1_ASAP7_75t_L g1825 ( 
.A1(n_1566),
.A2(n_1584),
.B(n_1492),
.Y(n_1825)
);

NOR2xp67_ASAP7_75t_L g1826 ( 
.A(n_1699),
.B(n_1461),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1496),
.B(n_1468),
.Y(n_1827)
);

INVx8_ASAP7_75t_L g1828 ( 
.A(n_1568),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1472),
.B(n_1538),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1497),
.B(n_1568),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1477),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1510),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1570),
.B(n_1655),
.Y(n_1833)
);

AND2x4_ASAP7_75t_L g1834 ( 
.A(n_1497),
.B(n_1557),
.Y(n_1834)
);

OAI21x1_ASAP7_75t_L g1835 ( 
.A1(n_1446),
.A2(n_1584),
.B(n_1483),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1523),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1594),
.Y(n_1837)
);

AND2x4_ASAP7_75t_L g1838 ( 
.A(n_1497),
.B(n_1557),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1611),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1629),
.Y(n_1840)
);

INVx1_ASAP7_75t_SL g1841 ( 
.A(n_1657),
.Y(n_1841)
);

AO31x2_ASAP7_75t_L g1842 ( 
.A1(n_1578),
.A2(n_1450),
.A3(n_1575),
.B(n_1514),
.Y(n_1842)
);

BUFx4f_ASAP7_75t_SL g1843 ( 
.A(n_1603),
.Y(n_1843)
);

OAI21x1_ASAP7_75t_L g1844 ( 
.A1(n_1691),
.A2(n_1561),
.B(n_1560),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_L g1845 ( 
.A(n_1486),
.B(n_1533),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1646),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1647),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1671),
.B(n_1495),
.Y(n_1848)
);

INVx1_ASAP7_75t_SL g1849 ( 
.A(n_1632),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1472),
.B(n_1552),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1517),
.B(n_1457),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1650),
.Y(n_1852)
);

BUFx2_ASAP7_75t_R g1853 ( 
.A(n_1460),
.Y(n_1853)
);

AOI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1569),
.A2(n_1551),
.B(n_1545),
.Y(n_1854)
);

OA21x2_ASAP7_75t_L g1855 ( 
.A1(n_1488),
.A2(n_1501),
.B(n_1567),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1567),
.B(n_1470),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1661),
.Y(n_1857)
);

INVx6_ASAP7_75t_L g1858 ( 
.A(n_1457),
.Y(n_1858)
);

AOI22x1_ASAP7_75t_L g1859 ( 
.A1(n_1503),
.A2(n_1564),
.B1(n_1541),
.B2(n_1577),
.Y(n_1859)
);

INVx3_ASAP7_75t_SL g1860 ( 
.A(n_1574),
.Y(n_1860)
);

NOR2xp67_ASAP7_75t_SL g1861 ( 
.A(n_1695),
.B(n_1443),
.Y(n_1861)
);

A2O1A1Ixp33_ASAP7_75t_L g1862 ( 
.A1(n_1464),
.A2(n_1450),
.B(n_1448),
.C(n_1444),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1476),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1589),
.B(n_1666),
.Y(n_1864)
);

AOI22x1_ASAP7_75t_L g1865 ( 
.A1(n_1556),
.A2(n_1572),
.B1(n_1516),
.B2(n_1563),
.Y(n_1865)
);

AO21x2_ASAP7_75t_L g1866 ( 
.A1(n_1453),
.A2(n_1572),
.B(n_1587),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1677),
.B(n_1580),
.Y(n_1867)
);

AO31x2_ASAP7_75t_L g1868 ( 
.A1(n_1454),
.A2(n_1489),
.A3(n_1563),
.B(n_1487),
.Y(n_1868)
);

AOI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1520),
.A2(n_1555),
.B1(n_1476),
.B2(n_1513),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1513),
.Y(n_1870)
);

AOI22xp5_ASAP7_75t_L g1871 ( 
.A1(n_1513),
.A2(n_1025),
.B1(n_933),
.B2(n_973),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1447),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1447),
.Y(n_1873)
);

NAND3xp33_ASAP7_75t_L g1874 ( 
.A(n_1573),
.B(n_1243),
.C(n_1667),
.Y(n_1874)
);

AND2x4_ASAP7_75t_L g1875 ( 
.A(n_1455),
.B(n_1614),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1524),
.B(n_865),
.Y(n_1876)
);

INVx1_ASAP7_75t_SL g1877 ( 
.A(n_1628),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1447),
.Y(n_1878)
);

OAI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1534),
.A2(n_1536),
.B(n_1268),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1524),
.B(n_865),
.Y(n_1880)
);

AO21x2_ASAP7_75t_L g1881 ( 
.A1(n_1586),
.A2(n_1546),
.B(n_1608),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1447),
.Y(n_1882)
);

NOR2xp67_ASAP7_75t_L g1883 ( 
.A(n_1455),
.B(n_1441),
.Y(n_1883)
);

AOI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1615),
.A2(n_1025),
.B1(n_933),
.B2(n_973),
.Y(n_1884)
);

NAND2x1p5_ASAP7_75t_L g1885 ( 
.A(n_1455),
.B(n_1614),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1447),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_SL g1887 ( 
.A(n_1521),
.B(n_1490),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1524),
.B(n_865),
.Y(n_1888)
);

AND2x4_ASAP7_75t_L g1889 ( 
.A(n_1455),
.B(n_1614),
.Y(n_1889)
);

AOI22xp33_ASAP7_75t_L g1890 ( 
.A1(n_1544),
.A2(n_1126),
.B1(n_1565),
.B2(n_1606),
.Y(n_1890)
);

INVxp67_ASAP7_75t_L g1891 ( 
.A(n_1876),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1702),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1704),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1706),
.Y(n_1894)
);

HB1xp67_ASAP7_75t_L g1895 ( 
.A(n_1762),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1712),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1713),
.Y(n_1897)
);

BUFx3_ASAP7_75t_L g1898 ( 
.A(n_1828),
.Y(n_1898)
);

OR2x6_ASAP7_75t_L g1899 ( 
.A(n_1811),
.B(n_1828),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1750),
.B(n_1747),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1735),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1774),
.B(n_1779),
.Y(n_1902)
);

HB1xp67_ASAP7_75t_SL g1903 ( 
.A(n_1785),
.Y(n_1903)
);

INVx3_ASAP7_75t_L g1904 ( 
.A(n_1828),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1836),
.B(n_1840),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1729),
.Y(n_1906)
);

CKINVDCx20_ASAP7_75t_R g1907 ( 
.A(n_1767),
.Y(n_1907)
);

BUFx2_ASAP7_75t_L g1908 ( 
.A(n_1781),
.Y(n_1908)
);

INVxp67_ASAP7_75t_L g1909 ( 
.A(n_1880),
.Y(n_1909)
);

AO21x1_ASAP7_75t_SL g1910 ( 
.A1(n_1716),
.A2(n_1812),
.B(n_1707),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1778),
.B(n_1780),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1836),
.B(n_1840),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1729),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1715),
.Y(n_1914)
);

HB1xp67_ASAP7_75t_L g1915 ( 
.A(n_1703),
.Y(n_1915)
);

AND2x4_ASAP7_75t_L g1916 ( 
.A(n_1830),
.B(n_1834),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1846),
.B(n_1852),
.Y(n_1917)
);

HB1xp67_ASAP7_75t_L g1918 ( 
.A(n_1703),
.Y(n_1918)
);

HB1xp67_ASAP7_75t_L g1919 ( 
.A(n_1740),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1846),
.B(n_1852),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1750),
.B(n_1764),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1888),
.B(n_1711),
.Y(n_1922)
);

BUFx8_ASAP7_75t_L g1923 ( 
.A(n_1772),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1857),
.B(n_1775),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1857),
.B(n_1775),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1708),
.B(n_1766),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1709),
.B(n_1884),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1717),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1719),
.B(n_1832),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1718),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1719),
.B(n_1837),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1721),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1726),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1732),
.Y(n_1934)
);

OR2x2_ASAP7_75t_L g1935 ( 
.A(n_1777),
.B(n_1817),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1736),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1705),
.B(n_1714),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1839),
.B(n_1847),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1738),
.Y(n_1939)
);

BUFx3_ASAP7_75t_L g1940 ( 
.A(n_1724),
.Y(n_1940)
);

HB1xp67_ASAP7_75t_L g1941 ( 
.A(n_1731),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1746),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1705),
.B(n_1871),
.Y(n_1943)
);

OAI21x1_ASAP7_75t_L g1944 ( 
.A1(n_1754),
.A2(n_1742),
.B(n_1753),
.Y(n_1944)
);

OAI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1862),
.A2(n_1874),
.B(n_1827),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1751),
.Y(n_1946)
);

AO21x2_ASAP7_75t_L g1947 ( 
.A1(n_1761),
.A2(n_1769),
.B(n_1757),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1737),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1760),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1872),
.Y(n_1950)
);

OAI21xp5_ASAP7_75t_L g1951 ( 
.A1(n_1862),
.A2(n_1854),
.B(n_1829),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1783),
.B(n_1784),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1873),
.Y(n_1953)
);

HB1xp67_ASAP7_75t_L g1954 ( 
.A(n_1877),
.Y(n_1954)
);

HB1xp67_ASAP7_75t_L g1955 ( 
.A(n_1734),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1878),
.Y(n_1956)
);

HB1xp67_ASAP7_75t_L g1957 ( 
.A(n_1748),
.Y(n_1957)
);

BUFx3_ASAP7_75t_L g1958 ( 
.A(n_1724),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1882),
.Y(n_1959)
);

CKINVDCx5p33_ASAP7_75t_R g1960 ( 
.A(n_1759),
.Y(n_1960)
);

OR2x6_ASAP7_75t_L g1961 ( 
.A(n_1811),
.B(n_1722),
.Y(n_1961)
);

HB1xp67_ASAP7_75t_L g1962 ( 
.A(n_1883),
.Y(n_1962)
);

OAI21x1_ASAP7_75t_SL g1963 ( 
.A1(n_1819),
.A2(n_1859),
.B(n_1720),
.Y(n_1963)
);

HB1xp67_ASAP7_75t_L g1964 ( 
.A(n_1787),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1886),
.Y(n_1965)
);

INVx2_ASAP7_75t_SL g1966 ( 
.A(n_1724),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1781),
.Y(n_1967)
);

INVx2_ASAP7_75t_SL g1968 ( 
.A(n_1875),
.Y(n_1968)
);

AND2x4_ASAP7_75t_L g1969 ( 
.A(n_1830),
.B(n_1834),
.Y(n_1969)
);

CKINVDCx14_ASAP7_75t_R g1970 ( 
.A(n_1759),
.Y(n_1970)
);

HB1xp67_ASAP7_75t_L g1971 ( 
.A(n_1811),
.Y(n_1971)
);

HB1xp67_ASAP7_75t_L g1972 ( 
.A(n_1728),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1765),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1770),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1792),
.Y(n_1975)
);

INVx3_ASAP7_75t_L g1976 ( 
.A(n_1875),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1800),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1821),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1890),
.B(n_1808),
.Y(n_1979)
);

BUFx2_ASAP7_75t_L g1980 ( 
.A(n_1792),
.Y(n_1980)
);

OR2x2_ASAP7_75t_L g1981 ( 
.A(n_1792),
.B(n_1810),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1831),
.Y(n_1982)
);

OR2x2_ASAP7_75t_L g1983 ( 
.A(n_1810),
.B(n_1801),
.Y(n_1983)
);

BUFx3_ASAP7_75t_L g1984 ( 
.A(n_1875),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1890),
.B(n_1804),
.Y(n_1985)
);

BUFx2_ASAP7_75t_L g1986 ( 
.A(n_1799),
.Y(n_1986)
);

OR2x2_ASAP7_75t_L g1987 ( 
.A(n_1856),
.B(n_1842),
.Y(n_1987)
);

AO21x2_ASAP7_75t_L g1988 ( 
.A1(n_1727),
.A2(n_1743),
.B(n_1879),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1870),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1863),
.Y(n_1990)
);

NOR2xp33_ASAP7_75t_L g1991 ( 
.A(n_1756),
.B(n_1853),
.Y(n_1991)
);

HB1xp67_ASAP7_75t_L g1992 ( 
.A(n_1752),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1809),
.B(n_1805),
.Y(n_1993)
);

AOI22xp33_ASAP7_75t_L g1994 ( 
.A1(n_1756),
.A2(n_1790),
.B1(n_1786),
.B2(n_1793),
.Y(n_1994)
);

AND2x4_ASAP7_75t_L g1995 ( 
.A(n_1838),
.B(n_1844),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1850),
.Y(n_1996)
);

AO21x2_ASAP7_75t_L g1997 ( 
.A1(n_1791),
.A2(n_1744),
.B(n_1869),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1739),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1739),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1885),
.Y(n_2000)
);

BUFx3_ASAP7_75t_L g2001 ( 
.A(n_1889),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1892),
.Y(n_2002)
);

BUFx2_ASAP7_75t_L g2003 ( 
.A(n_1995),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1893),
.Y(n_2004)
);

NAND3xp33_ASAP7_75t_L g2005 ( 
.A(n_1945),
.B(n_1848),
.C(n_1865),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1894),
.Y(n_2006)
);

INVxp67_ASAP7_75t_SL g2007 ( 
.A(n_1981),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1896),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1897),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1914),
.Y(n_2010)
);

CKINVDCx11_ASAP7_75t_R g2011 ( 
.A(n_1907),
.Y(n_2011)
);

AND2x4_ASAP7_75t_L g2012 ( 
.A(n_1995),
.B(n_1720),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1928),
.Y(n_2013)
);

HB1xp67_ASAP7_75t_L g2014 ( 
.A(n_1895),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1989),
.Y(n_2015)
);

NOR2x1_ASAP7_75t_SL g2016 ( 
.A(n_1899),
.B(n_1807),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1905),
.B(n_1868),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1926),
.B(n_1796),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1912),
.B(n_1868),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1930),
.Y(n_2020)
);

INVx4_ASAP7_75t_L g2021 ( 
.A(n_1899),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1932),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1926),
.B(n_1806),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1917),
.B(n_1868),
.Y(n_2024)
);

HB1xp67_ASAP7_75t_L g2025 ( 
.A(n_1972),
.Y(n_2025)
);

INVx1_ASAP7_75t_SL g2026 ( 
.A(n_1960),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1920),
.B(n_1868),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1989),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1911),
.B(n_1788),
.Y(n_2029)
);

BUFx3_ASAP7_75t_L g2030 ( 
.A(n_1898),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1911),
.B(n_1789),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1990),
.Y(n_2032)
);

AND2x4_ASAP7_75t_L g2033 ( 
.A(n_1995),
.B(n_1789),
.Y(n_2033)
);

OR2x2_ASAP7_75t_L g2034 ( 
.A(n_1983),
.B(n_1987),
.Y(n_2034)
);

INVx2_ASAP7_75t_SL g2035 ( 
.A(n_2001),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1911),
.B(n_1803),
.Y(n_2036)
);

AND2x4_ASAP7_75t_L g2037 ( 
.A(n_1961),
.B(n_1803),
.Y(n_2037)
);

INVx2_ASAP7_75t_SL g2038 ( 
.A(n_2001),
.Y(n_2038)
);

HB1xp67_ASAP7_75t_L g2039 ( 
.A(n_1919),
.Y(n_2039)
);

BUFx3_ASAP7_75t_L g2040 ( 
.A(n_1898),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1933),
.Y(n_2041)
);

AOI22xp33_ASAP7_75t_L g2042 ( 
.A1(n_1937),
.A2(n_1723),
.B1(n_1855),
.B2(n_1845),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1986),
.B(n_1924),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1983),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1934),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1936),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1986),
.B(n_1924),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1939),
.Y(n_2048)
);

NAND2xp33_ASAP7_75t_R g2049 ( 
.A(n_1960),
.B(n_1818),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1942),
.Y(n_2050)
);

INVx4_ASAP7_75t_L g2051 ( 
.A(n_1899),
.Y(n_2051)
);

AOI221xp5_ASAP7_75t_L g2052 ( 
.A1(n_1927),
.A2(n_1845),
.B1(n_1823),
.B2(n_1824),
.C(n_1815),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1902),
.B(n_1833),
.Y(n_2053)
);

BUFx2_ASAP7_75t_L g2054 ( 
.A(n_1908),
.Y(n_2054)
);

AOI22xp33_ASAP7_75t_L g2055 ( 
.A1(n_1943),
.A2(n_1855),
.B1(n_1861),
.B2(n_1867),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1902),
.B(n_1841),
.Y(n_2056)
);

OR2x2_ASAP7_75t_L g2057 ( 
.A(n_1987),
.B(n_1813),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1978),
.B(n_1842),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1921),
.B(n_1842),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_1925),
.B(n_1814),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1948),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_1925),
.B(n_1820),
.Y(n_2062)
);

OR2x2_ASAP7_75t_L g2063 ( 
.A(n_1915),
.B(n_1797),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_1967),
.B(n_1773),
.Y(n_2064)
);

HB1xp67_ASAP7_75t_L g2065 ( 
.A(n_1918),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_1967),
.B(n_1773),
.Y(n_2066)
);

NOR2xp33_ASAP7_75t_L g2067 ( 
.A(n_1922),
.B(n_1772),
.Y(n_2067)
);

BUFx2_ASAP7_75t_L g2068 ( 
.A(n_1908),
.Y(n_2068)
);

OR2x2_ASAP7_75t_L g2069 ( 
.A(n_1935),
.B(n_1881),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1946),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_1975),
.B(n_1881),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1949),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1950),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1953),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1900),
.B(n_1842),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1938),
.B(n_1866),
.Y(n_2076)
);

BUFx3_ASAP7_75t_L g2077 ( 
.A(n_1904),
.Y(n_2077)
);

CKINVDCx16_ASAP7_75t_R g2078 ( 
.A(n_1970),
.Y(n_2078)
);

OR2x2_ASAP7_75t_L g2079 ( 
.A(n_1935),
.B(n_1749),
.Y(n_2079)
);

BUFx3_ASAP7_75t_L g2080 ( 
.A(n_1904),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1956),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1959),
.Y(n_2082)
);

OA21x2_ASAP7_75t_L g2083 ( 
.A1(n_1944),
.A2(n_1835),
.B(n_1825),
.Y(n_2083)
);

HB1xp67_ASAP7_75t_L g2084 ( 
.A(n_1941),
.Y(n_2084)
);

AND2x4_ASAP7_75t_SL g2085 ( 
.A(n_1899),
.B(n_1758),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1952),
.B(n_1802),
.Y(n_2086)
);

NOR2xp33_ASAP7_75t_L g2087 ( 
.A(n_1996),
.B(n_1767),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_2059),
.B(n_1980),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_2061),
.Y(n_2089)
);

INVx2_ASAP7_75t_SL g2090 ( 
.A(n_2003),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2015),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2043),
.B(n_1980),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_2075),
.B(n_2044),
.Y(n_2093)
);

INVx2_ASAP7_75t_SL g2094 ( 
.A(n_2003),
.Y(n_2094)
);

INVx5_ASAP7_75t_L g2095 ( 
.A(n_2021),
.Y(n_2095)
);

NOR2xp33_ASAP7_75t_L g2096 ( 
.A(n_2087),
.B(n_1843),
.Y(n_2096)
);

AND2x4_ASAP7_75t_L g2097 ( 
.A(n_2012),
.B(n_2033),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2043),
.B(n_1906),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2015),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2028),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2028),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2032),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_2047),
.B(n_1913),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_2071),
.B(n_1947),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_2076),
.B(n_1947),
.Y(n_2105)
);

BUFx2_ASAP7_75t_L g2106 ( 
.A(n_2007),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2076),
.B(n_1947),
.Y(n_2107)
);

BUFx2_ASAP7_75t_L g2108 ( 
.A(n_2054),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2017),
.B(n_1988),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_2029),
.B(n_1988),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_2029),
.B(n_1988),
.Y(n_2111)
);

BUFx6f_ASAP7_75t_L g2112 ( 
.A(n_2083),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_2017),
.B(n_1910),
.Y(n_2113)
);

INVx1_ASAP7_75t_SL g2114 ( 
.A(n_2030),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2019),
.B(n_1910),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2058),
.B(n_1929),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2019),
.B(n_1997),
.Y(n_2117)
);

OR2x2_ASAP7_75t_L g2118 ( 
.A(n_2034),
.B(n_2069),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_2079),
.B(n_2024),
.Y(n_2119)
);

BUFx2_ASAP7_75t_L g2120 ( 
.A(n_2054),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_2024),
.B(n_1997),
.Y(n_2121)
);

AND2x4_ASAP7_75t_L g2122 ( 
.A(n_2012),
.B(n_1901),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2064),
.Y(n_2123)
);

HB1xp67_ASAP7_75t_L g2124 ( 
.A(n_2065),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2064),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2109),
.B(n_2027),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2124),
.B(n_2014),
.Y(n_2127)
);

OR2x2_ASAP7_75t_L g2128 ( 
.A(n_2118),
.B(n_2063),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2091),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_2089),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2091),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_2109),
.B(n_2027),
.Y(n_2132)
);

NAND2x1_ASAP7_75t_L g2133 ( 
.A(n_2090),
.B(n_1963),
.Y(n_2133)
);

OR2x2_ASAP7_75t_L g2134 ( 
.A(n_2118),
.B(n_2063),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2099),
.Y(n_2135)
);

INVx4_ASAP7_75t_L g2136 ( 
.A(n_2095),
.Y(n_2136)
);

INVx3_ASAP7_75t_L g2137 ( 
.A(n_2112),
.Y(n_2137)
);

AND2x4_ASAP7_75t_SL g2138 ( 
.A(n_2097),
.B(n_2021),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2105),
.B(n_2060),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_2124),
.B(n_2025),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2099),
.Y(n_2141)
);

INVx1_ASAP7_75t_SL g2142 ( 
.A(n_2114),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_2105),
.B(n_2060),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_2123),
.B(n_2084),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_2123),
.B(n_2039),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_2107),
.B(n_2062),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2100),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2125),
.B(n_2002),
.Y(n_2148)
);

OR2x2_ASAP7_75t_L g2149 ( 
.A(n_2119),
.B(n_2057),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_2107),
.B(n_2062),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2100),
.Y(n_2151)
);

AND2x4_ASAP7_75t_SL g2152 ( 
.A(n_2097),
.B(n_2021),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2125),
.B(n_2004),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2101),
.Y(n_2154)
);

OR2x2_ASAP7_75t_L g2155 ( 
.A(n_2119),
.B(n_2057),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_2110),
.B(n_2066),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2101),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_2110),
.B(n_2066),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2102),
.Y(n_2159)
);

AND2x4_ASAP7_75t_L g2160 ( 
.A(n_2122),
.B(n_2037),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_2110),
.B(n_2031),
.Y(n_2161)
);

NAND2xp33_ASAP7_75t_L g2162 ( 
.A(n_2114),
.B(n_1818),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2102),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2111),
.B(n_2031),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2111),
.B(n_2036),
.Y(n_2165)
);

OR2x6_ASAP7_75t_L g2166 ( 
.A(n_2106),
.B(n_2068),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2111),
.B(n_2036),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2145),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_2126),
.B(n_2093),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2144),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2129),
.Y(n_2171)
);

OR2x2_ASAP7_75t_L g2172 ( 
.A(n_2128),
.B(n_2088),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2156),
.B(n_2104),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_2126),
.B(n_2132),
.Y(n_2174)
);

NOR2x1_ASAP7_75t_L g2175 ( 
.A(n_2136),
.B(n_1907),
.Y(n_2175)
);

NAND2x1p5_ASAP7_75t_L g2176 ( 
.A(n_2136),
.B(n_2095),
.Y(n_2176)
);

OAI22xp5_ASAP7_75t_L g2177 ( 
.A1(n_2136),
.A2(n_2095),
.B1(n_1903),
.B2(n_2051),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2129),
.Y(n_2178)
);

O2A1O1Ixp5_ASAP7_75t_L g2179 ( 
.A1(n_2136),
.A2(n_1991),
.B(n_2067),
.C(n_2051),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_2130),
.Y(n_2180)
);

BUFx2_ASAP7_75t_L g2181 ( 
.A(n_2166),
.Y(n_2181)
);

OR2x2_ASAP7_75t_L g2182 ( 
.A(n_2128),
.B(n_2088),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_2156),
.B(n_2104),
.Y(n_2183)
);

OR2x2_ASAP7_75t_L g2184 ( 
.A(n_2134),
.B(n_2106),
.Y(n_2184)
);

NOR2xp33_ASAP7_75t_L g2185 ( 
.A(n_2127),
.B(n_2011),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2131),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2158),
.B(n_2104),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2131),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_2132),
.B(n_2158),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_2139),
.B(n_2117),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2135),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_2139),
.B(n_2143),
.Y(n_2192)
);

OR2x2_ASAP7_75t_L g2193 ( 
.A(n_2134),
.B(n_2140),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2143),
.B(n_2093),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2135),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2141),
.Y(n_2196)
);

AND2x4_ASAP7_75t_L g2197 ( 
.A(n_2166),
.B(n_2097),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2141),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_2146),
.B(n_2117),
.Y(n_2199)
);

INVx3_ASAP7_75t_L g2200 ( 
.A(n_2133),
.Y(n_2200)
);

INVxp67_ASAP7_75t_L g2201 ( 
.A(n_2142),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_2146),
.B(n_2121),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2147),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2147),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2190),
.B(n_2150),
.Y(n_2205)
);

INVx2_ASAP7_75t_SL g2206 ( 
.A(n_2175),
.Y(n_2206)
);

A2O1A1Ixp33_ASAP7_75t_L g2207 ( 
.A1(n_2179),
.A2(n_2162),
.B(n_2152),
.C(n_2138),
.Y(n_2207)
);

OAI22xp33_ASAP7_75t_L g2208 ( 
.A1(n_2176),
.A2(n_2166),
.B1(n_2095),
.B2(n_2133),
.Y(n_2208)
);

OR2x2_ASAP7_75t_L g2209 ( 
.A(n_2184),
.B(n_2149),
.Y(n_2209)
);

OAI221xp5_ASAP7_75t_L g2210 ( 
.A1(n_2181),
.A2(n_2200),
.B1(n_2176),
.B2(n_2201),
.C(n_2170),
.Y(n_2210)
);

INVxp67_ASAP7_75t_L g2211 ( 
.A(n_2185),
.Y(n_2211)
);

OAI31xp33_ASAP7_75t_L g2212 ( 
.A1(n_2176),
.A2(n_1962),
.A3(n_2040),
.B(n_2030),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2184),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2193),
.Y(n_2214)
);

OAI21xp33_ASAP7_75t_L g2215 ( 
.A1(n_2172),
.A2(n_2166),
.B(n_2115),
.Y(n_2215)
);

INVxp67_ASAP7_75t_L g2216 ( 
.A(n_2193),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_2173),
.B(n_2183),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_2190),
.B(n_2150),
.Y(n_2218)
);

NAND2xp33_ASAP7_75t_L g2219 ( 
.A(n_2177),
.B(n_2095),
.Y(n_2219)
);

AOI22xp5_ASAP7_75t_L g2220 ( 
.A1(n_2197),
.A2(n_2113),
.B1(n_2115),
.B2(n_2166),
.Y(n_2220)
);

OAI322xp33_ASAP7_75t_L g2221 ( 
.A1(n_2172),
.A2(n_2182),
.A3(n_2168),
.B1(n_2169),
.B2(n_2174),
.C1(n_2194),
.C2(n_2189),
.Y(n_2221)
);

NAND3xp33_ASAP7_75t_L g2222 ( 
.A(n_2181),
.B(n_2005),
.C(n_2055),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2202),
.B(n_2167),
.Y(n_2223)
);

AOI22xp5_ASAP7_75t_L g2224 ( 
.A1(n_2197),
.A2(n_2113),
.B1(n_2160),
.B2(n_2092),
.Y(n_2224)
);

OAI322xp33_ASAP7_75t_L g2225 ( 
.A1(n_2182),
.A2(n_2149),
.A3(n_2155),
.B1(n_2148),
.B2(n_2153),
.C1(n_2116),
.C2(n_1891),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2186),
.Y(n_2226)
);

AOI21xp33_ASAP7_75t_L g2227 ( 
.A1(n_2200),
.A2(n_1849),
.B(n_1909),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_2202),
.B(n_2161),
.Y(n_2228)
);

AND2x4_ASAP7_75t_L g2229 ( 
.A(n_2197),
.B(n_2160),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2186),
.Y(n_2230)
);

OAI33xp33_ASAP7_75t_L g2231 ( 
.A1(n_2199),
.A2(n_2155),
.A3(n_2116),
.B1(n_2056),
.B2(n_2053),
.B3(n_1979),
.Y(n_2231)
);

OR2x2_ASAP7_75t_L g2232 ( 
.A(n_2192),
.B(n_2161),
.Y(n_2232)
);

INVxp67_ASAP7_75t_L g2233 ( 
.A(n_2171),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2178),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2173),
.B(n_2183),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2188),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_2180),
.Y(n_2237)
);

INVxp67_ASAP7_75t_L g2238 ( 
.A(n_2211),
.Y(n_2238)
);

AND2x4_ASAP7_75t_L g2239 ( 
.A(n_2206),
.B(n_2200),
.Y(n_2239)
);

AOI22xp5_ASAP7_75t_L g2240 ( 
.A1(n_2231),
.A2(n_2187),
.B1(n_2192),
.B2(n_2160),
.Y(n_2240)
);

OAI21xp33_ASAP7_75t_L g2241 ( 
.A1(n_2215),
.A2(n_2187),
.B(n_2191),
.Y(n_2241)
);

OAI211xp5_ASAP7_75t_SL g2242 ( 
.A1(n_2210),
.A2(n_2011),
.B(n_2026),
.C(n_2042),
.Y(n_2242)
);

AOI322xp5_ASAP7_75t_L g2243 ( 
.A1(n_2216),
.A2(n_2164),
.A3(n_2165),
.B1(n_2167),
.B2(n_2092),
.C1(n_1955),
.C2(n_1957),
.Y(n_2243)
);

HB1xp67_ASAP7_75t_L g2244 ( 
.A(n_2233),
.Y(n_2244)
);

AND2x2_ASAP7_75t_L g2245 ( 
.A(n_2229),
.B(n_2164),
.Y(n_2245)
);

OAI21xp33_ASAP7_75t_SL g2246 ( 
.A1(n_2212),
.A2(n_2094),
.B(n_2090),
.Y(n_2246)
);

AOI221x1_ASAP7_75t_SL g2247 ( 
.A1(n_2214),
.A2(n_2023),
.B1(n_2018),
.B2(n_2096),
.C(n_1826),
.Y(n_2247)
);

OAI211xp5_ASAP7_75t_L g2248 ( 
.A1(n_2207),
.A2(n_1733),
.B(n_2040),
.C(n_1771),
.Y(n_2248)
);

OAI321xp33_ASAP7_75t_L g2249 ( 
.A1(n_2208),
.A2(n_2094),
.A3(n_2090),
.B1(n_2120),
.B2(n_2108),
.C(n_1951),
.Y(n_2249)
);

AOI221xp5_ASAP7_75t_L g2250 ( 
.A1(n_2221),
.A2(n_2196),
.B1(n_2203),
.B2(n_2198),
.C(n_2195),
.Y(n_2250)
);

AO21x1_ASAP7_75t_L g2251 ( 
.A1(n_2227),
.A2(n_2051),
.B(n_2138),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2226),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2213),
.B(n_2204),
.Y(n_2253)
);

AOI21xp5_ASAP7_75t_R g2254 ( 
.A1(n_2229),
.A2(n_1782),
.B(n_2078),
.Y(n_2254)
);

O2A1O1Ixp5_ASAP7_75t_L g2255 ( 
.A1(n_2225),
.A2(n_2180),
.B(n_2137),
.C(n_2154),
.Y(n_2255)
);

OAI221xp5_ASAP7_75t_L g2256 ( 
.A1(n_2220),
.A2(n_2120),
.B1(n_2108),
.B2(n_2094),
.C(n_1864),
.Y(n_2256)
);

OAI222xp33_ASAP7_75t_L g2257 ( 
.A1(n_2224),
.A2(n_2095),
.B1(n_2160),
.B2(n_2165),
.C1(n_2121),
.C2(n_2151),
.Y(n_2257)
);

OAI22xp5_ASAP7_75t_L g2258 ( 
.A1(n_2254),
.A2(n_2232),
.B1(n_2235),
.B2(n_2217),
.Y(n_2258)
);

AOI221xp5_ASAP7_75t_L g2259 ( 
.A1(n_2247),
.A2(n_2227),
.B1(n_2222),
.B2(n_2236),
.C(n_2234),
.Y(n_2259)
);

A2O1A1Ixp33_ASAP7_75t_L g2260 ( 
.A1(n_2246),
.A2(n_2219),
.B(n_2209),
.C(n_2152),
.Y(n_2260)
);

AOI22xp5_ASAP7_75t_L g2261 ( 
.A1(n_2248),
.A2(n_2217),
.B1(n_2235),
.B2(n_2230),
.Y(n_2261)
);

OAI221xp5_ASAP7_75t_SL g2262 ( 
.A1(n_2248),
.A2(n_1994),
.B1(n_2205),
.B2(n_2228),
.C(n_2223),
.Y(n_2262)
);

A2O1A1Ixp33_ASAP7_75t_L g2263 ( 
.A1(n_2255),
.A2(n_2152),
.B(n_2138),
.C(n_2218),
.Y(n_2263)
);

NOR2xp67_ASAP7_75t_L g2264 ( 
.A(n_2249),
.B(n_2095),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_SL g2265 ( 
.A(n_2251),
.B(n_2250),
.Y(n_2265)
);

AOI21xp5_ASAP7_75t_L g2266 ( 
.A1(n_2254),
.A2(n_2016),
.B(n_1887),
.Y(n_2266)
);

A2O1A1Ixp33_ASAP7_75t_L g2267 ( 
.A1(n_2241),
.A2(n_1710),
.B(n_1771),
.C(n_1904),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2253),
.Y(n_2268)
);

AOI221xp5_ASAP7_75t_L g2269 ( 
.A1(n_2238),
.A2(n_1954),
.B1(n_2237),
.B2(n_1964),
.C(n_2052),
.Y(n_2269)
);

OAI32xp33_ASAP7_75t_L g2270 ( 
.A1(n_2242),
.A2(n_1741),
.A3(n_1725),
.B1(n_2080),
.B2(n_2077),
.Y(n_2270)
);

OAI21xp33_ASAP7_75t_L g2271 ( 
.A1(n_2243),
.A2(n_2154),
.B(n_2151),
.Y(n_2271)
);

OAI22xp33_ASAP7_75t_L g2272 ( 
.A1(n_2240),
.A2(n_2080),
.B1(n_2077),
.B2(n_2038),
.Y(n_2272)
);

AOI21xp5_ASAP7_75t_L g2273 ( 
.A1(n_2257),
.A2(n_2016),
.B(n_1741),
.Y(n_2273)
);

NAND5xp2_ASAP7_75t_L g2274 ( 
.A(n_2256),
.B(n_1782),
.C(n_1929),
.D(n_1931),
.E(n_1885),
.Y(n_2274)
);

AOI211xp5_ASAP7_75t_L g2275 ( 
.A1(n_2244),
.A2(n_1860),
.B(n_1923),
.C(n_1985),
.Y(n_2275)
);

AOI221xp5_ASAP7_75t_L g2276 ( 
.A1(n_2239),
.A2(n_2006),
.B1(n_2010),
.B2(n_2009),
.C(n_2008),
.Y(n_2276)
);

AOI22xp5_ASAP7_75t_L g2277 ( 
.A1(n_2239),
.A2(n_2097),
.B1(n_1931),
.B2(n_2098),
.Y(n_2277)
);

NAND5xp2_ASAP7_75t_SL g2278 ( 
.A(n_2245),
.B(n_1923),
.C(n_2049),
.D(n_1725),
.E(n_1860),
.Y(n_2278)
);

NOR2x1_ASAP7_75t_L g2279 ( 
.A(n_2266),
.B(n_1798),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2268),
.Y(n_2280)
);

NOR4xp25_ASAP7_75t_L g2281 ( 
.A(n_2265),
.B(n_2252),
.C(n_1982),
.D(n_1973),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2261),
.Y(n_2282)
);

NAND4xp25_ASAP7_75t_L g2283 ( 
.A(n_2262),
.B(n_1993),
.C(n_1940),
.D(n_1984),
.Y(n_2283)
);

OAI211xp5_ASAP7_75t_L g2284 ( 
.A1(n_2270),
.A2(n_1798),
.B(n_1923),
.C(n_1822),
.Y(n_2284)
);

AOI221xp5_ASAP7_75t_L g2285 ( 
.A1(n_2272),
.A2(n_2072),
.B1(n_2070),
.B2(n_2081),
.C(n_2013),
.Y(n_2285)
);

NOR2xp33_ASAP7_75t_L g2286 ( 
.A(n_2258),
.B(n_1843),
.Y(n_2286)
);

AOI211xp5_ASAP7_75t_L g2287 ( 
.A1(n_2272),
.A2(n_1851),
.B(n_2022),
.C(n_2020),
.Y(n_2287)
);

NOR2x1_ASAP7_75t_L g2288 ( 
.A(n_2267),
.B(n_1998),
.Y(n_2288)
);

NAND3xp33_ASAP7_75t_L g2289 ( 
.A(n_2259),
.B(n_1794),
.C(n_1965),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_2260),
.B(n_2098),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2276),
.B(n_2157),
.Y(n_2291)
);

AOI221xp5_ASAP7_75t_L g2292 ( 
.A1(n_2271),
.A2(n_2082),
.B1(n_2045),
.B2(n_2046),
.C(n_2041),
.Y(n_2292)
);

AOI222xp33_ASAP7_75t_L g2293 ( 
.A1(n_2264),
.A2(n_2048),
.B1(n_2074),
.B2(n_2050),
.C1(n_2073),
.C2(n_1974),
.Y(n_2293)
);

NOR2x1_ASAP7_75t_L g2294 ( 
.A(n_2284),
.B(n_2273),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2286),
.B(n_2277),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2282),
.B(n_2269),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2281),
.B(n_2275),
.Y(n_2297)
);

NAND3xp33_ASAP7_75t_L g2298 ( 
.A(n_2283),
.B(n_2263),
.C(n_1795),
.Y(n_2298)
);

NOR3x1_ASAP7_75t_L g2299 ( 
.A(n_2289),
.B(n_2278),
.C(n_2274),
.Y(n_2299)
);

NOR3xp33_ASAP7_75t_L g2300 ( 
.A(n_2279),
.B(n_1763),
.C(n_1755),
.Y(n_2300)
);

NAND4xp25_ASAP7_75t_L g2301 ( 
.A(n_2293),
.B(n_1958),
.C(n_1984),
.D(n_1940),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_2290),
.B(n_2103),
.Y(n_2302)
);

AND2x2_ASAP7_75t_SL g2303 ( 
.A(n_2285),
.B(n_2085),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2280),
.Y(n_2304)
);

NOR2x1_ASAP7_75t_SL g2305 ( 
.A(n_2291),
.B(n_1999),
.Y(n_2305)
);

NOR3xp33_ASAP7_75t_L g2306 ( 
.A(n_2288),
.B(n_1763),
.C(n_1755),
.Y(n_2306)
);

NAND2x1p5_ASAP7_75t_L g2307 ( 
.A(n_2287),
.B(n_1730),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2304),
.Y(n_2308)
);

OR2x2_ASAP7_75t_L g2309 ( 
.A(n_2296),
.B(n_2157),
.Y(n_2309)
);

NOR2x1_ASAP7_75t_L g2310 ( 
.A(n_2294),
.B(n_2297),
.Y(n_2310)
);

NOR2x1p5_ASAP7_75t_L g2311 ( 
.A(n_2304),
.B(n_2292),
.Y(n_2311)
);

OAI31xp33_ASAP7_75t_SL g2312 ( 
.A1(n_2298),
.A2(n_2000),
.A3(n_1916),
.B(n_1969),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_2295),
.B(n_2159),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2307),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2302),
.B(n_2159),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_2305),
.Y(n_2316)
);

NOR2x1_ASAP7_75t_L g2317 ( 
.A(n_2301),
.B(n_1776),
.Y(n_2317)
);

NAND3xp33_ASAP7_75t_SL g2318 ( 
.A(n_2314),
.B(n_2300),
.C(n_2299),
.Y(n_2318)
);

XNOR2x1_ASAP7_75t_SL g2319 ( 
.A(n_2308),
.B(n_2310),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2313),
.Y(n_2320)
);

OR2x6_ASAP7_75t_L g2321 ( 
.A(n_2316),
.B(n_1858),
.Y(n_2321)
);

OR2x6_ASAP7_75t_L g2322 ( 
.A(n_2317),
.B(n_1858),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2311),
.B(n_2303),
.Y(n_2323)
);

OAI22xp5_ASAP7_75t_L g2324 ( 
.A1(n_2309),
.A2(n_2306),
.B1(n_2086),
.B2(n_2163),
.Y(n_2324)
);

NOR2xp67_ASAP7_75t_SL g2325 ( 
.A(n_2315),
.B(n_1858),
.Y(n_2325)
);

AND2x4_ASAP7_75t_L g2326 ( 
.A(n_2317),
.B(n_1992),
.Y(n_2326)
);

XNOR2xp5_ASAP7_75t_L g2327 ( 
.A(n_2319),
.B(n_2312),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2320),
.Y(n_2328)
);

A2O1A1Ixp33_ASAP7_75t_L g2329 ( 
.A1(n_2323),
.A2(n_1971),
.B(n_1977),
.C(n_1952),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2324),
.Y(n_2330)
);

NOR2xp33_ASAP7_75t_L g2331 ( 
.A(n_2318),
.B(n_2137),
.Y(n_2331)
);

AOI22xp5_ASAP7_75t_L g2332 ( 
.A1(n_2321),
.A2(n_1966),
.B1(n_1968),
.B2(n_1976),
.Y(n_2332)
);

OAI22x1_ASAP7_75t_SL g2333 ( 
.A1(n_2325),
.A2(n_1745),
.B1(n_1968),
.B2(n_1966),
.Y(n_2333)
);

OAI21x1_ASAP7_75t_SL g2334 ( 
.A1(n_2327),
.A2(n_2322),
.B(n_2326),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2328),
.Y(n_2335)
);

OAI22xp5_ASAP7_75t_L g2336 ( 
.A1(n_2331),
.A2(n_2038),
.B1(n_2035),
.B2(n_2137),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2335),
.B(n_2330),
.Y(n_2337)
);

BUFx2_ASAP7_75t_L g2338 ( 
.A(n_2337),
.Y(n_2338)
);

AOI222xp33_ASAP7_75t_L g2339 ( 
.A1(n_2338),
.A2(n_2334),
.B1(n_2333),
.B2(n_2329),
.C1(n_2336),
.C2(n_1776),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2339),
.B(n_2332),
.Y(n_2340)
);

OAI21xp5_ASAP7_75t_L g2341 ( 
.A1(n_2340),
.A2(n_1768),
.B(n_1816),
.Y(n_2341)
);


endmodule