module fake_jpeg_25444_n_271 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_271);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_271;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_3),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_38),
.B(n_41),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_22),
.B(n_18),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_28),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_20),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_47),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_49),
.B(n_2),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_38),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_50),
.B(n_52),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_45),
.B(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_51),
.B(n_58),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_47),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_29),
.B1(n_19),
.B2(n_22),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_53),
.A2(n_64),
.B1(n_72),
.B2(n_32),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_21),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_21),
.Y(n_59)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_19),
.B1(n_29),
.B2(n_33),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_61),
.A2(n_32),
.B1(n_4),
.B2(n_6),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_18),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_65),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_19),
.B1(n_18),
.B2(n_33),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_28),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_34),
.Y(n_66)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_39),
.B(n_20),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_46),
.B(n_44),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_20),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_70),
.Y(n_94)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_23),
.B1(n_26),
.B2(n_24),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_43),
.B(n_35),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_0),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_43),
.A2(n_35),
.B1(n_24),
.B2(n_26),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_75),
.A2(n_23),
.B1(n_17),
.B2(n_27),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_17),
.B(n_1),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_71),
.B(n_30),
.C(n_51),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_77),
.B(n_95),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_78),
.A2(n_87),
.B(n_67),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_83),
.Y(n_117)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_50),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_31),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_90),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_49),
.A2(n_44),
.B1(n_32),
.B2(n_31),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_106),
.Y(n_121)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_97),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_100),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_67),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_102),
.Y(n_128)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_101),
.Y(n_115)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_108),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_67),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_104),
.B(n_105),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_2),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_16),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_111),
.A2(n_95),
.B1(n_105),
.B2(n_93),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_52),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_120),
.C(n_88),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_94),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_69),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_55),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_135),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_107),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_126),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_7),
.B(n_8),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_127),
.A2(n_7),
.B(n_8),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_100),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_130),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_103),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_133),
.Y(n_155)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_55),
.Y(n_135)
);

AOI22x1_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_81),
.B1(n_80),
.B2(n_90),
.Y(n_138)
);

OA22x2_ASAP7_75t_L g174 ( 
.A1(n_138),
.A2(n_116),
.B1(n_69),
.B2(n_112),
.Y(n_174)
);

NOR3xp33_ASAP7_75t_SL g139 ( 
.A(n_137),
.B(n_87),
.C(n_85),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_139),
.B(n_147),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_121),
.A2(n_83),
.B1(n_80),
.B2(n_98),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_140),
.A2(n_145),
.B1(n_151),
.B2(n_161),
.Y(n_168)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_141),
.B(n_142),
.Y(n_166)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_144),
.B(n_148),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_121),
.A2(n_60),
.B1(n_91),
.B2(n_110),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_126),
.B(n_92),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_150),
.B(n_153),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_77),
.B1(n_105),
.B2(n_109),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_158),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_163),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_119),
.B(n_96),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_160),
.B(n_130),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_111),
.A2(n_60),
.B1(n_54),
.B2(n_86),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_60),
.B1(n_54),
.B2(n_57),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_141),
.B1(n_144),
.B2(n_161),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_114),
.B(n_69),
.C(n_16),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_137),
.C(n_158),
.Y(n_175)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_149),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_146),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_167),
.B(n_170),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_155),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_175),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_181),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_120),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_184),
.C(n_190),
.Y(n_194)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_185),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_123),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_182),
.A2(n_113),
.B1(n_124),
.B2(n_9),
.Y(n_200)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_188),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_123),
.C(n_133),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_127),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_187),
.Y(n_210)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_162),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_138),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_139),
.B(n_164),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_132),
.C(n_118),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_188),
.A2(n_138),
.B1(n_148),
.B2(n_153),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_191),
.A2(n_200),
.B1(n_183),
.B2(n_179),
.Y(n_215)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_193),
.Y(n_214)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_198),
.Y(n_219)
);

AOI322xp5_ASAP7_75t_L g198 ( 
.A1(n_173),
.A2(n_159),
.A3(n_151),
.B1(n_145),
.B2(n_154),
.C1(n_112),
.C2(n_134),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_170),
.A2(n_132),
.B(n_118),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_199),
.A2(n_206),
.B1(n_180),
.B2(n_185),
.Y(n_220)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_169),
.Y(n_203)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_203),
.Y(n_212)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_187),
.A2(n_113),
.B1(n_124),
.B2(n_9),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_7),
.C(n_8),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_175),
.C(n_178),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_202),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_210),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_215),
.A2(n_224),
.B1(n_225),
.B2(n_205),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_193),
.Y(n_228)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_199),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_218),
.Y(n_230)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_220),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_208),
.A2(n_168),
.B1(n_176),
.B2(n_174),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_191),
.A2(n_168),
.B1(n_174),
.B2(n_177),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_227),
.Y(n_237)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_231),
.Y(n_242)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_212),
.B(n_195),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_232),
.B(n_227),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_223),
.A2(n_209),
.B1(n_197),
.B2(n_207),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_233),
.A2(n_235),
.B1(n_219),
.B2(n_226),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_194),
.C(n_202),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_238),
.C(n_240),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_174),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_192),
.C(n_211),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_215),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_210),
.C(n_196),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_230),
.A2(n_217),
.B(n_225),
.Y(n_241)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_241),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_243),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_245),
.B(n_247),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_246),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_236),
.B(n_201),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_229),
.A2(n_201),
.B(n_218),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_250),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_238),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_240),
.B(n_10),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_245),
.A2(n_233),
.B1(n_237),
.B2(n_234),
.Y(n_251)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_251),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_256),
.A2(n_254),
.B(n_252),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_260),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_244),
.C(n_242),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_239),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_255),
.Y(n_265)
);

AOI21x1_ASAP7_75t_L g262 ( 
.A1(n_253),
.A2(n_249),
.B(n_244),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_262),
.A2(n_256),
.B(n_11),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_261),
.Y(n_264)
);

O2A1O1Ixp33_ASAP7_75t_SL g267 ( 
.A1(n_264),
.A2(n_265),
.B(n_266),
.C(n_259),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_267),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_263),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_269),
.A2(n_268),
.B(n_11),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_271)
);


endmodule