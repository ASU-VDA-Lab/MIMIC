module fake_jpeg_19461_n_318 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_318);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_10),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx2_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_11),
.B(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_35),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g34 ( 
.A(n_14),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_35),
.B1(n_32),
.B2(n_25),
.Y(n_41)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_36),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_47),
.B1(n_34),
.B2(n_30),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_22),
.B1(n_20),
.B2(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_55),
.Y(n_71)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_47),
.A2(n_25),
.B1(n_34),
.B2(n_35),
.Y(n_51)
);

AO22x1_ASAP7_75t_SL g78 ( 
.A1(n_51),
.A2(n_54),
.B1(n_32),
.B2(n_41),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_52),
.B(n_57),
.Y(n_69)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_47),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_46),
.B(n_11),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_59),
.Y(n_73)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_60),
.Y(n_67)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_61),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_54),
.A2(n_34),
.B1(n_40),
.B2(n_35),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_63),
.A2(n_72),
.B1(n_78),
.B2(n_39),
.Y(n_88)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_54),
.A2(n_34),
.B1(n_40),
.B2(n_32),
.Y(n_72)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_46),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_42),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_52),
.C(n_54),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_85),
.C(n_90),
.Y(n_118)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_95),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_69),
.B(n_57),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_87),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_84),
.B(n_90),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_54),
.C(n_38),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

OAI32xp33_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_38),
.A3(n_39),
.B1(n_30),
.B2(n_20),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_78),
.B1(n_76),
.B2(n_61),
.Y(n_104)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_89),
.A2(n_65),
.B1(n_64),
.B2(n_75),
.Y(n_116)
);

FAx1_ASAP7_75t_SL g90 ( 
.A(n_71),
.B(n_25),
.CI(n_40),
.CON(n_90),
.SN(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_22),
.B(n_60),
.C(n_59),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_93),
.Y(n_99)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_70),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_63),
.B1(n_72),
.B2(n_78),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_106),
.B1(n_90),
.B2(n_65),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_78),
.B(n_70),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_101),
.A2(n_103),
.B(n_107),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_79),
.A2(n_69),
.B(n_70),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_104),
.A2(n_112),
.B1(n_65),
.B2(n_89),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_80),
.A2(n_78),
.B1(n_43),
.B2(n_49),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_66),
.B(n_67),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_92),
.A2(n_66),
.B(n_67),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_108),
.A2(n_27),
.B(n_45),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_93),
.B(n_22),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_27),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_86),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_119),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_43),
.B1(n_49),
.B2(n_65),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_67),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_114),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_83),
.B(n_75),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_53),
.B1(n_96),
.B2(n_28),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_118),
.B(n_27),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_74),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_89),
.Y(n_121)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_121),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_90),
.C(n_92),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_143),
.C(n_147),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_123),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_124),
.A2(n_131),
.B1(n_141),
.B2(n_102),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_129),
.B1(n_130),
.B2(n_137),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_111),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_127),
.B(n_138),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_101),
.A2(n_43),
.B1(n_82),
.B2(n_91),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_104),
.A2(n_91),
.B1(n_64),
.B2(n_75),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_68),
.B1(n_58),
.B2(n_56),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_119),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_139),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_96),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_134),
.A2(n_0),
.B(n_1),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_28),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_150),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_99),
.A2(n_28),
.B1(n_96),
.B2(n_20),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_11),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_100),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_98),
.A2(n_44),
.B1(n_26),
.B2(n_29),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_97),
.B(n_16),
.Y(n_142)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_27),
.C(n_45),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_99),
.A2(n_44),
.B1(n_23),
.B2(n_24),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_110),
.B1(n_117),
.B2(n_120),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_115),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_21),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_138),
.A2(n_108),
.B1(n_105),
.B2(n_114),
.Y(n_153)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_109),
.C(n_105),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_164),
.C(n_146),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_135),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_157),
.B(n_171),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_158),
.B(n_131),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_128),
.A2(n_117),
.B1(n_102),
.B2(n_115),
.Y(n_159)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_159),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_162),
.A2(n_163),
.B1(n_166),
.B2(n_173),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_125),
.A2(n_109),
.B1(n_44),
.B2(n_36),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_122),
.C(n_143),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_130),
.A2(n_31),
.B1(n_36),
.B2(n_29),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_167),
.Y(n_188)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_126),
.Y(n_171)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_124),
.A2(n_23),
.B1(n_21),
.B2(n_18),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_176),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_165),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_185),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_128),
.Y(n_183)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_174),
.B(n_161),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_175),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_195),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_190),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_154),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_129),
.B1(n_140),
.B2(n_145),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_191),
.A2(n_196),
.B1(n_187),
.B2(n_197),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_146),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_198),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_150),
.C(n_127),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_204),
.C(n_189),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_170),
.A2(n_144),
.B(n_139),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_180),
.A2(n_134),
.B1(n_137),
.B2(n_141),
.Y(n_196)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_167),
.A2(n_179),
.B(n_152),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_152),
.B(n_126),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_199),
.A2(n_169),
.B(n_165),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_201),
.B(n_203),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_149),
.C(n_45),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_201),
.A2(n_184),
.B1(n_206),
.B2(n_177),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_207),
.A2(n_214),
.B1(n_222),
.B2(n_227),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_202),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_211),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_188),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_199),
.A2(n_177),
.B1(n_160),
.B2(n_173),
.Y(n_214)
);

FAx1_ASAP7_75t_SL g216 ( 
.A(n_193),
.B(n_155),
.CI(n_163),
.CON(n_216),
.SN(n_216)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_225),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_156),
.C(n_166),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_31),
.C(n_29),
.Y(n_246)
);

OA21x2_ASAP7_75t_L g221 ( 
.A1(n_200),
.A2(n_160),
.B(n_178),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_230),
.B1(n_10),
.B2(n_9),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_199),
.A2(n_156),
.B1(n_123),
.B2(n_2),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_224),
.A2(n_228),
.B1(n_209),
.B2(n_221),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_27),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_226),
.B(n_205),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_187),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_191),
.A2(n_23),
.B1(n_21),
.B2(n_18),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_27),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_36),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_181),
.A2(n_18),
.B1(n_19),
.B2(n_24),
.Y(n_230)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_215),
.B(n_196),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_244),
.Y(n_255)
);

FAx1_ASAP7_75t_SL g237 ( 
.A(n_215),
.B(n_203),
.CI(n_182),
.CON(n_237),
.SN(n_237)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_243),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_227),
.A2(n_213),
.B1(n_222),
.B2(n_220),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_238),
.A2(n_241),
.B1(n_242),
.B2(n_9),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_208),
.A2(n_192),
.B(n_19),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_239),
.A2(n_236),
.B(n_242),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_218),
.A2(n_214),
.B1(n_212),
.B2(n_207),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_221),
.A2(n_19),
.B1(n_45),
.B2(n_12),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_217),
.A2(n_12),
.B1(n_15),
.B2(n_16),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_247),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_246),
.B(n_249),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_16),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_9),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_31),
.C(n_29),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_225),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_16),
.Y(n_256)
);

OAI221xp5_ASAP7_75t_L g251 ( 
.A1(n_244),
.A2(n_219),
.B1(n_216),
.B2(n_229),
.C(n_228),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_251),
.A2(n_1),
.B(n_3),
.Y(n_280)
);

FAx1_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_224),
.CI(n_31),
.CON(n_252),
.SN(n_252)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_262),
.Y(n_271)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_253),
.B(n_259),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_246),
.Y(n_254)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_254),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_245),
.Y(n_273)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_15),
.Y(n_259)
);

INVxp67_ASAP7_75t_SL g260 ( 
.A(n_243),
.Y(n_260)
);

INVx11_ASAP7_75t_L g268 ( 
.A(n_260),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_233),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_247),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_266),
.B(n_237),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_269),
.A2(n_274),
.B(n_276),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_26),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_232),
.B(n_250),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_275),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_258),
.A2(n_234),
.B(n_249),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_12),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_26),
.C(n_17),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_15),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_252),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_279),
.A2(n_280),
.B1(n_3),
.B2(n_4),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_261),
.C(n_255),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_282),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_253),
.C(n_254),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_252),
.Y(n_283)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_283),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_287),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_26),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_291),
.C(n_292),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_290),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_12),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_12),
.Y(n_292)
);

AOI21x1_ASAP7_75t_L g293 ( 
.A1(n_268),
.A2(n_3),
.B(n_4),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_293),
.A2(n_272),
.B1(n_5),
.B2(n_6),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_278),
.C(n_279),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_301),
.Y(n_306)
);

AOI21xp33_ASAP7_75t_L g304 ( 
.A1(n_300),
.A2(n_303),
.B(n_4),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_289),
.A2(n_268),
.B1(n_17),
.B2(n_13),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_17),
.C(n_14),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_5),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_283),
.A2(n_288),
.B(n_292),
.Y(n_303)
);

AO21x1_ASAP7_75t_L g311 ( 
.A1(n_304),
.A2(n_307),
.B(n_308),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_17),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_295),
.C(n_296),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_297),
.A2(n_14),
.B(n_6),
.Y(n_307)
);

AOI21xp33_ASAP7_75t_L g309 ( 
.A1(n_306),
.A2(n_295),
.B(n_298),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_309),
.A2(n_300),
.B(n_6),
.Y(n_312)
);

AO221x1_ASAP7_75t_L g313 ( 
.A1(n_310),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_313),
.C(n_311),
.Y(n_314)
);

MAJx2_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_5),
.C(n_7),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_7),
.C(n_8),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_8),
.C(n_314),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_8),
.Y(n_318)
);


endmodule