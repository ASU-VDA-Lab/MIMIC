module real_jpeg_32721_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_0),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_0),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_1),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_1),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_1),
.B(n_308),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_1),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_1),
.B(n_396),
.Y(n_395)
);

AND2x2_ASAP7_75t_SL g436 ( 
.A(n_1),
.B(n_437),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_2),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_2),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_2),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_2),
.B(n_43),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_2),
.B(n_103),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_2),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_2),
.B(n_100),
.Y(n_154)
);

AND2x4_ASAP7_75t_SL g184 ( 
.A(n_2),
.B(n_185),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_3),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_3),
.B(n_116),
.Y(n_115)
);

AND2x4_ASAP7_75t_L g140 ( 
.A(n_3),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_3),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_3),
.B(n_172),
.Y(n_171)
);

NAND2xp33_ASAP7_75t_R g219 ( 
.A(n_3),
.B(n_220),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_4),
.A2(n_19),
.B(n_482),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_4),
.B(n_483),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_5),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_5),
.B(n_132),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_5),
.A2(n_216),
.B(n_218),
.Y(n_215)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_5),
.Y(n_279)
);

NAND2x1_ASAP7_75t_SL g310 ( 
.A(n_5),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_5),
.B(n_216),
.Y(n_338)
);

AND2x2_ASAP7_75t_SL g419 ( 
.A(n_5),
.B(n_420),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_5),
.B(n_449),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_6),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_6),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_7),
.Y(n_278)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_8),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_8),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_9),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_9),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_9),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_9),
.B(n_179),
.Y(n_178)
);

AND2x2_ASAP7_75t_SL g226 ( 
.A(n_9),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_9),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_9),
.B(n_270),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_10),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_10),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_10),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_12),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_12),
.B(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g229 ( 
.A(n_12),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_12),
.B(n_98),
.Y(n_239)
);

AND2x2_ASAP7_75t_SL g280 ( 
.A(n_12),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_12),
.B(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_12),
.B(n_374),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_12),
.B(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_13),
.Y(n_106)
);

INVx4_ASAP7_75t_L g403 ( 
.A(n_13),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_14),
.B(n_43),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_14),
.B(n_172),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_14),
.B(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_14),
.B(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_14),
.B(n_440),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_14),
.B(n_453),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_14),
.B(n_458),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_15),
.Y(n_483)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_16),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_16),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_17),
.B(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_17),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_17),
.B(n_58),
.Y(n_70)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_17),
.B(n_82),
.Y(n_81)
);

AND2x4_ASAP7_75t_SL g110 ( 
.A(n_17),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_17),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_17),
.B(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_17),
.B(n_43),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_191),
.Y(n_19)
);

NAND2xp33_ASAP7_75t_R g20 ( 
.A(n_21),
.B(n_190),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_160),
.Y(n_21)
);

NAND2x1p5_ASAP7_75t_L g190 ( 
.A(n_22),
.B(n_160),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_93),
.C(n_119),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_24),
.B(n_94),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_66),
.Y(n_24)
);

INVxp33_ASAP7_75t_L g162 ( 
.A(n_25),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_40),
.C(n_50),
.Y(n_25)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_26),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_36),
.B2(n_39),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_33),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

MAJx2_ASAP7_75t_L g86 ( 
.A(n_30),
.B(n_36),
.C(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_32),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_32),
.Y(n_132)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_32),
.Y(n_181)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_33),
.B(n_96),
.Y(n_95)
);

XOR2x2_ASAP7_75t_L g365 ( 
.A(n_33),
.B(n_147),
.Y(n_365)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_35),
.Y(n_228)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_35),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_35),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_36),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_46),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_36),
.B(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_36),
.A2(n_39),
.B1(n_373),
.B2(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_38),
.Y(n_148)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_38),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_39),
.B(n_373),
.Y(n_372)
);

XOR2x1_ASAP7_75t_L g208 ( 
.A(n_40),
.B(n_50),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_45),
.B(n_49),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_41),
.A2(n_42),
.B1(n_46),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_46),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_46),
.B(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_46),
.A2(n_136),
.B1(n_268),
.B2(n_269),
.Y(n_304)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_49),
.Y(n_330)
);

XNOR2x1_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_51),
.A2(n_118),
.B1(n_236),
.B2(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22x1_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_60),
.B1(n_64),
.B2(n_65),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_55),
.Y(n_64)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_59),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_60),
.Y(n_65)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_63),
.Y(n_185)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_63),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_65),
.C(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_85),
.B1(n_91),
.B2(n_92),
.Y(n_66)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_77),
.C(n_80),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_68),
.B(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_71),
.C(n_75),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_69),
.A2(n_70),
.B1(n_75),
.B2(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_69),
.A2(n_70),
.B1(n_171),
.B2(n_174),
.Y(n_170)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVxp67_ASAP7_75t_SL g123 ( 
.A(n_71),
.Y(n_123)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx5_ASAP7_75t_L g442 ( 
.A(n_73),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_76),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_77),
.A2(n_80),
.B1(n_81),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_77),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_80),
.A2(n_81),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_80),
.B(n_86),
.C(n_90),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_82),
.Y(n_173)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_84),
.Y(n_217)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_87),
.B(n_102),
.C(n_107),
.Y(n_189)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_91),
.B(n_162),
.C(n_163),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_92),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_108),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_95),
.B(n_109),
.C(n_117),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_101),
.B1(n_102),
.B2(n_107),
.Y(n_96)
);

INVxp67_ASAP7_75t_SL g107 ( 
.A(n_97),
.Y(n_107)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_100),
.Y(n_329)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_101),
.A2(n_102),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_101),
.A2(n_102),
.B1(n_274),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

MAJx2_ASAP7_75t_L g273 ( 
.A(n_102),
.B(n_274),
.C(n_280),
.Y(n_273)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_106),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_117),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_110),
.B(n_113),
.C(n_188),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_113),
.A2(n_133),
.B1(n_289),
.B2(n_291),
.Y(n_288)
);

INVxp33_ASAP7_75t_L g188 ( 
.A(n_115),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_118),
.B(n_183),
.C(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_119),
.B(n_196),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_137),
.C(n_155),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_120),
.A2(n_121),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.C(n_134),
.Y(n_121)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_122),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_126),
.B(n_134),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.C(n_133),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_127),
.A2(n_128),
.B1(n_131),
.B2(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_131),
.Y(n_290)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_132),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_137),
.A2(n_156),
.B1(n_157),
.B2(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_137),
.Y(n_203)
);

MAJx2_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_149),
.C(n_153),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_138),
.A2(n_139),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.C(n_147),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_140),
.B(n_143),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_147),
.B(n_213),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_148),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_149),
.A2(n_150),
.B1(n_153),
.B2(n_154),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_150),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_151),
.Y(n_238)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_152),
.Y(n_437)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_176),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_175),
.Y(n_169)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_171),
.Y(n_174)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_186),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_182),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_183),
.B(n_334),
.Y(n_333)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);

OA21x2_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_292),
.B(n_473),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_244),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

INVxp33_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_195),
.B(n_198),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_195),
.B(n_198),
.Y(n_481)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_204),
.C(n_209),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_200),
.A2(n_205),
.B1(n_206),
.B2(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_200),
.Y(n_248)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_247),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_209),
.B(n_247),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_232),
.C(n_240),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_211),
.B(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_214),
.C(n_221),
.Y(n_211)
);

XNOR2x1_ASAP7_75t_L g346 ( 
.A(n_212),
.B(n_347),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_214),
.A2(n_215),
.B1(n_221),
.B2(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NOR2xp67_ASAP7_75t_SL g336 ( 
.A(n_215),
.B(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_219),
.B(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_221),
.Y(n_348)
);

MAJx2_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_226),
.C(n_229),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_222),
.A2(n_223),
.B1(n_226),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_226),
.Y(n_265)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_264),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_231),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_241),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.C(n_239),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_235),
.Y(n_287)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_236),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_237),
.B(n_239),
.Y(n_286)
);

INVxp33_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_242),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_245),
.A2(n_475),
.B(n_481),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_249),
.B(n_250),
.Y(n_245)
);

NAND3xp33_ASAP7_75t_L g476 ( 
.A(n_246),
.B(n_249),
.C(n_250),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_256),
.C(n_260),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_253),
.A2(n_254),
.B1(n_257),
.B2(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVxp67_ASAP7_75t_SL g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_257),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_261),
.B(n_353),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_285),
.C(n_288),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_262),
.B(n_342),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_266),
.C(n_273),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_263),
.B(n_298),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_266),
.A2(n_267),
.B1(n_273),
.B2(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_272),
.Y(n_461)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_273),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_274),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_279),
.Y(n_274)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_278),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_279),
.B(n_400),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_280),
.B(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_285),
.B(n_288),
.Y(n_342)
);

XOR2x2_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_289),
.Y(n_291)
);

NAND3xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_349),
.C(n_355),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_340),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_294),
.B(n_340),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_300),
.C(n_316),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_296),
.A2(n_297),
.B1(n_318),
.B2(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_300),
.B(n_358),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g360 ( 
.A(n_300),
.B(n_358),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_304),
.C(n_305),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_301),
.B(n_363),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_304),
.B(n_306),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_310),
.C(n_315),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_307),
.B(n_310),
.Y(n_406)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx3_ASAP7_75t_SL g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_315),
.B(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_318),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_331),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_319),
.B(n_336),
.C(n_345),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_324),
.C(n_330),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_320),
.A2(n_321),
.B1(n_324),
.B2(n_325),
.Y(n_379)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_326),
.B(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_330),
.B(n_379),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_333),
.B1(n_336),
.B2(n_339),
.Y(n_331)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_332),
.Y(n_345)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_336),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_343),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_341),
.B(n_344),
.C(n_346),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_346),
.Y(n_343)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_350),
.A2(n_478),
.B(n_479),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g479 ( 
.A(n_351),
.B(n_352),
.Y(n_479)
);

OAI21x1_ASAP7_75t_SL g355 ( 
.A1(n_356),
.A2(n_380),
.B(n_472),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_360),
.B(n_361),
.Y(n_356)
);

NAND3xp33_ASAP7_75t_L g472 ( 
.A(n_357),
.B(n_360),
.C(n_361),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_364),
.C(n_377),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_362),
.B(n_408),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_364),
.B(n_378),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.C(n_372),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_365),
.A2(n_366),
.B1(n_367),
.B2(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_365),
.Y(n_386)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_372),
.B(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_373),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_409),
.B(n_471),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_407),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_382),
.B(n_407),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_387),
.C(n_404),
.Y(n_382)
);

INVxp33_ASAP7_75t_SL g383 ( 
.A(n_384),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_384),
.B(n_427),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_387),
.A2(n_388),
.B1(n_405),
.B2(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_394),
.C(n_399),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_389),
.A2(n_390),
.B1(n_394),
.B2(n_395),
.Y(n_414)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_399),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_402),
.Y(n_454)
);

INVx4_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_405),
.Y(n_428)
);

OAI21x1_ASAP7_75t_SL g409 ( 
.A1(n_410),
.A2(n_429),
.B(n_470),
.Y(n_409)
);

NOR2xp67_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_426),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_411),
.B(n_426),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_415),
.C(n_418),
.Y(n_411)
);

XNOR2x2_ASAP7_75t_L g466 ( 
.A(n_412),
.B(n_467),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_414),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_415),
.A2(n_416),
.B1(n_418),
.B2(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_418),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_423),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_419),
.B(n_423),
.Y(n_433)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

AOI21x1_ASAP7_75t_L g429 ( 
.A1(n_430),
.A2(n_464),
.B(n_469),
.Y(n_429)
);

OAI21x1_ASAP7_75t_L g430 ( 
.A1(n_431),
.A2(n_450),
.B(n_463),
.Y(n_430)
);

NOR2x1_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_443),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_432),
.B(n_443),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_434),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_433),
.B(n_436),
.C(n_438),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_435),
.A2(n_436),
.B1(n_438),
.B2(n_439),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_448),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_444),
.B(n_448),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_444),
.B(n_457),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx4_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_451),
.A2(n_456),
.B(n_462),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_455),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_452),
.B(n_455),
.Y(n_462)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_466),
.Y(n_464)
);

NOR2xp67_ASAP7_75t_L g469 ( 
.A(n_465),
.B(n_466),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_474),
.A2(n_477),
.B(n_480),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_476),
.Y(n_474)
);


endmodule