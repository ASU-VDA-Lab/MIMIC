module fake_aes_12647_n_653 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_653);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_653;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_466;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g85 ( .A(n_57), .Y(n_85) );
BUFx10_ASAP7_75t_L g86 ( .A(n_64), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_14), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_34), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_31), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_82), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_73), .Y(n_91) );
BUFx2_ASAP7_75t_L g92 ( .A(n_49), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_58), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_79), .Y(n_94) );
BUFx6f_ASAP7_75t_L g95 ( .A(n_74), .Y(n_95) );
INVx1_ASAP7_75t_SL g96 ( .A(n_81), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_42), .Y(n_97) );
BUFx5_ASAP7_75t_L g98 ( .A(n_19), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_54), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_60), .Y(n_100) );
INVx1_ASAP7_75t_SL g101 ( .A(n_8), .Y(n_101) );
BUFx6f_ASAP7_75t_L g102 ( .A(n_66), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_76), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_25), .B(n_63), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_72), .Y(n_105) );
BUFx10_ASAP7_75t_L g106 ( .A(n_46), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_53), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_40), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_32), .Y(n_109) );
INVx1_ASAP7_75t_SL g110 ( .A(n_28), .Y(n_110) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_61), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_52), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_24), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_44), .Y(n_114) );
INVxp67_ASAP7_75t_L g115 ( .A(n_62), .Y(n_115) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_77), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_80), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_29), .Y(n_118) );
INVxp33_ASAP7_75t_SL g119 ( .A(n_22), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_27), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_13), .Y(n_121) );
BUFx2_ASAP7_75t_L g122 ( .A(n_48), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_14), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_70), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_26), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_2), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_67), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_43), .Y(n_128) );
BUFx12f_ASAP7_75t_L g129 ( .A(n_86), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_98), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_98), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_98), .Y(n_132) );
HB1xp67_ASAP7_75t_L g133 ( .A(n_121), .Y(n_133) );
AND2x4_ASAP7_75t_L g134 ( .A(n_126), .B(n_0), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_92), .B(n_0), .Y(n_135) );
BUFx8_ASAP7_75t_L g136 ( .A(n_122), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_98), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_116), .Y(n_138) );
INVx6_ASAP7_75t_L g139 ( .A(n_86), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_86), .B(n_1), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_95), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_98), .Y(n_142) );
BUFx2_ASAP7_75t_L g143 ( .A(n_98), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_95), .Y(n_144) );
BUFx2_ASAP7_75t_L g145 ( .A(n_98), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_87), .B(n_1), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_95), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_85), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_134), .Y(n_149) );
OAI22xp33_ASAP7_75t_SL g150 ( .A1(n_140), .A2(n_119), .B1(n_101), .B2(n_123), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_141), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_141), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_139), .B(n_115), .Y(n_153) );
AOI22xp33_ASAP7_75t_L g154 ( .A1(n_134), .A2(n_126), .B1(n_119), .B2(n_112), .Y(n_154) );
BUFx10_ASAP7_75t_L g155 ( .A(n_139), .Y(n_155) );
AO22x2_ASAP7_75t_L g156 ( .A1(n_134), .A2(n_85), .B1(n_125), .B2(n_118), .Y(n_156) );
AOI22xp5_ASAP7_75t_L g157 ( .A1(n_135), .A2(n_88), .B1(n_94), .B2(n_124), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_134), .B(n_89), .Y(n_158) );
NAND3xp33_ASAP7_75t_L g159 ( .A(n_135), .B(n_88), .C(n_94), .Y(n_159) );
BUFx10_ASAP7_75t_L g160 ( .A(n_139), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_141), .Y(n_161) );
BUFx2_ASAP7_75t_L g162 ( .A(n_136), .Y(n_162) );
BUFx4f_ASAP7_75t_L g163 ( .A(n_143), .Y(n_163) );
BUFx3_ASAP7_75t_L g164 ( .A(n_143), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_133), .B(n_106), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_129), .B(n_106), .Y(n_166) );
AND2x4_ASAP7_75t_L g167 ( .A(n_145), .B(n_90), .Y(n_167) );
OR2x2_ASAP7_75t_L g168 ( .A(n_138), .B(n_108), .Y(n_168) );
INVx5_ASAP7_75t_L g169 ( .A(n_141), .Y(n_169) );
INVx2_ASAP7_75t_SL g170 ( .A(n_139), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_141), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_130), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_130), .Y(n_173) );
OR2x2_ASAP7_75t_L g174 ( .A(n_146), .B(n_108), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_137), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_141), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_137), .Y(n_177) );
INVx3_ASAP7_75t_L g178 ( .A(n_148), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_172), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_163), .B(n_136), .Y(n_180) );
INVx2_ASAP7_75t_SL g181 ( .A(n_156), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_163), .B(n_136), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_156), .A2(n_167), .B1(n_158), .B2(n_149), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_167), .B(n_145), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_149), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_163), .B(n_136), .Y(n_186) );
OR2x6_ASAP7_75t_L g187 ( .A(n_162), .B(n_129), .Y(n_187) );
AND2x6_ASAP7_75t_SL g188 ( .A(n_165), .B(n_91), .Y(n_188) );
BUFx8_ASAP7_75t_L g189 ( .A(n_162), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_149), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_172), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_167), .B(n_114), .Y(n_192) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_174), .Y(n_193) );
AND2x4_ASAP7_75t_L g194 ( .A(n_167), .B(n_148), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_174), .B(n_114), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_156), .A2(n_131), .B1(n_132), .B2(n_142), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_173), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_165), .B(n_106), .Y(n_198) );
OR2x4_ASAP7_75t_L g199 ( .A(n_168), .B(n_93), .Y(n_199) );
BUFx3_ASAP7_75t_L g200 ( .A(n_164), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_173), .Y(n_201) );
AND2x6_ASAP7_75t_SL g202 ( .A(n_153), .B(n_97), .Y(n_202) );
OR2x2_ASAP7_75t_L g203 ( .A(n_157), .B(n_120), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_163), .B(n_120), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_168), .B(n_124), .Y(n_205) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_156), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_175), .Y(n_207) );
AND2x4_ASAP7_75t_SL g208 ( .A(n_155), .B(n_100), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_164), .B(n_131), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_164), .B(n_132), .Y(n_210) );
INVx2_ASAP7_75t_SL g211 ( .A(n_156), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_158), .A2(n_142), .B(n_117), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_155), .B(n_99), .Y(n_213) );
INVx2_ASAP7_75t_SL g214 ( .A(n_155), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_158), .B(n_103), .Y(n_215) );
OAI22xp5_ASAP7_75t_SL g216 ( .A1(n_154), .A2(n_109), .B1(n_113), .B2(n_128), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_155), .B(n_127), .Y(n_217) );
OR2x2_ASAP7_75t_L g218 ( .A(n_159), .B(n_2), .Y(n_218) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_183), .A2(n_149), .B(n_158), .C(n_178), .Y(n_219) );
BUFx2_ASAP7_75t_L g220 ( .A(n_189), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_193), .B(n_150), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_189), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_SL g223 ( .A1(n_181), .A2(n_177), .B(n_175), .C(n_170), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_183), .B(n_200), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_209), .A2(n_177), .B(n_170), .Y(n_225) );
OAI321xp33_ASAP7_75t_L g226 ( .A1(n_216), .A2(n_107), .A3(n_105), .B1(n_147), .B2(n_144), .C(n_95), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_198), .A2(n_166), .B1(n_160), .B2(n_178), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_206), .A2(n_178), .B(n_96), .C(n_110), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_200), .Y(n_229) );
INVx3_ASAP7_75t_L g230 ( .A(n_179), .Y(n_230) );
NAND2x1p5_ASAP7_75t_L g231 ( .A(n_181), .B(n_178), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_212), .A2(n_210), .B(n_185), .Y(n_232) );
OAI22xp33_ASAP7_75t_L g233 ( .A1(n_187), .A2(n_160), .B1(n_111), .B2(n_102), .Y(n_233) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_185), .A2(n_104), .B(n_102), .C(n_111), .Y(n_234) );
OAI21x1_ASAP7_75t_L g235 ( .A1(n_190), .A2(n_176), .B(n_171), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_184), .B(n_160), .Y(n_236) );
OAI21xp5_ASAP7_75t_L g237 ( .A1(n_190), .A2(n_176), .B(n_171), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_211), .B(n_160), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_194), .B(n_3), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_192), .A2(n_176), .B(n_171), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_194), .B(n_3), .Y(n_241) );
AOI21x1_ASAP7_75t_L g242 ( .A1(n_204), .A2(n_161), .B(n_152), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_211), .A2(n_161), .B(n_152), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_194), .B(n_4), .Y(n_244) );
OAI21xp5_ASAP7_75t_L g245 ( .A1(n_179), .A2(n_161), .B(n_152), .Y(n_245) );
OR2x2_ASAP7_75t_L g246 ( .A(n_203), .B(n_4), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_215), .A2(n_151), .B(n_169), .Y(n_247) );
OA22x2_ASAP7_75t_L g248 ( .A1(n_216), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_198), .B(n_5), .Y(n_249) );
INVx5_ASAP7_75t_L g250 ( .A(n_187), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_195), .A2(n_151), .B(n_169), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_203), .B(n_6), .Y(n_252) );
OAI21xp5_ASAP7_75t_L g253 ( .A1(n_191), .A2(n_151), .B(n_169), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_232), .A2(n_191), .B(n_197), .Y(n_254) );
AO21x1_ASAP7_75t_L g255 ( .A1(n_228), .A2(n_218), .B(n_180), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_232), .A2(n_207), .B(n_201), .Y(n_256) );
AO31x2_ASAP7_75t_L g257 ( .A1(n_234), .A2(n_197), .A3(n_207), .B(n_201), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_239), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_243), .A2(n_196), .B(n_182), .Y(n_259) );
OAI21x1_ASAP7_75t_L g260 ( .A1(n_235), .A2(n_186), .B(n_217), .Y(n_260) );
OR2x6_ASAP7_75t_L g261 ( .A(n_220), .B(n_187), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_243), .A2(n_240), .B(n_223), .Y(n_262) );
OR2x2_ASAP7_75t_L g263 ( .A(n_246), .B(n_187), .Y(n_263) );
INVx1_ASAP7_75t_SL g264 ( .A(n_222), .Y(n_264) );
OAI21x1_ASAP7_75t_L g265 ( .A1(n_242), .A2(n_213), .B(n_218), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_SL g266 ( .A1(n_233), .A2(n_214), .B(n_205), .C(n_199), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_225), .A2(n_199), .B(n_214), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_241), .Y(n_268) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_250), .Y(n_269) );
BUFx2_ASAP7_75t_L g270 ( .A(n_250), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_230), .Y(n_271) );
OA21x2_ASAP7_75t_L g272 ( .A1(n_245), .A2(n_199), .B(n_102), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_251), .A2(n_208), .B(n_169), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_252), .A2(n_189), .B1(n_208), .B2(n_188), .Y(n_274) );
O2A1O1Ixp5_ASAP7_75t_L g275 ( .A1(n_238), .A2(n_202), .B(n_188), .C(n_111), .Y(n_275) );
A2O1A1Ixp33_ASAP7_75t_L g276 ( .A1(n_219), .A2(n_202), .B(n_111), .C(n_102), .Y(n_276) );
OAI22x1_ASAP7_75t_L g277 ( .A1(n_250), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_277) );
OAI21xp5_ASAP7_75t_L g278 ( .A1(n_247), .A2(n_169), .B(n_147), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_258), .B(n_224), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g280 ( .A1(n_268), .A2(n_248), .B1(n_221), .B2(n_249), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_271), .Y(n_281) );
AND2x4_ASAP7_75t_L g282 ( .A(n_270), .B(n_250), .Y(n_282) );
OAI21x1_ASAP7_75t_L g283 ( .A1(n_262), .A2(n_237), .B(n_253), .Y(n_283) );
AO31x2_ASAP7_75t_L g284 ( .A1(n_254), .A2(n_244), .A3(n_226), .B(n_248), .Y(n_284) );
AO31x2_ASAP7_75t_L g285 ( .A1(n_254), .A2(n_236), .A3(n_147), .B(n_144), .Y(n_285) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_269), .Y(n_286) );
OAI21xp5_ASAP7_75t_SL g287 ( .A1(n_274), .A2(n_263), .B(n_276), .Y(n_287) );
AO21x2_ASAP7_75t_L g288 ( .A1(n_262), .A2(n_227), .B(n_147), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_267), .B(n_230), .Y(n_289) );
BUFx2_ASAP7_75t_L g290 ( .A(n_261), .Y(n_290) );
AO21x2_ASAP7_75t_L g291 ( .A1(n_256), .A2(n_147), .B(n_144), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_272), .B(n_231), .Y(n_292) );
A2O1A1Ixp33_ASAP7_75t_L g293 ( .A1(n_267), .A2(n_229), .B(n_147), .C(n_144), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_261), .B(n_229), .Y(n_294) );
OA21x2_ASAP7_75t_L g295 ( .A1(n_256), .A2(n_144), .B(n_231), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_257), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_272), .B(n_229), .Y(n_297) );
INVx2_ASAP7_75t_SL g298 ( .A(n_261), .Y(n_298) );
INVx4_ASAP7_75t_SL g299 ( .A(n_257), .Y(n_299) );
AO21x2_ASAP7_75t_L g300 ( .A1(n_259), .A2(n_144), .B(n_10), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_259), .B(n_9), .Y(n_301) );
AOI21x1_ASAP7_75t_L g302 ( .A1(n_301), .A2(n_255), .B(n_265), .Y(n_302) );
BUFx8_ASAP7_75t_L g303 ( .A(n_290), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_296), .Y(n_304) );
OA21x2_ASAP7_75t_L g305 ( .A1(n_293), .A2(n_278), .B(n_260), .Y(n_305) );
BUFx2_ASAP7_75t_L g306 ( .A(n_295), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_296), .B(n_257), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_291), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_280), .B(n_277), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_285), .Y(n_310) );
OA21x2_ASAP7_75t_L g311 ( .A1(n_293), .A2(n_273), .B(n_275), .Y(n_311) );
INVx3_ASAP7_75t_L g312 ( .A(n_295), .Y(n_312) );
AO21x2_ASAP7_75t_L g313 ( .A1(n_301), .A2(n_266), .B(n_273), .Y(n_313) );
BUFx3_ASAP7_75t_L g314 ( .A(n_295), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_285), .Y(n_315) );
AO21x2_ASAP7_75t_L g316 ( .A1(n_300), .A2(n_10), .B(n_11), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_291), .Y(n_317) );
INVx3_ASAP7_75t_L g318 ( .A(n_295), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_285), .Y(n_319) );
AO21x2_ASAP7_75t_L g320 ( .A1(n_300), .A2(n_11), .B(n_12), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_285), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_285), .Y(n_322) );
BUFx2_ASAP7_75t_L g323 ( .A(n_295), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_285), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_280), .B(n_12), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_285), .Y(n_326) );
INVxp33_ASAP7_75t_L g327 ( .A(n_286), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_289), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_292), .B(n_13), .Y(n_329) );
OR2x6_ASAP7_75t_L g330 ( .A(n_292), .B(n_289), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_304), .Y(n_331) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_314), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_330), .B(n_299), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_308), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_309), .B(n_279), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_308), .Y(n_336) );
AO21x2_ASAP7_75t_L g337 ( .A1(n_310), .A2(n_300), .B(n_291), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_304), .B(n_300), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_304), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_309), .B(n_279), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_306), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_310), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_330), .B(n_299), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_310), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_330), .B(n_299), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_315), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_330), .B(n_287), .Y(n_347) );
AO21x2_ASAP7_75t_L g348 ( .A1(n_315), .A2(n_291), .B(n_288), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_315), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_303), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_330), .B(n_287), .Y(n_351) );
INVx3_ASAP7_75t_L g352 ( .A(n_314), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_314), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_319), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_319), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_308), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_330), .B(n_299), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_330), .B(n_299), .Y(n_358) );
INVx3_ASAP7_75t_L g359 ( .A(n_314), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_330), .B(n_299), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_306), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_319), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_307), .B(n_288), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_307), .B(n_288), .Y(n_364) );
AND2x4_ASAP7_75t_SL g365 ( .A(n_329), .B(n_282), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_321), .Y(n_366) );
AND2x4_ASAP7_75t_L g367 ( .A(n_312), .B(n_297), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_308), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_307), .B(n_288), .Y(n_369) );
INVx4_ASAP7_75t_L g370 ( .A(n_306), .Y(n_370) );
INVx2_ASAP7_75t_SL g371 ( .A(n_312), .Y(n_371) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_323), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_317), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_321), .B(n_297), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_328), .B(n_323), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_317), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_321), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_317), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_374), .B(n_323), .Y(n_379) );
AND2x4_ASAP7_75t_SL g380 ( .A(n_370), .B(n_329), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_335), .B(n_329), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_374), .B(n_312), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_334), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_375), .B(n_327), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_331), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_363), .B(n_312), .Y(n_386) );
AND2x4_ASAP7_75t_L g387 ( .A(n_333), .B(n_312), .Y(n_387) );
NAND2x1p5_ASAP7_75t_L g388 ( .A(n_370), .B(n_290), .Y(n_388) );
NOR2x1_ASAP7_75t_L g389 ( .A(n_370), .B(n_316), .Y(n_389) );
NOR2x1_ASAP7_75t_L g390 ( .A(n_370), .B(n_316), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_335), .B(n_309), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_331), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_363), .B(n_318), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_363), .B(n_318), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_364), .B(n_318), .Y(n_395) );
BUFx2_ASAP7_75t_L g396 ( .A(n_350), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_339), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_340), .B(n_325), .Y(n_398) );
NAND2x1p5_ASAP7_75t_L g399 ( .A(n_370), .B(n_298), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_364), .B(n_318), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_365), .B(n_325), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_342), .Y(n_402) );
AND2x4_ASAP7_75t_L g403 ( .A(n_333), .B(n_318), .Y(n_403) );
INVx1_ASAP7_75t_SL g404 ( .A(n_365), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_344), .Y(n_405) );
INVx2_ASAP7_75t_SL g406 ( .A(n_332), .Y(n_406) );
BUFx3_ASAP7_75t_L g407 ( .A(n_365), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_375), .B(n_318), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_346), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_361), .Y(n_410) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_361), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_346), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_349), .B(n_328), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_349), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_354), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_354), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_355), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_355), .Y(n_418) );
NAND3xp33_ASAP7_75t_L g419 ( .A(n_362), .B(n_326), .C(n_324), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_371), .B(n_322), .Y(n_420) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_372), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_362), .B(n_324), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_334), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_369), .B(n_326), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_334), .Y(n_425) );
AND2x4_ASAP7_75t_L g426 ( .A(n_333), .B(n_343), .Y(n_426) );
BUFx2_ASAP7_75t_L g427 ( .A(n_353), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_366), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_366), .B(n_326), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_341), .B(n_317), .Y(n_430) );
BUFx3_ASAP7_75t_L g431 ( .A(n_352), .Y(n_431) );
BUFx2_ASAP7_75t_L g432 ( .A(n_341), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_377), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_347), .B(n_316), .Y(n_434) );
INVxp67_ASAP7_75t_L g435 ( .A(n_377), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_338), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_369), .B(n_316), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_347), .B(n_316), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_351), .B(n_320), .Y(n_439) );
NAND3xp33_ASAP7_75t_SL g440 ( .A(n_396), .B(n_264), .C(n_388), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_427), .Y(n_441) );
OR2x6_ASAP7_75t_L g442 ( .A(n_407), .B(n_352), .Y(n_442) );
NAND3xp33_ASAP7_75t_L g443 ( .A(n_389), .B(n_338), .C(n_303), .Y(n_443) );
CKINVDCx16_ASAP7_75t_R g444 ( .A(n_407), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_380), .B(n_343), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_436), .B(n_338), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_424), .B(n_359), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_406), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_424), .B(n_359), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_391), .B(n_371), .Y(n_450) );
NOR2xp33_ASAP7_75t_SL g451 ( .A(n_380), .B(n_359), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_437), .B(n_371), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_406), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_379), .B(n_359), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_379), .B(n_336), .Y(n_455) );
NOR2x1_ASAP7_75t_L g456 ( .A(n_419), .B(n_320), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_384), .B(n_298), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_408), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_385), .Y(n_459) );
NOR2xp67_ASAP7_75t_R g460 ( .A(n_431), .B(n_336), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_392), .Y(n_461) );
AND3x2_ASAP7_75t_L g462 ( .A(n_432), .B(n_357), .C(n_358), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_397), .Y(n_463) );
INVxp67_ASAP7_75t_L g464 ( .A(n_410), .Y(n_464) );
INVx2_ASAP7_75t_SL g465 ( .A(n_404), .Y(n_465) );
NOR2x1_ASAP7_75t_L g466 ( .A(n_390), .B(n_320), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_381), .B(n_356), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_426), .B(n_343), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_402), .Y(n_469) );
AND2x4_ASAP7_75t_SL g470 ( .A(n_426), .B(n_282), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_405), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_409), .Y(n_472) );
OR2x6_ASAP7_75t_L g473 ( .A(n_399), .B(n_345), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_412), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_383), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_382), .B(n_367), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_414), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_415), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_416), .B(n_356), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_417), .B(n_356), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_398), .B(n_15), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_401), .B(n_15), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_418), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_428), .Y(n_484) );
INVx1_ASAP7_75t_SL g485 ( .A(n_431), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_433), .B(n_368), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_386), .B(n_358), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_435), .B(n_368), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_393), .B(n_367), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_422), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_429), .B(n_373), .Y(n_491) );
INVxp67_ASAP7_75t_L g492 ( .A(n_411), .Y(n_492) );
OR2x6_ASAP7_75t_L g493 ( .A(n_399), .B(n_360), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_394), .B(n_373), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_394), .B(n_360), .Y(n_495) );
AND2x4_ASAP7_75t_L g496 ( .A(n_387), .B(n_367), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_413), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_395), .B(n_373), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_411), .Y(n_499) );
NAND2x1_ASAP7_75t_SL g500 ( .A(n_421), .B(n_367), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_395), .B(n_376), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_423), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_400), .B(n_376), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_400), .B(n_367), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_420), .A2(n_292), .B(n_311), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_421), .Y(n_506) );
INVx2_ASAP7_75t_SL g507 ( .A(n_444), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_490), .B(n_438), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_442), .B(n_387), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_459), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_455), .B(n_430), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_452), .B(n_434), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_461), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_487), .B(n_403), .Y(n_514) );
OAI21xp33_ASAP7_75t_L g515 ( .A1(n_440), .A2(n_439), .B(n_388), .Y(n_515) );
NAND4xp25_ASAP7_75t_L g516 ( .A(n_481), .B(n_294), .C(n_420), .D(n_403), .Y(n_516) );
INVx1_ASAP7_75t_SL g517 ( .A(n_485), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_463), .Y(n_518) );
INVx1_ASAP7_75t_SL g519 ( .A(n_485), .Y(n_519) );
INVx2_ASAP7_75t_SL g520 ( .A(n_470), .Y(n_520) );
NOR2xp67_ASAP7_75t_L g521 ( .A(n_443), .B(n_425), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_497), .B(n_378), .Y(n_522) );
INVx2_ASAP7_75t_SL g523 ( .A(n_465), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_447), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_469), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_499), .B(n_337), .Y(n_526) );
INVxp67_ASAP7_75t_SL g527 ( .A(n_453), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_494), .B(n_378), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_506), .B(n_378), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_464), .B(n_320), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_471), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_498), .B(n_348), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_472), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_451), .A2(n_320), .B1(n_303), .B2(n_282), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_501), .B(n_348), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_449), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_503), .B(n_348), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_458), .B(n_337), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_474), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_495), .B(n_337), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_477), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_478), .Y(n_542) );
NOR2x1_ASAP7_75t_L g543 ( .A(n_443), .B(n_311), .Y(n_543) );
NAND3xp33_ASAP7_75t_L g544 ( .A(n_456), .B(n_303), .C(n_311), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_454), .B(n_313), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_482), .B(n_468), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_483), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_484), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_475), .Y(n_549) );
OR2x6_ASAP7_75t_L g550 ( .A(n_473), .B(n_297), .Y(n_550) );
NOR2x1_ASAP7_75t_SL g551 ( .A(n_473), .B(n_313), .Y(n_551) );
INVxp67_ASAP7_75t_L g552 ( .A(n_441), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_492), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_479), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_442), .B(n_313), .Y(n_555) );
INVx2_ASAP7_75t_SL g556 ( .A(n_473), .Y(n_556) );
NAND2xp33_ASAP7_75t_L g557 ( .A(n_445), .B(n_294), .Y(n_557) );
INVxp67_ASAP7_75t_L g558 ( .A(n_460), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_476), .B(n_16), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_500), .Y(n_560) );
OAI21xp5_ASAP7_75t_L g561 ( .A1(n_466), .A2(n_311), .B(n_282), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_448), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_479), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_480), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_480), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_554), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_514), .B(n_496), .Y(n_567) );
A2O1A1Ixp33_ASAP7_75t_L g568 ( .A1(n_515), .A2(n_505), .B(n_504), .C(n_489), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_563), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_564), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_565), .Y(n_571) );
AO22x1_ASAP7_75t_L g572 ( .A1(n_507), .A2(n_460), .B1(n_462), .B2(n_303), .Y(n_572) );
OAI21xp5_ASAP7_75t_SL g573 ( .A1(n_516), .A2(n_457), .B(n_282), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_550), .A2(n_493), .B1(n_442), .B2(n_450), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_553), .B(n_446), .Y(n_575) );
OAI21xp33_ASAP7_75t_L g576 ( .A1(n_515), .A2(n_446), .B(n_467), .Y(n_576) );
NOR4xp25_ASAP7_75t_SL g577 ( .A(n_527), .B(n_493), .C(n_303), .D(n_488), .Y(n_577) );
NOR2x1p5_ASAP7_75t_L g578 ( .A(n_516), .B(n_491), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_549), .Y(n_579) );
NAND4xp25_ASAP7_75t_L g580 ( .A(n_559), .B(n_294), .C(n_491), .D(n_486), .Y(n_580) );
OAI21xp5_ASAP7_75t_L g581 ( .A1(n_521), .A2(n_493), .B(n_486), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_557), .A2(n_502), .B1(n_311), .B2(n_305), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_510), .Y(n_583) );
XOR2x2_ASAP7_75t_L g584 ( .A(n_546), .B(n_16), .Y(n_584) );
INVx1_ASAP7_75t_SL g585 ( .A(n_517), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_513), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_511), .B(n_305), .Y(n_587) );
CKINVDCx16_ASAP7_75t_R g588 ( .A(n_520), .Y(n_588) );
AOI22xp33_ASAP7_75t_SL g589 ( .A1(n_556), .A2(n_305), .B1(n_281), .B2(n_283), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_518), .Y(n_590) );
AOI21xp33_ASAP7_75t_L g591 ( .A1(n_530), .A2(n_17), .B(n_18), .Y(n_591) );
INVxp67_ASAP7_75t_SL g592 ( .A(n_562), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_540), .B(n_302), .Y(n_593) );
OAI221xp5_ASAP7_75t_L g594 ( .A1(n_521), .A2(n_17), .B1(n_18), .B2(n_20), .C(n_21), .Y(n_594) );
AO22x1_ASAP7_75t_L g595 ( .A1(n_560), .A2(n_20), .B1(n_21), .B2(n_284), .Y(n_595) );
CKINVDCx16_ASAP7_75t_R g596 ( .A(n_523), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_517), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_560), .B(n_284), .Y(n_598) );
OAI21xp5_ASAP7_75t_SL g599 ( .A1(n_558), .A2(n_284), .B(n_23), .Y(n_599) );
OAI21xp5_ASAP7_75t_L g600 ( .A1(n_573), .A2(n_534), .B(n_519), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_573), .A2(n_534), .B1(n_519), .B2(n_509), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_596), .A2(n_509), .B1(n_552), .B2(n_508), .Y(n_602) );
AO221x1_ASAP7_75t_L g603 ( .A1(n_574), .A2(n_536), .B1(n_524), .B2(n_531), .C(n_539), .Y(n_603) );
AOI21xp33_ASAP7_75t_L g604 ( .A1(n_594), .A2(n_526), .B(n_544), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g605 ( .A1(n_572), .A2(n_551), .B(n_522), .Y(n_605) );
NAND3xp33_ASAP7_75t_L g606 ( .A(n_568), .B(n_544), .C(n_526), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_580), .A2(n_555), .B1(n_532), .B2(n_535), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_588), .A2(n_537), .B1(n_512), .B2(n_545), .Y(n_608) );
OAI221xp5_ASAP7_75t_L g609 ( .A1(n_576), .A2(n_581), .B1(n_580), .B2(n_599), .C(n_584), .Y(n_609) );
OAI221xp5_ASAP7_75t_L g610 ( .A1(n_581), .A2(n_543), .B1(n_525), .B2(n_548), .C(n_547), .Y(n_610) );
OAI31xp33_ASAP7_75t_SL g611 ( .A1(n_592), .A2(n_555), .A3(n_561), .B(n_542), .Y(n_611) );
AOI221x1_ASAP7_75t_SL g612 ( .A1(n_591), .A2(n_541), .B1(n_533), .B2(n_529), .C(n_561), .Y(n_612) );
OAI221xp5_ASAP7_75t_L g613 ( .A1(n_599), .A2(n_538), .B1(n_528), .B2(n_35), .C(n_36), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_566), .Y(n_614) );
AOI32xp33_ASAP7_75t_L g615 ( .A1(n_585), .A2(n_30), .A3(n_33), .B1(n_37), .B2(n_38), .Y(n_615) );
O2A1O1Ixp33_ASAP7_75t_L g616 ( .A1(n_585), .A2(n_39), .B(n_41), .C(n_45), .Y(n_616) );
INVxp67_ASAP7_75t_L g617 ( .A(n_597), .Y(n_617) );
INVx2_ASAP7_75t_SL g618 ( .A(n_567), .Y(n_618) );
OAI22xp33_ASAP7_75t_L g619 ( .A1(n_587), .A2(n_47), .B1(n_50), .B2(n_51), .Y(n_619) );
OAI221xp5_ASAP7_75t_L g620 ( .A1(n_575), .A2(n_55), .B1(n_56), .B2(n_59), .C(n_65), .Y(n_620) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_577), .A2(n_68), .B(n_69), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_569), .B(n_71), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g623 ( .A1(n_595), .A2(n_75), .B(n_78), .Y(n_623) );
OAI221xp5_ASAP7_75t_L g624 ( .A1(n_589), .A2(n_83), .B1(n_84), .B2(n_593), .C(n_571), .Y(n_624) );
AOI21xp5_ASAP7_75t_L g625 ( .A1(n_598), .A2(n_570), .B(n_579), .Y(n_625) );
OAI211xp5_ASAP7_75t_SL g626 ( .A1(n_582), .A2(n_586), .B(n_583), .C(n_590), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_573), .A2(n_580), .B1(n_568), .B2(n_576), .C(n_591), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_578), .B(n_566), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_585), .B(n_567), .Y(n_629) );
AND2x4_ASAP7_75t_L g630 ( .A(n_629), .B(n_618), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_602), .B(n_628), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_614), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_612), .B(n_627), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_612), .B(n_607), .Y(n_634) );
NAND4xp25_ASAP7_75t_L g635 ( .A(n_609), .B(n_611), .C(n_601), .D(n_600), .Y(n_635) );
NOR4xp25_ASAP7_75t_L g636 ( .A(n_606), .B(n_626), .C(n_610), .D(n_608), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_630), .B(n_603), .Y(n_637) );
NAND4xp25_ASAP7_75t_L g638 ( .A(n_633), .B(n_623), .C(n_624), .D(n_615), .Y(n_638) );
NAND3xp33_ASAP7_75t_SL g639 ( .A(n_636), .B(n_616), .C(n_621), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g640 ( .A(n_635), .B(n_620), .C(n_604), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_637), .B(n_631), .Y(n_641) );
AND2x4_ASAP7_75t_L g642 ( .A(n_640), .B(n_632), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_639), .B(n_634), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_643), .B(n_638), .Y(n_644) );
NOR3xp33_ASAP7_75t_SL g645 ( .A(n_642), .B(n_613), .C(n_619), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_644), .Y(n_646) );
INVx3_ASAP7_75t_L g647 ( .A(n_645), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_647), .A2(n_641), .B1(n_642), .B2(n_617), .Y(n_648) );
INVx2_ASAP7_75t_SL g649 ( .A(n_646), .Y(n_649) );
OAI21xp5_ASAP7_75t_L g650 ( .A1(n_648), .A2(n_647), .B(n_646), .Y(n_650) );
OAI21xp5_ASAP7_75t_SL g651 ( .A1(n_650), .A2(n_647), .B(n_649), .Y(n_651) );
AO21x2_ASAP7_75t_L g652 ( .A1(n_651), .A2(n_647), .B(n_605), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_652), .A2(n_625), .B(n_622), .Y(n_653) );
endmodule