module fake_jpeg_27745_n_201 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_201);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_36),
.Y(n_49)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_0),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_37),
.A2(n_30),
.B1(n_22),
.B2(n_27),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_55),
.B1(n_60),
.B2(n_19),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_41),
.Y(n_70)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_30),
.B1(n_27),
.B2(n_22),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_48),
.A2(n_58),
.B1(n_59),
.B2(n_53),
.Y(n_81)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_52),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_32),
.A2(n_15),
.B1(n_29),
.B2(n_28),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_54),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_33),
.A2(n_25),
.B1(n_19),
.B2(n_20),
.Y(n_55)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_41),
.Y(n_80)
);

AO22x2_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_31),
.B1(n_24),
.B2(n_23),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_19),
.B1(n_20),
.B2(n_25),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_49),
.B(n_36),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_71),
.Y(n_97)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_63),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_31),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_43),
.Y(n_86)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_75),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_0),
.C(n_1),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_77),
.Y(n_101)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_46),
.B(n_45),
.C(n_44),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_52),
.B(n_50),
.C(n_21),
.Y(n_91)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_47),
.B1(n_43),
.B2(n_57),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_58),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_98),
.C(n_79),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_58),
.B1(n_53),
.B2(n_45),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_83),
.A2(n_84),
.B1(n_89),
.B2(n_93),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_75),
.A2(n_59),
.B1(n_44),
.B2(n_47),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_86),
.B(n_96),
.Y(n_115)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_50),
.B1(n_25),
.B2(n_20),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_68),
.A2(n_50),
.B1(n_24),
.B2(n_31),
.Y(n_96)
);

MAJx2_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_24),
.C(n_1),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_29),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_102),
.B(n_15),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_24),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_73),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_64),
.Y(n_104)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_64),
.Y(n_105)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_100),
.A2(n_78),
.B(n_70),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_107),
.A2(n_118),
.B(n_122),
.Y(n_132)
);

MAJx2_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_98),
.C(n_94),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_117),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_110),
.B(n_112),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_113),
.B(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_73),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_77),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_67),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_121),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_71),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_120),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_61),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_63),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_129),
.C(n_115),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_94),
.B(n_101),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_127),
.B(n_134),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_95),
.B(n_93),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_95),
.C(n_89),
.Y(n_129)
);

OAI22x1_ASAP7_75t_L g130 ( 
.A1(n_111),
.A2(n_96),
.B1(n_74),
.B2(n_52),
.Y(n_130)
);

AOI22x1_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_28),
.B1(n_26),
.B2(n_17),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_88),
.B1(n_90),
.B2(n_85),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_133),
.A2(n_114),
.B1(n_115),
.B2(n_117),
.Y(n_145)
);

NAND2x1_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_88),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_111),
.A2(n_74),
.B(n_52),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_135),
.A2(n_2),
.B(n_3),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_0),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_151),
.Y(n_156)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_145),
.A2(n_148),
.B1(n_149),
.B2(n_154),
.Y(n_167)
);

OAI32xp33_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_118),
.A3(n_113),
.B1(n_106),
.B2(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_112),
.B1(n_90),
.B2(n_85),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_26),
.C(n_17),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_124),
.C(n_131),
.Y(n_165)
);

AOI221xp5_ASAP7_75t_L g151 ( 
.A1(n_126),
.A2(n_16),
.B1(n_2),
.B2(n_3),
.C(n_5),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_153),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_16),
.B1(n_3),
.B2(n_5),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_155),
.A2(n_132),
.B(n_130),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_127),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_147),
.A2(n_155),
.B(n_146),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_164),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_147),
.A2(n_135),
.B(n_134),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_150),
.C(n_128),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_136),
.B1(n_149),
.B2(n_140),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_174),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_174),
.C(n_175),
.Y(n_180)
);

XNOR2x1_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_128),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_172),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_149),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_139),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_163),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_181),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_182),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_172),
.B(n_160),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_165),
.C(n_166),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_171),
.B(n_156),
.Y(n_183)
);

OAI221xp5_ASAP7_75t_L g189 ( 
.A1(n_183),
.A2(n_156),
.B1(n_137),
.B2(n_7),
.C(n_8),
.Y(n_189)
);

AO21x1_ASAP7_75t_L g184 ( 
.A1(n_178),
.A2(n_161),
.B(n_159),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_184),
.A2(n_187),
.B(n_189),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_180),
.A2(n_170),
.B(n_159),
.Y(n_187)
);

NAND4xp25_ASAP7_75t_SL g188 ( 
.A(n_177),
.B(n_137),
.C(n_173),
.D(n_7),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_185),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_2),
.C(n_6),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_190),
.B(n_192),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_185),
.B(n_6),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_10),
.C(n_11),
.Y(n_196)
);

NOR3xp33_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_8),
.C(n_9),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_13),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_196),
.B(n_13),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_197),
.A2(n_198),
.B(n_194),
.Y(n_199)
);

OAI21x1_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_13),
.B(n_14),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_14),
.C(n_196),
.Y(n_201)
);


endmodule