module fake_netlist_5_1702_n_1708 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1708);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1708;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_150;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1556;
wire n_1384;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_152;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_151;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1689;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g150 ( 
.A(n_15),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_112),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_34),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_7),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_43),
.Y(n_155)
);

BUFx10_ASAP7_75t_L g156 ( 
.A(n_67),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_136),
.Y(n_157)
);

INVx4_ASAP7_75t_R g158 ( 
.A(n_57),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_30),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_52),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_105),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_135),
.Y(n_162)
);

BUFx2_ASAP7_75t_SL g163 ( 
.A(n_23),
.Y(n_163)
);

INVxp33_ASAP7_75t_SL g164 ( 
.A(n_40),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_20),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_31),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_30),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_10),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_120),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_5),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_81),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_4),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_88),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_62),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_87),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_134),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_60),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_123),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_52),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_45),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_41),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_61),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_99),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_95),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_66),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_145),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_75),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_124),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_10),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_31),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_5),
.Y(n_192)
);

BUFx10_ASAP7_75t_L g193 ( 
.A(n_118),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_114),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_21),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_51),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_24),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_101),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_96),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_100),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_69),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_129),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_144),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_26),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_127),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_43),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_12),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_107),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_139),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_9),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_58),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_68),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_6),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_0),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_74),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_17),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_133),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_59),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_48),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_79),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_115),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_103),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_130),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_148),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_51),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_21),
.Y(n_226)
);

INVxp67_ASAP7_75t_SL g227 ( 
.A(n_40),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_54),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_140),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_27),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_63),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_20),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_27),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_91),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_11),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_84),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_131),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_147),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_149),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_92),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_29),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_80),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_2),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_38),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_29),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_121),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_76),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_1),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_128),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_14),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_73),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_0),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_102),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_11),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_26),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_34),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_4),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_12),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_13),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_38),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_15),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_90),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_19),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_78),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_65),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_64),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_82),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_9),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_1),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_49),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_24),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_56),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_48),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_25),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_25),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_85),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_23),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_44),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_7),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_110),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_28),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_14),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_47),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_111),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_17),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_32),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_45),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_106),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_18),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_2),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_44),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_70),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_72),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_19),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_109),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_6),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_143),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_104),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_36),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_93),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_138),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_256),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_256),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_256),
.Y(n_304)
);

BUFx6f_ASAP7_75t_SL g305 ( 
.A(n_156),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_256),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_171),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_256),
.Y(n_308)
);

NOR2xp67_ASAP7_75t_L g309 ( 
.A(n_214),
.B(n_3),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_151),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_157),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_201),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_256),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_273),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_273),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_273),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_201),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_159),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_173),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_273),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_273),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_273),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_289),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_289),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_154),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_271),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_289),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g328 ( 
.A(n_230),
.B(n_3),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_161),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_219),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_289),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_289),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_212),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_265),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_289),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_175),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_214),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_298),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_258),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_162),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_160),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_258),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_169),
.Y(n_343)
);

INVxp33_ASAP7_75t_L g344 ( 
.A(n_150),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_269),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_269),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_281),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_281),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_282),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_156),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_282),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_174),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_176),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_178),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_287),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_287),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_182),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_183),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_271),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_186),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_271),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_150),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_152),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_152),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_164),
.B(n_8),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_155),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_187),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_153),
.B(n_8),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_175),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_188),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_259),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_194),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_302),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_359),
.B(n_177),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_308),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_359),
.B(n_177),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_308),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_316),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_316),
.Y(n_379)
);

AND2x4_ASAP7_75t_L g380 ( 
.A(n_302),
.B(n_239),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_303),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_303),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_304),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_368),
.B(n_185),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_304),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_306),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_306),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_312),
.B(n_247),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_313),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_313),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_314),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_314),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_315),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_315),
.Y(n_394)
);

CKINVDCx6p67_ASAP7_75t_R g395 ( 
.A(n_305),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_320),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_320),
.B(n_247),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_321),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_321),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_322),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_322),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_361),
.B(n_239),
.Y(n_402)
);

INVx5_ASAP7_75t_L g403 ( 
.A(n_342),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_323),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_323),
.B(n_153),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_324),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_324),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_327),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_361),
.B(n_184),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_327),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_326),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_331),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_331),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_371),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_332),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_332),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_335),
.B(n_184),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_335),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_342),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_337),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_337),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_339),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_326),
.B(n_190),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_339),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_345),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_345),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_346),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_346),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_341),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_347),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_347),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_348),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_336),
.B(n_190),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_369),
.B(n_198),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_348),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_325),
.Y(n_436)
);

INVx4_ASAP7_75t_L g437 ( 
.A(n_349),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_380),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_429),
.B(n_310),
.Y(n_439)
);

NAND2xp33_ASAP7_75t_R g440 ( 
.A(n_411),
.B(n_311),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_414),
.B(n_350),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_429),
.B(n_329),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_414),
.B(n_350),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_419),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_414),
.B(n_433),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_433),
.A2(n_317),
.B1(n_309),
.B2(n_365),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_411),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_417),
.Y(n_448)
);

NAND2xp33_ASAP7_75t_L g449 ( 
.A(n_384),
.B(n_185),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_395),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_417),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_417),
.Y(n_452)
);

INVx4_ASAP7_75t_SL g453 ( 
.A(n_417),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_417),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_R g455 ( 
.A(n_436),
.B(n_13),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_L g456 ( 
.A1(n_433),
.A2(n_309),
.B1(n_168),
.B2(n_291),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_419),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_411),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_429),
.B(n_340),
.Y(n_459)
);

NAND3xp33_ASAP7_75t_L g460 ( 
.A(n_388),
.B(n_352),
.C(n_343),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_433),
.B(n_353),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_411),
.B(n_357),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_419),
.Y(n_463)
);

NAND3xp33_ASAP7_75t_L g464 ( 
.A(n_388),
.B(n_370),
.C(n_360),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_388),
.B(n_372),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_436),
.A2(n_328),
.B1(n_227),
.B2(n_299),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_417),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_433),
.B(n_237),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_380),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_434),
.B(n_380),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_417),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_419),
.Y(n_472)
);

INVx5_ASAP7_75t_L g473 ( 
.A(n_383),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_434),
.B(n_301),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_419),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_434),
.A2(n_168),
.B1(n_155),
.B2(n_195),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_436),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_384),
.A2(n_250),
.B1(n_204),
.B2(n_207),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_423),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_417),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_423),
.Y(n_481)
);

OR2x6_ASAP7_75t_L g482 ( 
.A(n_423),
.B(n_163),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_434),
.B(n_199),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_381),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_383),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_423),
.B(n_354),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_383),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_423),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_380),
.B(n_200),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_381),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_384),
.B(n_358),
.Y(n_491)
);

OAI21xp33_ASAP7_75t_SL g492 ( 
.A1(n_409),
.A2(n_405),
.B(n_376),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_373),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_373),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_373),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_373),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_374),
.B(n_367),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_374),
.B(n_318),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_381),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_374),
.B(n_330),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_374),
.B(n_307),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_374),
.B(n_156),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_409),
.B(n_349),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_382),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_376),
.B(n_305),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_376),
.B(n_156),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_409),
.B(n_351),
.Y(n_507)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_380),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_381),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_381),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_382),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_385),
.Y(n_512)
);

BUFx10_ASAP7_75t_L g513 ( 
.A(n_380),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_376),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_382),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_382),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_380),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_387),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_387),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_387),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_376),
.B(n_193),
.Y(n_521)
);

AND3x2_ASAP7_75t_L g522 ( 
.A(n_402),
.B(n_277),
.C(n_222),
.Y(n_522)
);

INVx4_ASAP7_75t_L g523 ( 
.A(n_380),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_387),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_394),
.Y(n_525)
);

BUFx4f_ASAP7_75t_L g526 ( 
.A(n_395),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_402),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_394),
.Y(n_528)
);

NAND2xp33_ASAP7_75t_L g529 ( 
.A(n_409),
.B(n_185),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_383),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_394),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_402),
.Y(n_532)
);

INVxp67_ASAP7_75t_SL g533 ( 
.A(n_397),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_402),
.B(n_205),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_402),
.B(n_208),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_409),
.B(n_193),
.Y(n_536)
);

AND3x2_ASAP7_75t_L g537 ( 
.A(n_421),
.B(n_202),
.C(n_198),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_385),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_383),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_394),
.Y(n_540)
);

BUFx10_ASAP7_75t_L g541 ( 
.A(n_395),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_383),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_395),
.B(n_305),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_401),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_437),
.B(n_193),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_401),
.Y(n_546)
);

OR2x6_ASAP7_75t_L g547 ( 
.A(n_405),
.B(n_163),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_421),
.B(n_351),
.Y(n_548)
);

INVx1_ASAP7_75t_SL g549 ( 
.A(n_395),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_385),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_401),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_385),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_385),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_401),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_408),
.B(n_211),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_437),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_386),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_421),
.B(n_355),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_421),
.B(n_422),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_408),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_422),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_386),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_408),
.B(n_217),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_408),
.B(n_218),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_386),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_410),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_410),
.Y(n_567)
);

BUFx4f_ASAP7_75t_L g568 ( 
.A(n_383),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_437),
.B(n_344),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_386),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_405),
.B(n_362),
.Y(n_571)
);

INVxp33_ASAP7_75t_SL g572 ( 
.A(n_397),
.Y(n_572)
);

INVxp67_ASAP7_75t_SL g573 ( 
.A(n_397),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_410),
.Y(n_574)
);

BUFx6f_ASAP7_75t_SL g575 ( 
.A(n_437),
.Y(n_575)
);

OR2x6_ASAP7_75t_L g576 ( 
.A(n_437),
.B(n_189),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_422),
.Y(n_577)
);

AND2x2_ASAP7_75t_SL g578 ( 
.A(n_437),
.B(n_185),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_422),
.B(n_355),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_410),
.B(n_220),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_386),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_437),
.B(n_193),
.Y(n_582)
);

NAND2xp33_ASAP7_75t_SL g583 ( 
.A(n_437),
.B(n_165),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_389),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_533),
.B(n_573),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_572),
.B(n_415),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_572),
.B(n_166),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_532),
.B(n_362),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_527),
.B(n_415),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_492),
.B(n_185),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_444),
.Y(n_591)
);

INVxp67_ASAP7_75t_SL g592 ( 
.A(n_532),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_527),
.B(n_415),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_491),
.A2(n_319),
.B1(n_333),
.B2(n_334),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_444),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_492),
.B(n_452),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_438),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_452),
.B(n_185),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_438),
.Y(n_599)
);

OR2x2_ASAP7_75t_L g600 ( 
.A(n_447),
.B(n_363),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_514),
.B(n_488),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_479),
.B(n_167),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_445),
.B(n_338),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_452),
.B(n_229),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_445),
.B(n_363),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_559),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_481),
.B(n_461),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_561),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_488),
.B(n_415),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_452),
.B(n_229),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_448),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_569),
.B(n_416),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_440),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_577),
.B(n_416),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_577),
.B(n_416),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_460),
.B(n_170),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_447),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_578),
.B(n_416),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_578),
.B(n_427),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_452),
.B(n_229),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_458),
.Y(n_621)
);

NAND2x1p5_ASAP7_75t_L g622 ( 
.A(n_526),
.B(n_469),
.Y(n_622)
);

INVx8_ASAP7_75t_L g623 ( 
.A(n_482),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_578),
.B(n_427),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_470),
.B(n_427),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_559),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_493),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_540),
.B(n_544),
.Y(n_628)
);

NOR2x1p5_ASAP7_75t_L g629 ( 
.A(n_450),
.B(n_172),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_503),
.B(n_364),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_457),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_497),
.A2(n_223),
.B1(n_224),
.B2(n_228),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_560),
.B(n_427),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_457),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_451),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_503),
.B(n_364),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_471),
.B(n_229),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_501),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_446),
.A2(n_253),
.B1(n_231),
.B2(n_221),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_463),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_458),
.Y(n_641)
);

OAI22x1_ASAP7_75t_R g642 ( 
.A1(n_455),
.A2(n_245),
.B1(n_248),
.B2(n_244),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_451),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_501),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_454),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_477),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_464),
.B(n_179),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_498),
.B(n_180),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_463),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_454),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_560),
.B(n_427),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_449),
.A2(n_263),
.B1(n_255),
.B2(n_296),
.Y(n_652)
);

OA21x2_ASAP7_75t_L g653 ( 
.A1(n_493),
.A2(n_399),
.B(n_389),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g654 ( 
.A1(n_468),
.A2(n_231),
.B1(n_221),
.B2(n_215),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_471),
.B(n_229),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_500),
.B(n_181),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_465),
.B(n_192),
.Y(n_657)
);

BUFx2_ASAP7_75t_L g658 ( 
.A(n_477),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_471),
.B(n_229),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_471),
.B(n_234),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_469),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_507),
.B(n_427),
.Y(n_662)
);

INVxp67_ASAP7_75t_SL g663 ( 
.A(n_542),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_449),
.A2(n_547),
.B1(n_571),
.B2(n_476),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_441),
.B(n_366),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_439),
.B(n_196),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_467),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_467),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_474),
.A2(n_267),
.B1(n_236),
.B2(n_238),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_517),
.B(n_366),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_480),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_571),
.B(n_390),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_480),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_517),
.B(n_202),
.Y(n_674)
);

O2A1O1Ixp33_ASAP7_75t_L g675 ( 
.A1(n_483),
.A2(n_189),
.B(n_263),
.C(n_255),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_494),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_472),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_534),
.B(n_535),
.Y(n_678)
);

INVx8_ASAP7_75t_L g679 ( 
.A(n_482),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_471),
.B(n_240),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_442),
.B(n_197),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_508),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_462),
.B(n_206),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_459),
.B(n_210),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_482),
.B(n_216),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_494),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_513),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_495),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_450),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_508),
.B(n_242),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_482),
.B(n_486),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_495),
.Y(n_692)
);

NAND2xp33_ASAP7_75t_L g693 ( 
.A(n_489),
.B(n_246),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_508),
.B(n_523),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_496),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_523),
.B(n_249),
.Y(n_696)
);

AO221x1_ASAP7_75t_L g697 ( 
.A1(n_485),
.A2(n_296),
.B1(n_195),
.B2(n_191),
.C(n_291),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_523),
.Y(n_698)
);

NAND3xp33_ASAP7_75t_L g699 ( 
.A(n_478),
.B(n_260),
.C(n_225),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_556),
.B(n_251),
.Y(n_700)
);

INVxp33_ASAP7_75t_L g701 ( 
.A(n_443),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_555),
.B(n_390),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_513),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_526),
.B(n_513),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_496),
.Y(n_705)
);

INVx4_ASAP7_75t_L g706 ( 
.A(n_453),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_504),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_504),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_563),
.B(n_564),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_547),
.A2(n_209),
.B1(n_203),
.B2(n_215),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_511),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_541),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_576),
.B(n_203),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_511),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_548),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_472),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_526),
.B(n_262),
.Y(n_717)
);

INVxp33_ASAP7_75t_L g718 ( 
.A(n_478),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_453),
.B(n_264),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_580),
.B(n_390),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_547),
.B(n_226),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_541),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_515),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_515),
.B(n_516),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_475),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_547),
.B(n_232),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_453),
.B(n_272),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_516),
.B(n_390),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_518),
.B(n_390),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_518),
.Y(n_730)
);

OAI22xp33_ASAP7_75t_L g731 ( 
.A1(n_466),
.A2(n_191),
.B1(n_213),
.B2(n_286),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_519),
.B(n_390),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_519),
.B(n_391),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_520),
.B(n_391),
.Y(n_734)
);

O2A1O1Ixp33_ASAP7_75t_L g735 ( 
.A1(n_529),
.A2(n_213),
.B(n_286),
.C(n_428),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_520),
.B(n_391),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_524),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_524),
.B(n_391),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_542),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_466),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_475),
.Y(n_741)
);

OR2x6_ASAP7_75t_L g742 ( 
.A(n_502),
.B(n_506),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_484),
.Y(n_743)
);

NOR2x1p5_ASAP7_75t_L g744 ( 
.A(n_455),
.B(n_233),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_525),
.B(n_391),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_525),
.B(n_391),
.Y(n_746)
);

HB1xp67_ASAP7_75t_L g747 ( 
.A(n_521),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_528),
.B(n_391),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_528),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_453),
.B(n_276),
.Y(n_750)
);

O2A1O1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_639),
.A2(n_536),
.B(n_582),
.C(n_545),
.Y(n_751)
);

OAI21xp5_ASAP7_75t_L g752 ( 
.A1(n_619),
.A2(n_568),
.B(n_546),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_L g753 ( 
.A1(n_585),
.A2(n_529),
.B(n_568),
.Y(n_753)
);

OAI21xp5_ASAP7_75t_L g754 ( 
.A1(n_624),
.A2(n_568),
.B(n_546),
.Y(n_754)
);

NOR2xp67_ASAP7_75t_L g755 ( 
.A(n_689),
.B(n_543),
.Y(n_755)
);

INVx6_ASAP7_75t_L g756 ( 
.A(n_623),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_607),
.B(n_505),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_718),
.A2(n_576),
.B1(n_583),
.B2(n_456),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_596),
.A2(n_551),
.B(n_531),
.Y(n_759)
);

A2O1A1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_666),
.A2(n_549),
.B(n_209),
.C(n_253),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_607),
.B(n_531),
.Y(n_761)
);

A2O1A1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_666),
.A2(n_681),
.B(n_683),
.C(n_678),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_606),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_683),
.B(n_522),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_596),
.A2(n_625),
.B(n_682),
.Y(n_765)
);

A2O1A1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_657),
.A2(n_266),
.B(n_284),
.C(n_300),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_715),
.B(n_554),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_691),
.A2(n_709),
.B1(n_647),
.B2(n_616),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_715),
.B(n_554),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_597),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_682),
.A2(n_487),
.B(n_485),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_597),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_698),
.A2(n_487),
.B(n_485),
.Y(n_773)
);

INVx4_ASAP7_75t_L g774 ( 
.A(n_597),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_626),
.B(n_566),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_613),
.Y(n_776)
);

AOI21xp33_ASAP7_75t_L g777 ( 
.A1(n_657),
.A2(n_576),
.B(n_297),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_627),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_601),
.B(n_567),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_611),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_586),
.B(n_567),
.Y(n_781)
);

O2A1O1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_654),
.A2(n_576),
.B(n_574),
.C(n_297),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_605),
.B(n_574),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_592),
.B(n_548),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_664),
.B(n_558),
.Y(n_785)
);

AOI21x1_ASAP7_75t_L g786 ( 
.A1(n_690),
.A2(n_584),
.B(n_581),
.Y(n_786)
);

INVx1_ASAP7_75t_SL g787 ( 
.A(n_658),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_587),
.B(n_541),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_664),
.B(n_558),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_670),
.B(n_579),
.Y(n_790)
);

O2A1O1Ixp33_ASAP7_75t_L g791 ( 
.A1(n_590),
.A2(n_584),
.B(n_581),
.C(n_484),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_694),
.A2(n_530),
.B(n_487),
.Y(n_792)
);

OAI21xp5_ASAP7_75t_L g793 ( 
.A1(n_618),
.A2(n_490),
.B(n_570),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_670),
.B(n_530),
.Y(n_794)
);

BUFx12f_ASAP7_75t_L g795 ( 
.A(n_646),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_588),
.B(n_539),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_694),
.A2(n_539),
.B(n_570),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_663),
.A2(n_550),
.B(n_565),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_588),
.B(n_490),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_617),
.Y(n_800)
);

INVxp67_ASAP7_75t_L g801 ( 
.A(n_600),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_702),
.A2(n_550),
.B(n_565),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_635),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_602),
.B(n_356),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_643),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_645),
.B(n_499),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_720),
.A2(n_510),
.B(n_562),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_687),
.B(n_280),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_650),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_662),
.A2(n_509),
.B(n_557),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_667),
.B(n_499),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_668),
.B(n_512),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_671),
.B(n_512),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_673),
.B(n_538),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_687),
.B(n_288),
.Y(n_815)
);

O2A1O1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_590),
.A2(n_553),
.B(n_552),
.C(n_538),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_707),
.Y(n_817)
);

O2A1O1Ixp5_ASAP7_75t_L g818 ( 
.A1(n_690),
.A2(n_553),
.B(n_552),
.C(n_428),
.Y(n_818)
);

NAND2x1p5_ASAP7_75t_L g819 ( 
.A(n_706),
.B(n_542),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_602),
.B(n_356),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_672),
.A2(n_391),
.B(n_392),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_708),
.Y(n_822)
);

A2O1A1Ixp33_ASAP7_75t_L g823 ( 
.A1(n_616),
.A2(n_428),
.B(n_430),
.C(n_292),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_628),
.A2(n_542),
.B(n_473),
.Y(n_824)
);

HB1xp67_ASAP7_75t_L g825 ( 
.A(n_621),
.Y(n_825)
);

AOI21x1_ASAP7_75t_L g826 ( 
.A1(n_696),
.A2(n_389),
.B(n_407),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_661),
.A2(n_575),
.B1(n_295),
.B2(n_293),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_599),
.B(n_630),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_703),
.A2(n_542),
.B(n_473),
.Y(n_829)
);

NOR2xp67_ASAP7_75t_L g830 ( 
.A(n_594),
.B(n_53),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_630),
.B(n_636),
.Y(n_831)
);

AO21x1_ASAP7_75t_L g832 ( 
.A1(n_647),
.A2(n_428),
.B(n_430),
.Y(n_832)
);

OAI21xp5_ASAP7_75t_L g833 ( 
.A1(n_612),
.A2(n_413),
.B(n_393),
.Y(n_833)
);

O2A1O1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_710),
.A2(n_430),
.B(n_407),
.C(n_399),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_636),
.B(n_430),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_SL g836 ( 
.A(n_603),
.B(n_638),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_708),
.Y(n_837)
);

AOI21x1_ASAP7_75t_L g838 ( 
.A1(n_696),
.A2(n_406),
.B(n_400),
.Y(n_838)
);

INVx4_ASAP7_75t_L g839 ( 
.A(n_597),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_633),
.A2(n_375),
.B(n_377),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_641),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_687),
.B(n_235),
.Y(n_842)
);

NOR2xp67_ASAP7_75t_L g843 ( 
.A(n_747),
.B(n_55),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_651),
.A2(n_375),
.B(n_377),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_676),
.B(n_537),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_686),
.B(n_392),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_687),
.B(n_241),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_704),
.A2(n_378),
.B(n_379),
.Y(n_848)
);

INVx4_ASAP7_75t_L g849 ( 
.A(n_706),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_688),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_L g851 ( 
.A1(n_661),
.A2(n_252),
.B1(n_243),
.B2(n_257),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_692),
.B(n_392),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_608),
.B(n_254),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_695),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_705),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_704),
.A2(n_375),
.B(n_377),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_711),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_665),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_714),
.B(n_392),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_589),
.A2(n_379),
.B(n_378),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_593),
.A2(n_379),
.B(n_378),
.Y(n_861)
);

AO22x1_ASAP7_75t_L g862 ( 
.A1(n_701),
.A2(n_684),
.B1(n_691),
.B2(n_721),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_723),
.B(n_392),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_684),
.B(n_261),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_730),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_737),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_728),
.A2(n_413),
.B(n_393),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_749),
.B(n_392),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_648),
.B(n_656),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_724),
.A2(n_379),
.B(n_378),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_609),
.A2(n_379),
.B(n_378),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_599),
.B(n_420),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_729),
.A2(n_393),
.B(n_392),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_660),
.A2(n_418),
.B(n_400),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_674),
.B(n_420),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_653),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_740),
.B(n_268),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_648),
.B(n_270),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_653),
.Y(n_879)
);

AO22x1_ASAP7_75t_L g880 ( 
.A1(n_721),
.A2(n_278),
.B1(n_275),
.B2(n_274),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_653),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_669),
.B(n_656),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_660),
.A2(n_404),
.B(n_418),
.Y(n_883)
);

NOR2xp67_ASAP7_75t_L g884 ( 
.A(n_632),
.B(n_699),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_685),
.B(n_712),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_622),
.A2(n_283),
.B1(n_294),
.B2(n_290),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_680),
.A2(n_404),
.B(n_389),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_732),
.Y(n_888)
);

AND3x1_ASAP7_75t_SL g889 ( 
.A(n_744),
.B(n_279),
.C(n_285),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_680),
.A2(n_406),
.B(n_389),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_591),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_685),
.B(n_431),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_713),
.B(n_393),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_726),
.B(n_742),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_742),
.B(n_712),
.Y(n_895)
);

AND2x2_ASAP7_75t_SL g896 ( 
.A(n_652),
.B(n_158),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_733),
.A2(n_738),
.B(n_748),
.Y(n_897)
);

NOR2x1_ASAP7_75t_L g898 ( 
.A(n_722),
.B(n_392),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_742),
.B(n_420),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_622),
.A2(n_393),
.B1(n_413),
.B2(n_431),
.Y(n_900)
);

NAND2x1p5_ASAP7_75t_L g901 ( 
.A(n_739),
.B(n_473),
.Y(n_901)
);

AOI21x1_ASAP7_75t_L g902 ( 
.A1(n_700),
.A2(n_407),
.B(n_404),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_713),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_734),
.A2(n_407),
.B(n_418),
.Y(n_904)
);

OR2x6_ASAP7_75t_L g905 ( 
.A(n_623),
.B(n_431),
.Y(n_905)
);

NAND2x1_ASAP7_75t_L g906 ( 
.A(n_739),
.B(n_158),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_644),
.B(n_16),
.Y(n_907)
);

AO21x1_ASAP7_75t_L g908 ( 
.A1(n_700),
.A2(n_399),
.B(n_400),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_629),
.B(n_431),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_722),
.B(n_432),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_652),
.A2(n_393),
.B1(n_413),
.B2(n_420),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_623),
.B(n_431),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_736),
.A2(n_407),
.B(n_418),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_739),
.B(n_432),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_745),
.A2(n_400),
.B(n_404),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_679),
.B(n_424),
.Y(n_916)
);

O2A1O1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_731),
.A2(n_418),
.B(n_399),
.C(n_400),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_679),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_739),
.B(n_432),
.Y(n_919)
);

OR2x6_ASAP7_75t_L g920 ( 
.A(n_679),
.B(n_435),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_746),
.A2(n_404),
.B(n_406),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_614),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_598),
.A2(n_406),
.B(n_399),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_675),
.B(n_425),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_869),
.B(n_757),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_765),
.A2(n_750),
.B(n_719),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_762),
.B(n_615),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_765),
.A2(n_750),
.B(n_719),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_768),
.B(n_731),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_778),
.Y(n_930)
);

NAND2x1p5_ASAP7_75t_L g931 ( 
.A(n_849),
.B(n_598),
.Y(n_931)
);

AND2x6_ASAP7_75t_L g932 ( 
.A(n_876),
.B(n_743),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_SL g933 ( 
.A1(n_882),
.A2(n_717),
.B(n_727),
.C(n_604),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_787),
.B(n_604),
.Y(n_934)
);

INVx4_ASAP7_75t_L g935 ( 
.A(n_770),
.Y(n_935)
);

OR2x2_ASAP7_75t_L g936 ( 
.A(n_801),
.B(n_610),
.Y(n_936)
);

AO22x1_ASAP7_75t_L g937 ( 
.A1(n_788),
.A2(n_642),
.B1(n_697),
.B2(n_716),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_753),
.A2(n_727),
.B(n_620),
.Y(n_938)
);

INVxp67_ASAP7_75t_L g939 ( 
.A(n_800),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_877),
.B(n_610),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_SL g941 ( 
.A(n_896),
.B(n_735),
.Y(n_941)
);

NOR2x1_ASAP7_75t_SL g942 ( 
.A(n_849),
.B(n_770),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_858),
.B(n_620),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_828),
.B(n_741),
.Y(n_944)
);

NAND2x1p5_ASAP7_75t_L g945 ( 
.A(n_774),
.B(n_637),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_753),
.A2(n_637),
.B(n_655),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_817),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_825),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_770),
.Y(n_949)
);

O2A1O1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_864),
.A2(n_693),
.B(n_655),
.C(n_659),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_804),
.B(n_725),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_761),
.A2(n_659),
.B1(n_677),
.B2(n_649),
.Y(n_952)
);

O2A1O1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_766),
.A2(n_640),
.B(n_634),
.C(n_631),
.Y(n_953)
);

INVx1_ASAP7_75t_SL g954 ( 
.A(n_831),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_820),
.B(n_595),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_772),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_784),
.A2(n_473),
.B(n_403),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_R g958 ( 
.A(n_776),
.B(n_98),
.Y(n_958)
);

INVx3_ASAP7_75t_SL g959 ( 
.A(n_841),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_795),
.Y(n_960)
);

NOR3xp33_ASAP7_75t_L g961 ( 
.A(n_862),
.B(n_424),
.C(n_426),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_828),
.B(n_432),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_781),
.B(n_435),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_790),
.A2(n_473),
.B(n_403),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_878),
.B(n_16),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_772),
.Y(n_966)
);

OR2x2_ASAP7_75t_L g967 ( 
.A(n_903),
.B(n_435),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_895),
.Y(n_968)
);

INVx4_ASAP7_75t_L g969 ( 
.A(n_772),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_822),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_764),
.B(n_18),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_783),
.A2(n_403),
.B(n_393),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_918),
.B(n_435),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_794),
.A2(n_796),
.B(n_751),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_779),
.B(n_435),
.Y(n_975)
);

AOI221xp5_ASAP7_75t_L g976 ( 
.A1(n_907),
.A2(n_426),
.B1(n_425),
.B2(n_424),
.C(n_420),
.Y(n_976)
);

AOI21x1_ASAP7_75t_L g977 ( 
.A1(n_786),
.A2(n_838),
.B(n_826),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_837),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_799),
.A2(n_403),
.B(n_413),
.Y(n_979)
);

INVxp67_ASAP7_75t_L g980 ( 
.A(n_836),
.Y(n_980)
);

BUFx12f_ASAP7_75t_L g981 ( 
.A(n_756),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_884),
.B(n_432),
.Y(n_982)
);

INVx4_ASAP7_75t_L g983 ( 
.A(n_756),
.Y(n_983)
);

O2A1O1Ixp5_ASAP7_75t_L g984 ( 
.A1(n_777),
.A2(n_426),
.B(n_425),
.C(n_424),
.Y(n_984)
);

BUFx2_ASAP7_75t_L g985 ( 
.A(n_895),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_752),
.A2(n_403),
.B(n_413),
.Y(n_986)
);

INVx1_ASAP7_75t_SL g987 ( 
.A(n_892),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_894),
.B(n_22),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_888),
.B(n_426),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_754),
.A2(n_403),
.B(n_413),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_780),
.B(n_803),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_805),
.B(n_426),
.Y(n_992)
);

AOI21xp33_ASAP7_75t_L g993 ( 
.A1(n_785),
.A2(n_424),
.B(n_28),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_789),
.A2(n_403),
.B(n_412),
.Y(n_994)
);

OA22x2_ASAP7_75t_L g995 ( 
.A1(n_853),
.A2(n_22),
.B1(n_32),
.B2(n_33),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_759),
.A2(n_403),
.B(n_412),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_756),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_885),
.B(n_33),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_905),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_763),
.B(n_432),
.Y(n_1000)
);

INVx5_ASAP7_75t_L g1001 ( 
.A(n_905),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_905),
.Y(n_1002)
);

AO21x1_ASAP7_75t_L g1003 ( 
.A1(n_897),
.A2(n_782),
.B(n_874),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_809),
.B(n_850),
.Y(n_1004)
);

INVx4_ASAP7_75t_L g1005 ( 
.A(n_774),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_922),
.B(n_886),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_854),
.Y(n_1007)
);

INVxp67_ASAP7_75t_L g1008 ( 
.A(n_851),
.Y(n_1008)
);

INVx2_ASAP7_75t_SL g1009 ( 
.A(n_909),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_857),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_775),
.A2(n_403),
.B(n_412),
.Y(n_1011)
);

A2O1A1Ixp33_ASAP7_75t_SL g1012 ( 
.A1(n_758),
.A2(n_94),
.B(n_146),
.C(n_141),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_891),
.Y(n_1013)
);

INVxp67_ASAP7_75t_SL g1014 ( 
.A(n_875),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_755),
.B(n_432),
.Y(n_1015)
);

O2A1O1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_760),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_899),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_875),
.A2(n_432),
.B1(n_412),
.B2(n_398),
.Y(n_1018)
);

BUFx2_ASAP7_75t_L g1019 ( 
.A(n_899),
.Y(n_1019)
);

OR2x4_ASAP7_75t_L g1020 ( 
.A(n_845),
.B(n_855),
.Y(n_1020)
);

BUFx3_ASAP7_75t_L g1021 ( 
.A(n_912),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_916),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_SL g1023 ( 
.A1(n_865),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_843),
.A2(n_432),
.B(n_412),
.C(n_398),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_866),
.A2(n_769),
.B1(n_767),
.B2(n_835),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_922),
.B(n_432),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_879),
.A2(n_432),
.B1(n_412),
.B2(n_398),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_920),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_922),
.B(n_39),
.Y(n_1029)
);

AOI221x1_ASAP7_75t_L g1030 ( 
.A1(n_823),
.A2(n_432),
.B1(n_412),
.B2(n_398),
.C(n_396),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_880),
.B(n_41),
.Y(n_1031)
);

CKINVDCx16_ASAP7_75t_R g1032 ( 
.A(n_920),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_872),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_830),
.B(n_412),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_829),
.A2(n_403),
.B(n_412),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_806),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_897),
.A2(n_403),
.B(n_412),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_793),
.A2(n_403),
.B(n_412),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_818),
.A2(n_398),
.B(n_396),
.C(n_383),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_881),
.B(n_398),
.Y(n_1040)
);

OR2x6_ASAP7_75t_L g1041 ( 
.A(n_920),
.B(n_398),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_872),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_811),
.A2(n_398),
.B1(n_396),
.B2(n_383),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_839),
.B(n_398),
.Y(n_1044)
);

CKINVDCx16_ASAP7_75t_R g1045 ( 
.A(n_839),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_842),
.B(n_42),
.Y(n_1046)
);

NAND2xp33_ASAP7_75t_R g1047 ( 
.A(n_924),
.B(n_893),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_824),
.A2(n_771),
.B(n_773),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_847),
.B(n_398),
.Y(n_1049)
);

INVx4_ASAP7_75t_L g1050 ( 
.A(n_819),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_808),
.A2(n_42),
.B(n_46),
.C(n_47),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_898),
.B(n_46),
.Y(n_1052)
);

NAND3xp33_ASAP7_75t_SL g1053 ( 
.A(n_815),
.B(n_49),
.C(n_50),
.Y(n_1053)
);

INVx5_ASAP7_75t_L g1054 ( 
.A(n_819),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_812),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_813),
.Y(n_1056)
);

BUFx4f_ASAP7_75t_SL g1057 ( 
.A(n_910),
.Y(n_1057)
);

OR2x2_ASAP7_75t_L g1058 ( 
.A(n_814),
.B(n_50),
.Y(n_1058)
);

NOR2x1_ASAP7_75t_R g1059 ( 
.A(n_889),
.B(n_398),
.Y(n_1059)
);

HB1xp67_ASAP7_75t_L g1060 ( 
.A(n_906),
.Y(n_1060)
);

AOI221xp5_ASAP7_75t_L g1061 ( 
.A1(n_827),
.A2(n_396),
.B1(n_383),
.B2(n_83),
.C(n_86),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_846),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_940),
.A2(n_816),
.B(n_791),
.C(n_810),
.Y(n_1063)
);

AO31x2_ASAP7_75t_L g1064 ( 
.A1(n_1030),
.A2(n_832),
.A3(n_1003),
.B(n_908),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_925),
.B(n_868),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_987),
.B(n_954),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_980),
.B(n_852),
.Y(n_1067)
);

OA21x2_ASAP7_75t_L g1068 ( 
.A1(n_974),
.A2(n_928),
.B(n_926),
.Y(n_1068)
);

AO31x2_ASAP7_75t_L g1069 ( 
.A1(n_1039),
.A2(n_887),
.A3(n_874),
.B(n_883),
.Y(n_1069)
);

INVxp67_ASAP7_75t_L g1070 ( 
.A(n_948),
.Y(n_1070)
);

OR2x2_ASAP7_75t_L g1071 ( 
.A(n_954),
.B(n_1022),
.Y(n_1071)
);

BUFx8_ASAP7_75t_L g1072 ( 
.A(n_981),
.Y(n_1072)
);

INVx2_ASAP7_75t_SL g1073 ( 
.A(n_959),
.Y(n_1073)
);

BUFx10_ASAP7_75t_L g1074 ( 
.A(n_1020),
.Y(n_1074)
);

NAND3xp33_ASAP7_75t_L g1075 ( 
.A(n_965),
.B(n_883),
.C(n_887),
.Y(n_1075)
);

AOI21x1_ASAP7_75t_L g1076 ( 
.A1(n_977),
.A2(n_902),
.B(n_890),
.Y(n_1076)
);

OR2x6_ASAP7_75t_SL g1077 ( 
.A(n_997),
.B(n_863),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_968),
.Y(n_1078)
);

BUFx12f_ASAP7_75t_L g1079 ( 
.A(n_960),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_SL g1080 ( 
.A1(n_1016),
.A2(n_917),
.B(n_890),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_987),
.B(n_1036),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_991),
.Y(n_1082)
);

AO22x2_ASAP7_75t_L g1083 ( 
.A1(n_929),
.A2(n_900),
.B1(n_856),
.B2(n_848),
.Y(n_1083)
);

NAND3xp33_ASAP7_75t_L g1084 ( 
.A(n_971),
.B(n_834),
.C(n_921),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_927),
.A2(n_807),
.B(n_802),
.Y(n_1085)
);

AOI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_1006),
.A2(n_859),
.B1(n_919),
.B2(n_914),
.Y(n_1086)
);

AO21x1_ASAP7_75t_L g1087 ( 
.A1(n_941),
.A2(n_848),
.B(n_856),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_1021),
.B(n_821),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_SL g1089 ( 
.A1(n_927),
.A2(n_833),
.B(n_901),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1004),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_933),
.A2(n_798),
.B(n_797),
.Y(n_1091)
);

OAI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_941),
.A2(n_792),
.B1(n_911),
.B2(n_873),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_998),
.A2(n_904),
.B(n_921),
.C(n_915),
.Y(n_1093)
);

NAND2xp33_ASAP7_75t_SL g1094 ( 
.A(n_958),
.B(n_867),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_938),
.A2(n_870),
.B(n_860),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_947),
.Y(n_1096)
);

HB1xp67_ASAP7_75t_L g1097 ( 
.A(n_939),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_1008),
.A2(n_915),
.B1(n_913),
.B2(n_904),
.Y(n_1098)
);

OA21x2_ASAP7_75t_L g1099 ( 
.A1(n_946),
.A2(n_984),
.B(n_1048),
.Y(n_1099)
);

O2A1O1Ixp33_ASAP7_75t_SL g1100 ( 
.A1(n_1012),
.A2(n_913),
.B(n_923),
.C(n_871),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_1037),
.A2(n_840),
.B(n_844),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_978),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_988),
.A2(n_871),
.B(n_861),
.C(n_840),
.Y(n_1103)
);

AO22x2_ASAP7_75t_L g1104 ( 
.A1(n_1053),
.A2(n_923),
.B1(n_77),
.B2(n_89),
.Y(n_1104)
);

AO31x2_ASAP7_75t_L g1105 ( 
.A1(n_1024),
.A2(n_71),
.A3(n_97),
.B(n_108),
.Y(n_1105)
);

O2A1O1Ixp5_ASAP7_75t_L g1106 ( 
.A1(n_937),
.A2(n_113),
.B(n_116),
.C(n_119),
.Y(n_1106)
);

AO31x2_ASAP7_75t_L g1107 ( 
.A1(n_1025),
.A2(n_122),
.A3(n_125),
.B(n_126),
.Y(n_1107)
);

O2A1O1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_1031),
.A2(n_132),
.B(n_137),
.C(n_383),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1056),
.B(n_383),
.Y(n_1109)
);

NAND3xp33_ASAP7_75t_SL g1110 ( 
.A(n_1051),
.B(n_396),
.C(n_1023),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_951),
.A2(n_396),
.B(n_955),
.Y(n_1111)
);

INVx5_ASAP7_75t_L g1112 ( 
.A(n_1041),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_950),
.A2(n_396),
.B(n_943),
.C(n_1061),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_993),
.A2(n_396),
.B(n_934),
.C(n_1029),
.Y(n_1114)
);

OA21x2_ASAP7_75t_L g1115 ( 
.A1(n_993),
.A2(n_396),
.B(n_986),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_963),
.A2(n_396),
.B(n_1025),
.Y(n_1116)
);

AND2x6_ASAP7_75t_L g1117 ( 
.A(n_999),
.B(n_396),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_985),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_1055),
.A2(n_1009),
.B(n_1058),
.C(n_1046),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_930),
.Y(n_1120)
);

OA21x2_ASAP7_75t_L g1121 ( 
.A1(n_990),
.A2(n_1038),
.B(n_975),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_1020),
.B(n_1019),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_936),
.A2(n_1017),
.B(n_1042),
.C(n_982),
.Y(n_1123)
);

NOR2xp67_ASAP7_75t_L g1124 ( 
.A(n_1007),
.B(n_1010),
.Y(n_1124)
);

AOI221x1_ASAP7_75t_L g1125 ( 
.A1(n_961),
.A2(n_952),
.B1(n_994),
.B2(n_1052),
.C(n_975),
.Y(n_1125)
);

AO32x2_ASAP7_75t_L g1126 ( 
.A1(n_952),
.A2(n_1027),
.A3(n_1047),
.B1(n_1043),
.B2(n_969),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_949),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1014),
.B(n_1062),
.Y(n_1128)
);

OAI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_995),
.A2(n_1032),
.B1(n_1057),
.B2(n_1045),
.Y(n_1129)
);

AO31x2_ASAP7_75t_L g1130 ( 
.A1(n_1027),
.A2(n_1040),
.A3(n_989),
.B(n_1043),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_1033),
.B(n_1013),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_989),
.A2(n_1054),
.B(n_1034),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1054),
.A2(n_942),
.B(n_1026),
.Y(n_1133)
);

INVx5_ASAP7_75t_L g1134 ( 
.A(n_1041),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1054),
.A2(n_931),
.B(n_953),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1000),
.A2(n_996),
.B(n_964),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1001),
.A2(n_1054),
.B1(n_983),
.B2(n_931),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_967),
.B(n_970),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_SL g1139 ( 
.A1(n_995),
.A2(n_1001),
.B1(n_1028),
.B2(n_1002),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_944),
.B(n_973),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_979),
.A2(n_957),
.B(n_992),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1049),
.A2(n_972),
.B(n_945),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_945),
.A2(n_1015),
.B(n_1001),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1035),
.A2(n_1011),
.B(n_1044),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_SL g1145 ( 
.A(n_1005),
.B(n_1001),
.Y(n_1145)
);

O2A1O1Ixp33_ASAP7_75t_SL g1146 ( 
.A1(n_962),
.A2(n_1060),
.B(n_956),
.C(n_976),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_973),
.A2(n_956),
.B(n_1028),
.C(n_1002),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_999),
.A2(n_1028),
.B1(n_1002),
.B2(n_1050),
.Y(n_1148)
);

AND2x2_ASAP7_75t_SL g1149 ( 
.A(n_999),
.B(n_1005),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_932),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1059),
.A2(n_1018),
.B(n_932),
.C(n_969),
.Y(n_1151)
);

AO31x2_ASAP7_75t_L g1152 ( 
.A1(n_935),
.A2(n_932),
.A3(n_966),
.B(n_832),
.Y(n_1152)
);

NAND4xp25_ASAP7_75t_L g1153 ( 
.A(n_966),
.B(n_932),
.C(n_330),
.D(n_318),
.Y(n_1153)
);

INVxp67_ASAP7_75t_SL g1154 ( 
.A(n_966),
.Y(n_1154)
);

CKINVDCx11_ASAP7_75t_R g1155 ( 
.A(n_959),
.Y(n_1155)
);

O2A1O1Ixp33_ASAP7_75t_SL g1156 ( 
.A1(n_929),
.A2(n_762),
.B(n_882),
.C(n_1012),
.Y(n_1156)
);

NAND3xp33_ASAP7_75t_L g1157 ( 
.A(n_965),
.B(n_683),
.C(n_681),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_981),
.Y(n_1158)
);

OAI21xp33_ASAP7_75t_SL g1159 ( 
.A1(n_929),
.A2(n_896),
.B(n_768),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_940),
.A2(n_762),
.B(n_768),
.C(n_869),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_926),
.A2(n_762),
.B(n_698),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_981),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_926),
.A2(n_762),
.B(n_698),
.Y(n_1163)
);

OR2x2_ASAP7_75t_L g1164 ( 
.A(n_954),
.B(n_644),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_991),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_926),
.A2(n_762),
.B(n_698),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_925),
.B(n_607),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_991),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_925),
.B(n_607),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_940),
.A2(n_762),
.B(n_768),
.C(n_869),
.Y(n_1170)
);

NAND3x1_ASAP7_75t_L g1171 ( 
.A(n_971),
.B(n_594),
.C(n_1031),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_926),
.A2(n_762),
.B(n_698),
.Y(n_1172)
);

O2A1O1Ixp33_ASAP7_75t_SL g1173 ( 
.A1(n_929),
.A2(n_762),
.B(n_882),
.C(n_1012),
.Y(n_1173)
);

OAI22x1_ASAP7_75t_L g1174 ( 
.A1(n_929),
.A2(n_768),
.B1(n_971),
.B2(n_988),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_925),
.B(n_607),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_925),
.B(n_603),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_940),
.A2(n_762),
.B(n_768),
.C(n_869),
.Y(n_1177)
);

AO31x2_ASAP7_75t_L g1178 ( 
.A1(n_1030),
.A2(n_832),
.A3(n_1003),
.B(n_762),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_925),
.B(n_307),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_926),
.A2(n_762),
.B(n_698),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_948),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_940),
.A2(n_762),
.B(n_768),
.C(n_869),
.Y(n_1182)
);

AOI221xp5_ASAP7_75t_SL g1183 ( 
.A1(n_929),
.A2(n_965),
.B1(n_639),
.B2(n_683),
.C(n_762),
.Y(n_1183)
);

AO32x2_ASAP7_75t_L g1184 ( 
.A1(n_1025),
.A2(n_639),
.A3(n_952),
.B1(n_710),
.B2(n_654),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_926),
.A2(n_762),
.B(n_698),
.Y(n_1185)
);

NAND3xp33_ASAP7_75t_L g1186 ( 
.A(n_965),
.B(n_683),
.C(n_681),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_977),
.A2(n_1048),
.B(n_786),
.Y(n_1187)
);

NOR2x1_ASAP7_75t_L g1188 ( 
.A(n_983),
.B(n_712),
.Y(n_1188)
);

AOI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_929),
.A2(n_869),
.B1(n_836),
.B2(n_613),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_926),
.A2(n_762),
.B(n_698),
.Y(n_1190)
);

AO31x2_ASAP7_75t_L g1191 ( 
.A1(n_1030),
.A2(n_832),
.A3(n_1003),
.B(n_762),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_925),
.B(n_607),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_SL g1193 ( 
.A1(n_971),
.A2(n_414),
.B(n_594),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1167),
.A2(n_1175),
.B1(n_1169),
.B2(n_1192),
.Y(n_1194)
);

BUFx12f_ASAP7_75t_L g1195 ( 
.A(n_1155),
.Y(n_1195)
);

INVx2_ASAP7_75t_SL g1196 ( 
.A(n_1072),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1160),
.B(n_1170),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_1072),
.Y(n_1198)
);

INVx2_ASAP7_75t_SL g1199 ( 
.A(n_1162),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_1118),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1102),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1157),
.A2(n_1186),
.B1(n_1174),
.B2(n_1179),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_1162),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1176),
.A2(n_1159),
.B1(n_1110),
.B2(n_1189),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1129),
.A2(n_1104),
.B1(n_1153),
.B2(n_1164),
.Y(n_1205)
);

AOI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1171),
.A2(n_1193),
.B1(n_1183),
.B2(n_1067),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_1162),
.Y(n_1207)
);

NAND2x1p5_ASAP7_75t_L g1208 ( 
.A(n_1112),
.B(n_1134),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1104),
.A2(n_1094),
.B1(n_1088),
.B2(n_1139),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1161),
.A2(n_1172),
.B(n_1163),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1122),
.A2(n_1084),
.B1(n_1065),
.B2(n_1140),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1120),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_SL g1213 ( 
.A1(n_1082),
.A2(n_1168),
.B1(n_1165),
.B2(n_1090),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1177),
.B(n_1182),
.Y(n_1214)
);

BUFx2_ASAP7_75t_L g1215 ( 
.A(n_1181),
.Y(n_1215)
);

HB1xp67_ASAP7_75t_L g1216 ( 
.A(n_1071),
.Y(n_1216)
);

INVx8_ASAP7_75t_L g1217 ( 
.A(n_1117),
.Y(n_1217)
);

CKINVDCx6p67_ASAP7_75t_R g1218 ( 
.A(n_1079),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1081),
.B(n_1114),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_1073),
.Y(n_1220)
);

BUFx2_ASAP7_75t_L g1221 ( 
.A(n_1078),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_SL g1222 ( 
.A1(n_1108),
.A2(n_1119),
.B(n_1113),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_SL g1223 ( 
.A1(n_1112),
.A2(n_1134),
.B1(n_1145),
.B2(n_1149),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1112),
.A2(n_1134),
.B1(n_1066),
.B2(n_1128),
.Y(n_1224)
);

CKINVDCx11_ASAP7_75t_R g1225 ( 
.A(n_1077),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_SL g1226 ( 
.A1(n_1074),
.A2(n_1080),
.B1(n_1075),
.B2(n_1097),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1156),
.B(n_1173),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1138),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1074),
.A2(n_1131),
.B1(n_1092),
.B2(n_1070),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_SL g1230 ( 
.A1(n_1137),
.A2(n_1083),
.B1(n_1190),
.B2(n_1166),
.Y(n_1230)
);

OAI21xp33_ASAP7_75t_L g1231 ( 
.A1(n_1123),
.A2(n_1086),
.B(n_1093),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1124),
.A2(n_1142),
.B1(n_1087),
.B2(n_1150),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1158),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1148),
.A2(n_1188),
.B1(n_1147),
.B2(n_1154),
.Y(n_1234)
);

CKINVDCx20_ASAP7_75t_R g1235 ( 
.A(n_1127),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1098),
.A2(n_1111),
.B1(n_1180),
.B2(n_1185),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1109),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1152),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1117),
.Y(n_1239)
);

CKINVDCx11_ASAP7_75t_R g1240 ( 
.A(n_1106),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1089),
.A2(n_1151),
.B1(n_1063),
.B2(n_1135),
.Y(n_1241)
);

OAI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1125),
.A2(n_1143),
.B1(n_1133),
.B2(n_1132),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1117),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1116),
.B(n_1191),
.Y(n_1244)
);

OR2x2_ASAP7_75t_L g1245 ( 
.A(n_1152),
.B(n_1191),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1068),
.A2(n_1121),
.B1(n_1115),
.B2(n_1141),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1117),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1101),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_SL g1249 ( 
.A1(n_1184),
.A2(n_1115),
.B1(n_1121),
.B2(n_1099),
.Y(n_1249)
);

NAND2x1p5_ASAP7_75t_L g1250 ( 
.A(n_1144),
.B(n_1136),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_SL g1251 ( 
.A1(n_1184),
.A2(n_1126),
.B1(n_1099),
.B2(n_1107),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_SL g1252 ( 
.A1(n_1126),
.A2(n_1107),
.B1(n_1091),
.B2(n_1085),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1126),
.Y(n_1253)
);

CKINVDCx20_ASAP7_75t_R g1254 ( 
.A(n_1095),
.Y(n_1254)
);

OAI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1146),
.A2(n_1076),
.B1(n_1107),
.B2(n_1105),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1105),
.B(n_1191),
.Y(n_1256)
);

CKINVDCx11_ASAP7_75t_R g1257 ( 
.A(n_1105),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1103),
.A2(n_1100),
.B(n_1187),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1178),
.A2(n_1130),
.B1(n_1064),
.B2(n_1069),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_1069),
.Y(n_1260)
);

BUFx8_ASAP7_75t_SL g1261 ( 
.A(n_1064),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1130),
.A2(n_1186),
.B1(n_1157),
.B2(n_1174),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1176),
.B(n_603),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_SL g1264 ( 
.A1(n_1157),
.A2(n_869),
.B1(n_1186),
.B2(n_683),
.Y(n_1264)
);

CKINVDCx6p67_ASAP7_75t_R g1265 ( 
.A(n_1155),
.Y(n_1265)
);

INVxp67_ASAP7_75t_SL g1266 ( 
.A(n_1066),
.Y(n_1266)
);

INVx1_ASAP7_75t_SL g1267 ( 
.A(n_1164),
.Y(n_1267)
);

INVx6_ASAP7_75t_L g1268 ( 
.A(n_1072),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1157),
.A2(n_1186),
.B1(n_1174),
.B2(n_869),
.Y(n_1269)
);

BUFx12f_ASAP7_75t_L g1270 ( 
.A(n_1155),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1096),
.Y(n_1271)
);

INVx2_ASAP7_75t_SL g1272 ( 
.A(n_1072),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_1072),
.Y(n_1273)
);

INVx4_ASAP7_75t_L g1274 ( 
.A(n_1162),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1167),
.A2(n_1169),
.B1(n_1192),
.B2(n_1175),
.Y(n_1275)
);

AOI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1171),
.A2(n_836),
.B1(n_1193),
.B2(n_869),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_SL g1277 ( 
.A1(n_1157),
.A2(n_869),
.B1(n_1186),
.B2(n_683),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_SL g1278 ( 
.A1(n_1157),
.A2(n_869),
.B1(n_1186),
.B2(n_683),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_SL g1279 ( 
.A1(n_1157),
.A2(n_414),
.B1(n_995),
.B2(n_1186),
.Y(n_1279)
);

BUFx10_ASAP7_75t_L g1280 ( 
.A(n_1162),
.Y(n_1280)
);

BUFx12f_ASAP7_75t_L g1281 ( 
.A(n_1155),
.Y(n_1281)
);

INVx6_ASAP7_75t_L g1282 ( 
.A(n_1072),
.Y(n_1282)
);

INVx4_ASAP7_75t_L g1283 ( 
.A(n_1162),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_1117),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1167),
.B(n_925),
.Y(n_1285)
);

OAI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1193),
.A2(n_1157),
.B1(n_1186),
.B2(n_718),
.Y(n_1286)
);

CKINVDCx11_ASAP7_75t_R g1287 ( 
.A(n_1155),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1118),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1096),
.Y(n_1289)
);

OAI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1193),
.A2(n_1157),
.B1(n_1186),
.B2(n_718),
.Y(n_1290)
);

INVx2_ASAP7_75t_SL g1291 ( 
.A(n_1072),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_SL g1292 ( 
.A1(n_1157),
.A2(n_414),
.B1(n_995),
.B2(n_1186),
.Y(n_1292)
);

BUFx12f_ASAP7_75t_L g1293 ( 
.A(n_1155),
.Y(n_1293)
);

INVx4_ASAP7_75t_L g1294 ( 
.A(n_1162),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1157),
.A2(n_1186),
.B1(n_1174),
.B2(n_869),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1072),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1072),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1167),
.A2(n_1169),
.B1(n_1192),
.B2(n_1175),
.Y(n_1298)
);

OAI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1193),
.A2(n_1157),
.B1(n_1186),
.B2(n_718),
.Y(n_1299)
);

BUFx4_ASAP7_75t_SL g1300 ( 
.A(n_1118),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1157),
.A2(n_1186),
.B1(n_1174),
.B2(n_869),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_SL g1302 ( 
.A1(n_1157),
.A2(n_414),
.B1(n_995),
.B2(n_1186),
.Y(n_1302)
);

INVx1_ASAP7_75t_SL g1303 ( 
.A(n_1164),
.Y(n_1303)
);

INVx5_ASAP7_75t_L g1304 ( 
.A(n_1112),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1157),
.A2(n_1186),
.B1(n_1174),
.B2(n_869),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1157),
.A2(n_1186),
.B1(n_1174),
.B2(n_869),
.Y(n_1306)
);

INVx3_ASAP7_75t_L g1307 ( 
.A(n_1117),
.Y(n_1307)
);

INVx6_ASAP7_75t_L g1308 ( 
.A(n_1072),
.Y(n_1308)
);

BUFx3_ASAP7_75t_L g1309 ( 
.A(n_1072),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1096),
.Y(n_1310)
);

AOI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1171),
.A2(n_836),
.B1(n_1193),
.B2(n_869),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1167),
.A2(n_1169),
.B1(n_1192),
.B2(n_1175),
.Y(n_1312)
);

BUFx4f_ASAP7_75t_SL g1313 ( 
.A(n_1195),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1266),
.B(n_1194),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1254),
.B(n_1238),
.Y(n_1315)
);

NAND2x1p5_ASAP7_75t_L g1316 ( 
.A(n_1260),
.B(n_1304),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_1245),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1258),
.A2(n_1210),
.B(n_1250),
.Y(n_1318)
);

AO21x2_ASAP7_75t_L g1319 ( 
.A1(n_1255),
.A2(n_1258),
.B(n_1210),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_1250),
.Y(n_1320)
);

OR2x6_ASAP7_75t_L g1321 ( 
.A(n_1241),
.B(n_1248),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1256),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1253),
.B(n_1262),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1244),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1304),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1201),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1224),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1271),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1259),
.B(n_1251),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1246),
.A2(n_1236),
.B(n_1241),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1251),
.B(n_1289),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1310),
.Y(n_1332)
);

AND2x2_ASAP7_75t_SL g1333 ( 
.A(n_1197),
.B(n_1214),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1213),
.B(n_1197),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1227),
.Y(n_1335)
);

BUFx2_ASAP7_75t_L g1336 ( 
.A(n_1261),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1249),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1212),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1213),
.B(n_1214),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1231),
.Y(n_1340)
);

OR2x2_ASAP7_75t_L g1341 ( 
.A(n_1219),
.B(n_1216),
.Y(n_1341)
);

OA21x2_ASAP7_75t_L g1342 ( 
.A1(n_1222),
.A2(n_1232),
.B(n_1209),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1224),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1252),
.Y(n_1344)
);

OAI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1264),
.A2(n_1278),
.B(n_1277),
.Y(n_1345)
);

AO31x2_ASAP7_75t_L g1346 ( 
.A1(n_1237),
.A2(n_1219),
.A3(n_1252),
.B(n_1312),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1257),
.Y(n_1347)
);

AOI222xp33_ASAP7_75t_L g1348 ( 
.A1(n_1194),
.A2(n_1312),
.B1(n_1275),
.B2(n_1298),
.C1(n_1285),
.C2(n_1286),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1242),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1230),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1208),
.A2(n_1284),
.B(n_1307),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1230),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1267),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1206),
.B(n_1202),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1226),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1226),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1303),
.Y(n_1357)
);

CKINVDCx6p67_ASAP7_75t_R g1358 ( 
.A(n_1270),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1275),
.B(n_1298),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1228),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1234),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1263),
.B(n_1311),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1211),
.B(n_1285),
.Y(n_1363)
);

AO21x2_ASAP7_75t_L g1364 ( 
.A1(n_1290),
.A2(n_1299),
.B(n_1276),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1269),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1240),
.A2(n_1204),
.B1(n_1306),
.B2(n_1305),
.Y(n_1366)
);

AO21x2_ASAP7_75t_L g1367 ( 
.A1(n_1295),
.A2(n_1301),
.B(n_1292),
.Y(n_1367)
);

AOI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1215),
.A2(n_1221),
.B(n_1223),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1247),
.A2(n_1307),
.B(n_1284),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1279),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1279),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1292),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1302),
.B(n_1205),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1302),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1243),
.B(n_1229),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_SL g1376 ( 
.A1(n_1268),
.A2(n_1308),
.B1(n_1282),
.B2(n_1223),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1217),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1288),
.B(n_1220),
.Y(n_1378)
);

INVx2_ASAP7_75t_SL g1379 ( 
.A(n_1280),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1239),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1225),
.B(n_1203),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1203),
.Y(n_1382)
);

CKINVDCx6p67_ASAP7_75t_R g1383 ( 
.A(n_1281),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1203),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1207),
.Y(n_1385)
);

AOI222xp33_ASAP7_75t_L g1386 ( 
.A1(n_1268),
.A2(n_1308),
.B1(n_1282),
.B2(n_1287),
.C1(n_1297),
.C2(n_1309),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1207),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1274),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1274),
.B(n_1294),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1199),
.B(n_1294),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1283),
.Y(n_1391)
);

A2O1A1Ixp33_ASAP7_75t_SL g1392 ( 
.A1(n_1345),
.A2(n_1280),
.B(n_1308),
.C(n_1282),
.Y(n_1392)
);

A2O1A1Ixp33_ASAP7_75t_SL g1393 ( 
.A1(n_1345),
.A2(n_1340),
.B(n_1374),
.C(n_1372),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1318),
.A2(n_1268),
.B(n_1218),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1314),
.B(n_1233),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1315),
.B(n_1235),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_1358),
.Y(n_1397)
);

AOI221xp5_ASAP7_75t_L g1398 ( 
.A1(n_1373),
.A2(n_1196),
.B1(n_1296),
.B2(n_1291),
.C(n_1273),
.Y(n_1398)
);

OA21x2_ASAP7_75t_L g1399 ( 
.A1(n_1318),
.A2(n_1272),
.B(n_1198),
.Y(n_1399)
);

AOI221xp5_ASAP7_75t_L g1400 ( 
.A1(n_1373),
.A2(n_1200),
.B1(n_1300),
.B2(n_1265),
.C(n_1293),
.Y(n_1400)
);

O2A1O1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1359),
.A2(n_1348),
.B(n_1340),
.C(n_1354),
.Y(n_1401)
);

A2O1A1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1333),
.A2(n_1359),
.B(n_1354),
.C(n_1350),
.Y(n_1402)
);

AND4x1_ASAP7_75t_L g1403 ( 
.A(n_1386),
.B(n_1348),
.C(n_1366),
.D(n_1381),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1341),
.B(n_1314),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_1363),
.B(n_1361),
.Y(n_1405)
);

O2A1O1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1370),
.A2(n_1372),
.B(n_1374),
.C(n_1371),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1315),
.B(n_1347),
.Y(n_1407)
);

A2O1A1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1333),
.A2(n_1350),
.B(n_1352),
.C(n_1349),
.Y(n_1408)
);

A2O1A1Ixp33_ASAP7_75t_L g1409 ( 
.A1(n_1333),
.A2(n_1352),
.B(n_1349),
.C(n_1339),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1315),
.B(n_1347),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1331),
.B(n_1329),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1353),
.B(n_1357),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1361),
.A2(n_1362),
.B(n_1330),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1334),
.B(n_1339),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1336),
.A2(n_1371),
.B1(n_1370),
.B2(n_1347),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1334),
.B(n_1360),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1330),
.A2(n_1365),
.B(n_1342),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1358),
.Y(n_1418)
);

AOI221xp5_ASAP7_75t_L g1419 ( 
.A1(n_1365),
.A2(n_1356),
.B1(n_1355),
.B2(n_1364),
.C(n_1344),
.Y(n_1419)
);

AOI221xp5_ASAP7_75t_L g1420 ( 
.A1(n_1355),
.A2(n_1356),
.B1(n_1364),
.B2(n_1344),
.C(n_1367),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1331),
.B(n_1329),
.Y(n_1421)
);

NOR2x1_ASAP7_75t_SL g1422 ( 
.A(n_1368),
.B(n_1335),
.Y(n_1422)
);

AOI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1368),
.A2(n_1337),
.B(n_1327),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1319),
.A2(n_1321),
.B(n_1342),
.Y(n_1424)
);

NOR3xp33_ASAP7_75t_SL g1425 ( 
.A(n_1376),
.B(n_1380),
.C(n_1377),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1337),
.B(n_1323),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1369),
.A2(n_1351),
.B(n_1316),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1323),
.B(n_1327),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1322),
.B(n_1332),
.Y(n_1429)
);

INVx3_ASAP7_75t_L g1430 ( 
.A(n_1369),
.Y(n_1430)
);

BUFx4f_ASAP7_75t_SL g1431 ( 
.A(n_1358),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1364),
.A2(n_1367),
.B1(n_1342),
.B2(n_1376),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1343),
.B(n_1317),
.Y(n_1433)
);

AND2x2_ASAP7_75t_SL g1434 ( 
.A(n_1342),
.B(n_1343),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1322),
.B(n_1326),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1322),
.B(n_1351),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1326),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1360),
.B(n_1328),
.Y(n_1438)
);

INVx4_ASAP7_75t_L g1439 ( 
.A(n_1325),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_SL g1440 ( 
.A(n_1402),
.B(n_1375),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1429),
.B(n_1346),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1429),
.B(n_1346),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1436),
.B(n_1346),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1433),
.B(n_1404),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1436),
.B(n_1346),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1402),
.A2(n_1336),
.B1(n_1342),
.B2(n_1375),
.Y(n_1446)
);

INVx4_ASAP7_75t_L g1447 ( 
.A(n_1439),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1435),
.B(n_1346),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1430),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1435),
.B(n_1346),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1427),
.B(n_1320),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1437),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1437),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1432),
.A2(n_1364),
.B1(n_1367),
.B2(n_1375),
.Y(n_1454)
);

BUFx6f_ASAP7_75t_L g1455 ( 
.A(n_1394),
.Y(n_1455)
);

CKINVDCx20_ASAP7_75t_R g1456 ( 
.A(n_1431),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1424),
.B(n_1434),
.Y(n_1457)
);

NAND3xp33_ASAP7_75t_L g1458 ( 
.A(n_1403),
.B(n_1386),
.C(n_1338),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1434),
.B(n_1319),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1411),
.B(n_1319),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1411),
.B(n_1319),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1421),
.B(n_1324),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1405),
.B(n_1380),
.Y(n_1463)
);

NAND3xp33_ASAP7_75t_L g1464 ( 
.A(n_1458),
.B(n_1419),
.C(n_1432),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1458),
.A2(n_1367),
.B1(n_1420),
.B2(n_1413),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1452),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1460),
.B(n_1416),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1452),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1450),
.B(n_1412),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_1455),
.Y(n_1470)
);

AOI211xp5_ASAP7_75t_SL g1471 ( 
.A1(n_1446),
.A2(n_1408),
.B(n_1409),
.C(n_1415),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1443),
.B(n_1426),
.Y(n_1472)
);

NAND2x1_ASAP7_75t_L g1473 ( 
.A(n_1455),
.B(n_1399),
.Y(n_1473)
);

BUFx2_ASAP7_75t_L g1474 ( 
.A(n_1451),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1452),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1450),
.B(n_1417),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1460),
.B(n_1428),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1443),
.B(n_1426),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1443),
.B(n_1399),
.Y(n_1479)
);

AO21x2_ASAP7_75t_L g1480 ( 
.A1(n_1454),
.A2(n_1422),
.B(n_1423),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1453),
.Y(n_1481)
);

BUFx6f_ASAP7_75t_L g1482 ( 
.A(n_1455),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1446),
.A2(n_1409),
.B(n_1408),
.Y(n_1483)
);

O2A1O1Ixp5_ASAP7_75t_L g1484 ( 
.A1(n_1440),
.A2(n_1392),
.B(n_1393),
.C(n_1395),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1449),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1453),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1453),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_SL g1488 ( 
.A1(n_1459),
.A2(n_1414),
.B1(n_1396),
.B2(n_1375),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1451),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1445),
.B(n_1399),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1460),
.B(n_1438),
.Y(n_1491)
);

BUFx2_ASAP7_75t_L g1492 ( 
.A(n_1451),
.Y(n_1492)
);

NAND3xp33_ASAP7_75t_SL g1493 ( 
.A(n_1454),
.B(n_1393),
.C(n_1401),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1463),
.B(n_1407),
.Y(n_1494)
);

BUFx3_ASAP7_75t_L g1495 ( 
.A(n_1455),
.Y(n_1495)
);

BUFx3_ASAP7_75t_L g1496 ( 
.A(n_1455),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_R g1497 ( 
.A(n_1456),
.B(n_1397),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1470),
.Y(n_1498)
);

INVx1_ASAP7_75t_SL g1499 ( 
.A(n_1497),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1470),
.B(n_1451),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1474),
.B(n_1457),
.Y(n_1501)
);

OAI21xp33_ASAP7_75t_L g1502 ( 
.A1(n_1493),
.A2(n_1440),
.B(n_1457),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1467),
.B(n_1461),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1466),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1466),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1468),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1474),
.B(n_1457),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1467),
.B(n_1461),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1474),
.B(n_1459),
.Y(n_1509)
);

NOR3xp33_ASAP7_75t_L g1510 ( 
.A(n_1493),
.B(n_1392),
.C(n_1400),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1489),
.B(n_1459),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1468),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1475),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1475),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1472),
.B(n_1461),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1481),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1472),
.B(n_1448),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1485),
.Y(n_1518)
);

BUFx2_ASAP7_75t_L g1519 ( 
.A(n_1470),
.Y(n_1519)
);

AND2x4_ASAP7_75t_SL g1520 ( 
.A(n_1482),
.B(n_1447),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1489),
.B(n_1441),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1464),
.A2(n_1410),
.B1(n_1463),
.B2(n_1398),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1489),
.B(n_1441),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1481),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1469),
.B(n_1462),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1472),
.B(n_1448),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1486),
.Y(n_1527)
);

NAND2x1p5_ASAP7_75t_L g1528 ( 
.A(n_1473),
.B(n_1455),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1478),
.B(n_1448),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1486),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1492),
.B(n_1442),
.Y(n_1531)
);

INVx2_ASAP7_75t_SL g1532 ( 
.A(n_1482),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1469),
.B(n_1462),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1476),
.B(n_1444),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1476),
.B(n_1444),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1487),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1478),
.B(n_1442),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1502),
.B(n_1494),
.Y(n_1538)
);

OAI22xp33_ASAP7_75t_R g1539 ( 
.A1(n_1499),
.A2(n_1476),
.B1(n_1464),
.B2(n_1471),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1512),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1518),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1512),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1534),
.B(n_1469),
.Y(n_1543)
);

OAI32xp33_ASAP7_75t_L g1544 ( 
.A1(n_1510),
.A2(n_1465),
.A3(n_1471),
.B1(n_1495),
.B2(n_1496),
.Y(n_1544)
);

AOI21xp5_ASAP7_75t_L g1545 ( 
.A1(n_1502),
.A2(n_1483),
.B(n_1484),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1517),
.B(n_1479),
.Y(n_1546)
);

NAND3xp33_ASAP7_75t_SL g1547 ( 
.A(n_1510),
.B(n_1483),
.C(n_1484),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1517),
.B(n_1526),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1504),
.Y(n_1549)
);

INVxp67_ASAP7_75t_SL g1550 ( 
.A(n_1534),
.Y(n_1550)
);

OAI31xp33_ASAP7_75t_SL g1551 ( 
.A1(n_1499),
.A2(n_1488),
.A3(n_1494),
.B(n_1479),
.Y(n_1551)
);

INVx3_ASAP7_75t_L g1552 ( 
.A(n_1520),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1518),
.Y(n_1553)
);

NAND2x1_ASAP7_75t_L g1554 ( 
.A(n_1498),
.B(n_1482),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1522),
.B(n_1477),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1526),
.B(n_1479),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1535),
.B(n_1477),
.Y(n_1557)
);

BUFx6f_ASAP7_75t_L g1558 ( 
.A(n_1532),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1504),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1505),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1535),
.B(n_1383),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1503),
.B(n_1465),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1503),
.B(n_1478),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1525),
.B(n_1491),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1508),
.B(n_1491),
.Y(n_1565)
);

NAND4xp25_ASAP7_75t_L g1566 ( 
.A(n_1501),
.B(n_1406),
.C(n_1488),
.D(n_1495),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1505),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1520),
.B(n_1470),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1529),
.B(n_1490),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1506),
.Y(n_1570)
);

NOR2x1p5_ASAP7_75t_L g1571 ( 
.A(n_1525),
.B(n_1383),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1498),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1529),
.B(n_1537),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1506),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1537),
.B(n_1490),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1508),
.B(n_1533),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1513),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1513),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1518),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1549),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1550),
.B(n_1533),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1558),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1557),
.B(n_1536),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1543),
.B(n_1536),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1572),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1540),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1545),
.B(n_1515),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1549),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1538),
.B(n_1515),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1548),
.B(n_1521),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1559),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1555),
.B(n_1501),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1559),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1560),
.Y(n_1594)
);

OAI21xp33_ASAP7_75t_L g1595 ( 
.A1(n_1547),
.A2(n_1507),
.B(n_1501),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1548),
.B(n_1521),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1562),
.B(n_1507),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1573),
.B(n_1521),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1561),
.B(n_1507),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1551),
.B(n_1509),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1573),
.B(n_1523),
.Y(n_1601)
);

AOI21xp33_ASAP7_75t_L g1602 ( 
.A1(n_1544),
.A2(n_1554),
.B(n_1552),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1560),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1544),
.B(n_1397),
.Y(n_1604)
);

NOR2x1_ASAP7_75t_SL g1605 ( 
.A(n_1543),
.B(n_1480),
.Y(n_1605)
);

NAND4xp25_ASAP7_75t_L g1606 ( 
.A(n_1566),
.B(n_1519),
.C(n_1381),
.D(n_1511),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1577),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1552),
.B(n_1523),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1552),
.B(n_1520),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1558),
.Y(n_1610)
);

NAND2x1p5_ASAP7_75t_L g1611 ( 
.A(n_1554),
.B(n_1473),
.Y(n_1611)
);

AO22x1_ASAP7_75t_L g1612 ( 
.A1(n_1539),
.A2(n_1568),
.B1(n_1418),
.B2(n_1542),
.Y(n_1612)
);

AOI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1539),
.A2(n_1480),
.B1(n_1425),
.B2(n_1490),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1564),
.B(n_1514),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1604),
.A2(n_1571),
.B1(n_1480),
.B2(n_1568),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1585),
.Y(n_1616)
);

OAI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1604),
.A2(n_1568),
.B1(n_1564),
.B2(n_1563),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1587),
.B(n_1565),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1580),
.Y(n_1619)
);

OAI222xp33_ASAP7_75t_L g1620 ( 
.A1(n_1600),
.A2(n_1528),
.B1(n_1576),
.B2(n_1473),
.C1(n_1519),
.C2(n_1509),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1586),
.B(n_1567),
.Y(n_1621)
);

OA22x2_ASAP7_75t_L g1622 ( 
.A1(n_1613),
.A2(n_1532),
.B1(n_1570),
.B2(n_1574),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1592),
.B(n_1546),
.Y(n_1623)
);

OAI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1606),
.A2(n_1482),
.B1(n_1528),
.B2(n_1496),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1595),
.B(n_1546),
.Y(n_1625)
);

OAI21xp33_ASAP7_75t_L g1626 ( 
.A1(n_1597),
.A2(n_1511),
.B(n_1509),
.Y(n_1626)
);

AOI22x1_ASAP7_75t_L g1627 ( 
.A1(n_1609),
.A2(n_1418),
.B1(n_1528),
.B2(n_1558),
.Y(n_1627)
);

OAI32xp33_ASAP7_75t_L g1628 ( 
.A1(n_1602),
.A2(n_1528),
.A3(n_1496),
.B1(n_1495),
.B2(n_1511),
.Y(n_1628)
);

AOI221xp5_ASAP7_75t_L g1629 ( 
.A1(n_1612),
.A2(n_1589),
.B1(n_1591),
.B2(n_1593),
.C(n_1588),
.Y(n_1629)
);

INVxp67_ASAP7_75t_L g1630 ( 
.A(n_1609),
.Y(n_1630)
);

INVxp67_ASAP7_75t_L g1631 ( 
.A(n_1609),
.Y(n_1631)
);

OAI21xp33_ASAP7_75t_L g1632 ( 
.A1(n_1599),
.A2(n_1578),
.B(n_1577),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_SL g1633 ( 
.A(n_1608),
.B(n_1313),
.Y(n_1633)
);

XOR2x2_ASAP7_75t_L g1634 ( 
.A(n_1608),
.B(n_1497),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1581),
.B(n_1558),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1594),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1590),
.Y(n_1637)
);

AOI221xp5_ASAP7_75t_L g1638 ( 
.A1(n_1603),
.A2(n_1578),
.B1(n_1480),
.B2(n_1482),
.C(n_1495),
.Y(n_1638)
);

AOI21xp33_ASAP7_75t_L g1639 ( 
.A1(n_1582),
.A2(n_1480),
.B(n_1532),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1630),
.B(n_1590),
.Y(n_1640)
);

AOI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1629),
.A2(n_1633),
.B1(n_1622),
.B2(n_1617),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1622),
.A2(n_1607),
.B1(n_1610),
.B2(n_1582),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1616),
.B(n_1596),
.Y(n_1643)
);

O2A1O1Ixp5_ASAP7_75t_L g1644 ( 
.A1(n_1628),
.A2(n_1610),
.B(n_1581),
.C(n_1584),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1631),
.B(n_1596),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1634),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1637),
.Y(n_1647)
);

AOI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1629),
.A2(n_1605),
.B(n_1611),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1625),
.B(n_1583),
.Y(n_1649)
);

NAND2x1p5_ASAP7_75t_L g1650 ( 
.A(n_1627),
.B(n_1383),
.Y(n_1650)
);

OAI21xp33_ASAP7_75t_SL g1651 ( 
.A1(n_1638),
.A2(n_1601),
.B(n_1598),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1619),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1636),
.Y(n_1653)
);

OAI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1615),
.A2(n_1611),
.B(n_1583),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1618),
.B(n_1456),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1621),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1632),
.B(n_1598),
.Y(n_1657)
);

OR4x1_ASAP7_75t_L g1658 ( 
.A(n_1635),
.B(n_1379),
.C(n_1382),
.D(n_1516),
.Y(n_1658)
);

INVxp67_ASAP7_75t_L g1659 ( 
.A(n_1647),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1646),
.A2(n_1626),
.B1(n_1638),
.B2(n_1623),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1645),
.B(n_1601),
.Y(n_1661)
);

BUFx2_ASAP7_75t_L g1662 ( 
.A(n_1645),
.Y(n_1662)
);

NOR2x1_ASAP7_75t_L g1663 ( 
.A(n_1646),
.B(n_1620),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1647),
.Y(n_1664)
);

INVxp67_ASAP7_75t_SL g1665 ( 
.A(n_1643),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1640),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1652),
.Y(n_1667)
);

OAI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1641),
.A2(n_1611),
.B1(n_1624),
.B2(n_1482),
.Y(n_1668)
);

AOI211xp5_ASAP7_75t_L g1669 ( 
.A1(n_1668),
.A2(n_1648),
.B(n_1654),
.C(n_1656),
.Y(n_1669)
);

O2A1O1Ixp33_ASAP7_75t_L g1670 ( 
.A1(n_1663),
.A2(n_1644),
.B(n_1653),
.C(n_1642),
.Y(n_1670)
);

NAND4xp25_ASAP7_75t_L g1671 ( 
.A(n_1660),
.B(n_1655),
.C(n_1642),
.D(n_1649),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1662),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1661),
.Y(n_1673)
);

NAND4xp25_ASAP7_75t_L g1674 ( 
.A(n_1666),
.B(n_1655),
.C(n_1657),
.D(n_1639),
.Y(n_1674)
);

NOR2x1_ASAP7_75t_L g1675 ( 
.A(n_1664),
.B(n_1558),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1659),
.Y(n_1676)
);

NAND3xp33_ASAP7_75t_L g1677 ( 
.A(n_1659),
.B(n_1651),
.C(n_1614),
.Y(n_1677)
);

OAI221xp5_ASAP7_75t_L g1678 ( 
.A1(n_1670),
.A2(n_1650),
.B1(n_1665),
.B2(n_1667),
.C(n_1614),
.Y(n_1678)
);

OAI221xp5_ASAP7_75t_L g1679 ( 
.A1(n_1671),
.A2(n_1650),
.B1(n_1584),
.B2(n_1496),
.C(n_1482),
.Y(n_1679)
);

OAI21xp33_ASAP7_75t_L g1680 ( 
.A1(n_1674),
.A2(n_1541),
.B(n_1579),
.Y(n_1680)
);

AO21x1_ASAP7_75t_L g1681 ( 
.A1(n_1669),
.A2(n_1658),
.B(n_1579),
.Y(n_1681)
);

OAI211xp5_ASAP7_75t_L g1682 ( 
.A1(n_1677),
.A2(n_1672),
.B(n_1676),
.C(n_1675),
.Y(n_1682)
);

AOI21x1_ASAP7_75t_L g1683 ( 
.A1(n_1682),
.A2(n_1673),
.B(n_1553),
.Y(n_1683)
);

INVxp33_ASAP7_75t_L g1684 ( 
.A(n_1678),
.Y(n_1684)
);

O2A1O1Ixp5_ASAP7_75t_SL g1685 ( 
.A1(n_1679),
.A2(n_1658),
.B(n_1514),
.C(n_1516),
.Y(n_1685)
);

AOI221xp5_ASAP7_75t_L g1686 ( 
.A1(n_1680),
.A2(n_1482),
.B1(n_1541),
.B2(n_1553),
.C(n_1556),
.Y(n_1686)
);

OAI211xp5_ASAP7_75t_L g1687 ( 
.A1(n_1681),
.A2(n_1378),
.B(n_1379),
.C(n_1492),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1678),
.A2(n_1500),
.B(n_1569),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1683),
.Y(n_1689)
);

AND2x4_ASAP7_75t_L g1690 ( 
.A(n_1688),
.B(n_1500),
.Y(n_1690)
);

NAND4xp75_ASAP7_75t_L g1691 ( 
.A(n_1684),
.B(n_1379),
.C(n_1390),
.D(n_1556),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1687),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1686),
.B(n_1500),
.Y(n_1693)
);

OAI211xp5_ASAP7_75t_SL g1694 ( 
.A1(n_1689),
.A2(n_1685),
.B(n_1382),
.C(n_1377),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_SL g1695 ( 
.A(n_1692),
.B(n_1500),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1691),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1696),
.B(n_1690),
.Y(n_1697)
);

AOI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1697),
.A2(n_1695),
.B1(n_1690),
.B2(n_1691),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1698),
.Y(n_1699)
);

CKINVDCx16_ASAP7_75t_R g1700 ( 
.A(n_1699),
.Y(n_1700)
);

AOI221xp5_ASAP7_75t_L g1701 ( 
.A1(n_1700),
.A2(n_1694),
.B1(n_1693),
.B2(n_1530),
.C(n_1524),
.Y(n_1701)
);

AOI22xp33_ASAP7_75t_SL g1702 ( 
.A1(n_1701),
.A2(n_1575),
.B1(n_1569),
.B2(n_1492),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1701),
.A2(n_1575),
.B(n_1389),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1702),
.A2(n_1531),
.B1(n_1523),
.B2(n_1389),
.Y(n_1704)
);

OAI21x1_ASAP7_75t_SL g1705 ( 
.A1(n_1703),
.A2(n_1388),
.B(n_1391),
.Y(n_1705)
);

OAI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1704),
.A2(n_1530),
.B1(n_1527),
.B2(n_1524),
.Y(n_1706)
);

AOI221xp5_ASAP7_75t_L g1707 ( 
.A1(n_1706),
.A2(n_1705),
.B1(n_1527),
.B2(n_1390),
.C(n_1531),
.Y(n_1707)
);

AOI211xp5_ASAP7_75t_L g1708 ( 
.A1(n_1707),
.A2(n_1385),
.B(n_1384),
.C(n_1387),
.Y(n_1708)
);


endmodule