module fake_jpeg_15755_n_62 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_62);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_62;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_7),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_0),
.B(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_17),
.B(n_18),
.Y(n_23)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_13),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_20),
.B(n_13),
.Y(n_25)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_14),
.Y(n_24)
);

NOR2x1_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_18),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_8),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_16),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_30),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_22),
.A2(n_21),
.B1(n_8),
.B2(n_12),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_23),
.A2(n_16),
.B1(n_12),
.B2(n_11),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_15),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_19),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_26),
.A2(n_10),
.B(n_11),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_10),
.B(n_15),
.Y(n_40)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_33),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_29),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_44),
.A2(n_46),
.B(n_47),
.Y(n_50)
);

XOR2x2_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_31),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_32),
.B1(n_34),
.B2(n_19),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_SL g52 ( 
.A1(n_48),
.A2(n_37),
.B(n_36),
.C(n_15),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_45),
.A2(n_34),
.B1(n_40),
.B2(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

AO22x1_ASAP7_75t_SL g51 ( 
.A1(n_46),
.A2(n_41),
.B1(n_14),
.B2(n_19),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_51),
.A2(n_52),
.B1(n_43),
.B2(n_15),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_48),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_0),
.C(n_2),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_55),
.A2(n_52),
.B1(n_44),
.B2(n_15),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_56),
.B(n_3),
.Y(n_59)
);

MAJx2_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_53),
.C(n_54),
.Y(n_58)
);

BUFx24_ASAP7_75t_SL g60 ( 
.A(n_58),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_59),
.B1(n_5),
.B2(n_6),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_5),
.Y(n_62)
);


endmodule