module fake_jpeg_21904_n_132 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx2_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_10),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_30),
.B(n_33),
.Y(n_53)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_23),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_15),
.B1(n_25),
.B2(n_21),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_3),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_36),
.B(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_27),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_17),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_29),
.B(n_19),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_54),
.Y(n_64)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_50),
.A2(n_27),
.B1(n_40),
.B2(n_6),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_25),
.Y(n_51)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_16),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_35),
.B(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_57),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_27),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_31),
.A2(n_27),
.B(n_17),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_4),
.B(n_5),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_28),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_11),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_24),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_81),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_33),
.C(n_39),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_74),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_67),
.B(n_79),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g68 ( 
.A1(n_49),
.A2(n_10),
.B(n_13),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_68),
.A2(n_71),
.B(n_73),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_40),
.B(n_5),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_6),
.C(n_7),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_78),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_6),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_50),
.A2(n_11),
.B1(n_58),
.B2(n_45),
.Y(n_81)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_64),
.B(n_57),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_71),
.C(n_79),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_64),
.B(n_42),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_92),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_53),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_66),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_93),
.A2(n_88),
.B(n_86),
.Y(n_99)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_72),
.Y(n_104)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_56),
.C(n_42),
.Y(n_95)
);

AOI21xp33_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_72),
.B(n_60),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_99),
.C(n_101),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_55),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_81),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_69),
.C(n_74),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_105),
.C(n_82),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_88),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_86),
.B(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_114),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_113),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_99),
.B(n_86),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_98),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_91),
.B1(n_85),
.B2(n_89),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_70),
.B1(n_87),
.B2(n_56),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_105),
.C(n_103),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_83),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_104),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_112),
.A2(n_101),
.B1(n_106),
.B2(n_102),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_115),
.A2(n_47),
.B1(n_62),
.B2(n_100),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_118),
.C(n_111),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_69),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_117),
.C(n_116),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_111),
.Y(n_122)
);

OAI21x1_ASAP7_75t_SL g126 ( 
.A1(n_122),
.A2(n_123),
.B(n_115),
.Y(n_126)
);

OAI21x1_ASAP7_75t_L g123 ( 
.A1(n_120),
.A2(n_73),
.B(n_109),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_125),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_127),
.C(n_121),
.Y(n_129)
);

AOI322xp5_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_130),
.A3(n_48),
.B1(n_77),
.B2(n_127),
.C1(n_124),
.C2(n_119),
.Y(n_131)
);

OAI31xp33_ASAP7_75t_L g130 ( 
.A1(n_128),
.A2(n_122),
.A3(n_77),
.B(n_76),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_48),
.Y(n_132)
);


endmodule