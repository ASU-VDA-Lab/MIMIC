module fake_jpeg_65_n_158 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_158);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

NOR2xp67_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_55),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_60),
.B(n_45),
.Y(n_71)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_60),
.A2(n_58),
.B1(n_56),
.B2(n_55),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_63),
.A2(n_41),
.B1(n_59),
.B2(n_43),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_59),
.A2(n_41),
.B1(n_53),
.B2(n_52),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_71),
.Y(n_78)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_48),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_70),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_76),
.B(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_72),
.B1(n_50),
.B2(n_46),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_70),
.Y(n_80)
);

BUFx8_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_87),
.Y(n_93)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_51),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_1),
.Y(n_101)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_61),
.C(n_62),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_20),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_81),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_94),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_74),
.A2(n_62),
.B1(n_88),
.B2(n_85),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_92),
.A2(n_95),
.B1(n_39),
.B2(n_36),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_81),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_47),
.B(n_72),
.Y(n_96)
);

NOR2x1_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_78),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_72),
.B1(n_50),
.B2(n_49),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_100),
.B1(n_78),
.B2(n_3),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_84),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_103),
.Y(n_112)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_96),
.A2(n_87),
.B1(n_78),
.B2(n_22),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_106),
.Y(n_128)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_109),
.A2(n_113),
.B1(n_99),
.B2(n_9),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_2),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_116),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_24),
.B1(n_38),
.B2(n_37),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_115),
.B1(n_8),
.B2(n_9),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_102),
.B(n_4),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_34),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_121),
.C(n_100),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_6),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_119),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_90),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_120),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_32),
.C(n_31),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_126),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_113),
.B1(n_112),
.B2(n_121),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_30),
.B(n_28),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_125),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_108),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_127),
.B(n_131),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_107),
.A2(n_10),
.B(n_11),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_129),
.A2(n_105),
.B(n_15),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_27),
.C(n_26),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_134),
.Y(n_138)
);

AO221x1_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_25),
.C(n_13),
.Y(n_134)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_141),
.B(n_142),
.C(n_129),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_140),
.B(n_128),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_143),
.B(n_144),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_128),
.C(n_122),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_146),
.C(n_136),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_130),
.C(n_134),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_149),
.B(n_150),
.C(n_135),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_137),
.C(n_142),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_152),
.A2(n_126),
.B1(n_148),
.B2(n_133),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_123),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_12),
.B(n_15),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_16),
.C(n_17),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_17),
.B(n_18),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_18),
.Y(n_158)
);


endmodule