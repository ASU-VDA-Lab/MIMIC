module fake_netlist_5_463_n_431 (n_10, n_24, n_61, n_75, n_65, n_74, n_57, n_37, n_31, n_13, n_66, n_60, n_16, n_43, n_0, n_58, n_9, n_69, n_18, n_42, n_22, n_1, n_45, n_46, n_21, n_38, n_4, n_35, n_73, n_17, n_19, n_30, n_5, n_33, n_14, n_23, n_29, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_62, n_71, n_59, n_26, n_55, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_36, n_76, n_27, n_64, n_28, n_70, n_68, n_72, n_32, n_41, n_56, n_51, n_63, n_11, n_7, n_15, n_48, n_50, n_52, n_431);

input n_10;
input n_24;
input n_61;
input n_75;
input n_65;
input n_74;
input n_57;
input n_37;
input n_31;
input n_13;
input n_66;
input n_60;
input n_16;
input n_43;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_42;
input n_22;
input n_1;
input n_45;
input n_46;
input n_21;
input n_38;
input n_4;
input n_35;
input n_73;
input n_17;
input n_19;
input n_30;
input n_5;
input n_33;
input n_14;
input n_23;
input n_29;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_62;
input n_71;
input n_59;
input n_26;
input n_55;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_36;
input n_76;
input n_27;
input n_64;
input n_28;
input n_70;
input n_68;
input n_72;
input n_32;
input n_41;
input n_56;
input n_51;
input n_63;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;

output n_431;

wire n_137;
wire n_294;
wire n_318;
wire n_419;
wire n_380;
wire n_82;
wire n_194;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_124;
wire n_86;
wire n_146;
wire n_136;
wire n_315;
wire n_268;
wire n_408;
wire n_376;
wire n_127;
wire n_235;
wire n_226;
wire n_353;
wire n_351;
wire n_367;
wire n_397;
wire n_111;
wire n_155;
wire n_116;
wire n_423;
wire n_284;
wire n_245;
wire n_139;
wire n_105;
wire n_280;
wire n_378;
wire n_382;
wire n_254;
wire n_302;
wire n_265;
wire n_293;
wire n_372;
wire n_244;
wire n_173;
wire n_198;
wire n_247;
wire n_314;
wire n_368;
wire n_321;
wire n_292;
wire n_100;
wire n_417;
wire n_212;
wire n_385;
wire n_119;
wire n_275;
wire n_252;
wire n_295;
wire n_133;
wire n_330;
wire n_147;
wire n_373;
wire n_307;
wire n_87;
wire n_150;
wire n_106;
wire n_209;
wire n_259;
wire n_375;
wire n_301;
wire n_93;
wire n_186;
wire n_134;
wire n_191;
wire n_171;
wire n_153;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_260;
wire n_298;
wire n_320;
wire n_286;
wire n_122;
wire n_282;
wire n_331;
wire n_406;
wire n_325;
wire n_132;
wire n_90;
wire n_101;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_371;
wire n_152;
wire n_317;
wire n_323;
wire n_195;
wire n_356;
wire n_227;
wire n_271;
wire n_94;
wire n_335;
wire n_123;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_297;
wire n_156;
wire n_225;
wire n_377;
wire n_219;
wire n_157;
wire n_131;
wire n_192;
wire n_223;
wire n_392;
wire n_158;
wire n_138;
wire n_264;
wire n_109;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_95;
wire n_185;
wire n_183;
wire n_243;
wire n_398;
wire n_396;
wire n_347;
wire n_169;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_290;
wire n_221;
wire n_178;
wire n_386;
wire n_287;
wire n_344;
wire n_422;
wire n_104;
wire n_415;
wire n_141;
wire n_355;
wire n_336;
wire n_145;
wire n_337;
wire n_430;
wire n_313;
wire n_88;
wire n_216;
wire n_168;
wire n_395;
wire n_164;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_328;
wire n_140;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_241;
wire n_357;
wire n_184;
wire n_78;
wire n_144;
wire n_114;
wire n_96;
wire n_165;
wire n_213;
wire n_129;
wire n_342;
wire n_98;
wire n_361;
wire n_363;
wire n_413;
wire n_402;
wire n_197;
wire n_107;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_384;
wire n_80;
wire n_277;
wire n_92;
wire n_338;
wire n_149;
wire n_333;
wire n_309;
wire n_84;
wire n_130;
wire n_322;
wire n_258;
wire n_79;
wire n_151;
wire n_306;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_112;
wire n_85;
wire n_239;
wire n_420;
wire n_310;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_102;
wire n_77;
wire n_161;
wire n_273;
wire n_349;
wire n_270;
wire n_230;
wire n_81;
wire n_118;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_172;
wire n_206;
wire n_217;
wire n_312;
wire n_429;
wire n_345;
wire n_210;
wire n_365;
wire n_91;
wire n_176;
wire n_182;
wire n_143;
wire n_83;
wire n_354;
wire n_237;
wire n_425;
wire n_407;
wire n_180;
wire n_340;
wire n_207;
wire n_346;
wire n_393;
wire n_229;
wire n_108;
wire n_177;
wire n_403;
wire n_421;
wire n_405;
wire n_359;
wire n_117;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_113;
wire n_246;
wire n_179;
wire n_125;
wire n_410;
wire n_269;
wire n_128;
wire n_285;
wire n_412;
wire n_120;
wire n_232;
wire n_327;
wire n_135;
wire n_126;
wire n_202;
wire n_266;
wire n_272;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_426;
wire n_409;
wire n_154;
wire n_148;
wire n_300;
wire n_159;
wire n_334;
wire n_391;
wire n_175;
wire n_262;
wire n_238;
wire n_99;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_121;
wire n_242;
wire n_360;
wire n_200;
wire n_162;
wire n_222;
wire n_89;
wire n_115;
wire n_324;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_103;
wire n_348;
wire n_97;
wire n_166;
wire n_424;
wire n_256;
wire n_305;
wire n_278;
wire n_110;

INVx1_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

NOR2xp67_ASAP7_75t_L g79 ( 
.A(n_37),
.B(n_52),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_71),
.Y(n_80)
);

CKINVDCx5p33_ASAP7_75t_R g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_16),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_64),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_23),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

CKINVDCx5p33_ASAP7_75t_R g89 ( 
.A(n_3),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_49),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVxp67_ASAP7_75t_SL g93 ( 
.A(n_13),
.Y(n_93)
);

CKINVDCx5p33_ASAP7_75t_R g94 ( 
.A(n_8),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_43),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_20),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_29),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_63),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_4),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g103 ( 
.A(n_7),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_6),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_4),
.Y(n_106)
);

NOR2xp67_ASAP7_75t_L g107 ( 
.A(n_60),
.B(n_18),
.Y(n_107)
);

CKINVDCx5p33_ASAP7_75t_R g108 ( 
.A(n_57),
.Y(n_108)
);

CKINVDCx5p33_ASAP7_75t_R g109 ( 
.A(n_31),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_39),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_3),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_56),
.Y(n_115)
);

BUFx10_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_2),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_11),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_28),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_32),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_14),
.Y(n_121)
);

AND2x4_ASAP7_75t_L g122 ( 
.A(n_25),
.B(n_26),
.Y(n_122)
);

NOR2xp67_ASAP7_75t_L g123 ( 
.A(n_15),
.B(n_41),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_10),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_50),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_8),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_51),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_46),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_48),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_30),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_44),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_14),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_21),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_13),
.Y(n_137)
);

BUFx8_ASAP7_75t_SL g138 ( 
.A(n_66),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_35),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_72),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_7),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_12),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_0),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_1),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_1),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_19),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_137),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_143),
.Y(n_149)
);

AND2x4_ASAP7_75t_L g150 ( 
.A(n_102),
.B(n_36),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_95),
.B(n_5),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_9),
.B1(n_12),
.B2(n_17),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_27),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_112),
.Y(n_157)
);

AND2x4_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_42),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_92),
.B(n_67),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_104),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

AND2x4_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_69),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_125),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_118),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

AND2x4_ASAP7_75t_L g169 ( 
.A(n_122),
.B(n_75),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_141),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_116),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_121),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_77),
.Y(n_174)
);

BUFx8_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_127),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_78),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_86),
.A2(n_126),
.B1(n_94),
.B2(n_103),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_82),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_89),
.Y(n_180)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_87),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_83),
.Y(n_182)
);

OAI21x1_ASAP7_75t_L g183 ( 
.A1(n_84),
.A2(n_147),
.B(n_113),
.Y(n_183)
);

AND2x6_ASAP7_75t_L g184 ( 
.A(n_88),
.B(n_97),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_90),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_106),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_99),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_145),
.A2(n_146),
.B1(n_134),
.B2(n_93),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_105),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_123),
.B(n_117),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_110),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_111),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_128),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_129),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_100),
.B(n_135),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_130),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_80),
.A2(n_115),
.B1(n_140),
.B2(n_91),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_132),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_136),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_87),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_81),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_80),
.A2(n_115),
.B1(n_85),
.B2(n_91),
.Y(n_202)
);

AND2x4_ASAP7_75t_L g203 ( 
.A(n_79),
.B(n_107),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_85),
.A2(n_133),
.B1(n_131),
.B2(n_108),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_96),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_98),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_109),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_157),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g209 ( 
.A(n_203),
.Y(n_209)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_157),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_200),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_154),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_149),
.Y(n_213)
);

AND2x4_ASAP7_75t_L g214 ( 
.A(n_158),
.B(n_119),
.Y(n_214)
);

OR2x6_ASAP7_75t_L g215 ( 
.A(n_165),
.B(n_138),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_120),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_156),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_139),
.Y(n_218)
);

OR2x6_ASAP7_75t_L g219 ( 
.A(n_165),
.B(n_152),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_151),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_178),
.A2(n_204),
.B1(n_188),
.B2(n_190),
.Y(n_221)
);

INVxp33_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_168),
.B(n_171),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_158),
.B(n_164),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_171),
.B(n_207),
.Y(n_225)
);

NAND3xp33_ASAP7_75t_L g226 ( 
.A(n_170),
.B(n_193),
.C(n_185),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_157),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_160),
.Y(n_228)
);

AND2x4_ASAP7_75t_L g229 ( 
.A(n_158),
.B(n_164),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_160),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_207),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_166),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_166),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_181),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_164),
.B(n_169),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_169),
.A2(n_186),
.B1(n_180),
.B2(n_155),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_166),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_172),
.Y(n_238)
);

BUFx4f_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_206),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_206),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_180),
.B(n_186),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_172),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_174),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_153),
.Y(n_245)
);

AND2x4_ASAP7_75t_L g246 ( 
.A(n_150),
.B(n_183),
.Y(n_246)
);

NAND2xp33_ASAP7_75t_SL g247 ( 
.A(n_161),
.B(n_173),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_245),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_216),
.B(n_182),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_184),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_224),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_228),
.Y(n_254)
);

BUFx8_ASAP7_75t_L g255 ( 
.A(n_212),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_199),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_233),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_211),
.B(n_197),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_184),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_198),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_220),
.A2(n_184),
.B1(n_175),
.B2(n_187),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_242),
.Y(n_262)
);

INVxp33_ASAP7_75t_L g263 ( 
.A(n_220),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_213),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_237),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_225),
.B(n_192),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_218),
.B(n_191),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_237),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_209),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_231),
.B(n_194),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_177),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_210),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_L g274 ( 
.A1(n_221),
.A2(n_176),
.B1(n_163),
.B2(n_159),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_208),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_240),
.B(n_223),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_236),
.B(n_179),
.Y(n_277)
);

INVx8_ASAP7_75t_L g278 ( 
.A(n_215),
.Y(n_278)
);

NOR2xp67_ASAP7_75t_L g279 ( 
.A(n_226),
.B(n_189),
.Y(n_279)
);

AND2x4_ASAP7_75t_L g280 ( 
.A(n_234),
.B(n_167),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_246),
.B(n_177),
.Y(n_281)
);

OR2x6_ASAP7_75t_L g282 ( 
.A(n_215),
.B(n_162),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_209),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_253),
.A2(n_214),
.B1(n_219),
.B2(n_239),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_253),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_247),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_247),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_251),
.Y(n_288)
);

AND2x4_ASAP7_75t_L g289 ( 
.A(n_250),
.B(n_219),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_248),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_280),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_265),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_260),
.B(n_230),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_277),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_255),
.B(n_148),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_148),
.Y(n_296)
);

A2O1A1Ixp33_ASAP7_75t_L g297 ( 
.A1(n_259),
.A2(n_281),
.B(n_256),
.C(n_252),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_258),
.B(n_208),
.Y(n_299)
);

AND2x4_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_217),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_249),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_267),
.B(n_196),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_254),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_261),
.B(n_238),
.Y(n_304)
);

OR2x6_ASAP7_75t_L g305 ( 
.A(n_278),
.B(n_282),
.Y(n_305)
);

AO32x1_ASAP7_75t_L g306 ( 
.A1(n_257),
.A2(n_264),
.A3(n_275),
.B1(n_269),
.B2(n_266),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_273),
.B(n_232),
.Y(n_307)
);

NOR2xp67_ASAP7_75t_L g308 ( 
.A(n_278),
.B(n_238),
.Y(n_308)
);

BUFx4f_ASAP7_75t_L g309 ( 
.A(n_278),
.Y(n_309)
);

NAND2x1p5_ASAP7_75t_L g310 ( 
.A(n_262),
.B(n_244),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_276),
.B(n_235),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_283),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_287),
.B(n_294),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_301),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_284),
.A2(n_302),
.B1(n_297),
.B2(n_299),
.Y(n_315)
);

CKINVDCx6p67_ASAP7_75t_R g316 ( 
.A(n_305),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_303),
.Y(n_317)
);

NAND2x1p5_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_291),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_292),
.Y(n_319)
);

AO21x2_ASAP7_75t_L g320 ( 
.A1(n_304),
.A2(n_307),
.B(n_293),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_300),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_298),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_289),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_298),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_290),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_296),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_305),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_306),
.A2(n_309),
.B(n_295),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_309),
.B(n_306),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_301),
.Y(n_330)
);

AOI221xp5_ASAP7_75t_L g331 ( 
.A1(n_286),
.A2(n_263),
.B1(n_220),
.B2(n_274),
.C(n_195),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_301),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_283),
.B(n_263),
.Y(n_333)
);

NAND3x1_ASAP7_75t_L g334 ( 
.A(n_296),
.B(n_202),
.C(n_197),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_301),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_311),
.B(n_285),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_309),
.B(n_80),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_311),
.B(n_285),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_288),
.Y(n_339)
);

AND2x4_ASAP7_75t_L g340 ( 
.A(n_298),
.B(n_308),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_298),
.B(n_262),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_288),
.B(n_263),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_301),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_301),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_301),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_301),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_342),
.B(n_339),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_317),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_315),
.A2(n_313),
.B(n_336),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_338),
.B(n_331),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_335),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_323),
.Y(n_352)
);

OR2x2_ASAP7_75t_L g353 ( 
.A(n_312),
.B(n_333),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_343),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_344),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_314),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_316),
.Y(n_357)
);

AND2x6_ASAP7_75t_L g358 ( 
.A(n_329),
.B(n_322),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_330),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_332),
.Y(n_360)
);

AND2x4_ASAP7_75t_L g361 ( 
.A(n_340),
.B(n_327),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_345),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_346),
.B(n_319),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_327),
.Y(n_364)
);

CKINVDCx11_ASAP7_75t_R g365 ( 
.A(n_324),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_324),
.B(n_337),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_321),
.B(n_326),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_365),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_348),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_350),
.B(n_320),
.Y(n_370)
);

OR2x6_ASAP7_75t_L g371 ( 
.A(n_349),
.B(n_328),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_347),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_347),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_351),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_354),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_355),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_363),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_356),
.Y(n_378)
);

OR2x2_ASAP7_75t_L g379 ( 
.A(n_353),
.B(n_318),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_359),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_361),
.B(n_340),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_360),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_352),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_353),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_366),
.B(n_325),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_362),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_373),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_379),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g389 ( 
.A(n_379),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_370),
.B(n_371),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_381),
.B(n_361),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_377),
.B(n_358),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_369),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_385),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_390),
.B(n_385),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_390),
.B(n_384),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_390),
.B(n_375),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_393),
.Y(n_398)
);

NAND4xp25_ASAP7_75t_L g399 ( 
.A(n_387),
.B(n_372),
.C(n_367),
.D(n_374),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_386),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_393),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_388),
.B(n_386),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_388),
.B(n_382),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_389),
.B(n_383),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_396),
.B(n_389),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_396),
.B(n_394),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_399),
.A2(n_334),
.B1(n_391),
.B2(n_381),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_400),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_398),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_395),
.B(n_394),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_401),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g412 ( 
.A(n_406),
.B(n_395),
.Y(n_412)
);

INVx2_ASAP7_75t_SL g413 ( 
.A(n_410),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_407),
.B(n_404),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_411),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_414),
.B(n_408),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_413),
.B(n_408),
.Y(n_417)
);

O2A1O1Ixp5_ASAP7_75t_L g418 ( 
.A1(n_415),
.A2(n_405),
.B(n_409),
.C(n_402),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_417),
.B(n_357),
.Y(n_419)
);

OAI211xp5_ASAP7_75t_SL g420 ( 
.A1(n_419),
.A2(n_416),
.B(n_418),
.C(n_412),
.Y(n_420)
);

NOR3xp33_ASAP7_75t_L g421 ( 
.A(n_420),
.B(n_368),
.C(n_365),
.Y(n_421)
);

NAND4xp25_ASAP7_75t_L g422 ( 
.A(n_421),
.B(n_368),
.C(n_364),
.D(n_403),
.Y(n_422)
);

NOR2x1_ASAP7_75t_L g423 ( 
.A(n_422),
.B(n_357),
.Y(n_423)
);

NAND3xp33_ASAP7_75t_L g424 ( 
.A(n_422),
.B(n_364),
.C(n_392),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_423),
.B(n_397),
.Y(n_425)
);

NOR2xp67_ASAP7_75t_L g426 ( 
.A(n_425),
.B(n_424),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_426),
.B(n_397),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_427),
.A2(n_361),
.B(n_381),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_428),
.B(n_376),
.Y(n_429)
);

AOI21xp33_ASAP7_75t_L g430 ( 
.A1(n_429),
.A2(n_341),
.B(n_382),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_430),
.A2(n_381),
.B1(n_380),
.B2(n_378),
.Y(n_431)
);


endmodule