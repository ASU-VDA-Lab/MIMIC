module fake_jpeg_9137_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_40),
.Y(n_67)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_46),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_18),
.B(n_0),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_55),
.B(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_20),
.B1(n_35),
.B2(n_30),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_57),
.A2(n_43),
.B1(n_35),
.B2(n_47),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_17),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_58),
.B(n_60),
.Y(n_95)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_39),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_70),
.B(n_80),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_72),
.Y(n_106)
);

AO22x2_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_38),
.B1(n_47),
.B2(n_41),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_41),
.B1(n_66),
.B2(n_52),
.Y(n_103)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_76),
.Y(n_110)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_78),
.Y(n_120)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_18),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_82),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_50),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_53),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_89),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_84),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_86),
.Y(n_125)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_91),
.A2(n_94),
.B1(n_66),
.B2(n_30),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_92),
.A2(n_24),
.B1(n_20),
.B2(n_22),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_50),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_97),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_62),
.A2(n_30),
.B1(n_24),
.B2(n_20),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_62),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_31),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_31),
.Y(n_113)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_101),
.B(n_104),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_76),
.B1(n_74),
.B2(n_91),
.Y(n_133)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

OAI22x1_ASAP7_75t_L g151 ( 
.A1(n_105),
.A2(n_23),
.B1(n_36),
.B2(n_26),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_111),
.B(n_112),
.Y(n_156)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_114),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_61),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_116),
.A2(n_87),
.B1(n_71),
.B2(n_25),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_70),
.B(n_48),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_84),
.B(n_86),
.Y(n_137)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_127),
.B1(n_128),
.B2(n_81),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_80),
.B(n_17),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_121),
.B(n_123),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_80),
.B(n_28),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_70),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_129),
.B(n_130),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_73),
.B(n_24),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_142),
.B(n_153),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_133),
.A2(n_138),
.B1(n_151),
.B2(n_102),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_134),
.B(n_122),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_137),
.A2(n_144),
.B(n_147),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_83),
.B1(n_87),
.B2(n_90),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_139),
.A2(n_148),
.B1(n_157),
.B2(n_125),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_128),
.A2(n_83),
.B1(n_75),
.B2(n_42),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_102),
.B1(n_100),
.B2(n_124),
.Y(n_173)
);

BUFx8_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_126),
.A2(n_25),
.B(n_34),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_SL g144 ( 
.A1(n_114),
.A2(n_88),
.B(n_85),
.C(n_98),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_150),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_118),
.A2(n_113),
.B(n_101),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_116),
.A2(n_78),
.B1(n_71),
.B2(n_34),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_117),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_31),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_154),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_106),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_29),
.Y(n_154)
);

OAI32xp33_ASAP7_75t_L g155 ( 
.A1(n_106),
.A2(n_23),
.A3(n_32),
.B1(n_36),
.B2(n_26),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_124),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_103),
.A2(n_28),
.B1(n_32),
.B2(n_37),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_158),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_161),
.A2(n_173),
.B1(n_186),
.B2(n_184),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_164),
.B(n_166),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_154),
.A2(n_109),
.B(n_123),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_165),
.A2(n_172),
.B(n_177),
.Y(n_222)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_167),
.A2(n_187),
.B1(n_188),
.B2(n_143),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_168),
.B(n_192),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_121),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_181),
.C(n_182),
.Y(n_199)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_175),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

OA21x2_ASAP7_75t_L g172 ( 
.A1(n_129),
.A2(n_122),
.B(n_125),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_135),
.B(n_111),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_137),
.A2(n_142),
.B(n_153),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_134),
.B(n_100),
.Y(n_180)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_115),
.C(n_104),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_131),
.B(n_112),
.C(n_108),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_130),
.B(n_33),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_189),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_139),
.A2(n_23),
.B(n_32),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_186),
.A2(n_21),
.B(n_158),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_157),
.A2(n_108),
.B1(n_33),
.B2(n_29),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_151),
.A2(n_33),
.B1(n_29),
.B2(n_23),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_144),
.B(n_33),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_191),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_144),
.B(n_33),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_149),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_190),
.A2(n_143),
.B1(n_136),
.B2(n_141),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_194),
.A2(n_220),
.B1(n_187),
.B2(n_172),
.Y(n_226)
);

AO22x1_ASAP7_75t_L g196 ( 
.A1(n_189),
.A2(n_191),
.B1(n_172),
.B2(n_176),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_182),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_197),
.A2(n_208),
.B1(n_183),
.B2(n_188),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_29),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_204),
.C(n_213),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_203),
.A2(n_212),
.B1(n_216),
.B2(n_165),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_141),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_159),
.A2(n_21),
.B(n_1),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_3),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_180),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_209),
.B(n_210),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_175),
.B(n_158),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_159),
.A2(n_9),
.B1(n_10),
.B2(n_15),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_170),
.B(n_158),
.C(n_21),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_21),
.C(n_1),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_217),
.C(n_3),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_173),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_0),
.C(n_2),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_167),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_219),
.A2(n_171),
.B1(n_162),
.B2(n_166),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_168),
.A2(n_178),
.B1(n_162),
.B2(n_172),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_163),
.B(n_9),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_221),
.B(n_10),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_223),
.A2(n_233),
.B1(n_247),
.B2(n_202),
.Y(n_254)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_193),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_227),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_225),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_226),
.A2(n_231),
.B1(n_232),
.B2(n_238),
.Y(n_262)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_193),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_206),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_228),
.B(n_230),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_169),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_235),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_194),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_218),
.A2(n_192),
.B1(n_163),
.B2(n_160),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_3),
.Y(n_234)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_234),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_9),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_198),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_239),
.A2(n_208),
.B(n_196),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_241),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_198),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_199),
.B(n_7),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_248),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_205),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_195),
.B(n_4),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_246),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_199),
.B(n_4),
.C(n_5),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_217),
.C(n_222),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_220),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_218),
.A2(n_5),
.B1(n_6),
.B2(n_12),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_6),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_258),
.C(n_266),
.Y(n_283)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_222),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_256),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_214),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_228),
.A2(n_215),
.B1(n_201),
.B2(n_196),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_257),
.A2(n_227),
.B(n_224),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_213),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_260),
.A2(n_223),
.B(n_237),
.Y(n_281)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_261),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_233),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_239),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_203),
.Y(n_266)
);

FAx1_ASAP7_75t_SL g267 ( 
.A(n_241),
.B(n_219),
.CI(n_212),
.CON(n_267),
.SN(n_267)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_267),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_245),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_270),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_226),
.B(n_6),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_252),
.Y(n_272)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_272),
.Y(n_296)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_269),
.Y(n_273)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_273),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_274),
.Y(n_295)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_277),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_265),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_262),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_280),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_270),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_282),
.Y(n_288)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_257),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_248),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_235),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_253),
.C(n_250),
.Y(n_290)
);

XOR2x2_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_264),
.Y(n_289)
);

OAI21x1_ASAP7_75t_L g311 ( 
.A1(n_289),
.A2(n_250),
.B(n_12),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_300),
.C(n_275),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_255),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_249),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_274),
.A2(n_251),
.B1(n_263),
.B2(n_267),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_294),
.A2(n_301),
.B1(n_302),
.B2(n_13),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_272),
.A2(n_247),
.B1(n_256),
.B2(n_258),
.Y(n_297)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_297),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_271),
.C(n_287),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_249),
.C(n_285),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_278),
.A2(n_244),
.B1(n_234),
.B2(n_243),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_281),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_283),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_306),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_308),
.C(n_312),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_307),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_286),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_273),
.C(n_286),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_276),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_309),
.Y(n_321)
);

NOR2xp67_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_284),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_311),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_12),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_313),
.A2(n_302),
.B1(n_296),
.B2(n_298),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_15),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_14),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_317),
.B(n_322),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_314),
.A2(n_291),
.B(n_295),
.Y(n_318)
);

A2O1A1Ixp33_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_312),
.B(n_305),
.C(n_304),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_315),
.A2(n_297),
.B1(n_288),
.B2(n_15),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_324),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_326),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_14),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_5),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_328),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_321),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_329),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_319),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_332),
.A2(n_331),
.B(n_329),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_335),
.Y(n_336)
);

BUFx24_ASAP7_75t_SL g337 ( 
.A(n_336),
.Y(n_337)
);

OA21x2_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_334),
.B(n_330),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_333),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_316),
.B(n_331),
.Y(n_340)
);


endmodule