module fake_netlist_1_5059_n_44 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_44);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_44;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_25;
wire n_30;
wire n_26;
wire n_16;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
INVx1_ASAP7_75t_L g16 ( .A(n_6), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_8), .Y(n_17) );
BUFx3_ASAP7_75t_L g18 ( .A(n_14), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_3), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_4), .Y(n_20) );
AND2x4_ASAP7_75t_L g21 ( .A(n_11), .B(n_2), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_7), .Y(n_22) );
NOR2xp33_ASAP7_75t_L g23 ( .A(n_17), .B(n_0), .Y(n_23) );
BUFx3_ASAP7_75t_L g24 ( .A(n_18), .Y(n_24) );
AND3x2_ASAP7_75t_SL g25 ( .A(n_20), .B(n_0), .C(n_1), .Y(n_25) );
INVx8_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
INVx2_ASAP7_75t_L g27 ( .A(n_24), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_26), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
NAND2xp5_ASAP7_75t_L g31 ( .A(n_28), .B(n_23), .Y(n_31) );
AND2x2_ASAP7_75t_L g32 ( .A(n_30), .B(n_29), .Y(n_32) );
AOI22xp33_ASAP7_75t_L g33 ( .A1(n_30), .A2(n_21), .B1(n_19), .B2(n_22), .Y(n_33) );
INVxp33_ASAP7_75t_SL g34 ( .A(n_32), .Y(n_34) );
OAI221xp5_ASAP7_75t_SL g35 ( .A1(n_33), .A2(n_31), .B1(n_16), .B2(n_22), .C(n_25), .Y(n_35) );
AOI211xp5_ASAP7_75t_L g36 ( .A1(n_32), .A2(n_16), .B(n_21), .C(n_20), .Y(n_36) );
NOR3xp33_ASAP7_75t_L g37 ( .A(n_35), .B(n_17), .C(n_21), .Y(n_37) );
NAND2xp5_ASAP7_75t_L g38 ( .A(n_34), .B(n_1), .Y(n_38) );
INVx1_ASAP7_75t_L g39 ( .A(n_36), .Y(n_39) );
OAI22xp5_ASAP7_75t_L g40 ( .A1(n_39), .A2(n_18), .B1(n_3), .B2(n_4), .Y(n_40) );
AOI31xp33_ASAP7_75t_L g41 ( .A1(n_38), .A2(n_2), .A3(n_5), .B(n_6), .Y(n_41) );
INVx1_ASAP7_75t_L g42 ( .A(n_41), .Y(n_42) );
OAI22xp5_ASAP7_75t_L g43 ( .A1(n_40), .A2(n_37), .B1(n_7), .B2(n_5), .Y(n_43) );
AOI322xp5_ASAP7_75t_L g44 ( .A1(n_42), .A2(n_9), .A3(n_10), .B1(n_12), .B2(n_13), .C1(n_15), .C2(n_43), .Y(n_44) );
endmodule