module fake_jpeg_27016_n_138 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_138);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_138;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx4f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g30 ( 
.A(n_20),
.Y(n_30)
);

CKINVDCx6p67_ASAP7_75t_R g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_35),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_36),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_41)
);

NAND3xp33_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_10),
.C(n_9),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_38),
.B(n_39),
.Y(n_52)
);

NAND3xp33_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_10),
.C(n_8),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_32),
.A2(n_27),
.B1(n_13),
.B2(n_16),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_14),
.B1(n_16),
.B2(n_21),
.Y(n_46)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_32),
.B1(n_30),
.B2(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_14),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_35),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_13),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_61),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_47),
.Y(n_54)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_22),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_64),
.Y(n_72)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_60),
.A2(n_62),
.B1(n_45),
.B2(n_43),
.Y(n_75)
);

AO22x1_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_30),
.B1(n_32),
.B2(n_28),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g71 ( 
.A(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_66),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_22),
.Y(n_66)
);

A2O1A1O1Ixp25_ASAP7_75t_L g70 ( 
.A1(n_56),
.A2(n_45),
.B(n_30),
.C(n_31),
.D(n_14),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_70),
.A2(n_62),
.B(n_60),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_25),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_80),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_78),
.B1(n_82),
.B2(n_31),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_45),
.B1(n_28),
.B2(n_42),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_18),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_21),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_50),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_53),
.A2(n_28),
.B1(n_42),
.B2(n_29),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_77),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_88),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_52),
.B(n_50),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_84),
.A2(n_89),
.B(n_82),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_78),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_69),
.A2(n_64),
.B1(n_60),
.B2(n_59),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_90),
.B1(n_93),
.B2(n_67),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_57),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_60),
.B1(n_63),
.B2(n_55),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_95),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_75),
.A2(n_62),
.B1(n_54),
.B2(n_29),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_94),
.A2(n_79),
.B1(n_67),
.B2(n_71),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_71),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_81),
.C(n_76),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_100),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_86),
.B(n_76),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_102),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_70),
.B(n_79),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_99),
.A2(n_106),
.B(n_19),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_68),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_103),
.A2(n_91),
.B(n_19),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_105),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_18),
.B(n_25),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_107),
.Y(n_120)
);

A2O1A1O1Ixp25_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_93),
.B(n_94),
.C(n_24),
.D(n_92),
.Y(n_109)
);

OAI322xp33_ASAP7_75t_L g117 ( 
.A1(n_109),
.A2(n_114),
.A3(n_33),
.B1(n_35),
.B2(n_23),
.C1(n_104),
.C2(n_105),
.Y(n_117)
);

MAJx2_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_114),
.C(n_109),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_101),
.Y(n_112)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

A2O1A1O1Ixp25_ASAP7_75t_L g114 ( 
.A1(n_106),
.A2(n_35),
.B(n_33),
.C(n_23),
.D(n_15),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_117),
.A2(n_121),
.B(n_108),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_111),
.A2(n_96),
.B1(n_33),
.B2(n_2),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_119),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_124),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_125),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_116),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_115),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_0),
.B(n_1),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_125),
.A2(n_121),
.B1(n_115),
.B2(n_2),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_129),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_128),
.A2(n_0),
.B(n_2),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_133),
.Y(n_135)
);

OAI21x1_ASAP7_75t_L g133 ( 
.A1(n_130),
.A2(n_3),
.B(n_4),
.Y(n_133)
);

BUFx24_ASAP7_75t_SL g134 ( 
.A(n_131),
.Y(n_134)
);

MAJx2_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_127),
.C(n_4),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_5),
.B1(n_135),
.B2(n_126),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_5),
.Y(n_138)
);


endmodule