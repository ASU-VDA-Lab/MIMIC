module fake_netlist_1_5026_n_637 (n_117, n_44, n_133, n_149, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_125, n_9, n_10, n_130, n_103, n_19, n_87, n_137, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_146, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_46, n_31, n_58, n_122, n_138, n_126, n_118, n_32, n_0, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_75, n_105, n_159, n_72, n_136, n_43, n_76, n_89, n_68, n_144, n_27, n_53, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_3, n_18, n_110, n_66, n_134, n_1, n_82, n_106, n_15, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_637);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_125;
input n_9;
input n_10;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_146;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_118;
input n_32;
input n_0;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_75;
input n_105;
input n_159;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_68;
input n_144;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_82;
input n_106;
input n_15;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_637;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_612;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_202;
wire n_386;
wire n_432;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_599;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_529;
wire n_455;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_178;
wire n_616;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_438;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_524;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_187;
wire n_375;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_44), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_153), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_48), .Y(n_163) );
CKINVDCx16_ASAP7_75t_R g164 ( .A(n_130), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_95), .Y(n_165) );
BUFx2_ASAP7_75t_L g166 ( .A(n_57), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_21), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_135), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_113), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_77), .Y(n_170) );
INVx2_ASAP7_75t_SL g171 ( .A(n_53), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_119), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_157), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_107), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_37), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_123), .Y(n_176) );
BUFx2_ASAP7_75t_L g177 ( .A(n_42), .Y(n_177) );
INVxp67_ASAP7_75t_L g178 ( .A(n_1), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_116), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_150), .Y(n_180) );
BUFx5_ASAP7_75t_L g181 ( .A(n_9), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_15), .Y(n_182) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_97), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_122), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_78), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_8), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_0), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_29), .Y(n_188) );
NOR2xp67_ASAP7_75t_L g189 ( .A(n_17), .B(n_38), .Y(n_189) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_136), .Y(n_190) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_59), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_143), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g193 ( .A(n_80), .Y(n_193) );
BUFx3_ASAP7_75t_L g194 ( .A(n_34), .Y(n_194) );
OR2x2_ASAP7_75t_L g195 ( .A(n_159), .B(n_22), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_108), .Y(n_196) );
BUFx2_ASAP7_75t_L g197 ( .A(n_12), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_117), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_131), .Y(n_199) );
INVx1_ASAP7_75t_SL g200 ( .A(n_7), .Y(n_200) );
BUFx2_ASAP7_75t_SL g201 ( .A(n_127), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_109), .Y(n_202) );
INVxp67_ASAP7_75t_SL g203 ( .A(n_58), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_133), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_118), .Y(n_205) );
CKINVDCx14_ASAP7_75t_R g206 ( .A(n_132), .Y(n_206) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_124), .Y(n_207) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_46), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_102), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_79), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_129), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_146), .Y(n_212) );
INVxp67_ASAP7_75t_SL g213 ( .A(n_86), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_134), .Y(n_214) );
INVx1_ASAP7_75t_SL g215 ( .A(n_74), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_2), .Y(n_216) );
INVx1_ASAP7_75t_SL g217 ( .A(n_41), .Y(n_217) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_126), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_138), .Y(n_219) );
CKINVDCx16_ASAP7_75t_R g220 ( .A(n_18), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_114), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_111), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_151), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_147), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_28), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_112), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_1), .Y(n_227) );
INVxp67_ASAP7_75t_L g228 ( .A(n_67), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_101), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_125), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_137), .Y(n_231) );
INVx1_ASAP7_75t_SL g232 ( .A(n_87), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_39), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_92), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_96), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_62), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_121), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_89), .Y(n_238) );
CKINVDCx16_ASAP7_75t_R g239 ( .A(n_81), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_56), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_47), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_16), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_24), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_141), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_35), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_140), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_139), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_55), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_43), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_73), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_152), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_142), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_128), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_63), .Y(n_254) );
NOR2xp67_ASAP7_75t_L g255 ( .A(n_149), .B(n_20), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_13), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_110), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_19), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_75), .Y(n_259) );
NOR2xp67_ASAP7_75t_L g260 ( .A(n_144), .B(n_120), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_115), .Y(n_261) );
INVx1_ASAP7_75t_SL g262 ( .A(n_85), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_160), .Y(n_263) );
INVxp67_ASAP7_75t_L g264 ( .A(n_227), .Y(n_264) );
AND2x4_ASAP7_75t_L g265 ( .A(n_166), .B(n_0), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_177), .B(n_2), .Y(n_266) );
BUFx6f_ASAP7_75t_L g267 ( .A(n_168), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_167), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_181), .Y(n_269) );
INVx5_ASAP7_75t_L g270 ( .A(n_168), .Y(n_270) );
OA21x2_ASAP7_75t_L g271 ( .A1(n_170), .A2(n_106), .B(n_156), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_197), .B(n_3), .Y(n_272) );
BUFx12f_ASAP7_75t_L g273 ( .A(n_187), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_165), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_181), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_168), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_207), .B(n_171), .Y(n_277) );
OA21x2_ASAP7_75t_L g278 ( .A1(n_173), .A2(n_105), .B(n_155), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_181), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_178), .B(n_3), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_175), .Y(n_281) );
AND2x4_ASAP7_75t_L g282 ( .A(n_194), .B(n_4), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_164), .B(n_4), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_220), .A2(n_5), .B1(n_6), .B2(n_10), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_181), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_176), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_269), .Y(n_287) );
BUFx2_ASAP7_75t_L g288 ( .A(n_273), .Y(n_288) );
OAI22xp33_ASAP7_75t_L g289 ( .A1(n_284), .A2(n_216), .B1(n_239), .B2(n_193), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_275), .Y(n_290) );
INVx1_ASAP7_75t_SL g291 ( .A(n_283), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_279), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_277), .B(n_206), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_285), .Y(n_294) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_264), .B(n_228), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_281), .B(n_161), .Y(n_296) );
INVx3_ASAP7_75t_L g297 ( .A(n_282), .Y(n_297) );
OAI22xp5_ASAP7_75t_SL g298 ( .A1(n_274), .A2(n_174), .B1(n_186), .B2(n_213), .Y(n_298) );
INVx4_ASAP7_75t_L g299 ( .A(n_265), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_268), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_268), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_286), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_300), .B(n_283), .Y(n_303) );
OAI22xp33_ASAP7_75t_L g304 ( .A1(n_291), .A2(n_280), .B1(n_266), .B2(n_272), .Y(n_304) );
BUFx2_ASAP7_75t_L g305 ( .A(n_288), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_293), .B(n_200), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_299), .B(n_163), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_302), .B(n_169), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_301), .B(n_172), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_296), .B(n_179), .Y(n_310) );
NOR2xp67_ASAP7_75t_L g311 ( .A(n_299), .B(n_270), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_297), .B(n_180), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_297), .Y(n_313) );
AND2x2_ASAP7_75t_SL g314 ( .A(n_298), .B(n_271), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g315 ( .A1(n_290), .A2(n_201), .B1(n_188), .B2(n_196), .Y(n_315) );
NAND2xp5_ASAP7_75t_SL g316 ( .A(n_295), .B(n_183), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_304), .B(n_289), .Y(n_317) );
INVxp67_ASAP7_75t_L g318 ( .A(n_305), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_313), .Y(n_319) );
AO21x2_ASAP7_75t_L g320 ( .A1(n_303), .A2(n_198), .B(n_182), .Y(n_320) );
CKINVDCx8_ASAP7_75t_R g321 ( .A(n_306), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_303), .B(n_292), .Y(n_322) );
OR2x2_ASAP7_75t_L g323 ( .A(n_316), .B(n_287), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_309), .A2(n_294), .B(n_278), .Y(n_324) );
BUFx2_ASAP7_75t_L g325 ( .A(n_308), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_312), .B(n_215), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_314), .Y(n_327) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_310), .A2(n_278), .B(n_271), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_307), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_315), .B(n_203), .Y(n_330) );
A2O1A1Ixp33_ASAP7_75t_L g331 ( .A1(n_317), .A2(n_311), .B(n_233), .C(n_252), .Y(n_331) );
OAI21x1_ASAP7_75t_L g332 ( .A1(n_328), .A2(n_195), .B(n_199), .Y(n_332) );
OA22x2_ASAP7_75t_L g333 ( .A1(n_318), .A2(n_263), .B1(n_184), .B2(n_261), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_322), .B(n_214), .Y(n_334) );
AOI21xp5_ASAP7_75t_SL g335 ( .A1(n_320), .A2(n_222), .B(n_219), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_325), .B(n_224), .Y(n_336) );
INVxp67_ASAP7_75t_L g337 ( .A(n_320), .Y(n_337) );
OAI21x1_ASAP7_75t_L g338 ( .A1(n_324), .A2(n_238), .B(n_235), .Y(n_338) );
NOR2x1_ASAP7_75t_SL g339 ( .A(n_323), .B(n_241), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g340 ( .A1(n_327), .A2(n_246), .B1(n_244), .B2(n_247), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_330), .B(n_249), .Y(n_341) );
OAI21x1_ASAP7_75t_L g342 ( .A1(n_329), .A2(n_254), .B(n_253), .Y(n_342) );
OAI21x1_ASAP7_75t_L g343 ( .A1(n_330), .A2(n_185), .B(n_162), .Y(n_343) );
INVx6_ASAP7_75t_L g344 ( .A(n_321), .Y(n_344) );
OAI21xp5_ASAP7_75t_L g345 ( .A1(n_326), .A2(n_255), .B(n_189), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_319), .A2(n_209), .B(n_192), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_322), .B(n_190), .Y(n_347) );
OAI21x1_ASAP7_75t_L g348 ( .A1(n_328), .A2(n_229), .B(n_225), .Y(n_348) );
BUFx12f_ASAP7_75t_L g349 ( .A(n_323), .Y(n_349) );
CKINVDCx20_ASAP7_75t_R g350 ( .A(n_318), .Y(n_350) );
OAI21x1_ASAP7_75t_L g351 ( .A1(n_328), .A2(n_258), .B(n_230), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_343), .Y(n_352) );
AO21x2_ASAP7_75t_L g353 ( .A1(n_348), .A2(n_260), .B(n_181), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_332), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_342), .Y(n_355) );
AO21x2_ASAP7_75t_L g356 ( .A1(n_351), .A2(n_243), .B(n_218), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_334), .Y(n_357) );
INVx3_ASAP7_75t_L g358 ( .A(n_344), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_341), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_336), .Y(n_360) );
NOR2x1_ASAP7_75t_L g361 ( .A(n_350), .B(n_217), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_331), .B(n_191), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_344), .Y(n_363) );
OAI21x1_ASAP7_75t_L g364 ( .A1(n_338), .A2(n_243), .B(n_218), .Y(n_364) );
OAI21x1_ASAP7_75t_L g365 ( .A1(n_335), .A2(n_243), .B(n_218), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_339), .Y(n_366) );
NOR2x1_ASAP7_75t_R g367 ( .A(n_349), .B(n_202), .Y(n_367) );
OAI21x1_ASAP7_75t_L g368 ( .A1(n_346), .A2(n_11), .B(n_14), .Y(n_368) );
BUFx2_ASAP7_75t_SL g369 ( .A(n_333), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_337), .Y(n_370) );
OAI21x1_ASAP7_75t_SL g371 ( .A1(n_345), .A2(n_340), .B(n_347), .Y(n_371) );
OR2x6_ASAP7_75t_L g372 ( .A(n_344), .B(n_267), .Y(n_372) );
BUFx12f_ASAP7_75t_L g373 ( .A(n_344), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_336), .B(n_232), .Y(n_374) );
INVx1_ASAP7_75t_SL g375 ( .A(n_350), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_334), .Y(n_376) );
OR2x6_ASAP7_75t_L g377 ( .A(n_344), .B(n_267), .Y(n_377) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_334), .A2(n_262), .B1(n_204), .B2(n_237), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_343), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_334), .Y(n_380) );
INVx6_ASAP7_75t_L g381 ( .A(n_344), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_334), .Y(n_382) );
NAND2xp5_ASAP7_75t_SL g383 ( .A(n_350), .B(n_205), .Y(n_383) );
BUFx2_ASAP7_75t_L g384 ( .A(n_350), .Y(n_384) );
OAI21x1_ASAP7_75t_L g385 ( .A1(n_348), .A2(n_23), .B(n_25), .Y(n_385) );
NAND2x1p5_ASAP7_75t_L g386 ( .A(n_350), .B(n_270), .Y(n_386) );
OAI21x1_ASAP7_75t_L g387 ( .A1(n_348), .A2(n_26), .B(n_27), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_334), .Y(n_388) );
OAI21xp5_ASAP7_75t_L g389 ( .A1(n_337), .A2(n_240), .B(n_210), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_334), .A2(n_242), .B1(n_211), .B2(n_259), .Y(n_390) );
OAI21x1_ASAP7_75t_SL g391 ( .A1(n_339), .A2(n_30), .B(n_31), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_336), .B(n_208), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_374), .B(n_212), .Y(n_393) );
INVx1_ASAP7_75t_SL g394 ( .A(n_375), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_360), .B(n_221), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_370), .Y(n_396) );
BUFx2_ASAP7_75t_L g397 ( .A(n_384), .Y(n_397) );
A2O1A1Ixp33_ASAP7_75t_L g398 ( .A1(n_366), .A2(n_248), .B(n_226), .C(n_257), .Y(n_398) );
AO21x2_ASAP7_75t_L g399 ( .A1(n_371), .A2(n_276), .B(n_270), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_357), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_355), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_376), .B(n_223), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_380), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_382), .Y(n_404) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_372), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_388), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_359), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_369), .Y(n_408) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_384), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_369), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_372), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_354), .Y(n_412) );
OAI21x1_ASAP7_75t_L g413 ( .A1(n_364), .A2(n_276), .B(n_33), .Y(n_413) );
NOR3xp33_ASAP7_75t_L g414 ( .A(n_361), .B(n_256), .C(n_251), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_377), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_377), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_391), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_391), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_352), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_379), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_353), .Y(n_421) );
INVx2_ASAP7_75t_SL g422 ( .A(n_373), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_371), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_368), .Y(n_424) );
OAI21x1_ASAP7_75t_L g425 ( .A1(n_385), .A2(n_387), .B(n_365), .Y(n_425) );
OAI21x1_ASAP7_75t_L g426 ( .A1(n_356), .A2(n_32), .B(n_36), .Y(n_426) );
AO21x2_ASAP7_75t_L g427 ( .A1(n_389), .A2(n_250), .B(n_245), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_362), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_386), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_392), .Y(n_430) );
OA21x2_ASAP7_75t_L g431 ( .A1(n_378), .A2(n_236), .B(n_234), .Y(n_431) );
BUFx2_ASAP7_75t_SL g432 ( .A(n_358), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_381), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_381), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_363), .B(n_231), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_383), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_367), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_390), .B(n_40), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_360), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_384), .Y(n_440) );
BUFx2_ASAP7_75t_L g441 ( .A(n_384), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_370), .Y(n_442) );
BUFx2_ASAP7_75t_L g443 ( .A(n_384), .Y(n_443) );
OAI21xp33_ASAP7_75t_SL g444 ( .A1(n_366), .A2(n_45), .B(n_49), .Y(n_444) );
BUFx12f_ASAP7_75t_L g445 ( .A(n_363), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_370), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_370), .Y(n_447) );
INVx3_ASAP7_75t_L g448 ( .A(n_366), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_360), .B(n_158), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_374), .B(n_50), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_370), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_374), .B(n_51), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_370), .Y(n_453) );
INVx3_ASAP7_75t_L g454 ( .A(n_448), .Y(n_454) );
NOR2x1_ASAP7_75t_L g455 ( .A(n_448), .B(n_52), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_407), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_403), .B(n_154), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_400), .Y(n_458) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_396), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_439), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_396), .B(n_54), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_430), .B(n_60), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_404), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_430), .B(n_61), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_447), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_406), .B(n_64), .Y(n_466) );
AND2x2_ASAP7_75t_SL g467 ( .A(n_405), .B(n_65), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_447), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_453), .Y(n_469) );
INVx3_ASAP7_75t_L g470 ( .A(n_405), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_442), .B(n_66), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_453), .Y(n_472) );
BUFx2_ASAP7_75t_L g473 ( .A(n_405), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_446), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g475 ( .A(n_445), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_451), .Y(n_476) );
INVx3_ASAP7_75t_L g477 ( .A(n_408), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_401), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_401), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_397), .A2(n_68), .B1(n_69), .B2(n_70), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_395), .B(n_71), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_420), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_409), .B(n_72), .Y(n_483) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_433), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_440), .B(n_441), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_412), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_420), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_443), .B(n_76), .Y(n_488) );
INVxp67_ASAP7_75t_R g489 ( .A(n_437), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_419), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_410), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_428), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_428), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_423), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_421), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_429), .Y(n_496) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_429), .Y(n_497) );
INVx2_ASAP7_75t_SL g498 ( .A(n_422), .Y(n_498) );
BUFx2_ASAP7_75t_L g499 ( .A(n_411), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_417), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_394), .B(n_148), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_449), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_415), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_416), .Y(n_504) );
NAND2x1p5_ASAP7_75t_SL g505 ( .A(n_450), .B(n_452), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_436), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_434), .B(n_82), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_432), .B(n_145), .Y(n_508) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_399), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_418), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_498), .B(n_435), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_474), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_459), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_463), .B(n_393), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_465), .B(n_414), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_485), .B(n_431), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_469), .Y(n_517) );
AND2x4_ASAP7_75t_L g518 ( .A(n_496), .B(n_438), .Y(n_518) );
AND2x4_ASAP7_75t_L g519 ( .A(n_497), .B(n_427), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_460), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_456), .B(n_431), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_468), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_472), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_506), .B(n_402), .Y(n_524) );
BUFx2_ASAP7_75t_L g525 ( .A(n_477), .Y(n_525) );
OR2x6_ASAP7_75t_L g526 ( .A(n_508), .B(n_426), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_458), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_476), .B(n_424), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_478), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_492), .B(n_444), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_477), .B(n_425), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_499), .B(n_398), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_493), .B(n_413), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_504), .B(n_83), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_503), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_475), .B(n_84), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_454), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_467), .A2(n_88), .B1(n_90), .B2(n_91), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_479), .B(n_93), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_486), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_484), .B(n_94), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_454), .B(n_98), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_482), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_473), .B(n_99), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_482), .B(n_100), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_487), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_487), .Y(n_547) );
BUFx3_ASAP7_75t_L g548 ( .A(n_484), .Y(n_548) );
INVx3_ASAP7_75t_L g549 ( .A(n_470), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_484), .B(n_103), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_491), .B(n_104), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_490), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_552), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_543), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_546), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_525), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_525), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_513), .B(n_495), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_517), .B(n_495), .Y(n_559) );
NOR2xp67_ASAP7_75t_L g560 ( .A(n_538), .B(n_501), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_516), .B(n_490), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_512), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_520), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_535), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_519), .B(n_470), .Y(n_565) );
INVx3_ASAP7_75t_L g566 ( .A(n_531), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_522), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_540), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_527), .B(n_500), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_537), .B(n_510), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_523), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_529), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_547), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_518), .B(n_500), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_528), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_548), .B(n_489), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_521), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_514), .B(n_494), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_524), .B(n_505), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_563), .Y(n_580) );
NAND2x1_ASAP7_75t_SL g581 ( .A(n_560), .B(n_511), .Y(n_581) );
AND2x4_ASAP7_75t_L g582 ( .A(n_566), .B(n_531), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_574), .B(n_549), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_564), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_567), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_571), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_561), .B(n_532), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_575), .B(n_494), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_578), .B(n_530), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_558), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_579), .B(n_515), .Y(n_591) );
NOR2x1_ASAP7_75t_L g592 ( .A(n_576), .B(n_534), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_562), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_559), .Y(n_594) );
AND3x2_ASAP7_75t_L g595 ( .A(n_570), .B(n_536), .C(n_542), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_568), .Y(n_596) );
OAI32xp33_ASAP7_75t_L g597 ( .A1(n_591), .A2(n_566), .A3(n_565), .B1(n_557), .B2(n_556), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_580), .Y(n_598) );
INVxp67_ASAP7_75t_L g599 ( .A(n_592), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_584), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_590), .B(n_577), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_589), .B(n_572), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_585), .Y(n_603) );
OAI33xp33_ASAP7_75t_L g604 ( .A1(n_594), .A2(n_573), .A3(n_569), .B1(n_555), .B2(n_554), .B3(n_457), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_587), .B(n_554), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_586), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_602), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_599), .B(n_593), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_605), .B(n_596), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_601), .Y(n_610) );
INVxp33_ASAP7_75t_L g611 ( .A(n_598), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_600), .Y(n_612) );
AOI221xp5_ASAP7_75t_L g613 ( .A1(n_611), .A2(n_604), .B1(n_597), .B2(n_603), .C(n_606), .Y(n_613) );
AOI211xp5_ASAP7_75t_SL g614 ( .A1(n_608), .A2(n_595), .B(n_488), .C(n_581), .Y(n_614) );
NOR2xp33_ASAP7_75t_SL g615 ( .A(n_607), .B(n_583), .Y(n_615) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_610), .A2(n_612), .B1(n_609), .B2(n_582), .C(n_555), .Y(n_616) );
NOR4xp25_ASAP7_75t_L g617 ( .A(n_613), .B(n_616), .C(n_483), .D(n_464), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_614), .B(n_588), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_615), .A2(n_582), .B1(n_542), .B2(n_526), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_618), .Y(n_620) );
NOR2x1_ASAP7_75t_SL g621 ( .A(n_617), .B(n_526), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_620), .B(n_621), .Y(n_622) );
XNOR2xp5_ASAP7_75t_L g623 ( .A(n_620), .B(n_619), .Y(n_623) );
XNOR2x1_ASAP7_75t_L g624 ( .A(n_623), .B(n_481), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g625 ( .A(n_622), .B(n_455), .Y(n_625) );
BUFx10_ASAP7_75t_L g626 ( .A(n_624), .Y(n_626) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_625), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_627), .B(n_462), .Y(n_628) );
NOR2xp33_ASAP7_75t_SL g629 ( .A(n_626), .B(n_544), .Y(n_629) );
NAND2xp67_ASAP7_75t_L g630 ( .A(n_628), .B(n_507), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_629), .A2(n_502), .B1(n_480), .B2(n_461), .Y(n_631) );
OAI21xp5_ASAP7_75t_L g632 ( .A1(n_631), .A2(n_541), .B(n_466), .Y(n_632) );
OAI21xp5_ASAP7_75t_L g633 ( .A1(n_630), .A2(n_551), .B(n_545), .Y(n_633) );
OAI21x1_ASAP7_75t_SL g634 ( .A1(n_633), .A2(n_539), .B(n_533), .Y(n_634) );
OR2x6_ASAP7_75t_L g635 ( .A(n_634), .B(n_632), .Y(n_635) );
OR2x6_ASAP7_75t_L g636 ( .A(n_635), .B(n_550), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_636), .A2(n_553), .B1(n_509), .B2(n_471), .Y(n_637) );
endmodule