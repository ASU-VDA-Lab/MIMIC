module real_aes_17761_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1095;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1301;
wire n_728;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1648;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_733;
wire n_402;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1620;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_1524;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1605;
wire n_1056;
wire n_1592;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1619;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1617;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1584;
wire n_1277;
wire n_1049;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_1280;
wire n_394;
wire n_729;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_0), .A2(n_53), .B1(n_459), .B2(n_788), .Y(n_787) );
INVxp67_ASAP7_75t_SL g816 ( .A(n_0), .Y(n_816) );
INVx1_ASAP7_75t_L g947 ( .A(n_1), .Y(n_947) );
INVx1_ASAP7_75t_L g327 ( .A(n_2), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_2), .B(n_337), .Y(n_352) );
AND2x2_ASAP7_75t_L g1564 ( .A(n_2), .B(n_444), .Y(n_1564) );
AND2x2_ASAP7_75t_L g1572 ( .A(n_2), .B(n_226), .Y(n_1572) );
INVx1_ASAP7_75t_L g617 ( .A(n_3), .Y(n_617) );
INVx1_ASAP7_75t_L g855 ( .A(n_4), .Y(n_855) );
OAI22xp5_ASAP7_75t_SL g870 ( .A1(n_5), .A2(n_202), .B1(n_472), .B2(n_539), .Y(n_870) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_5), .A2(n_202), .B1(n_874), .B2(n_875), .Y(n_873) );
INVx1_ASAP7_75t_L g1127 ( .A(n_6), .Y(n_1127) );
INVx1_ASAP7_75t_L g842 ( .A(n_7), .Y(n_842) );
CKINVDCx5p33_ASAP7_75t_R g686 ( .A(n_8), .Y(n_686) );
INVx1_ASAP7_75t_L g763 ( .A(n_9), .Y(n_763) );
OAI22xp33_ASAP7_75t_L g871 ( .A1(n_10), .A2(n_139), .B1(n_329), .B2(n_544), .Y(n_871) );
OAI22xp33_ASAP7_75t_L g881 ( .A1(n_10), .A2(n_139), .B1(n_523), .B2(n_608), .Y(n_881) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_11), .A2(n_41), .B1(n_481), .B2(n_523), .Y(n_522) );
OAI22xp33_ASAP7_75t_L g543 ( .A1(n_11), .A2(n_41), .B1(n_329), .B2(n_544), .Y(n_543) );
CKINVDCx5p33_ASAP7_75t_R g1005 ( .A(n_12), .Y(n_1005) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_13), .A2(n_281), .B1(n_539), .B2(n_594), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_13), .A2(n_281), .B1(n_507), .B2(n_509), .Y(n_661) );
INVx2_ASAP7_75t_L g398 ( .A(n_14), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g1325 ( .A1(n_15), .A2(n_19), .B1(n_1309), .B2(n_1316), .Y(n_1325) );
INVx1_ASAP7_75t_L g1173 ( .A(n_16), .Y(n_1173) );
CKINVDCx5p33_ASAP7_75t_R g1550 ( .A(n_17), .Y(n_1550) );
INVx1_ASAP7_75t_L g1169 ( .A(n_18), .Y(n_1169) );
XNOR2xp5_ASAP7_75t_L g751 ( .A(n_19), .B(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g370 ( .A(n_20), .Y(n_370) );
INVx1_ASAP7_75t_L g1236 ( .A(n_21), .Y(n_1236) );
INVx1_ASAP7_75t_L g915 ( .A(n_22), .Y(n_915) );
INVx1_ASAP7_75t_L g1122 ( .A(n_23), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g1269 ( .A1(n_24), .A2(n_166), .B1(n_1270), .B2(n_1272), .Y(n_1269) );
AOI22xp33_ASAP7_75t_SL g1292 ( .A1(n_24), .A2(n_124), .B1(n_1208), .B2(n_1293), .Y(n_1292) );
AOI221xp5_ASAP7_75t_L g1150 ( .A1(n_25), .A2(n_80), .B1(n_695), .B2(n_1151), .C(n_1154), .Y(n_1150) );
AOI22xp33_ASAP7_75t_L g1205 ( .A1(n_25), .A2(n_39), .B1(n_1206), .B2(n_1208), .Y(n_1205) );
INVx1_ASAP7_75t_L g354 ( .A(n_26), .Y(n_354) );
OAI211xp5_ASAP7_75t_L g447 ( .A1(n_27), .A2(n_448), .B(n_452), .C(n_464), .Y(n_447) );
INVx1_ASAP7_75t_L g505 ( .A(n_27), .Y(n_505) );
INVx1_ASAP7_75t_L g1050 ( .A(n_28), .Y(n_1050) );
OAI221xp5_ASAP7_75t_L g968 ( .A1(n_29), .A2(n_79), .B1(n_508), .B2(n_969), .C(n_971), .Y(n_968) );
INVx1_ASAP7_75t_L g992 ( .A(n_29), .Y(n_992) );
OAI22xp5_ASAP7_75t_L g1105 ( .A1(n_30), .A2(n_284), .B1(n_994), .B2(n_1034), .Y(n_1105) );
OAI22xp33_ASAP7_75t_L g1115 ( .A1(n_30), .A2(n_284), .B1(n_508), .B2(n_511), .Y(n_1115) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_31), .Y(n_322) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_31), .B(n_320), .Y(n_1310) );
AOI22xp33_ASAP7_75t_L g1378 ( .A1(n_32), .A2(n_177), .B1(n_1309), .B2(n_1365), .Y(n_1378) );
OAI22xp33_ASAP7_75t_SL g593 ( .A1(n_33), .A2(n_156), .B1(n_539), .B2(n_594), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_33), .A2(n_156), .B1(n_507), .B2(n_598), .Y(n_597) );
OAI222xp33_ASAP7_75t_L g1262 ( .A1(n_34), .A2(n_186), .B1(n_303), .B2(n_819), .C1(n_820), .C2(n_1263), .Y(n_1262) );
OAI222xp33_ASAP7_75t_L g1298 ( .A1(n_34), .A2(n_186), .B1(n_303), .B2(n_459), .C1(n_625), .C2(n_788), .Y(n_1298) );
CKINVDCx5p33_ASAP7_75t_R g1622 ( .A(n_35), .Y(n_1622) );
INVx1_ASAP7_75t_L g867 ( .A(n_36), .Y(n_867) );
INVx1_ASAP7_75t_L g722 ( .A(n_37), .Y(n_722) );
INVxp67_ASAP7_75t_SL g786 ( .A(n_38), .Y(n_786) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_38), .A2(n_53), .B1(n_819), .B2(n_820), .Y(n_818) );
AOI221xp5_ASAP7_75t_L g1157 ( .A1(n_39), .A2(n_67), .B1(n_695), .B2(n_1151), .C(n_1158), .Y(n_1157) );
INVx1_ASAP7_75t_L g904 ( .A(n_40), .Y(n_904) );
OAI22xp33_ASAP7_75t_L g1106 ( .A1(n_42), .A2(n_240), .B1(n_441), .B2(n_899), .Y(n_1106) );
OAI22xp33_ASAP7_75t_SL g1108 ( .A1(n_42), .A2(n_240), .B1(n_483), .B2(n_1109), .Y(n_1108) );
OAI22xp5_ASAP7_75t_L g1532 ( .A1(n_43), .A2(n_1533), .B1(n_1537), .B2(n_1540), .Y(n_1532) );
INVx1_ASAP7_75t_L g1575 ( .A(n_43), .Y(n_1575) );
INVx1_ASAP7_75t_L g549 ( .A(n_44), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g1363 ( .A1(n_45), .A2(n_193), .B1(n_1316), .B2(n_1319), .Y(n_1363) );
AOI22xp5_ASAP7_75t_L g1334 ( .A1(n_46), .A2(n_298), .B1(n_1309), .B2(n_1313), .Y(n_1334) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_47), .Y(n_334) );
INVx1_ASAP7_75t_L g1163 ( .A(n_48), .Y(n_1163) );
AOI22xp33_ASAP7_75t_SL g1197 ( .A1(n_48), .A2(n_232), .B1(n_1198), .B2(n_1199), .Y(n_1197) );
INVx1_ASAP7_75t_L g950 ( .A(n_49), .Y(n_950) );
AOI22xp5_ASAP7_75t_L g1364 ( .A1(n_50), .A2(n_276), .B1(n_1309), .B2(n_1365), .Y(n_1364) );
INVx1_ASAP7_75t_L g1539 ( .A(n_51), .Y(n_1539) );
AOI22xp33_ASAP7_75t_L g1588 ( .A1(n_51), .A2(n_59), .B1(n_792), .B2(n_807), .Y(n_1588) );
AOI22xp5_ASAP7_75t_L g1315 ( .A1(n_52), .A2(n_111), .B1(n_1316), .B2(n_1319), .Y(n_1315) );
INVx1_ASAP7_75t_L g852 ( .A(n_54), .Y(n_852) );
INVx1_ASAP7_75t_L g1244 ( .A(n_55), .Y(n_1244) );
NAND2xp5_ASAP7_75t_L g973 ( .A(n_56), .B(n_500), .Y(n_973) );
INVxp67_ASAP7_75t_SL g989 ( .A(n_56), .Y(n_989) );
OAI211xp5_ASAP7_75t_SL g524 ( .A1(n_57), .A2(n_489), .B(n_492), .C(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g537 ( .A(n_57), .Y(n_537) );
OAI211xp5_ASAP7_75t_L g887 ( .A1(n_58), .A2(n_603), .B(n_663), .C(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g896 ( .A(n_58), .Y(n_896) );
AOI221xp5_ASAP7_75t_L g1525 ( .A1(n_59), .A2(n_300), .B1(n_1526), .B2(n_1527), .C(n_1528), .Y(n_1525) );
OAI22xp33_ASAP7_75t_L g528 ( .A1(n_60), .A2(n_162), .B1(n_507), .B2(n_509), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_60), .A2(n_162), .B1(n_539), .B2(n_540), .Y(n_538) );
INVx1_ASAP7_75t_L g850 ( .A(n_61), .Y(n_850) );
INVx1_ASAP7_75t_L g790 ( .A(n_62), .Y(n_790) );
INVx1_ASAP7_75t_L g1126 ( .A(n_63), .Y(n_1126) );
OAI22xp33_ASAP7_75t_L g742 ( .A1(n_64), .A2(n_267), .B1(n_329), .B2(n_544), .Y(n_742) );
OAI22xp33_ASAP7_75t_L g744 ( .A1(n_64), .A2(n_267), .B1(n_523), .B2(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g463 ( .A(n_65), .Y(n_463) );
OAI211xp5_ASAP7_75t_L g488 ( .A1(n_65), .A2(n_489), .B(n_492), .C(n_496), .Y(n_488) );
OAI22xp33_ASAP7_75t_L g978 ( .A1(n_66), .A2(n_171), .B1(n_483), .B2(n_979), .Y(n_978) );
INVxp67_ASAP7_75t_SL g991 ( .A(n_66), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g1200 ( .A1(n_67), .A2(n_80), .B1(n_1201), .B2(n_1203), .Y(n_1200) );
INVx1_ASAP7_75t_L g914 ( .A(n_68), .Y(n_914) );
CKINVDCx5p33_ASAP7_75t_R g1017 ( .A(n_69), .Y(n_1017) );
INVx1_ASAP7_75t_L g795 ( .A(n_70), .Y(n_795) );
INVx1_ASAP7_75t_L g910 ( .A(n_71), .Y(n_910) );
INVx1_ASAP7_75t_L g563 ( .A(n_72), .Y(n_563) );
CKINVDCx5p33_ASAP7_75t_R g1063 ( .A(n_73), .Y(n_1063) );
OAI211xp5_ASAP7_75t_L g1100 ( .A1(n_74), .A2(n_983), .B(n_1101), .C(n_1102), .Y(n_1100) );
INVx1_ASAP7_75t_L g1112 ( .A(n_74), .Y(n_1112) );
INVx1_ASAP7_75t_L g781 ( .A(n_75), .Y(n_781) );
INVx1_ASAP7_75t_L g949 ( .A(n_76), .Y(n_949) );
INVx1_ASAP7_75t_L g637 ( .A(n_77), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g1341 ( .A1(n_78), .A2(n_306), .B1(n_1316), .B2(n_1319), .Y(n_1341) );
OAI22xp33_ASAP7_75t_L g995 ( .A1(n_79), .A2(n_171), .B1(n_441), .B2(n_899), .Y(n_995) );
OAI22xp5_ASAP7_75t_L g1166 ( .A1(n_81), .A2(n_179), .B1(n_483), .B2(n_508), .Y(n_1166) );
INVx1_ASAP7_75t_L g1179 ( .A(n_81), .Y(n_1179) );
INVx1_ASAP7_75t_L g377 ( .A(n_82), .Y(n_377) );
INVx1_ASAP7_75t_L g1083 ( .A(n_83), .Y(n_1083) );
OAI211xp5_ASAP7_75t_L g1089 ( .A1(n_83), .A2(n_436), .B(n_603), .C(n_1090), .Y(n_1089) );
OAI22xp5_ASAP7_75t_L g1028 ( .A1(n_84), .A2(n_239), .B1(n_899), .B2(n_994), .Y(n_1028) );
OAI22xp5_ASAP7_75t_SL g1037 ( .A1(n_84), .A2(n_119), .B1(n_483), .B2(n_511), .Y(n_1037) );
INVx1_ASAP7_75t_L g562 ( .A(n_85), .Y(n_562) );
INVx1_ASAP7_75t_L g977 ( .A(n_86), .Y(n_977) );
INVx1_ASAP7_75t_L g890 ( .A(n_87), .Y(n_890) );
OAI211xp5_ASAP7_75t_L g893 ( .A1(n_87), .A2(n_653), .B(n_894), .C(n_895), .Y(n_893) );
CKINVDCx5p33_ASAP7_75t_R g1031 ( .A(n_88), .Y(n_1031) );
INVx1_ASAP7_75t_L g1130 ( .A(n_89), .Y(n_1130) );
CKINVDCx5p33_ASAP7_75t_R g1003 ( .A(n_90), .Y(n_1003) );
OAI22xp33_ASAP7_75t_L g440 ( .A1(n_91), .A2(n_149), .B1(n_329), .B2(n_441), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_91), .A2(n_149), .B1(n_481), .B2(n_484), .Y(n_480) );
INVx1_ASAP7_75t_L g1174 ( .A(n_92), .Y(n_1174) );
XNOR2xp5_ASAP7_75t_L g1610 ( .A(n_93), .B(n_1611), .Y(n_1610) );
AOI22xp5_ASAP7_75t_SL g1342 ( .A1(n_94), .A2(n_200), .B1(n_1309), .B2(n_1313), .Y(n_1342) );
INVx1_ASAP7_75t_L g765 ( .A(n_95), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_95), .A2(n_259), .B1(n_806), .B2(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g909 ( .A(n_96), .Y(n_909) );
CKINVDCx5p33_ASAP7_75t_R g1625 ( .A(n_97), .Y(n_1625) );
CKINVDCx5p33_ASAP7_75t_R g1013 ( .A(n_98), .Y(n_1013) );
OAI22xp33_ASAP7_75t_L g1553 ( .A1(n_99), .A2(n_133), .B1(n_1554), .B2(n_1556), .Y(n_1553) );
OAI22xp5_ASAP7_75t_L g1589 ( .A1(n_99), .A2(n_258), .B1(n_1590), .B2(n_1597), .Y(n_1589) );
INVx1_ASAP7_75t_L g1104 ( .A(n_100), .Y(n_1104) );
INVx1_ASAP7_75t_L g728 ( .A(n_101), .Y(n_728) );
OAI211xp5_ASAP7_75t_L g1079 ( .A1(n_102), .A2(n_578), .B(n_983), .C(n_1080), .Y(n_1079) );
INVx1_ASAP7_75t_L g1091 ( .A(n_102), .Y(n_1091) );
INVx1_ASAP7_75t_L g320 ( .A(n_103), .Y(n_320) );
INVx1_ASAP7_75t_L g845 ( .A(n_104), .Y(n_845) );
INVx1_ASAP7_75t_L g777 ( .A(n_105), .Y(n_777) );
INVx1_ASAP7_75t_L g1535 ( .A(n_106), .Y(n_1535) );
AOI22xp33_ASAP7_75t_L g1585 ( .A1(n_106), .A2(n_300), .B1(n_792), .B2(n_1576), .Y(n_1585) );
OAI22xp33_ASAP7_75t_L g1085 ( .A1(n_107), .A2(n_263), .B1(n_471), .B2(n_544), .Y(n_1085) );
OAI22xp33_ASAP7_75t_L g1092 ( .A1(n_107), .A2(n_145), .B1(n_508), .B2(n_511), .Y(n_1092) );
AOI22xp5_ASAP7_75t_L g1338 ( .A1(n_108), .A2(n_289), .B1(n_1313), .B2(n_1319), .Y(n_1338) );
INVx1_ASAP7_75t_L g591 ( .A(n_109), .Y(n_591) );
INVx1_ASAP7_75t_L g716 ( .A(n_110), .Y(n_716) );
INVx1_ASAP7_75t_L g761 ( .A(n_112), .Y(n_761) );
INVx1_ASAP7_75t_L g622 ( .A(n_113), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g1260 ( .A1(n_114), .A2(n_228), .B1(n_979), .B2(n_1261), .Y(n_1260) );
OAI22xp5_ASAP7_75t_L g1297 ( .A1(n_114), .A2(n_228), .B1(n_470), .B2(n_797), .Y(n_1297) );
CKINVDCx5p33_ASAP7_75t_R g1530 ( .A(n_115), .Y(n_1530) );
INVx1_ASAP7_75t_L g889 ( .A(n_116), .Y(n_889) );
INVx1_ASAP7_75t_L g1239 ( .A(n_117), .Y(n_1239) );
OAI22xp33_ASAP7_75t_SL g1033 ( .A1(n_118), .A2(n_119), .B1(n_441), .B2(n_1034), .Y(n_1033) );
OAI22xp5_ASAP7_75t_L g1041 ( .A1(n_118), .A2(n_123), .B1(n_1042), .B2(n_1043), .Y(n_1041) );
INVx1_ASAP7_75t_L g567 ( .A(n_120), .Y(n_567) );
INVx1_ASAP7_75t_L g1242 ( .A(n_121), .Y(n_1242) );
CKINVDCx5p33_ASAP7_75t_R g682 ( .A(n_122), .Y(n_682) );
INVx1_ASAP7_75t_L g1032 ( .A(n_123), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g1276 ( .A1(n_124), .A2(n_256), .B1(n_1151), .B2(n_1277), .Y(n_1276) );
INVx1_ASAP7_75t_L g907 ( .A(n_125), .Y(n_907) );
INVx1_ASAP7_75t_L g1240 ( .A(n_126), .Y(n_1240) );
AOI31xp33_ASAP7_75t_L g1142 ( .A1(n_127), .A2(n_1143), .A3(n_1165), .B(n_1177), .Y(n_1142) );
NAND2xp33_ASAP7_75t_SL g1193 ( .A(n_127), .B(n_1194), .Y(n_1193) );
INVxp67_ASAP7_75t_SL g1211 ( .A(n_127), .Y(n_1211) );
INVx1_ASAP7_75t_L g357 ( .A(n_128), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g685 ( .A(n_129), .Y(n_685) );
CKINVDCx5p33_ASAP7_75t_R g1623 ( .A(n_130), .Y(n_1623) );
OAI22xp33_ASAP7_75t_L g1638 ( .A1(n_131), .A2(n_173), .B1(n_544), .B2(n_1034), .Y(n_1638) );
OAI22xp33_ASAP7_75t_L g1644 ( .A1(n_131), .A2(n_165), .B1(n_508), .B2(n_511), .Y(n_1644) );
CKINVDCx5p33_ASAP7_75t_R g1616 ( .A(n_132), .Y(n_1616) );
INVx1_ASAP7_75t_L g1581 ( .A(n_133), .Y(n_1581) );
OAI22xp33_ASAP7_75t_L g891 ( .A1(n_134), .A2(n_148), .B1(n_608), .B2(n_610), .Y(n_891) );
OAI22xp33_ASAP7_75t_L g898 ( .A1(n_134), .A2(n_148), .B1(n_544), .B2(n_899), .Y(n_898) );
OAI211xp5_ASAP7_75t_L g589 ( .A1(n_135), .A2(n_531), .B(n_534), .C(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g606 ( .A(n_135), .Y(n_606) );
CKINVDCx5p33_ASAP7_75t_R g1009 ( .A(n_136), .Y(n_1009) );
INVx1_ASAP7_75t_L g592 ( .A(n_137), .Y(n_592) );
OAI211xp5_ASAP7_75t_L g600 ( .A1(n_137), .A2(n_601), .B(n_603), .C(n_604), .Y(n_600) );
INVx1_ASAP7_75t_L g555 ( .A(n_138), .Y(n_555) );
INVx1_ASAP7_75t_L g526 ( .A(n_140), .Y(n_526) );
INVx1_ASAP7_75t_L g379 ( .A(n_141), .Y(n_379) );
INVx1_ASAP7_75t_L g619 ( .A(n_142), .Y(n_619) );
OAI211xp5_ASAP7_75t_L g735 ( .A1(n_143), .A2(n_533), .B(n_534), .C(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g749 ( .A(n_143), .Y(n_749) );
INVx1_ASAP7_75t_L g737 ( .A(n_144), .Y(n_737) );
OAI22xp33_ASAP7_75t_L g1084 ( .A1(n_145), .A2(n_242), .B1(n_542), .B2(n_899), .Y(n_1084) );
INVx1_ASAP7_75t_L g1636 ( .A(n_146), .Y(n_1636) );
OAI211xp5_ASAP7_75t_L g1641 ( .A1(n_146), .A2(n_436), .B(n_603), .C(n_1642), .Y(n_1641) );
CKINVDCx5p33_ASAP7_75t_R g1055 ( .A(n_147), .Y(n_1055) );
INVx1_ASAP7_75t_L g946 ( .A(n_150), .Y(n_946) );
OAI211xp5_ASAP7_75t_SL g865 ( .A1(n_151), .A2(n_448), .B(n_534), .C(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g880 ( .A(n_151), .Y(n_880) );
INVx1_ASAP7_75t_L g1237 ( .A(n_152), .Y(n_1237) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_153), .A2(n_255), .B1(n_539), .B2(n_594), .Y(n_741) );
OAI22xp33_ASAP7_75t_L g750 ( .A1(n_153), .A2(n_255), .B1(n_507), .B2(n_598), .Y(n_750) );
INVx1_ASAP7_75t_L g906 ( .A(n_154), .Y(n_906) );
OAI211xp5_ASAP7_75t_L g1633 ( .A1(n_155), .A2(n_578), .B(n_983), .C(n_1634), .Y(n_1633) );
INVx1_ASAP7_75t_L g1643 ( .A(n_155), .Y(n_1643) );
INVx1_ASAP7_75t_L g1547 ( .A(n_157), .Y(n_1547) );
INVx1_ASAP7_75t_L g1375 ( .A(n_158), .Y(n_1375) );
AOI22xp5_ASAP7_75t_SL g1308 ( .A1(n_159), .A2(n_167), .B1(n_1309), .B2(n_1313), .Y(n_1308) );
INVx1_ASAP7_75t_L g636 ( .A(n_160), .Y(n_636) );
INVx1_ASAP7_75t_L g727 ( .A(n_161), .Y(n_727) );
OAI22xp33_ASAP7_75t_L g1637 ( .A1(n_163), .A2(n_165), .B1(n_542), .B2(n_899), .Y(n_1637) );
OAI22xp33_ASAP7_75t_L g1640 ( .A1(n_163), .A2(n_173), .B1(n_483), .B2(n_969), .Y(n_1640) );
INVx1_ASAP7_75t_L g527 ( .A(n_164), .Y(n_527) );
OAI211xp5_ASAP7_75t_L g530 ( .A1(n_164), .A2(n_531), .B(n_534), .C(n_535), .Y(n_530) );
AOI22xp33_ASAP7_75t_SL g1284 ( .A1(n_166), .A2(n_256), .B1(n_1285), .B2(n_1289), .Y(n_1284) );
INVx1_ASAP7_75t_L g711 ( .A(n_168), .Y(n_711) );
INVx1_ASAP7_75t_L g1233 ( .A(n_169), .Y(n_1233) );
INVx2_ASAP7_75t_L g1312 ( .A(n_170), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_170), .B(n_265), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_170), .B(n_1318), .Y(n_1320) );
AOI22xp5_ASAP7_75t_SL g1323 ( .A1(n_172), .A2(n_233), .B1(n_1319), .B2(n_1324), .Y(n_1323) );
CKINVDCx5p33_ASAP7_75t_R g1620 ( .A(n_174), .Y(n_1620) );
CKINVDCx5p33_ASAP7_75t_R g1012 ( .A(n_175), .Y(n_1012) );
INVx1_ASAP7_75t_L g551 ( .A(n_176), .Y(n_551) );
XNOR2xp5_ASAP7_75t_L g836 ( .A(n_178), .B(n_837), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g1183 ( .A1(n_179), .A2(n_247), .B1(n_994), .B2(n_1034), .Y(n_1183) );
AOI22xp5_ASAP7_75t_L g1330 ( .A1(n_180), .A2(n_285), .B1(n_1309), .B2(n_1324), .Y(n_1330) );
XOR2xp5_ASAP7_75t_L g931 ( .A(n_181), .B(n_932), .Y(n_931) );
AOI22xp5_ASAP7_75t_L g1333 ( .A1(n_181), .A2(n_235), .B1(n_1316), .B2(n_1319), .Y(n_1333) );
AOI22xp33_ASAP7_75t_L g1273 ( .A1(n_182), .A2(n_293), .B1(n_1267), .B2(n_1274), .Y(n_1273) );
AOI22xp33_ASAP7_75t_L g1291 ( .A1(n_182), .A2(n_222), .B1(n_1285), .B2(n_1289), .Y(n_1291) );
XNOR2x2_ASAP7_75t_L g344 ( .A(n_183), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g939 ( .A(n_184), .Y(n_939) );
INVx1_ASAP7_75t_L g1220 ( .A(n_185), .Y(n_1220) );
CKINVDCx5p33_ASAP7_75t_R g1061 ( .A(n_187), .Y(n_1061) );
INVx1_ASAP7_75t_L g1103 ( .A(n_188), .Y(n_1103) );
XOR2x2_ASAP7_75t_L g1097 ( .A(n_189), .B(n_1098), .Y(n_1097) );
AOI22xp5_ASAP7_75t_L g1339 ( .A1(n_189), .A2(n_248), .B1(n_1309), .B2(n_1316), .Y(n_1339) );
INVx1_ASAP7_75t_L g849 ( .A(n_190), .Y(n_849) );
CKINVDCx5p33_ASAP7_75t_R g655 ( .A(n_191), .Y(n_655) );
INVx1_ASAP7_75t_L g717 ( .A(n_192), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g886 ( .A1(n_194), .A2(n_211), .B1(n_507), .B2(n_875), .Y(n_886) );
OAI22xp5_ASAP7_75t_L g897 ( .A1(n_194), .A2(n_211), .B1(n_470), .B2(n_472), .Y(n_897) );
INVx1_ASAP7_75t_L g943 ( .A(n_195), .Y(n_943) );
OAI22xp33_ASAP7_75t_L g588 ( .A1(n_196), .A2(n_257), .B1(n_329), .B2(n_544), .Y(n_588) );
OAI22xp33_ASAP7_75t_L g607 ( .A1(n_196), .A2(n_257), .B1(n_608), .B2(n_610), .Y(n_607) );
INVx2_ASAP7_75t_L g397 ( .A(n_197), .Y(n_397) );
INVx1_ASAP7_75t_L g434 ( .A(n_197), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g1543 ( .A(n_197), .B(n_398), .Y(n_1543) );
CKINVDCx5p33_ASAP7_75t_R g1056 ( .A(n_198), .Y(n_1056) );
OAI22xp33_ASAP7_75t_L g1216 ( .A1(n_199), .A2(n_245), .B1(n_994), .B2(n_1034), .Y(n_1216) );
OAI22xp5_ASAP7_75t_SL g1223 ( .A1(n_199), .A2(n_220), .B1(n_483), .B2(n_508), .Y(n_1223) );
XOR2xp5_ASAP7_75t_L g1253 ( .A(n_201), .B(n_1254), .Y(n_1253) );
BUFx3_ASAP7_75t_L g404 ( .A(n_203), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g1066 ( .A(n_204), .Y(n_1066) );
CKINVDCx5p33_ASAP7_75t_R g683 ( .A(n_205), .Y(n_683) );
CKINVDCx5p33_ASAP7_75t_R g1626 ( .A(n_206), .Y(n_1626) );
XOR2xp5_ASAP7_75t_L g706 ( .A(n_207), .B(n_707), .Y(n_706) );
OAI221xp5_ASAP7_75t_L g1548 ( .A1(n_208), .A2(n_258), .B1(n_692), .B2(n_923), .C(n_1549), .Y(n_1548) );
OAI211xp5_ASAP7_75t_L g1565 ( .A1(n_208), .A2(n_1566), .B(n_1569), .C(n_1582), .Y(n_1565) );
AOI22xp33_ASAP7_75t_L g1266 ( .A1(n_209), .A2(n_222), .B1(n_1170), .B2(n_1267), .Y(n_1266) );
AOI22xp33_ASAP7_75t_L g1281 ( .A1(n_209), .A2(n_293), .B1(n_1282), .B2(n_1283), .Y(n_1281) );
CKINVDCx5p33_ASAP7_75t_R g1529 ( .A(n_210), .Y(n_1529) );
OA22x2_ASAP7_75t_L g883 ( .A1(n_212), .A2(n_884), .B1(n_927), .B2(n_928), .Y(n_883) );
INVxp67_ASAP7_75t_L g928 ( .A(n_212), .Y(n_928) );
AOI22xp5_ASAP7_75t_L g1329 ( .A1(n_212), .A2(n_243), .B1(n_1316), .B2(n_1319), .Y(n_1329) );
INVx1_ASAP7_75t_L g770 ( .A(n_213), .Y(n_770) );
INVx1_ASAP7_75t_L g657 ( .A(n_214), .Y(n_657) );
OAI211xp5_ASAP7_75t_L g662 ( .A1(n_214), .A2(n_603), .B(n_663), .C(n_666), .Y(n_662) );
INVx1_ASAP7_75t_L g712 ( .A(n_215), .Y(n_712) );
CKINVDCx5p33_ASAP7_75t_R g1619 ( .A(n_216), .Y(n_1619) );
CKINVDCx5p33_ASAP7_75t_R g1058 ( .A(n_217), .Y(n_1058) );
INVx1_ASAP7_75t_L g624 ( .A(n_218), .Y(n_624) );
INVx1_ASAP7_75t_L g1219 ( .A(n_219), .Y(n_1219) );
OAI22xp33_ASAP7_75t_L g1221 ( .A1(n_220), .A2(n_250), .B1(n_441), .B2(n_899), .Y(n_1221) );
CKINVDCx5p33_ASAP7_75t_R g680 ( .A(n_221), .Y(n_680) );
INVx1_ASAP7_75t_L g775 ( .A(n_223), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_223), .A2(n_266), .B1(n_804), .B2(n_806), .Y(n_803) );
XOR2xp5_ASAP7_75t_L g998 ( .A(n_224), .B(n_999), .Y(n_998) );
INVx1_ASAP7_75t_L g1123 ( .A(n_225), .Y(n_1123) );
BUFx3_ASAP7_75t_L g337 ( .A(n_226), .Y(n_337) );
INVx1_ASAP7_75t_L g444 ( .A(n_226), .Y(n_444) );
INVx1_ASAP7_75t_L g457 ( .A(n_227), .Y(n_457) );
XOR2x2_ASAP7_75t_L g519 ( .A(n_229), .B(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g937 ( .A(n_230), .Y(n_937) );
INVx1_ASAP7_75t_L g1119 ( .A(n_231), .Y(n_1119) );
AOI22xp5_ASAP7_75t_L g1144 ( .A1(n_232), .A2(n_253), .B1(n_1145), .B2(n_1146), .Y(n_1144) );
INVx1_ASAP7_75t_L g392 ( .A(n_234), .Y(n_392) );
INVx1_ASAP7_75t_L g1258 ( .A(n_236), .Y(n_1258) );
CKINVDCx5p33_ASAP7_75t_R g1538 ( .A(n_237), .Y(n_1538) );
OAI211xp5_ASAP7_75t_L g1217 ( .A1(n_238), .A2(n_625), .B(n_983), .C(n_1218), .Y(n_1217) );
INVx1_ASAP7_75t_L g1228 ( .A(n_238), .Y(n_1228) );
NOR2xp33_ASAP7_75t_L g1036 ( .A(n_239), .B(n_508), .Y(n_1036) );
CKINVDCx5p33_ASAP7_75t_R g1016 ( .A(n_241), .Y(n_1016) );
OAI22xp33_ASAP7_75t_L g1088 ( .A1(n_242), .A2(n_263), .B1(n_483), .B2(n_969), .Y(n_1088) );
XOR2x2_ASAP7_75t_L g585 ( .A(n_244), .B(n_586), .Y(n_585) );
OAI22xp33_ASAP7_75t_L g1229 ( .A1(n_245), .A2(n_250), .B1(n_511), .B2(n_969), .Y(n_1229) );
CKINVDCx5p33_ASAP7_75t_R g1617 ( .A(n_246), .Y(n_1617) );
OAI22xp5_ASAP7_75t_L g1175 ( .A1(n_247), .A2(n_286), .B1(n_511), .B2(n_969), .Y(n_1175) );
INVx1_ASAP7_75t_L g406 ( .A(n_249), .Y(n_406) );
INVx1_ASAP7_75t_L g412 ( .A(n_249), .Y(n_412) );
INVx1_ASAP7_75t_L g391 ( .A(n_251), .Y(n_391) );
INVx1_ASAP7_75t_L g365 ( .A(n_252), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g1204 ( .A1(n_253), .A2(n_288), .B1(n_1201), .B2(n_1203), .Y(n_1204) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_254), .A2(n_301), .B1(n_470), .B2(n_472), .Y(n_469) );
OAI22xp33_ASAP7_75t_L g506 ( .A1(n_254), .A2(n_301), .B1(n_507), .B2(n_509), .Y(n_506) );
INVx1_ASAP7_75t_L g773 ( .A(n_259), .Y(n_773) );
OAI22xp33_ASAP7_75t_L g659 ( .A1(n_260), .A2(n_262), .B1(n_329), .B2(n_544), .Y(n_659) );
OAI22xp33_ASAP7_75t_L g668 ( .A1(n_260), .A2(n_262), .B1(n_523), .B2(n_608), .Y(n_668) );
INVx1_ASAP7_75t_L g557 ( .A(n_261), .Y(n_557) );
INVx1_ASAP7_75t_L g941 ( .A(n_264), .Y(n_941) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_265), .B(n_1312), .Y(n_1311) );
INVx1_ASAP7_75t_L g1318 ( .A(n_265), .Y(n_1318) );
INVx1_ASAP7_75t_L g757 ( .A(n_266), .Y(n_757) );
INVx1_ASAP7_75t_L g1120 ( .A(n_268), .Y(n_1120) );
CKINVDCx5p33_ASAP7_75t_R g1059 ( .A(n_269), .Y(n_1059) );
CKINVDCx5p33_ASAP7_75t_R g672 ( .A(n_270), .Y(n_672) );
INVx1_ASAP7_75t_L g1257 ( .A(n_271), .Y(n_1257) );
INVx1_ASAP7_75t_L g1129 ( .A(n_272), .Y(n_1129) );
INVx1_ASAP7_75t_L g780 ( .A(n_273), .Y(n_780) );
INVx1_ASAP7_75t_L g1377 ( .A(n_274), .Y(n_1377) );
CKINVDCx5p33_ASAP7_75t_R g1635 ( .A(n_275), .Y(n_1635) );
OAI211xp5_ASAP7_75t_SL g1029 ( .A1(n_277), .A2(n_958), .B(n_983), .C(n_1030), .Y(n_1029) );
OAI211xp5_ASAP7_75t_SL g1038 ( .A1(n_277), .A2(n_492), .B(n_1039), .C(n_1040), .Y(n_1038) );
INVx1_ASAP7_75t_L g1234 ( .A(n_278), .Y(n_1234) );
INVx1_ASAP7_75t_L g868 ( .A(n_279), .Y(n_868) );
OAI211xp5_ASAP7_75t_SL g876 ( .A1(n_279), .A2(n_492), .B(n_877), .C(n_879), .Y(n_876) );
INVx1_ASAP7_75t_L g975 ( .A(n_280), .Y(n_975) );
XOR2x2_ASAP7_75t_L g1213 ( .A(n_282), .B(n_1214), .Y(n_1213) );
OAI211xp5_ASAP7_75t_L g652 ( .A1(n_283), .A2(n_533), .B(n_653), .C(n_654), .Y(n_652) );
INVx1_ASAP7_75t_L g667 ( .A(n_283), .Y(n_667) );
INVxp67_ASAP7_75t_SL g1181 ( .A(n_286), .Y(n_1181) );
INVx1_ASAP7_75t_L g738 ( .A(n_287), .Y(n_738) );
OAI211xp5_ASAP7_75t_L g747 ( .A1(n_287), .A2(n_602), .B(n_603), .C(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g1160 ( .A(n_288), .Y(n_1160) );
INVx1_ASAP7_75t_L g903 ( .A(n_290), .Y(n_903) );
CKINVDCx5p33_ASAP7_75t_R g674 ( .A(n_291), .Y(n_674) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_292), .Y(n_333) );
INVx1_ASAP7_75t_L g630 ( .A(n_294), .Y(n_630) );
CKINVDCx5p33_ASAP7_75t_R g1534 ( .A(n_295), .Y(n_1534) );
INVx1_ASAP7_75t_L g721 ( .A(n_296), .Y(n_721) );
CKINVDCx5p33_ASAP7_75t_R g677 ( .A(n_297), .Y(n_677) );
CKINVDCx5p33_ASAP7_75t_R g1082 ( .A(n_299), .Y(n_1082) );
CKINVDCx5p33_ASAP7_75t_R g1007 ( .A(n_302), .Y(n_1007) );
XOR2x2_ASAP7_75t_L g649 ( .A(n_304), .B(n_650), .Y(n_649) );
INVx2_ASAP7_75t_L g351 ( .A(n_305), .Y(n_351) );
INVx1_ASAP7_75t_L g387 ( .A(n_305), .Y(n_387) );
INVx1_ASAP7_75t_L g433 ( .A(n_305), .Y(n_433) );
INVx1_ASAP7_75t_L g1516 ( .A(n_306), .Y(n_1516) );
AOI22xp33_ASAP7_75t_L g1606 ( .A1(n_306), .A2(n_1607), .B1(n_1609), .B2(n_1645), .Y(n_1606) );
INVx1_ASAP7_75t_L g841 ( .A(n_307), .Y(n_841) );
INVx1_ASAP7_75t_L g844 ( .A(n_308), .Y(n_844) );
INVx1_ASAP7_75t_L g632 ( .A(n_309), .Y(n_632) );
INVx1_ASAP7_75t_L g566 ( .A(n_310), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g1067 ( .A(n_311), .Y(n_1067) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_338), .B(n_1301), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_323), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g1605 ( .A(n_317), .B(n_326), .Y(n_1605) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g1608 ( .A(n_319), .B(n_322), .Y(n_1608) );
INVx1_ASAP7_75t_L g1648 ( .A(n_319), .Y(n_1648) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g1650 ( .A(n_322), .B(n_1648), .Y(n_1650) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_328), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x4_ASAP7_75t_L g476 ( .A(n_326), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g382 ( .A(n_327), .B(n_337), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_328), .A2(n_442), .B1(n_780), .B2(n_781), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g1295 ( .A1(n_328), .A2(n_442), .B1(n_1257), .B2(n_1258), .Y(n_1295) );
AND2x4_ASAP7_75t_SL g1604 ( .A(n_328), .B(n_1605), .Y(n_1604) );
INVx3_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OR2x6_ASAP7_75t_L g329 ( .A(n_330), .B(n_335), .Y(n_329) );
OR2x6_ASAP7_75t_L g471 ( .A(n_330), .B(n_443), .Y(n_471) );
BUFx4f_ASAP7_75t_L g618 ( .A(n_330), .Y(n_618) );
OR2x2_ASAP7_75t_L g1034 ( .A(n_330), .B(n_443), .Y(n_1034) );
INVx1_ASAP7_75t_L g1138 ( .A(n_330), .Y(n_1138) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx4f_ASAP7_75t_L g356 ( .A(n_331), .Y(n_356) );
INVx3_ASAP7_75t_L g390 ( .A(n_331), .Y(n_390) );
INVx3_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx2_ASAP7_75t_L g363 ( .A(n_333), .Y(n_363) );
INVx2_ASAP7_75t_L g369 ( .A(n_333), .Y(n_369) );
NAND2x1_ASAP7_75t_L g372 ( .A(n_333), .B(n_334), .Y(n_372) );
AND2x2_ASAP7_75t_L g445 ( .A(n_333), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g462 ( .A(n_333), .Y(n_462) );
AND2x2_ASAP7_75t_L g468 ( .A(n_333), .B(n_334), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_334), .B(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g368 ( .A(n_334), .B(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g446 ( .A(n_334), .Y(n_446) );
BUFx2_ASAP7_75t_L g456 ( .A(n_334), .Y(n_456) );
INVx1_ASAP7_75t_L g794 ( .A(n_334), .Y(n_794) );
AND2x2_ASAP7_75t_L g808 ( .A(n_334), .B(n_363), .Y(n_808) );
OR2x6_ASAP7_75t_L g899 ( .A(n_335), .B(n_390), .Y(n_899) );
INVxp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g466 ( .A(n_336), .Y(n_466) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx2_ASAP7_75t_L g455 ( .A(n_337), .Y(n_455) );
AND2x4_ASAP7_75t_L g460 ( .A(n_337), .B(n_461), .Y(n_460) );
XNOR2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_1094), .Y(n_338) );
AOI22xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .B1(n_831), .B2(n_832), .Y(n_339) );
INVx2_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
XOR2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_582), .Y(n_341) );
OA21x2_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_518), .B(n_581), .Y(n_342) );
INVx2_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g581 ( .A(n_344), .B(n_519), .Y(n_581) );
NAND3xp33_ASAP7_75t_L g345 ( .A(n_346), .B(n_439), .C(n_479), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_347), .B(n_393), .Y(n_346) );
OAI33xp33_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_353), .A3(n_364), .B1(n_373), .B2(n_380), .B3(n_388), .Y(n_347) );
OAI33xp33_ASAP7_75t_L g568 ( .A1(n_348), .A2(n_569), .A3(n_572), .B1(n_577), .B2(n_579), .B3(n_580), .Y(n_568) );
OAI33xp33_ASAP7_75t_L g901 ( .A1(n_348), .A2(n_579), .A3(n_902), .B1(n_905), .B2(n_908), .B3(n_911), .Y(n_901) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g615 ( .A(n_349), .Y(n_615) );
INVx1_ASAP7_75t_L g675 ( .A(n_349), .Y(n_675) );
INVx2_ASAP7_75t_L g801 ( .A(n_349), .Y(n_801) );
INVx4_ASAP7_75t_L g1196 ( .A(n_349), .Y(n_1196) );
AND2x4_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
OR2x6_ASAP7_75t_L g951 ( .A(n_350), .B(n_952), .Y(n_951) );
OR2x2_ASAP7_75t_L g1018 ( .A(n_350), .B(n_952), .Y(n_1018) );
BUFx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g1156 ( .A(n_351), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1594 ( .A(n_351), .B(n_1572), .Y(n_1594) );
OAI22xp5_ASAP7_75t_SL g353 ( .A1(n_354), .A2(n_355), .B1(n_357), .B2(n_358), .Y(n_353) );
OAI22xp33_ASAP7_75t_L g399 ( .A1(n_354), .A2(n_377), .B1(n_400), .B2(n_407), .Y(n_399) );
INVx2_ASAP7_75t_SL g571 ( .A(n_355), .Y(n_571) );
INVx3_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_356), .Y(n_635) );
INVx4_ASAP7_75t_L g1070 ( .A(n_356), .Y(n_1070) );
OAI22xp33_ASAP7_75t_L g435 ( .A1(n_357), .A2(n_379), .B1(n_400), .B2(n_436), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_358), .A2(n_389), .B1(n_391), .B2(n_392), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_358), .A2(n_549), .B1(n_566), .B2(n_570), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_358), .A2(n_557), .B1(n_563), .B2(n_570), .Y(n_580) );
OAI22xp33_ASAP7_75t_L g671 ( .A1(n_358), .A2(n_672), .B1(n_673), .B2(n_674), .Y(n_671) );
OAI22xp33_ASAP7_75t_L g684 ( .A1(n_358), .A2(n_673), .B1(n_685), .B2(n_686), .Y(n_684) );
OAI22xp33_ASAP7_75t_L g840 ( .A1(n_358), .A2(n_389), .B1(n_841), .B2(n_842), .Y(n_840) );
INVx6_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx5_ASAP7_75t_L g620 ( .A(n_359), .Y(n_620) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g854 ( .A(n_360), .Y(n_854) );
INVx4_ASAP7_75t_L g956 ( .A(n_360), .Y(n_956) );
INVx2_ASAP7_75t_L g964 ( .A(n_360), .Y(n_964) );
INVx1_ASAP7_75t_L g1133 ( .A(n_360), .Y(n_1133) );
INVx2_ASAP7_75t_SL g1243 ( .A(n_360), .Y(n_1243) );
INVx8_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g474 ( .A(n_361), .B(n_455), .Y(n_474) );
OR2x2_ASAP7_75t_L g994 ( .A(n_361), .B(n_466), .Y(n_994) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_366), .B1(n_370), .B2(n_371), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_365), .A2(n_391), .B1(n_415), .B2(n_420), .Y(n_414) );
OAI221xp5_ASAP7_75t_L g802 ( .A1(n_366), .A2(n_533), .B1(n_763), .B2(n_770), .C(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g848 ( .A(n_366), .Y(n_848) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx2_ASAP7_75t_L g574 ( .A(n_367), .Y(n_574) );
INVx2_ASAP7_75t_L g1072 ( .A(n_367), .Y(n_1072) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx2_ASAP7_75t_L g376 ( .A(n_368), .Y(n_376) );
BUFx3_ASAP7_75t_L g629 ( .A(n_368), .Y(n_629) );
INVx1_ASAP7_75t_L g679 ( .A(n_368), .Y(n_679) );
BUFx2_ASAP7_75t_L g1075 ( .A(n_368), .Y(n_1075) );
AND2x2_ASAP7_75t_L g793 ( .A(n_369), .B(n_794), .Y(n_793) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_370), .A2(n_392), .B1(n_425), .B2(n_426), .Y(n_424) );
BUFx2_ASAP7_75t_SL g378 ( .A(n_371), .Y(n_378) );
BUFx3_ASAP7_75t_L g533 ( .A(n_371), .Y(n_533) );
INVx2_ASAP7_75t_SL g626 ( .A(n_371), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g1074 ( .A1(n_371), .A2(n_1056), .B1(n_1067), .B2(n_1075), .Y(n_1074) );
OAI22xp5_ASAP7_75t_L g1135 ( .A1(n_371), .A2(n_1022), .B1(n_1120), .B2(n_1130), .Y(n_1135) );
OR2x2_ASAP7_75t_L g1580 ( .A(n_371), .B(n_1578), .Y(n_1580) );
OAI22xp5_ASAP7_75t_L g1618 ( .A1(n_371), .A2(n_1072), .B1(n_1619), .B2(n_1620), .Y(n_1618) );
BUFx3_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_372), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_377), .B1(n_378), .B2(n_379), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g843 ( .A1(n_374), .A2(n_625), .B1(n_844), .B2(n_845), .Y(n_843) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx4_ASAP7_75t_L g623 ( .A(n_375), .Y(n_623) );
INVx4_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g846 ( .A1(n_378), .A2(n_847), .B1(n_849), .B2(n_850), .Y(n_846) );
OAI33xp33_ASAP7_75t_L g729 ( .A1(n_380), .A2(n_614), .A3(n_730), .B1(n_731), .B2(n_732), .B3(n_733), .Y(n_729) );
OAI33xp33_ASAP7_75t_L g839 ( .A1(n_380), .A2(n_614), .A3(n_840), .B1(n_843), .B2(n_846), .B3(n_851), .Y(n_839) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g579 ( .A(n_381), .Y(n_579) );
AOI33xp33_ASAP7_75t_L g1279 ( .A1(n_381), .A2(n_1280), .A3(n_1281), .B1(n_1284), .B2(n_1291), .B3(n_1292), .Y(n_1279) );
AND2x4_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
AND2x2_ASAP7_75t_SL g966 ( .A(n_382), .B(n_385), .Y(n_966) );
NAND2xp5_ASAP7_75t_L g1586 ( .A(n_382), .B(n_383), .Y(n_1586) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OR2x2_ASAP7_75t_L g395 ( .A(n_385), .B(n_396), .Y(n_395) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_385), .Y(n_517) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx2_ASAP7_75t_L g478 ( .A(n_386), .Y(n_478) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g851 ( .A1(n_389), .A2(n_852), .B1(n_853), .B2(n_855), .Y(n_851) );
BUFx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_SL g913 ( .A(n_390), .Y(n_913) );
BUFx3_ASAP7_75t_L g955 ( .A(n_390), .Y(n_955) );
BUFx6f_ASAP7_75t_L g962 ( .A(n_390), .Y(n_962) );
OAI33xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_399), .A3(n_414), .B1(n_424), .B2(n_428), .B3(n_435), .Y(n_393) );
OAI33xp33_ASAP7_75t_L g638 ( .A1(n_394), .A2(n_564), .A3(n_639), .B1(n_643), .B2(n_647), .B3(n_648), .Y(n_638) );
OAI33xp33_ASAP7_75t_L g709 ( .A1(n_394), .A2(n_710), .A3(n_715), .B1(n_718), .B2(n_723), .B3(n_726), .Y(n_709) );
BUFx4f_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx2_ASAP7_75t_L g547 ( .A(n_395), .Y(n_547) );
BUFx8_ASAP7_75t_L g688 ( .A(n_395), .Y(n_688) );
BUFx4f_ASAP7_75t_L g755 ( .A(n_395), .Y(n_755) );
NAND2xp33_ASAP7_75t_SL g396 ( .A(n_397), .B(n_398), .Y(n_396) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_397), .Y(n_515) );
AND3x4_ASAP7_75t_L g1155 ( .A(n_397), .B(n_500), .C(n_1156), .Y(n_1155) );
INVx1_ASAP7_75t_L g1524 ( .A(n_397), .Y(n_1524) );
AND2x2_ASAP7_75t_L g1531 ( .A(n_397), .B(n_500), .Y(n_1531) );
INVx3_ASAP7_75t_L g431 ( .A(n_398), .Y(n_431) );
BUFx3_ASAP7_75t_L g500 ( .A(n_398), .Y(n_500) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVxp67_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g691 ( .A(n_402), .Y(n_691) );
INVx1_ASAP7_75t_L g701 ( .A(n_402), .Y(n_701) );
BUFx3_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OR2x4_ASAP7_75t_L g483 ( .A(n_403), .B(n_431), .Y(n_483) );
OR2x4_ASAP7_75t_L g508 ( .A(n_403), .B(n_486), .Y(n_508) );
BUFx3_ASAP7_75t_L g550 ( .A(n_403), .Y(n_550) );
INVx2_ASAP7_75t_L g642 ( .A(n_403), .Y(n_642) );
BUFx4f_ASAP7_75t_L g936 ( .A(n_403), .Y(n_936) );
OR2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_404), .Y(n_413) );
INVx2_ASAP7_75t_L g419 ( .A(n_404), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_404), .B(n_412), .Y(n_423) );
AND2x4_ASAP7_75t_L g494 ( .A(n_404), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g1149 ( .A(n_405), .Y(n_1149) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVxp67_ASAP7_75t_L g418 ( .A(n_406), .Y(n_418) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx6f_ASAP7_75t_L g776 ( .A(n_409), .Y(n_776) );
OAI22xp5_ASAP7_75t_L g1015 ( .A1(n_409), .A2(n_936), .B1(n_1016), .B2(n_1017), .Y(n_1015) );
OAI22xp33_ASAP7_75t_L g1065 ( .A1(n_409), .A2(n_760), .B1(n_1066), .B2(n_1067), .Y(n_1065) );
OAI22xp33_ASAP7_75t_L g1128 ( .A1(n_409), .A2(n_936), .B1(n_1129), .B2(n_1130), .Y(n_1128) );
OAI22xp33_ASAP7_75t_L g1246 ( .A1(n_409), .A2(n_760), .B1(n_1233), .B2(n_1239), .Y(n_1246) );
OAI22xp33_ASAP7_75t_L g1631 ( .A1(n_409), .A2(n_760), .B1(n_1617), .B2(n_1623), .Y(n_1631) );
BUFx3_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx2_ASAP7_75t_L g438 ( .A(n_410), .Y(n_438) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_410), .Y(n_491) );
NAND2x1p5_ASAP7_75t_L g410 ( .A(n_411), .B(n_413), .Y(n_410) );
BUFx2_ASAP7_75t_L g504 ( .A(n_411), .Y(n_504) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g495 ( .A(n_412), .Y(n_495) );
BUFx2_ASAP7_75t_L g501 ( .A(n_413), .Y(n_501) );
INVx2_ASAP7_75t_L g1043 ( .A(n_413), .Y(n_1043) );
AND2x4_ASAP7_75t_L g1153 ( .A(n_413), .B(n_1046), .Y(n_1153) );
BUFx3_ASAP7_75t_L g556 ( .A(n_415), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_415), .A2(n_420), .B1(n_624), .B2(n_637), .Y(n_647) );
INVx8_ASAP7_75t_L g720 ( .A(n_415), .Y(n_720) );
INVx5_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_SL g425 ( .A(n_416), .Y(n_425) );
INVx3_ASAP7_75t_L g561 ( .A(n_416), .Y(n_561) );
INVx2_ASAP7_75t_SL g764 ( .A(n_416), .Y(n_764) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_417), .Y(n_487) );
BUFx8_ASAP7_75t_L g769 ( .A(n_417), .Y(n_769) );
INVx2_ASAP7_75t_L g925 ( .A(n_417), .Y(n_925) );
AND2x4_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
AND2x4_ASAP7_75t_L g1148 ( .A(n_419), .B(n_1149), .Y(n_1148) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_420), .A2(n_555), .B1(n_556), .B2(n_557), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_420), .A2(n_719), .B1(n_721), .B2(n_722), .Y(n_718) );
OAI22xp33_ASAP7_75t_L g919 ( .A1(n_420), .A2(n_906), .B1(n_914), .B2(n_920), .Y(n_919) );
CKINVDCx8_ASAP7_75t_R g420 ( .A(n_421), .Y(n_420) );
INVx3_ASAP7_75t_L g766 ( .A(n_421), .Y(n_766) );
INVx3_ASAP7_75t_L g1010 ( .A(n_421), .Y(n_1010) );
INVx3_ASAP7_75t_L g1014 ( .A(n_421), .Y(n_1014) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g772 ( .A(n_422), .Y(n_772) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx2_ASAP7_75t_L g427 ( .A(n_423), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_425), .A2(n_622), .B1(n_636), .B2(n_644), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g1011 ( .A1(n_425), .A2(n_1012), .B1(n_1013), .B2(n_1014), .Y(n_1011) );
OAI22xp5_ASAP7_75t_L g1630 ( .A1(n_425), .A2(n_766), .B1(n_1620), .B2(n_1626), .Y(n_1630) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_426), .A2(n_559), .B1(n_562), .B2(n_563), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g859 ( .A1(n_426), .A2(n_844), .B1(n_852), .B2(n_860), .Y(n_859) );
OAI22xp5_ASAP7_75t_L g861 ( .A1(n_426), .A2(n_845), .B1(n_855), .B2(n_862), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_426), .A2(n_907), .B1(n_915), .B2(n_923), .Y(n_922) );
BUFx3_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OR2x6_ASAP7_75t_L g511 ( .A(n_427), .B(n_431), .Y(n_511) );
INVx1_ASAP7_75t_L g646 ( .A(n_427), .Y(n_646) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_429), .Y(n_564) );
INVx2_ASAP7_75t_L g698 ( .A(n_429), .Y(n_698) );
INVx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx3_ASAP7_75t_L g725 ( .A(n_430), .Y(n_725) );
NAND3x1_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .C(n_434), .Y(n_430) );
INVx1_ASAP7_75t_L g486 ( .A(n_431), .Y(n_486) );
AND2x4_ASAP7_75t_L g493 ( .A(n_431), .B(n_494), .Y(n_493) );
NAND2x1p5_ASAP7_75t_L g952 ( .A(n_431), .B(n_434), .Y(n_952) );
AND2x4_ASAP7_75t_L g1523 ( .A(n_431), .B(n_1524), .Y(n_1523) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g1574 ( .A(n_433), .Y(n_1574) );
NAND2xp5_ASAP7_75t_L g1578 ( .A(n_433), .B(n_1564), .Y(n_1578) );
OAI22xp33_ASAP7_75t_L g565 ( .A1(n_436), .A2(n_550), .B1(n_566), .B2(n_567), .Y(n_565) );
OAI22xp33_ASAP7_75t_L g639 ( .A1(n_436), .A2(n_617), .B1(n_630), .B2(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g714 ( .A(n_438), .Y(n_714) );
INVx1_ASAP7_75t_L g878 ( .A(n_438), .Y(n_878) );
OR2x6_ASAP7_75t_L g1521 ( .A(n_438), .B(n_1522), .Y(n_1521) );
OAI221xp5_ASAP7_75t_L g1533 ( .A1(n_438), .A2(n_936), .B1(n_1534), .B2(n_1535), .C(n_1536), .Y(n_1533) );
OAI31xp33_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_447), .A3(n_469), .B(n_475), .Y(n_439) );
INVx4_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
CKINVDCx16_ASAP7_75t_R g544 ( .A(n_442), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g1178 ( .A1(n_442), .A2(n_1179), .B1(n_1180), .B2(n_1181), .Y(n_1178) );
AND2x4_ASAP7_75t_L g442 ( .A(n_443), .B(n_445), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
BUFx6f_ASAP7_75t_L g1202 ( .A(n_445), .Y(n_1202) );
INVx2_ASAP7_75t_L g1288 ( .A(n_445), .Y(n_1288) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_450), .A2(n_678), .B1(n_682), .B2(n_683), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_450), .A2(n_678), .B1(n_909), .B2(n_910), .Y(n_908) );
BUFx4f_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx4_ASAP7_75t_L g576 ( .A(n_451), .Y(n_576) );
BUFx4f_ASAP7_75t_L g631 ( .A(n_451), .Y(n_631) );
BUFx4f_ASAP7_75t_L g958 ( .A(n_451), .Y(n_958) );
BUFx6f_ASAP7_75t_L g960 ( .A(n_451), .Y(n_960) );
BUFx4f_ASAP7_75t_L g1023 ( .A(n_451), .Y(n_1023) );
OR2x6_ASAP7_75t_L g1600 ( .A(n_451), .B(n_1601), .Y(n_1600) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_457), .B1(n_458), .B2(n_463), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_453), .A2(n_867), .B1(n_868), .B2(n_869), .Y(n_866) );
BUFx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_454), .A2(n_460), .B1(n_591), .B2(n_592), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_454), .A2(n_737), .B1(n_738), .B2(n_739), .Y(n_736) );
INVx1_ASAP7_75t_L g788 ( .A(n_454), .Y(n_788) );
AOI22xp5_ASAP7_75t_L g1030 ( .A1(n_454), .A2(n_869), .B1(n_1031), .B2(n_1032), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_454), .A2(n_869), .B1(n_1103), .B2(n_1104), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g1218 ( .A1(n_454), .A2(n_869), .B1(n_1219), .B2(n_1220), .Y(n_1218) );
AND2x4_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
AND2x2_ASAP7_75t_L g536 ( .A(n_455), .B(n_456), .Y(n_536) );
AND2x2_ASAP7_75t_L g791 ( .A(n_455), .B(n_792), .Y(n_791) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_456), .B(n_466), .Y(n_1081) );
INVx1_ASAP7_75t_L g1596 ( .A(n_456), .Y(n_1596) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_457), .A2(n_497), .B1(n_502), .B2(n_505), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_458), .A2(n_526), .B1(n_536), .B2(n_537), .Y(n_535) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g656 ( .A(n_459), .Y(n_656) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g740 ( .A(n_460), .Y(n_740) );
BUFx3_ASAP7_75t_L g869 ( .A(n_460), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g1185 ( .A1(n_460), .A2(n_1081), .B1(n_1169), .B2(n_1173), .Y(n_1185) );
NAND2xp5_ASAP7_75t_L g1598 ( .A(n_461), .B(n_1572), .Y(n_1598) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g534 ( .A(n_465), .Y(n_534) );
INVx3_ASAP7_75t_L g653 ( .A(n_465), .Y(n_653) );
AOI211xp5_ASAP7_75t_L g782 ( .A1(n_465), .A2(n_783), .B(n_786), .C(n_787), .Y(n_782) );
NOR3xp33_ASAP7_75t_L g1296 ( .A(n_465), .B(n_1297), .C(n_1298), .Y(n_1296) );
AND2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
AND2x2_ASAP7_75t_L g984 ( .A(n_466), .B(n_985), .Y(n_984) );
BUFx6f_ASAP7_75t_L g785 ( .A(n_467), .Y(n_785) );
BUFx3_ASAP7_75t_L g988 ( .A(n_467), .Y(n_988) );
BUFx3_ASAP7_75t_L g1203 ( .A(n_467), .Y(n_1203) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g986 ( .A(n_468), .Y(n_986) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g539 ( .A(n_471), .Y(n_539) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g594 ( .A(n_473), .Y(n_594) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx2_ASAP7_75t_L g542 ( .A(n_474), .Y(n_542) );
INVx1_ASAP7_75t_L g798 ( .A(n_474), .Y(n_798) );
OAI31xp33_ASAP7_75t_L g529 ( .A1(n_475), .A2(n_530), .A3(n_538), .B(n_543), .Y(n_529) );
OAI31xp33_ASAP7_75t_SL g734 ( .A1(n_475), .A2(n_735), .A3(n_741), .B(n_742), .Y(n_734) );
OAI31xp33_ASAP7_75t_L g864 ( .A1(n_475), .A2(n_865), .A3(n_870), .B(n_871), .Y(n_864) );
BUFx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx2_ASAP7_75t_SL g595 ( .A(n_476), .Y(n_595) );
INVx1_ASAP7_75t_L g799 ( .A(n_476), .Y(n_799) );
OAI21xp5_ASAP7_75t_L g981 ( .A1(n_476), .A2(n_982), .B(n_995), .Y(n_981) );
OAI31xp33_ASAP7_75t_L g1027 ( .A1(n_476), .A2(n_1028), .A3(n_1029), .B(n_1033), .Y(n_1027) );
BUFx2_ASAP7_75t_L g1086 ( .A(n_476), .Y(n_1086) );
OAI31xp33_ASAP7_75t_L g1215 ( .A1(n_476), .A2(n_1216), .A3(n_1217), .B(n_1221), .Y(n_1215) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g1562 ( .A(n_478), .Y(n_1562) );
OR2x2_ASAP7_75t_L g1597 ( .A(n_478), .B(n_1598), .Y(n_1597) );
OAI31xp33_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_488), .A3(n_506), .B(n_512), .Y(n_479) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g609 ( .A(n_483), .Y(n_609) );
INVx1_ASAP7_75t_L g746 ( .A(n_483), .Y(n_746) );
INVx2_ASAP7_75t_SL g822 ( .A(n_483), .Y(n_822) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g523 ( .A(n_485), .Y(n_523) );
INVx1_ASAP7_75t_L g610 ( .A(n_485), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_485), .A2(n_780), .B1(n_781), .B2(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g1109 ( .A(n_485), .Y(n_1109) );
AOI22xp33_ASAP7_75t_L g1256 ( .A1(n_485), .A2(n_822), .B1(n_1257), .B2(n_1258), .Y(n_1256) );
AND2x4_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
AND2x2_ASAP7_75t_L g970 ( .A(n_486), .B(n_487), .Y(n_970) );
BUFx6f_ASAP7_75t_L g695 ( .A(n_487), .Y(n_695) );
INVx2_ASAP7_75t_L g697 ( .A(n_487), .Y(n_697) );
INVx2_ASAP7_75t_L g862 ( .A(n_487), .Y(n_862) );
BUFx6f_ASAP7_75t_L g921 ( .A(n_487), .Y(n_921) );
INVx2_ASAP7_75t_L g1008 ( .A(n_487), .Y(n_1008) );
OAI22xp33_ASAP7_75t_L g699 ( .A1(n_489), .A2(n_674), .B1(n_683), .B2(n_700), .Y(n_699) );
OAI22xp33_ASAP7_75t_L g726 ( .A1(n_489), .A2(n_640), .B1(n_727), .B2(n_728), .Y(n_726) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g602 ( .A(n_490), .Y(n_602) );
INVx2_ASAP7_75t_L g938 ( .A(n_490), .Y(n_938) );
INVx1_ASAP7_75t_L g1250 ( .A(n_490), .Y(n_1250) );
INVx1_ASAP7_75t_L g1263 ( .A(n_490), .Y(n_1263) );
INVx4_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx3_ASAP7_75t_L g553 ( .A(n_491), .Y(n_553) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_491), .Y(n_665) );
HB1xp67_ASAP7_75t_L g858 ( .A(n_491), .Y(n_858) );
OAI221xp5_ASAP7_75t_L g1528 ( .A1(n_491), .A2(n_862), .B1(n_1529), .B2(n_1530), .C(n_1531), .Y(n_1528) );
CKINVDCx8_ASAP7_75t_R g492 ( .A(n_493), .Y(n_492) );
CKINVDCx8_ASAP7_75t_R g603 ( .A(n_493), .Y(n_603) );
AOI211xp5_ASAP7_75t_L g815 ( .A1(n_493), .A2(n_816), .B(n_817), .C(n_818), .Y(n_815) );
NOR3xp33_ASAP7_75t_L g1259 ( .A(n_493), .B(n_1260), .C(n_1262), .Y(n_1259) );
BUFx3_ASAP7_75t_L g817 ( .A(n_494), .Y(n_817) );
BUFx2_ASAP7_75t_L g972 ( .A(n_494), .Y(n_972) );
BUFx2_ASAP7_75t_L g1145 ( .A(n_494), .Y(n_1145) );
INVx2_ASAP7_75t_L g1171 ( .A(n_494), .Y(n_1171) );
BUFx2_ASAP7_75t_L g1226 ( .A(n_494), .Y(n_1226) );
BUFx2_ASAP7_75t_L g1275 ( .A(n_494), .Y(n_1275) );
INVx1_ASAP7_75t_L g1046 ( .A(n_495), .Y(n_1046) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_497), .A2(n_502), .B1(n_526), .B2(n_527), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_497), .A2(n_502), .B1(n_867), .B2(n_880), .Y(n_879) );
BUFx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_501), .Y(n_498) );
AND2x4_ASAP7_75t_L g503 ( .A(n_499), .B(n_504), .Y(n_503) );
AND2x4_ASAP7_75t_L g605 ( .A(n_499), .B(n_501), .Y(n_605) );
AND2x4_ASAP7_75t_L g974 ( .A(n_499), .B(n_501), .Y(n_974) );
AND2x2_ASAP7_75t_L g976 ( .A(n_499), .B(n_504), .Y(n_976) );
INVx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_500), .B(n_1045), .Y(n_1044) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_503), .A2(n_591), .B1(n_605), .B2(n_606), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_503), .A2(n_605), .B1(n_655), .B2(n_667), .Y(n_666) );
AOI22xp33_ASAP7_75t_SL g748 ( .A1(n_503), .A2(n_605), .B1(n_737), .B2(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g820 ( .A(n_503), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_503), .A2(n_605), .B1(n_889), .B2(n_890), .Y(n_888) );
BUFx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_SL g824 ( .A(n_508), .Y(n_824) );
BUFx2_ASAP7_75t_L g874 ( .A(n_508), .Y(n_874) );
BUFx2_ASAP7_75t_L g1261 ( .A(n_508), .Y(n_1261) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g599 ( .A(n_511), .Y(n_599) );
INVx2_ASAP7_75t_L g825 ( .A(n_511), .Y(n_825) );
BUFx3_ASAP7_75t_L g875 ( .A(n_511), .Y(n_875) );
OAI31xp33_ASAP7_75t_L g521 ( .A1(n_512), .A2(n_522), .A3(n_524), .B(n_528), .Y(n_521) );
OAI31xp33_ASAP7_75t_L g872 ( .A1(n_512), .A2(n_873), .A3(n_876), .B(n_881), .Y(n_872) );
BUFx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_SL g513 ( .A(n_514), .B(n_516), .Y(n_513) );
AND2x2_ASAP7_75t_L g611 ( .A(n_514), .B(n_516), .Y(n_611) );
AND2x4_ASAP7_75t_L g827 ( .A(n_514), .B(n_516), .Y(n_827) );
AND2x2_ASAP7_75t_L g980 ( .A(n_514), .B(n_516), .Y(n_980) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_514), .B(n_516), .Y(n_1176) );
INVx1_ASAP7_75t_SL g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
NAND3xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_529), .C(n_545), .Y(n_520) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
OAI221xp5_ASAP7_75t_L g809 ( .A1(n_533), .A2(n_761), .B1(n_777), .B2(n_810), .C(n_812), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_536), .A2(n_655), .B1(n_656), .B2(n_657), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_536), .A2(n_656), .B1(n_889), .B2(n_896), .Y(n_895) );
AOI222xp33_ASAP7_75t_L g987 ( .A1(n_536), .A2(n_869), .B1(n_975), .B2(n_977), .C1(n_988), .C2(n_989), .Y(n_987) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_546), .B(n_568), .Y(n_545) );
OAI33xp33_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .A3(n_554), .B1(n_558), .B2(n_564), .B3(n_565), .Y(n_546) );
OAI33xp33_ASAP7_75t_L g856 ( .A1(n_547), .A2(n_564), .A3(n_857), .B1(n_859), .B2(n_861), .B3(n_863), .Y(n_856) );
OAI33xp33_ASAP7_75t_L g916 ( .A1(n_547), .A2(n_698), .A3(n_917), .B1(n_919), .B2(n_922), .B3(n_926), .Y(n_916) );
OAI33xp33_ASAP7_75t_L g934 ( .A1(n_547), .A2(n_935), .A3(n_940), .B1(n_944), .B2(n_948), .B3(n_951), .Y(n_934) );
OAI22xp33_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_550), .B1(n_551), .B2(n_552), .Y(n_548) );
OAI22xp33_ASAP7_75t_L g857 ( .A1(n_550), .A2(n_841), .B1(n_849), .B2(n_858), .Y(n_857) );
OAI22xp33_ASAP7_75t_L g863 ( .A1(n_550), .A2(n_713), .B1(n_842), .B2(n_850), .Y(n_863) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_551), .A2(n_567), .B1(n_573), .B2(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g692 ( .A(n_553), .Y(n_692) );
INVx3_ASAP7_75t_L g1004 ( .A(n_553), .Y(n_1004) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_555), .A2(n_562), .B1(n_573), .B2(n_575), .Y(n_572) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OAI22xp33_ASAP7_75t_SL g715 ( .A1(n_561), .A2(n_644), .B1(n_716), .B2(n_717), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g1247 ( .A1(n_561), .A2(n_1010), .B1(n_1236), .B2(n_1242), .Y(n_1247) );
OAI22xp5_ASAP7_75t_L g1537 ( .A1(n_561), .A2(n_766), .B1(n_1538), .B2(n_1539), .Y(n_1537) );
INVx1_ASAP7_75t_L g1278 ( .A(n_564), .Y(n_1278) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx4_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g578 ( .A(n_576), .Y(n_578) );
INVx1_ASAP7_75t_L g894 ( .A(n_576), .Y(n_894) );
INVx2_ASAP7_75t_L g1025 ( .A(n_576), .Y(n_1025) );
INVx2_ASAP7_75t_L g1073 ( .A(n_576), .Y(n_1073) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_578), .A2(n_677), .B1(n_678), .B2(n_680), .Y(n_676) );
OAI22xp33_ASAP7_75t_L g731 ( .A1(n_578), .A2(n_623), .B1(n_716), .B2(n_721), .Y(n_731) );
OAI33xp33_ASAP7_75t_L g613 ( .A1(n_579), .A2(n_614), .A3(n_616), .B1(n_621), .B2(n_627), .B3(n_633), .Y(n_613) );
OAI33xp33_ASAP7_75t_L g670 ( .A1(n_579), .A2(n_671), .A3(n_675), .B1(n_676), .B2(n_681), .B3(n_684), .Y(n_670) );
OAI22xp5_ASAP7_75t_SL g800 ( .A1(n_579), .A2(n_801), .B1(n_802), .B2(n_809), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_703), .B1(n_704), .B2(n_830), .Y(n_582) );
INVx1_ASAP7_75t_L g830 ( .A(n_583), .Y(n_830) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_585), .B1(n_649), .B2(n_702), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND3xp33_ASAP7_75t_L g586 ( .A(n_587), .B(n_596), .C(n_612), .Y(n_586) );
OAI31xp33_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .A3(n_593), .B(n_595), .Y(n_587) );
OAI31xp33_ASAP7_75t_L g651 ( .A1(n_595), .A2(n_652), .A3(n_658), .B(n_659), .Y(n_651) );
OAI31xp33_ASAP7_75t_L g892 ( .A1(n_595), .A2(n_893), .A3(n_897), .B(n_898), .Y(n_892) );
OAI31xp33_ASAP7_75t_SL g1099 ( .A1(n_595), .A2(n_1100), .A3(n_1105), .B(n_1106), .Y(n_1099) );
OAI31xp33_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_600), .A3(n_607), .B(n_611), .Y(n_596) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OAI22xp33_ASAP7_75t_L g648 ( .A1(n_602), .A2(n_619), .B1(n_632), .B2(n_640), .Y(n_648) );
NAND3xp33_ASAP7_75t_L g1110 ( .A(n_603), .B(n_1111), .C(n_1113), .Y(n_1110) );
NAND3xp33_ASAP7_75t_SL g1167 ( .A(n_603), .B(n_1168), .C(n_1172), .Y(n_1167) );
NAND3xp33_ASAP7_75t_SL g1224 ( .A(n_603), .B(n_1225), .C(n_1227), .Y(n_1224) );
INVx1_ASAP7_75t_L g819 ( .A(n_605), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_605), .A2(n_976), .B1(n_1103), .B2(n_1112), .Y(n_1111) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OAI31xp33_ASAP7_75t_L g660 ( .A1(n_611), .A2(n_661), .A3(n_662), .B(n_668), .Y(n_660) );
OAI31xp33_ASAP7_75t_L g743 ( .A1(n_611), .A2(n_744), .A3(n_747), .B(n_750), .Y(n_743) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_638), .Y(n_612) );
INVx1_ASAP7_75t_L g1280 ( .A(n_614), .Y(n_1280) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI33xp33_ASAP7_75t_L g1019 ( .A1(n_615), .A2(n_965), .A3(n_1020), .B1(n_1021), .B2(n_1024), .B3(n_1026), .Y(n_1019) );
OAI33xp33_ASAP7_75t_L g1231 ( .A1(n_615), .A2(n_1077), .A3(n_1232), .B1(n_1235), .B2(n_1238), .B3(n_1241), .Y(n_1231) );
OAI33xp33_ASAP7_75t_L g1614 ( .A1(n_615), .A2(n_1077), .A3(n_1615), .B1(n_1618), .B2(n_1621), .B3(n_1624), .Y(n_1614) );
OAI22xp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_618), .B1(n_619), .B2(n_620), .Y(n_616) );
OAI22xp33_ASAP7_75t_L g730 ( .A1(n_618), .A2(n_620), .B1(n_711), .B2(n_727), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_620), .A2(n_634), .B1(n_636), .B2(n_637), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_620), .A2(n_634), .B1(n_717), .B2(n_722), .Y(n_733) );
OAI22xp33_ASAP7_75t_L g902 ( .A1(n_620), .A2(n_673), .B1(n_903), .B2(n_904), .Y(n_902) );
OAI22xp5_ASAP7_75t_L g911 ( .A1(n_620), .A2(n_912), .B1(n_914), .B2(n_915), .Y(n_911) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_623), .B1(n_624), .B2(n_625), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_623), .A2(n_631), .B1(n_712), .B2(n_728), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g905 ( .A1(n_625), .A2(n_678), .B1(n_906), .B2(n_907), .Y(n_905) );
INVx5_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OAI22xp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_630), .B1(n_631), .B2(n_632), .Y(n_627) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g811 ( .A(n_629), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g957 ( .A1(n_629), .A2(n_941), .B1(n_946), .B2(n_958), .Y(n_957) );
OAI22xp5_ASAP7_75t_L g1024 ( .A1(n_629), .A2(n_1005), .B1(n_1017), .B2(n_1025), .Y(n_1024) );
OAI221xp5_ASAP7_75t_L g1584 ( .A1(n_629), .A2(n_1023), .B1(n_1530), .B2(n_1538), .C(n_1585), .Y(n_1584) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx3_ASAP7_75t_L g673 ( .A(n_635), .Y(n_673) );
OAI22xp33_ASAP7_75t_L g710 ( .A1(n_640), .A2(n_711), .B1(n_712), .B2(n_713), .Y(n_710) );
BUFx4f_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
INVx3_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_SL g760 ( .A(n_642), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_644), .A2(n_677), .B1(n_685), .B2(n_694), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_644), .A2(n_680), .B1(n_686), .B2(n_697), .Y(n_696) );
INVx3_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
BUFx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g1064 ( .A(n_646), .Y(n_1064) );
INVx1_ASAP7_75t_L g702 ( .A(n_649), .Y(n_702) );
NAND3xp33_ASAP7_75t_SL g650 ( .A(n_651), .B(n_660), .C(n_669), .Y(n_650) );
INVx2_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
OAI22xp33_ASAP7_75t_L g756 ( .A1(n_665), .A2(n_757), .B1(n_758), .B2(n_761), .Y(n_756) );
OAI22xp33_ASAP7_75t_L g926 ( .A1(n_665), .A2(n_690), .B1(n_904), .B2(n_910), .Y(n_926) );
OAI22xp33_ASAP7_75t_L g948 ( .A1(n_665), .A2(n_936), .B1(n_949), .B2(n_950), .Y(n_948) );
OAI22xp33_ASAP7_75t_L g1118 ( .A1(n_665), .A2(n_936), .B1(n_1119), .B2(n_1120), .Y(n_1118) );
OAI22xp33_ASAP7_75t_L g1628 ( .A1(n_665), .A2(n_760), .B1(n_1616), .B2(n_1622), .Y(n_1628) );
NOR2xp33_ASAP7_75t_SL g669 ( .A(n_670), .B(n_687), .Y(n_669) );
OAI22xp33_ASAP7_75t_L g689 ( .A1(n_672), .A2(n_682), .B1(n_690), .B2(n_692), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g959 ( .A1(n_678), .A2(n_939), .B1(n_950), .B2(n_960), .Y(n_959) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g1022 ( .A(n_679), .Y(n_1022) );
OAI33xp33_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_689), .A3(n_693), .B1(n_696), .B2(n_698), .B3(n_699), .Y(n_687) );
OAI22xp33_ASAP7_75t_L g917 ( .A1(n_690), .A2(n_903), .B1(n_909), .B2(n_918), .Y(n_917) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g860 ( .A(n_695), .Y(n_860) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_751), .B1(n_828), .B2(n_829), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
HB1xp67_ASAP7_75t_L g828 ( .A(n_706), .Y(n_828) );
NAND3xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_734), .C(n_743), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_709), .B(n_729), .Y(n_708) );
INVxp67_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
OAI33xp33_ASAP7_75t_L g753 ( .A1(n_723), .A2(n_754), .A3(n_756), .B1(n_762), .B2(n_767), .B3(n_774), .Y(n_753) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
BUFx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AOI22xp5_ASAP7_75t_L g1080 ( .A1(n_739), .A2(n_1081), .B1(n_1082), .B2(n_1083), .Y(n_1080) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g829 ( .A(n_751), .Y(n_829) );
NOR4xp25_ASAP7_75t_L g752 ( .A(n_753), .B(n_778), .C(n_800), .D(n_814), .Y(n_752) );
BUFx3_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
OAI33xp33_ASAP7_75t_L g1001 ( .A1(n_755), .A2(n_1002), .A3(n_1006), .B1(n_1011), .B2(n_1015), .B3(n_1018), .Y(n_1001) );
OAI33xp33_ASAP7_75t_L g1053 ( .A1(n_755), .A2(n_1018), .A3(n_1054), .B1(n_1057), .B2(n_1060), .B3(n_1065), .Y(n_1053) );
OAI33xp33_ASAP7_75t_L g1117 ( .A1(n_755), .A2(n_1018), .A3(n_1118), .B1(n_1121), .B2(n_1124), .B3(n_1128), .Y(n_1117) );
OAI33xp33_ASAP7_75t_L g1245 ( .A1(n_755), .A2(n_1018), .A3(n_1246), .B1(n_1247), .B2(n_1248), .B3(n_1249), .Y(n_1245) );
OAI33xp33_ASAP7_75t_L g1627 ( .A1(n_755), .A2(n_1018), .A3(n_1628), .B1(n_1629), .B2(n_1630), .B3(n_1631), .Y(n_1627) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx2_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
OAI22xp33_ASAP7_75t_L g774 ( .A1(n_760), .A2(n_775), .B1(n_776), .B2(n_777), .Y(n_774) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_764), .B1(n_765), .B2(n_766), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g944 ( .A1(n_766), .A2(n_945), .B1(n_946), .B2(n_947), .Y(n_944) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_770), .B1(n_771), .B2(n_773), .Y(n_767) );
INVx2_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
INVx3_ASAP7_75t_L g945 ( .A(n_769), .Y(n_945) );
INVx2_ASAP7_75t_SL g1125 ( .A(n_769), .Y(n_1125) );
OAI22xp5_ASAP7_75t_L g940 ( .A1(n_771), .A2(n_941), .B1(n_942), .B2(n_943), .Y(n_940) );
OAI22xp5_ASAP7_75t_L g1124 ( .A1(n_771), .A2(n_1125), .B1(n_1126), .B2(n_1127), .Y(n_1124) );
BUFx3_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
AOI31xp33_ASAP7_75t_SL g778 ( .A1(n_779), .A2(n_782), .A3(n_789), .B(n_799), .Y(n_778) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_791), .B1(n_795), .B2(n_796), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_790), .A2(n_795), .B1(n_824), .B2(n_825), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_791), .A2(n_991), .B1(n_992), .B2(n_993), .Y(n_990) );
BUFx6f_ASAP7_75t_L g813 ( .A(n_792), .Y(n_813) );
INVx3_ASAP7_75t_L g1207 ( .A(n_792), .Y(n_1207) );
BUFx6f_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx3_ASAP7_75t_L g805 ( .A(n_793), .Y(n_805) );
AND2x2_ASAP7_75t_L g1563 ( .A(n_793), .B(n_1564), .Y(n_1563) );
NAND2xp5_ASAP7_75t_L g1571 ( .A(n_793), .B(n_1572), .Y(n_1571) );
INVx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
AO21x1_ASAP7_75t_L g1177 ( .A1(n_799), .A2(n_1178), .B(n_1182), .Y(n_1177) );
AO21x1_ASAP7_75t_L g1294 ( .A1(n_799), .A2(n_1295), .B(n_1296), .Y(n_1294) );
OAI33xp33_ASAP7_75t_L g953 ( .A1(n_801), .A2(n_954), .A3(n_957), .B1(n_959), .B2(n_961), .B3(n_965), .Y(n_953) );
OAI33xp33_ASAP7_75t_L g1068 ( .A1(n_801), .A2(n_1069), .A3(n_1071), .B1(n_1074), .B2(n_1076), .B3(n_1077), .Y(n_1068) );
OAI33xp33_ASAP7_75t_L g1131 ( .A1(n_801), .A2(n_965), .A3(n_1132), .B1(n_1134), .B2(n_1135), .B3(n_1136), .Y(n_1131) );
OAI22xp5_ASAP7_75t_SL g1583 ( .A1(n_801), .A2(n_1584), .B1(n_1586), .B2(n_1587), .Y(n_1583) );
INVx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx2_ASAP7_75t_L g1198 ( .A(n_805), .Y(n_1198) );
INVx1_ASAP7_75t_L g1282 ( .A(n_805), .Y(n_1282) );
INVx2_ASAP7_75t_SL g1293 ( .A(n_805), .Y(n_1293) );
BUFx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
BUFx6f_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
BUFx3_ASAP7_75t_L g1199 ( .A(n_808), .Y(n_1199) );
INVx2_ASAP7_75t_L g1209 ( .A(n_808), .Y(n_1209) );
INVx3_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
AOI31xp33_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_821), .A3(n_823), .B(n_826), .Y(n_814) );
HB1xp67_ASAP7_75t_L g1114 ( .A(n_817), .Y(n_1114) );
INVx1_ASAP7_75t_L g1159 ( .A(n_817), .Y(n_1159) );
INVx2_ASAP7_75t_L g979 ( .A(n_825), .Y(n_979) );
AO21x1_ASAP7_75t_L g1255 ( .A1(n_826), .A2(n_1256), .B(n_1259), .Y(n_1255) );
CKINVDCx14_ASAP7_75t_R g826 ( .A(n_827), .Y(n_826) );
OAI31xp33_ASAP7_75t_L g885 ( .A1(n_827), .A2(n_886), .A3(n_887), .B(n_891), .Y(n_885) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
XOR2xp5_ASAP7_75t_L g832 ( .A(n_833), .B(n_929), .Y(n_832) );
INVx2_ASAP7_75t_SL g833 ( .A(n_834), .Y(n_833) );
OA22x2_ASAP7_75t_L g834 ( .A1(n_835), .A2(n_836), .B1(n_882), .B2(n_883), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
NAND3xp33_ASAP7_75t_L g837 ( .A(n_838), .B(n_864), .C(n_872), .Y(n_837) );
NOR2xp33_ASAP7_75t_SL g838 ( .A(n_839), .B(n_856), .Y(n_838) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
BUFx3_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
AOI22xp5_ASAP7_75t_L g1634 ( .A1(n_869), .A2(n_1081), .B1(n_1635), .B2(n_1636), .Y(n_1634) );
INVxp67_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g918 ( .A(n_878), .Y(n_918) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g927 ( .A(n_884), .Y(n_927) );
NAND3xp33_ASAP7_75t_L g884 ( .A(n_885), .B(n_892), .C(n_900), .Y(n_884) );
INVx1_ASAP7_75t_L g1180 ( .A(n_899), .Y(n_1180) );
NOR2xp33_ASAP7_75t_L g900 ( .A(n_901), .B(n_916), .Y(n_900) );
INVx2_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
INVx2_ASAP7_75t_SL g920 ( .A(n_921), .Y(n_920) );
INVx2_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
INVx2_ASAP7_75t_L g1062 ( .A(n_924), .Y(n_1062) );
INVx3_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
BUFx2_ASAP7_75t_L g942 ( .A(n_925), .Y(n_942) );
BUFx2_ASAP7_75t_L g1271 ( .A(n_925), .Y(n_1271) );
INVx1_ASAP7_75t_L g1277 ( .A(n_925), .Y(n_1277) );
XNOR2xp5_ASAP7_75t_L g929 ( .A(n_930), .B(n_996), .Y(n_929) );
HB1xp67_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
NAND3xp33_ASAP7_75t_L g932 ( .A(n_933), .B(n_967), .C(n_981), .Y(n_932) );
NOR2xp33_ASAP7_75t_L g933 ( .A(n_934), .B(n_953), .Y(n_933) );
OAI22xp33_ASAP7_75t_L g935 ( .A1(n_936), .A2(n_937), .B1(n_938), .B2(n_939), .Y(n_935) );
OAI22xp5_ASAP7_75t_L g1002 ( .A1(n_936), .A2(n_1003), .B1(n_1004), .B2(n_1005), .Y(n_1002) );
OAI22xp5_ASAP7_75t_L g1054 ( .A1(n_936), .A2(n_1004), .B1(n_1055), .B2(n_1056), .Y(n_1054) );
OAI22xp33_ASAP7_75t_L g1249 ( .A1(n_936), .A2(n_1234), .B1(n_1240), .B2(n_1250), .Y(n_1249) );
OAI22xp5_ASAP7_75t_L g954 ( .A1(n_937), .A2(n_949), .B1(n_955), .B2(n_956), .Y(n_954) );
OAI22xp5_ASAP7_75t_L g961 ( .A1(n_943), .A2(n_947), .B1(n_962), .B2(n_963), .Y(n_961) );
OAI22xp5_ASAP7_75t_L g1121 ( .A1(n_945), .A2(n_1064), .B1(n_1122), .B2(n_1123), .Y(n_1121) );
INVx1_ASAP7_75t_L g1164 ( .A(n_951), .Y(n_1164) );
INVx3_ASAP7_75t_L g1536 ( .A(n_952), .Y(n_1536) );
OAI22xp5_ASAP7_75t_L g1020 ( .A1(n_955), .A2(n_963), .B1(n_1003), .B2(n_1016), .Y(n_1020) );
OAI22xp5_ASAP7_75t_L g1026 ( .A1(n_955), .A2(n_956), .B1(n_1009), .B2(n_1013), .Y(n_1026) );
OAI22xp5_ASAP7_75t_L g1076 ( .A1(n_956), .A2(n_1059), .B1(n_1063), .B2(n_1070), .Y(n_1076) );
OAI22xp5_ASAP7_75t_L g1136 ( .A1(n_956), .A2(n_1123), .B1(n_1127), .B2(n_1137), .Y(n_1136) );
HB1xp67_ASAP7_75t_L g1101 ( .A(n_960), .Y(n_1101) );
OAI22xp5_ASAP7_75t_L g1235 ( .A1(n_960), .A2(n_1072), .B1(n_1236), .B2(n_1237), .Y(n_1235) );
OAI221xp5_ASAP7_75t_L g1587 ( .A1(n_960), .A2(n_1072), .B1(n_1529), .B2(n_1534), .C(n_1588), .Y(n_1587) );
OAI22xp5_ASAP7_75t_L g1621 ( .A1(n_960), .A2(n_1072), .B1(n_1622), .B2(n_1623), .Y(n_1621) );
OAI22xp5_ASAP7_75t_L g1069 ( .A1(n_963), .A2(n_1055), .B1(n_1066), .B2(n_1070), .Y(n_1069) );
OAI22xp5_ASAP7_75t_L g1232 ( .A1(n_963), .A2(n_1070), .B1(n_1233), .B2(n_1234), .Y(n_1232) );
OAI22xp5_ASAP7_75t_L g1624 ( .A1(n_963), .A2(n_1070), .B1(n_1625), .B2(n_1626), .Y(n_1624) );
BUFx6f_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
INVx2_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
INVx2_ASAP7_75t_L g1077 ( .A(n_966), .Y(n_1077) );
AOI33xp33_ASAP7_75t_L g1194 ( .A1(n_966), .A2(n_1195), .A3(n_1197), .B1(n_1200), .B2(n_1204), .B3(n_1205), .Y(n_1194) );
OAI21xp5_ASAP7_75t_L g967 ( .A1(n_968), .A2(n_978), .B(n_980), .Y(n_967) );
INVx2_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
AOI222xp33_ASAP7_75t_L g971 ( .A1(n_972), .A2(n_973), .B1(n_974), .B2(n_975), .C1(n_976), .C2(n_977), .Y(n_971) );
AOI22xp5_ASAP7_75t_L g1040 ( .A1(n_974), .A2(n_1031), .B1(n_1041), .B2(n_1044), .Y(n_1040) );
AOI22xp33_ASAP7_75t_SL g1090 ( .A1(n_974), .A2(n_976), .B1(n_1082), .B2(n_1091), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g1172 ( .A1(n_974), .A2(n_976), .B1(n_1173), .B2(n_1174), .Y(n_1172) );
AOI22xp33_ASAP7_75t_L g1227 ( .A1(n_974), .A2(n_976), .B1(n_1219), .B2(n_1228), .Y(n_1227) );
AOI22xp33_ASAP7_75t_SL g1642 ( .A1(n_974), .A2(n_976), .B1(n_1635), .B2(n_1643), .Y(n_1642) );
INVxp67_ASAP7_75t_L g1039 ( .A(n_976), .Y(n_1039) );
OAI31xp33_ASAP7_75t_SL g1035 ( .A1(n_980), .A2(n_1036), .A3(n_1037), .B(n_1038), .Y(n_1035) );
OAI31xp33_ASAP7_75t_SL g1087 ( .A1(n_980), .A2(n_1088), .A3(n_1089), .B(n_1092), .Y(n_1087) );
OAI31xp33_ASAP7_75t_L g1107 ( .A1(n_980), .A2(n_1108), .A3(n_1110), .B(n_1115), .Y(n_1107) );
OAI31xp33_ASAP7_75t_SL g1639 ( .A1(n_980), .A2(n_1640), .A3(n_1641), .B(n_1644), .Y(n_1639) );
NAND3xp33_ASAP7_75t_SL g982 ( .A(n_983), .B(n_987), .C(n_990), .Y(n_982) );
INVx2_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
INVx2_ASAP7_75t_L g1189 ( .A(n_984), .Y(n_1189) );
INVx1_ASAP7_75t_L g1188 ( .A(n_985), .Y(n_1188) );
INVx1_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
BUFx2_ASAP7_75t_L g1290 ( .A(n_986), .Y(n_1290) );
INVx1_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
AOI22xp5_ASAP7_75t_L g996 ( .A1(n_997), .A2(n_1047), .B1(n_1048), .B2(n_1093), .Y(n_996) );
INVx1_ASAP7_75t_L g1093 ( .A(n_997), .Y(n_1093) );
INVx1_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
NAND3xp33_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1027), .C(n_1035), .Y(n_999) );
NOR2xp33_ASAP7_75t_SL g1000 ( .A(n_1001), .B(n_1019), .Y(n_1000) );
OAI22xp5_ASAP7_75t_L g1006 ( .A1(n_1007), .A2(n_1008), .B1(n_1009), .B2(n_1010), .Y(n_1006) );
OAI22xp5_ASAP7_75t_L g1021 ( .A1(n_1007), .A2(n_1012), .B1(n_1022), .B2(n_1023), .Y(n_1021) );
OAI22xp5_ASAP7_75t_L g1057 ( .A1(n_1008), .A2(n_1010), .B1(n_1058), .B2(n_1059), .Y(n_1057) );
OAI22xp5_ASAP7_75t_L g1248 ( .A1(n_1008), .A2(n_1014), .B1(n_1237), .B2(n_1244), .Y(n_1248) );
OAI22xp5_ASAP7_75t_L g1629 ( .A1(n_1008), .A2(n_1010), .B1(n_1619), .B2(n_1625), .Y(n_1629) );
OAI22xp5_ASAP7_75t_L g1134 ( .A1(n_1022), .A2(n_1073), .B1(n_1122), .B2(n_1126), .Y(n_1134) );
OAI22xp5_ASAP7_75t_L g1238 ( .A1(n_1023), .A2(n_1072), .B1(n_1239), .B2(n_1240), .Y(n_1238) );
AND2x6_ASAP7_75t_L g1555 ( .A(n_1042), .B(n_1523), .Y(n_1555) );
INVx3_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1557 ( .A(n_1045), .B(n_1523), .Y(n_1557) );
INVx1_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
INVx1_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
HB1xp67_ASAP7_75t_L g1048 ( .A(n_1049), .Y(n_1048) );
XNOR2xp5_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1051), .Y(n_1049) );
AND3x1_ASAP7_75t_L g1051 ( .A(n_1052), .B(n_1078), .C(n_1087), .Y(n_1051) );
NOR2xp33_ASAP7_75t_SL g1052 ( .A(n_1053), .B(n_1068), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g1071 ( .A1(n_1058), .A2(n_1061), .B1(n_1072), .B2(n_1073), .Y(n_1071) );
OAI22xp5_ASAP7_75t_L g1060 ( .A1(n_1061), .A2(n_1062), .B1(n_1063), .B2(n_1064), .Y(n_1060) );
OAI22xp33_ASAP7_75t_L g1132 ( .A1(n_1070), .A2(n_1119), .B1(n_1129), .B2(n_1133), .Y(n_1132) );
OAI22xp5_ASAP7_75t_L g1241 ( .A1(n_1070), .A2(n_1242), .B1(n_1243), .B2(n_1244), .Y(n_1241) );
OAI22xp5_ASAP7_75t_L g1615 ( .A1(n_1070), .A2(n_1243), .B1(n_1616), .B2(n_1617), .Y(n_1615) );
OAI31xp33_ASAP7_75t_L g1078 ( .A1(n_1079), .A2(n_1084), .A3(n_1085), .B(n_1086), .Y(n_1078) );
OAI31xp33_ASAP7_75t_L g1632 ( .A1(n_1086), .A2(n_1633), .A3(n_1637), .B(n_1638), .Y(n_1632) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
XNOR2xp5_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1139), .Y(n_1095) );
INVx2_ASAP7_75t_SL g1096 ( .A(n_1097), .Y(n_1096) );
NAND3xp33_ASAP7_75t_L g1098 ( .A(n_1099), .B(n_1107), .C(n_1116), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g1113 ( .A(n_1104), .B(n_1114), .Y(n_1113) );
NOR2xp33_ASAP7_75t_L g1116 ( .A(n_1117), .B(n_1131), .Y(n_1116) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
AOI22xp5_ASAP7_75t_L g1139 ( .A1(n_1140), .A2(n_1251), .B1(n_1299), .B2(n_1300), .Y(n_1139) );
INVx2_ASAP7_75t_L g1300 ( .A(n_1140), .Y(n_1300) );
XNOR2x1_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1213), .Y(n_1140) );
OR2x2_ASAP7_75t_L g1141 ( .A(n_1142), .B(n_1190), .Y(n_1141) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1143), .Y(n_1192) );
AOI21xp5_ASAP7_75t_L g1143 ( .A1(n_1144), .A2(n_1150), .B(n_1157), .Y(n_1143) );
INVx2_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
INVx8_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
BUFx3_ASAP7_75t_L g1162 ( .A(n_1148), .Y(n_1162) );
BUFx3_ASAP7_75t_L g1527 ( .A(n_1148), .Y(n_1527) );
NAND2x1p5_ASAP7_75t_L g1546 ( .A(n_1148), .B(n_1523), .Y(n_1546) );
INVx2_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1152), .Y(n_1272) );
INVx5_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
BUFx12f_ASAP7_75t_L g1526 ( .A(n_1153), .Y(n_1526) );
AND2x4_ASAP7_75t_L g1541 ( .A(n_1153), .B(n_1542), .Y(n_1541) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
BUFx3_ASAP7_75t_L g1265 ( .A(n_1155), .Y(n_1265) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1156), .Y(n_1559) );
OAI221xp5_ASAP7_75t_L g1158 ( .A1(n_1159), .A2(n_1160), .B1(n_1161), .B2(n_1163), .C(n_1164), .Y(n_1158) );
INVx2_ASAP7_75t_L g1268 ( .A(n_1161), .Y(n_1268) );
INVx2_ASAP7_75t_SL g1161 ( .A(n_1162), .Y(n_1161) );
NAND2xp5_ASAP7_75t_L g1549 ( .A(n_1162), .B(n_1550), .Y(n_1549) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1165), .B(n_1177), .Y(n_1191) );
OAI31xp33_ASAP7_75t_SL g1165 ( .A1(n_1166), .A2(n_1167), .A3(n_1175), .B(n_1176), .Y(n_1165) );
NAND2xp5_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1170), .Y(n_1168) );
INVx2_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g1186 ( .A(n_1174), .B(n_1187), .Y(n_1186) );
OAI31xp33_ASAP7_75t_SL g1222 ( .A1(n_1176), .A2(n_1223), .A3(n_1224), .B(n_1229), .Y(n_1222) );
NOR2xp33_ASAP7_75t_L g1182 ( .A(n_1183), .B(n_1184), .Y(n_1182) );
NAND3xp33_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1186), .C(n_1189), .Y(n_1184) );
INVx2_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
OAI31xp33_ASAP7_75t_L g1190 ( .A1(n_1191), .A2(n_1192), .A3(n_1193), .B(n_1210), .Y(n_1190) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1194), .Y(n_1212) );
INVx2_ASAP7_75t_SL g1195 ( .A(n_1196), .Y(n_1195) );
HB1xp67_ASAP7_75t_L g1283 ( .A(n_1199), .Y(n_1283) );
BUFx6f_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1568 ( .A(n_1202), .B(n_1564), .Y(n_1568) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
INVx3_ASAP7_75t_L g1576 ( .A(n_1209), .Y(n_1576) );
NAND2xp5_ASAP7_75t_L g1210 ( .A(n_1211), .B(n_1212), .Y(n_1210) );
NAND3xp33_ASAP7_75t_SL g1214 ( .A(n_1215), .B(n_1222), .C(n_1230), .Y(n_1214) );
NAND2xp5_ASAP7_75t_L g1225 ( .A(n_1220), .B(n_1226), .Y(n_1225) );
NOR2xp33_ASAP7_75t_L g1230 ( .A(n_1231), .B(n_1245), .Y(n_1230) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1253), .Y(n_1252) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1253), .Y(n_1299) );
NAND4xp25_ASAP7_75t_SL g1254 ( .A(n_1255), .B(n_1264), .C(n_1279), .D(n_1294), .Y(n_1254) );
AOI33xp33_ASAP7_75t_L g1264 ( .A1(n_1265), .A2(n_1266), .A3(n_1269), .B1(n_1273), .B2(n_1276), .B3(n_1278), .Y(n_1264) );
BUFx2_ASAP7_75t_SL g1267 ( .A(n_1268), .Y(n_1267) );
INVx2_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
BUFx2_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
INVx2_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
INVx2_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
INVx2_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1290), .Y(n_1289) );
OAI221xp5_ASAP7_75t_SL g1301 ( .A1(n_1302), .A2(n_1512), .B1(n_1514), .B2(n_1602), .C(n_1606), .Y(n_1301) );
AND5x1_ASAP7_75t_L g1302 ( .A(n_1303), .B(n_1468), .C(n_1485), .D(n_1494), .E(n_1505), .Y(n_1302) );
OAI33xp33_ASAP7_75t_L g1303 ( .A1(n_1304), .A2(n_1396), .A3(n_1413), .B1(n_1422), .B2(n_1449), .B3(n_1463), .Y(n_1303) );
OAI211xp5_ASAP7_75t_SL g1304 ( .A1(n_1305), .A2(n_1326), .B(n_1343), .C(n_1386), .Y(n_1304) );
CKINVDCx5p33_ASAP7_75t_R g1403 ( .A(n_1305), .Y(n_1403) );
OR2x2_ASAP7_75t_L g1305 ( .A(n_1306), .B(n_1321), .Y(n_1305) );
AOI22xp33_ASAP7_75t_L g1352 ( .A1(n_1306), .A2(n_1353), .B1(n_1356), .B2(n_1359), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1359 ( .A(n_1306), .B(n_1360), .Y(n_1359) );
OR2x2_ASAP7_75t_L g1395 ( .A(n_1306), .B(n_1322), .Y(n_1395) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1306), .Y(n_1406) );
INVx2_ASAP7_75t_L g1424 ( .A(n_1306), .Y(n_1424) );
OR2x2_ASAP7_75t_L g1438 ( .A(n_1306), .B(n_1362), .Y(n_1438) );
AND2x2_ASAP7_75t_L g1484 ( .A(n_1306), .B(n_1361), .Y(n_1484) );
AND2x2_ASAP7_75t_L g1493 ( .A(n_1306), .B(n_1362), .Y(n_1493) );
INVx2_ASAP7_75t_L g1306 ( .A(n_1307), .Y(n_1306) );
OR2x2_ASAP7_75t_L g1345 ( .A(n_1307), .B(n_1321), .Y(n_1345) );
NAND2xp5_ASAP7_75t_L g1307 ( .A(n_1308), .B(n_1315), .Y(n_1307) );
AND2x6_ASAP7_75t_L g1309 ( .A(n_1310), .B(n_1311), .Y(n_1309) );
AND2x2_ASAP7_75t_L g1313 ( .A(n_1310), .B(n_1314), .Y(n_1313) );
AND2x4_ASAP7_75t_L g1316 ( .A(n_1310), .B(n_1317), .Y(n_1316) );
AND2x6_ASAP7_75t_L g1319 ( .A(n_1310), .B(n_1320), .Y(n_1319) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1310), .B(n_1314), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1365 ( .A(n_1310), .B(n_1314), .Y(n_1365) );
NAND2xp5_ASAP7_75t_L g1374 ( .A(n_1310), .B(n_1317), .Y(n_1374) );
AND2x2_ASAP7_75t_L g1317 ( .A(n_1312), .B(n_1318), .Y(n_1317) );
INVx2_ASAP7_75t_L g1376 ( .A(n_1319), .Y(n_1376) );
HB1xp67_ASAP7_75t_L g1647 ( .A(n_1320), .Y(n_1647) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1321), .Y(n_1367) );
NOR2xp33_ASAP7_75t_L g1481 ( .A(n_1321), .B(n_1408), .Y(n_1481) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1322), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g1322 ( .A(n_1323), .B(n_1325), .Y(n_1322) );
OR2x2_ASAP7_75t_L g1326 ( .A(n_1327), .B(n_1331), .Y(n_1326) );
NOR2xp33_ASAP7_75t_L g1353 ( .A(n_1327), .B(n_1354), .Y(n_1353) );
NAND2xp5_ASAP7_75t_L g1388 ( .A(n_1327), .B(n_1389), .Y(n_1388) );
AND2x2_ASAP7_75t_L g1421 ( .A(n_1327), .B(n_1403), .Y(n_1421) );
CKINVDCx5p33_ASAP7_75t_R g1448 ( .A(n_1327), .Y(n_1448) );
AND2x2_ASAP7_75t_L g1455 ( .A(n_1327), .B(n_1357), .Y(n_1455) );
NAND2xp5_ASAP7_75t_L g1464 ( .A(n_1327), .B(n_1370), .Y(n_1464) );
AND2x2_ASAP7_75t_L g1497 ( .A(n_1327), .B(n_1367), .Y(n_1497) );
INVx4_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
O2A1O1Ixp33_ASAP7_75t_L g1379 ( .A1(n_1328), .A2(n_1380), .B(n_1382), .C(n_1385), .Y(n_1379) );
AND2x2_ASAP7_75t_L g1383 ( .A(n_1328), .B(n_1384), .Y(n_1383) );
INVx4_ASAP7_75t_L g1399 ( .A(n_1328), .Y(n_1399) );
NOR2xp33_ASAP7_75t_L g1401 ( .A(n_1328), .B(n_1402), .Y(n_1401) );
OR2x2_ASAP7_75t_L g1405 ( .A(n_1328), .B(n_1349), .Y(n_1405) );
NAND2xp5_ASAP7_75t_L g1407 ( .A(n_1328), .B(n_1397), .Y(n_1407) );
NAND2xp5_ASAP7_75t_SL g1412 ( .A(n_1328), .B(n_1349), .Y(n_1412) );
NOR2xp33_ASAP7_75t_L g1419 ( .A(n_1328), .B(n_1350), .Y(n_1419) );
NOR3xp33_ASAP7_75t_L g1441 ( .A(n_1328), .B(n_1438), .C(n_1442), .Y(n_1441) );
AND2x2_ASAP7_75t_L g1492 ( .A(n_1328), .B(n_1391), .Y(n_1492) );
AND2x4_ASAP7_75t_SL g1328 ( .A(n_1329), .B(n_1330), .Y(n_1328) );
NOR2xp33_ASAP7_75t_L g1467 ( .A(n_1331), .B(n_1430), .Y(n_1467) );
OR2x2_ASAP7_75t_L g1331 ( .A(n_1332), .B(n_1335), .Y(n_1331) );
OR2x2_ASAP7_75t_L g1390 ( .A(n_1332), .B(n_1337), .Y(n_1390) );
OR2x2_ASAP7_75t_L g1435 ( .A(n_1332), .B(n_1436), .Y(n_1435) );
AND2x2_ASAP7_75t_L g1443 ( .A(n_1332), .B(n_1384), .Y(n_1443) );
NAND2xp5_ASAP7_75t_L g1509 ( .A(n_1332), .B(n_1419), .Y(n_1509) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1333), .B(n_1334), .Y(n_1332) );
AND2x2_ASAP7_75t_L g1349 ( .A(n_1333), .B(n_1334), .Y(n_1349) );
OR2x2_ASAP7_75t_L g1459 ( .A(n_1335), .B(n_1348), .Y(n_1459) );
NAND2xp5_ASAP7_75t_L g1506 ( .A(n_1335), .B(n_1507), .Y(n_1506) );
NAND2xp5_ASAP7_75t_L g1335 ( .A(n_1336), .B(n_1340), .Y(n_1335) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
OR2x2_ASAP7_75t_L g1350 ( .A(n_1337), .B(n_1340), .Y(n_1350) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1337), .Y(n_1355) );
AND2x2_ASAP7_75t_L g1370 ( .A(n_1337), .B(n_1340), .Y(n_1370) );
AND2x2_ASAP7_75t_L g1384 ( .A(n_1337), .B(n_1358), .Y(n_1384) );
NAND2xp5_ASAP7_75t_L g1428 ( .A(n_1337), .B(n_1349), .Y(n_1428) );
AND2x2_ASAP7_75t_L g1337 ( .A(n_1338), .B(n_1339), .Y(n_1337) );
INVx2_ASAP7_75t_L g1358 ( .A(n_1340), .Y(n_1358) );
NAND2x1p5_ASAP7_75t_L g1340 ( .A(n_1341), .B(n_1342), .Y(n_1340) );
AOI211xp5_ASAP7_75t_L g1343 ( .A1(n_1344), .A2(n_1346), .B(n_1351), .C(n_1379), .Y(n_1343) );
NAND2xp5_ASAP7_75t_L g1447 ( .A(n_1344), .B(n_1448), .Y(n_1447) );
CKINVDCx5p33_ASAP7_75t_R g1344 ( .A(n_1345), .Y(n_1344) );
OR2x2_ASAP7_75t_L g1511 ( .A(n_1345), .B(n_1361), .Y(n_1511) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1347), .Y(n_1346) );
NOR2xp33_ASAP7_75t_L g1439 ( .A(n_1347), .B(n_1393), .Y(n_1439) );
OR2x2_ASAP7_75t_L g1347 ( .A(n_1348), .B(n_1350), .Y(n_1347) );
NOR2xp33_ASAP7_75t_L g1357 ( .A(n_1348), .B(n_1358), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1391 ( .A(n_1348), .B(n_1384), .Y(n_1391) );
AND2x2_ASAP7_75t_L g1445 ( .A(n_1348), .B(n_1410), .Y(n_1445) );
A2O1A1Ixp33_ASAP7_75t_L g1505 ( .A1(n_1348), .A2(n_1506), .B(n_1508), .C(n_1510), .Y(n_1505) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1349), .Y(n_1348) );
OR2x2_ASAP7_75t_L g1354 ( .A(n_1349), .B(n_1355), .Y(n_1354) );
AND2x2_ASAP7_75t_L g1369 ( .A(n_1349), .B(n_1370), .Y(n_1369) );
AND2x2_ASAP7_75t_L g1381 ( .A(n_1349), .B(n_1355), .Y(n_1381) );
OR2x2_ASAP7_75t_L g1402 ( .A(n_1349), .B(n_1358), .Y(n_1402) );
AND2x2_ASAP7_75t_L g1478 ( .A(n_1349), .B(n_1358), .Y(n_1478) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1350), .Y(n_1410) );
OR2x2_ASAP7_75t_L g1471 ( .A(n_1350), .B(n_1405), .Y(n_1471) );
OAI221xp5_ASAP7_75t_SL g1351 ( .A1(n_1352), .A2(n_1361), .B1(n_1366), .B2(n_1368), .C(n_1371), .Y(n_1351) );
HB1xp67_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1359), .Y(n_1452) );
OR2x2_ASAP7_75t_L g1385 ( .A(n_1360), .B(n_1361), .Y(n_1385) );
INVx2_ASAP7_75t_L g1397 ( .A(n_1360), .Y(n_1397) );
OAI221xp5_ASAP7_75t_L g1413 ( .A1(n_1360), .A2(n_1406), .B1(n_1414), .B2(n_1418), .C(n_1420), .Y(n_1413) );
AND2x2_ASAP7_75t_L g1429 ( .A(n_1360), .B(n_1430), .Y(n_1429) );
AND2x2_ASAP7_75t_L g1457 ( .A(n_1360), .B(n_1399), .Y(n_1457) );
A2O1A1Ixp33_ASAP7_75t_L g1485 ( .A1(n_1360), .A2(n_1486), .B(n_1492), .C(n_1493), .Y(n_1485) );
OR2x2_ASAP7_75t_L g1366 ( .A(n_1361), .B(n_1367), .Y(n_1366) );
A2O1A1Ixp33_ASAP7_75t_L g1400 ( .A1(n_1361), .A2(n_1401), .B(n_1403), .C(n_1404), .Y(n_1400) );
CKINVDCx14_ASAP7_75t_R g1462 ( .A(n_1361), .Y(n_1462) );
INVx3_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1362), .Y(n_1394) );
AOI221xp5_ASAP7_75t_L g1468 ( .A1(n_1362), .A2(n_1397), .B1(n_1469), .B2(n_1472), .C(n_1479), .Y(n_1468) );
AND2x2_ASAP7_75t_L g1474 ( .A(n_1362), .B(n_1406), .Y(n_1474) );
OAI21xp33_ASAP7_75t_L g1479 ( .A1(n_1362), .A2(n_1480), .B(n_1482), .Y(n_1479) );
AND2x2_ASAP7_75t_L g1362 ( .A(n_1363), .B(n_1364), .Y(n_1362) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1367), .Y(n_1416) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
NAND2x1_ASAP7_75t_L g1398 ( .A(n_1369), .B(n_1399), .Y(n_1398) );
OAI21xp33_ASAP7_75t_L g1482 ( .A1(n_1369), .A2(n_1483), .B(n_1484), .Y(n_1482) );
OAI321xp33_ASAP7_75t_L g1404 ( .A1(n_1370), .A2(n_1380), .A3(n_1405), .B1(n_1406), .B2(n_1407), .C(n_1408), .Y(n_1404) );
INVx1_ASAP7_75t_L g1436 ( .A(n_1370), .Y(n_1436) );
OAI21xp5_ASAP7_75t_L g1444 ( .A1(n_1370), .A2(n_1445), .B(n_1446), .Y(n_1444) );
AND2x2_ASAP7_75t_L g1476 ( .A(n_1370), .B(n_1411), .Y(n_1476) );
AOI211xp5_ASAP7_75t_L g1453 ( .A1(n_1371), .A2(n_1454), .B(n_1455), .C(n_1456), .Y(n_1453) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
NAND2xp5_ASAP7_75t_L g1461 ( .A(n_1372), .B(n_1462), .Y(n_1461) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1373), .Y(n_1372) );
OAI221xp5_ASAP7_75t_L g1373 ( .A1(n_1374), .A2(n_1375), .B1(n_1376), .B2(n_1377), .C(n_1378), .Y(n_1373) );
CKINVDCx20_ASAP7_75t_R g1513 ( .A(n_1376), .Y(n_1513) );
NAND2xp5_ASAP7_75t_SL g1434 ( .A(n_1380), .B(n_1435), .Y(n_1434) );
O2A1O1Ixp33_ASAP7_75t_L g1449 ( .A1(n_1380), .A2(n_1450), .B(n_1453), .C(n_1460), .Y(n_1449) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1381), .Y(n_1380) );
NAND2xp5_ASAP7_75t_L g1420 ( .A(n_1381), .B(n_1421), .Y(n_1420) );
INVx1_ASAP7_75t_L g1382 ( .A(n_1383), .Y(n_1382) );
INVx1_ASAP7_75t_L g1507 ( .A(n_1384), .Y(n_1507) );
OAI322xp33_ASAP7_75t_L g1463 ( .A1(n_1385), .A2(n_1390), .A3(n_1394), .B1(n_1403), .B2(n_1464), .C1(n_1465), .C2(n_1466), .Y(n_1463) );
OAI21xp33_ASAP7_75t_L g1386 ( .A1(n_1387), .A2(n_1391), .B(n_1392), .Y(n_1386) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
INVxp67_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
NOR2xp33_ASAP7_75t_L g1417 ( .A(n_1390), .B(n_1399), .Y(n_1417) );
NAND2xp5_ASAP7_75t_L g1432 ( .A(n_1391), .B(n_1403), .Y(n_1432) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1391), .Y(n_1502) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
OR2x2_ASAP7_75t_L g1393 ( .A(n_1394), .B(n_1395), .Y(n_1393) );
NAND2xp5_ASAP7_75t_L g1496 ( .A(n_1394), .B(n_1497), .Y(n_1496) );
OAI21xp33_ASAP7_75t_L g1396 ( .A1(n_1397), .A2(n_1398), .B(n_1400), .Y(n_1396) );
OR2x2_ASAP7_75t_L g1465 ( .A(n_1397), .B(n_1438), .Y(n_1465) );
CKINVDCx5p33_ASAP7_75t_R g1430 ( .A(n_1399), .Y(n_1430) );
AND2x2_ASAP7_75t_L g1504 ( .A(n_1403), .B(n_1448), .Y(n_1504) );
NOR2xp33_ASAP7_75t_L g1425 ( .A(n_1406), .B(n_1426), .Y(n_1425) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1406), .Y(n_1454) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
AOI211xp5_ASAP7_75t_L g1423 ( .A1(n_1409), .A2(n_1424), .B(n_1425), .C(n_1431), .Y(n_1423) );
NAND2xp5_ASAP7_75t_L g1501 ( .A(n_1409), .B(n_1416), .Y(n_1501) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_1410), .B(n_1411), .Y(n_1409) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1412), .Y(n_1411) );
INVxp67_ASAP7_75t_L g1414 ( .A(n_1415), .Y(n_1414) );
AND2x2_ASAP7_75t_L g1415 ( .A(n_1416), .B(n_1417), .Y(n_1415) );
AND2x2_ASAP7_75t_L g1469 ( .A(n_1416), .B(n_1470), .Y(n_1469) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1419), .Y(n_1418) );
O2A1O1Ixp33_ASAP7_75t_L g1494 ( .A1(n_1421), .A2(n_1495), .B(n_1498), .C(n_1500), .Y(n_1494) );
NAND4xp25_ASAP7_75t_L g1422 ( .A(n_1423), .B(n_1433), .C(n_1440), .D(n_1444), .Y(n_1422) );
INVxp33_ASAP7_75t_L g1483 ( .A(n_1426), .Y(n_1483) );
NAND2xp5_ASAP7_75t_L g1426 ( .A(n_1427), .B(n_1429), .Y(n_1426) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
OR2x2_ASAP7_75t_L g1489 ( .A(n_1428), .B(n_1448), .Y(n_1489) );
AOI31xp33_ASAP7_75t_L g1433 ( .A1(n_1430), .A2(n_1434), .A3(n_1437), .B(n_1439), .Y(n_1433) );
NOR2xp33_ASAP7_75t_L g1451 ( .A(n_1430), .B(n_1452), .Y(n_1451) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1432), .Y(n_1431) );
CKINVDCx14_ASAP7_75t_R g1437 ( .A(n_1438), .Y(n_1437) );
OAI22xp5_ASAP7_75t_L g1472 ( .A1(n_1438), .A2(n_1473), .B1(n_1475), .B2(n_1477), .Y(n_1472) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1441), .Y(n_1440) );
AND2x2_ASAP7_75t_L g1499 ( .A(n_1442), .B(n_1491), .Y(n_1499) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1443), .Y(n_1442) );
INVx1_ASAP7_75t_L g1491 ( .A(n_1445), .Y(n_1491) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1447), .Y(n_1446) );
INVxp67_ASAP7_75t_SL g1450 ( .A(n_1451), .Y(n_1450) );
OAI22xp5_ASAP7_75t_L g1500 ( .A1(n_1454), .A2(n_1501), .B1(n_1502), .B2(n_1503), .Y(n_1500) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1455), .Y(n_1490) );
AND2x2_ASAP7_75t_L g1456 ( .A(n_1457), .B(n_1458), .Y(n_1456) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
INVx1_ASAP7_75t_L g1460 ( .A(n_1461), .Y(n_1460) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1467), .Y(n_1466) );
INVx1_ASAP7_75t_L g1470 ( .A(n_1471), .Y(n_1470) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1476), .Y(n_1475) );
CKINVDCx14_ASAP7_75t_R g1477 ( .A(n_1478), .Y(n_1477) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1481), .Y(n_1480) );
NAND2xp5_ASAP7_75t_L g1486 ( .A(n_1487), .B(n_1491), .Y(n_1486) );
INVxp67_ASAP7_75t_SL g1487 ( .A(n_1488), .Y(n_1487) );
NAND2xp5_ASAP7_75t_L g1488 ( .A(n_1489), .B(n_1490), .Y(n_1488) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
INVxp67_ASAP7_75t_L g1498 ( .A(n_1499), .Y(n_1498) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1504), .Y(n_1503) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1509), .Y(n_1508) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1511), .Y(n_1510) );
CKINVDCx20_ASAP7_75t_R g1512 ( .A(n_1513), .Y(n_1512) );
HB1xp67_ASAP7_75t_L g1514 ( .A(n_1515), .Y(n_1514) );
XNOR2x1_ASAP7_75t_L g1515 ( .A(n_1516), .B(n_1517), .Y(n_1515) );
OR2x2_ASAP7_75t_L g1517 ( .A(n_1518), .B(n_1565), .Y(n_1517) );
A2O1A1Ixp33_ASAP7_75t_L g1518 ( .A1(n_1519), .A2(n_1544), .B(n_1558), .C(n_1560), .Y(n_1518) );
NOR3xp33_ASAP7_75t_L g1519 ( .A(n_1520), .B(n_1525), .C(n_1532), .Y(n_1519) );
CKINVDCx5p33_ASAP7_75t_R g1520 ( .A(n_1521), .Y(n_1520) );
INVx1_ASAP7_75t_L g1522 ( .A(n_1523), .Y(n_1522) );
INVx3_ASAP7_75t_L g1540 ( .A(n_1541), .Y(n_1540) );
HB1xp67_ASAP7_75t_L g1552 ( .A(n_1542), .Y(n_1552) );
INVx1_ASAP7_75t_L g1542 ( .A(n_1543), .Y(n_1542) );
AOI221xp5_ASAP7_75t_L g1544 ( .A1(n_1545), .A2(n_1547), .B1(n_1548), .B2(n_1551), .C(n_1553), .Y(n_1544) );
INVx2_ASAP7_75t_L g1545 ( .A(n_1546), .Y(n_1545) );
AOI332xp33_ASAP7_75t_L g1569 ( .A1(n_1547), .A2(n_1570), .A3(n_1573), .B1(n_1575), .B2(n_1576), .B3(n_1577), .C1(n_1579), .C2(n_1581), .Y(n_1569) );
NAND2xp5_ASAP7_75t_L g1560 ( .A(n_1550), .B(n_1561), .Y(n_1560) );
BUFx2_ASAP7_75t_L g1551 ( .A(n_1552), .Y(n_1551) );
INVx4_ASAP7_75t_L g1554 ( .A(n_1555), .Y(n_1554) );
INVx2_ASAP7_75t_L g1556 ( .A(n_1557), .Y(n_1556) );
HB1xp67_ASAP7_75t_L g1558 ( .A(n_1559), .Y(n_1558) );
AND2x4_ASAP7_75t_L g1561 ( .A(n_1562), .B(n_1563), .Y(n_1561) );
AND2x4_ASAP7_75t_L g1567 ( .A(n_1562), .B(n_1568), .Y(n_1567) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1571), .Y(n_1570) );
INVx1_ASAP7_75t_L g1573 ( .A(n_1574), .Y(n_1573) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1578), .Y(n_1577) );
INVx2_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
NOR3xp33_ASAP7_75t_L g1582 ( .A(n_1583), .B(n_1589), .C(n_1599), .Y(n_1582) );
INVx2_ASAP7_75t_L g1590 ( .A(n_1591), .Y(n_1590) );
INVx2_ASAP7_75t_SL g1591 ( .A(n_1592), .Y(n_1591) );
NAND2x2_ASAP7_75t_L g1592 ( .A(n_1593), .B(n_1595), .Y(n_1592) );
INVx1_ASAP7_75t_L g1601 ( .A(n_1593), .Y(n_1601) );
INVx2_ASAP7_75t_L g1593 ( .A(n_1594), .Y(n_1593) );
INVx2_ASAP7_75t_SL g1595 ( .A(n_1596), .Y(n_1595) );
CKINVDCx5p33_ASAP7_75t_R g1599 ( .A(n_1600), .Y(n_1599) );
INVx1_ASAP7_75t_L g1602 ( .A(n_1603), .Y(n_1602) );
BUFx3_ASAP7_75t_L g1603 ( .A(n_1604), .Y(n_1603) );
BUFx3_ASAP7_75t_L g1607 ( .A(n_1608), .Y(n_1607) );
INVxp33_ASAP7_75t_SL g1609 ( .A(n_1610), .Y(n_1609) );
HB1xp67_ASAP7_75t_L g1611 ( .A(n_1612), .Y(n_1611) );
AND3x1_ASAP7_75t_L g1612 ( .A(n_1613), .B(n_1632), .C(n_1639), .Y(n_1612) );
NOR2xp33_ASAP7_75t_L g1613 ( .A(n_1614), .B(n_1627), .Y(n_1613) );
HB1xp67_ASAP7_75t_L g1645 ( .A(n_1646), .Y(n_1645) );
OAI21xp5_ASAP7_75t_L g1646 ( .A1(n_1647), .A2(n_1648), .B(n_1649), .Y(n_1646) );
INVx1_ASAP7_75t_L g1649 ( .A(n_1650), .Y(n_1649) );
endmodule