module fake_jpeg_13467_n_188 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_188);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_11),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_25),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_27),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_26),
.Y(n_64)
);

INVx11_ASAP7_75t_SL g65 ( 
.A(n_23),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_44),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_10),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_0),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_88),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_51),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_84),
.B(n_71),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_0),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_90),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_1),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_78),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_93),
.B(n_96),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_59),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_67),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_98),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_70),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_73),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_100),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_64),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_58),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_85),
.A2(n_71),
.B1(n_58),
.B2(n_52),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_52),
.B1(n_56),
.B2(n_76),
.Y(n_112)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_105),
.Y(n_108)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_111),
.Y(n_132)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_120),
.Y(n_136)
);

OA21x2_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_56),
.B(n_79),
.Y(n_115)
);

AO22x1_ASAP7_75t_L g149 ( 
.A1(n_115),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_149)
);

AOI22x1_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_80),
.B1(n_65),
.B2(n_53),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_2),
.B(n_3),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_92),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_117),
.B(n_118),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_62),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_102),
.B(n_72),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_119),
.Y(n_147)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_122),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_101),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_124),
.Y(n_135)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_2),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_60),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_126),
.B(n_8),
.Y(n_150)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_46),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_113),
.A2(n_80),
.B1(n_69),
.B2(n_68),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_113),
.A2(n_66),
.B1(n_65),
.B2(n_72),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_116),
.A2(n_74),
.B1(n_63),
.B2(n_75),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_119),
.A2(n_74),
.B(n_75),
.C(n_47),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_75),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_15),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_106),
.B(n_1),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_143),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_138),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_139),
.Y(n_157)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_115),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_146),
.B1(n_14),
.B2(n_15),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_110),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_115),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_149),
.A2(n_122),
.B(n_124),
.Y(n_152)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_127),
.B(n_119),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_153),
.B(n_164),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_154),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_148),
.A2(n_111),
.B1(n_32),
.B2(n_36),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_147),
.A2(n_13),
.B(n_14),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_160),
.Y(n_173)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_163),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_40),
.Y(n_163)
);

OAI32xp33_ASAP7_75t_L g164 ( 
.A1(n_132),
.A2(n_144),
.A3(n_149),
.B1(n_128),
.B2(n_135),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_165),
.A2(n_167),
.B1(n_146),
.B2(n_141),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_148),
.A2(n_16),
.B1(n_17),
.B2(n_20),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_166),
.A2(n_137),
.B1(n_136),
.B2(n_145),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_130),
.A2(n_16),
.B1(n_17),
.B2(n_24),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_159),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_168),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_170),
.A2(n_174),
.B1(n_163),
.B2(n_165),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_171),
.A2(n_155),
.B1(n_158),
.B2(n_153),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_161),
.A2(n_129),
.B1(n_131),
.B2(n_42),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_179),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_L g178 ( 
.A1(n_174),
.A2(n_161),
.B1(n_162),
.B2(n_157),
.Y(n_178)
);

OAI321xp33_ASAP7_75t_L g180 ( 
.A1(n_178),
.A2(n_172),
.A3(n_171),
.B1(n_175),
.B2(n_169),
.C(n_173),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_169),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_182),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_177),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_184),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_181),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_177),
.C(n_170),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_39),
.C(n_41),
.Y(n_188)
);


endmodule