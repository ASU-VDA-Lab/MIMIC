module fake_jpeg_21474_n_136 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_10),
.B(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_25),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_30),
.Y(n_44)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_15),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_15),
.B1(n_22),
.B2(n_20),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_42),
.B1(n_34),
.B2(n_2),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_21),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_31),
.A2(n_14),
.B1(n_22),
.B2(n_20),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_25),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_49),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_25),
.B(n_23),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_48),
.A2(n_13),
.B1(n_27),
.B2(n_17),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_25),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_27),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_19),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_51),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_17),
.B1(n_14),
.B2(n_13),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_41),
.B1(n_46),
.B2(n_39),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_54),
.B(n_58),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_19),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_56),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_26),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_59),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_34),
.Y(n_58)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_41),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_64),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

CKINVDCx11_ASAP7_75t_R g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_72),
.Y(n_82)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_37),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

NOR4xp25_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_54),
.C(n_58),
.D(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_40),
.Y(n_76)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_79),
.B1(n_39),
.B2(n_2),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_46),
.B(n_39),
.C(n_4),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_71),
.B(n_72),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_58),
.B(n_53),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_74),
.A2(n_61),
.B1(n_65),
.B2(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_76),
.B(n_10),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_89),
.B(n_91),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_65),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_67),
.Y(n_99)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_78),
.B(n_73),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_101),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_100),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_90),
.B(n_78),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_88),
.A2(n_69),
.B1(n_79),
.B2(n_77),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_79),
.B1(n_73),
.B2(n_92),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_104),
.B(n_82),
.Y(n_110)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_95),
.Y(n_106)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_99),
.C(n_98),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_111),
.Y(n_118)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_109),
.A2(n_60),
.B1(n_2),
.B2(n_4),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_8),
.B(n_81),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_86),
.C(n_85),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);

OAI321xp33_ASAP7_75t_L g117 ( 
.A1(n_113),
.A2(n_101),
.A3(n_94),
.B1(n_91),
.B2(n_71),
.C(n_81),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_117),
.A2(n_108),
.B(n_8),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_119),
.A2(n_120),
.B(n_0),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_107),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_123),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_114),
.A2(n_112),
.B(n_111),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_125),
.B(n_114),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_108),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_127),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_121),
.A2(n_115),
.B1(n_6),
.B2(n_7),
.Y(n_127)
);

BUFx24_ASAP7_75t_SL g130 ( 
.A(n_128),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_130),
.B(n_7),
.Y(n_134)
);

AO21x1_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_5),
.B(n_6),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_132),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_133),
.B(n_131),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_7),
.Y(n_136)
);


endmodule