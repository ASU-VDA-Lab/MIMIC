module fake_jpeg_8680_n_46 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_46);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_46;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_43;
wire n_37;
wire n_32;

INVx4_ASAP7_75t_SL g20 ( 
.A(n_18),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_17),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx6p67_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_25),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_28),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_1),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_1),
.C(n_3),
.Y(n_39)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_32),
.B(n_33),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_26),
.A2(n_8),
.B(n_2),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_39),
.C(n_13),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_42),
.A2(n_43),
.B(n_41),
.Y(n_44)
);

AOI322xp5_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_35),
.A3(n_37),
.B1(n_36),
.B2(n_34),
.C1(n_14),
.C2(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);


endmodule