module fake_netlist_5_2237_n_1739 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1739);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1739;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_152),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_31),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_85),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_111),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_87),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_17),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_43),
.Y(n_166)
);

BUFx10_ASAP7_75t_L g167 ( 
.A(n_65),
.Y(n_167)
);

BUFx10_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_47),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_12),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_139),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_45),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_39),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_19),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_17),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_53),
.Y(n_176)
);

CKINVDCx11_ASAP7_75t_R g177 ( 
.A(n_116),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_131),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_14),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_34),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_117),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_67),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_134),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_140),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_144),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_12),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_81),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_76),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_11),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_31),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_105),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_16),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_63),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_27),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_92),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_39),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_41),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_114),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_54),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_127),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_79),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_159),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_30),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_60),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_136),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_142),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_78),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_75),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_109),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_28),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_56),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_2),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_20),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_69),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_2),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_148),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_83),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_25),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_129),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_5),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_104),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_120),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_37),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_90),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_58),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_33),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_138),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_115),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_95),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_53),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_119),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_74),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_112),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_1),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_145),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_89),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_86),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_64),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_8),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_99),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_128),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_121),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_108),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_106),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_21),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_110),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_25),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_3),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_61),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_149),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_77),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_10),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_37),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_33),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_62),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_100),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_66),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_153),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_57),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_71),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_154),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_141),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_16),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_124),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_5),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_1),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_47),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_82),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_20),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_68),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_9),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_43),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_36),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_24),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_34),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_19),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_70),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_6),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_103),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_133),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_158),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_101),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_11),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_41),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_29),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_135),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_21),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_30),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_15),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_51),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_51),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_151),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_49),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_8),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_10),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_29),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_49),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_14),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_93),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_27),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_22),
.Y(n_301)
);

INVxp33_ASAP7_75t_L g302 ( 
.A(n_36),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_150),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_157),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_18),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_122),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_125),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_9),
.Y(n_308)
);

BUFx2_ASAP7_75t_SL g309 ( 
.A(n_6),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_24),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_22),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_73),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_97),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_126),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_13),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_192),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_192),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_192),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_180),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_206),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_183),
.Y(n_321)
);

INVxp33_ASAP7_75t_SL g322 ( 
.A(n_161),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_177),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_192),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_192),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_269),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_207),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_250),
.Y(n_328)
);

INVxp33_ASAP7_75t_SL g329 ( 
.A(n_161),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_259),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_269),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_286),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_298),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_246),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_269),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_269),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_269),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_163),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_199),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_202),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_218),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_204),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_219),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_218),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_205),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_209),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_266),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_226),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_266),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_297),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_288),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_297),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_226),
.Y(n_353)
);

INVxp33_ASAP7_75t_L g354 ( 
.A(n_302),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_245),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_219),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_214),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_245),
.Y(n_358)
);

INVxp33_ASAP7_75t_SL g359 ( 
.A(n_165),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_290),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_290),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_221),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_224),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_170),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_225),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_225),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_165),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_167),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_306),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_315),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_173),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_167),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_176),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_166),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_228),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_190),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_223),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_229),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_252),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_238),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_240),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_166),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_242),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_243),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_267),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_271),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_273),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_244),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_274),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_275),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_278),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_283),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_339),
.B(n_208),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_316),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_316),
.Y(n_395)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_334),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_317),
.B(n_306),
.Y(n_397)
);

AND2x6_ASAP7_75t_L g398 ( 
.A(n_334),
.B(n_246),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_334),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_340),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_317),
.Y(n_401)
);

AND2x4_ASAP7_75t_L g402 ( 
.A(n_318),
.B(n_164),
.Y(n_402)
);

AND2x4_ASAP7_75t_L g403 ( 
.A(n_318),
.B(n_164),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_342),
.B(n_237),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_324),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_324),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_325),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_325),
.B(n_237),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_345),
.B(n_255),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_357),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_326),
.B(n_331),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_374),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_326),
.Y(n_413)
);

NAND2xp33_ASAP7_75t_R g414 ( 
.A(n_322),
.B(n_160),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_362),
.B(n_255),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_331),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_335),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_335),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_363),
.B(n_261),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_336),
.B(n_261),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_336),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_337),
.Y(n_422)
);

NOR2x1_ASAP7_75t_L g423 ( 
.A(n_337),
.B(n_181),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_343),
.B(n_182),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_379),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_379),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_375),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_364),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_364),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_378),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_370),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_341),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_380),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_320),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_356),
.B(n_212),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_327),
.A2(n_294),
.B1(n_272),
.B2(n_296),
.Y(n_436)
);

NAND2xp33_ASAP7_75t_L g437 ( 
.A(n_383),
.B(n_169),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_341),
.Y(n_438)
);

CKINVDCx8_ASAP7_75t_R g439 ( 
.A(n_368),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_370),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_371),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_344),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_366),
.B(n_212),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_384),
.B(n_236),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_371),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_373),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_328),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_373),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_344),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_368),
.B(n_372),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_376),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_369),
.B(n_284),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_376),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_347),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_377),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_347),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_349),
.Y(n_457)
);

OA21x2_ASAP7_75t_L g458 ( 
.A1(n_349),
.A2(n_187),
.B(n_185),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_377),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_372),
.B(n_167),
.Y(n_460)
);

INVx4_ASAP7_75t_L g461 ( 
.A(n_388),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_350),
.Y(n_462)
);

AND2x6_ASAP7_75t_L g463 ( 
.A(n_343),
.B(n_246),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_354),
.B(n_168),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_338),
.B(n_188),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_397),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_394),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_397),
.B(n_343),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_411),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_394),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_393),
.B(n_319),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_399),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_412),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_399),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_395),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_395),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_444),
.B(n_321),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_435),
.B(n_365),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_407),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_399),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_404),
.B(n_321),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_409),
.B(n_365),
.Y(n_482)
);

AOI21x1_ASAP7_75t_L g483 ( 
.A1(n_405),
.A2(n_195),
.B(n_191),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_401),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_399),
.Y(n_485)
);

NOR2x1p5_ASAP7_75t_L g486 ( 
.A(n_461),
.B(n_323),
.Y(n_486)
);

INVx8_ASAP7_75t_L g487 ( 
.A(n_463),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_415),
.B(n_365),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_411),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_436),
.B(n_330),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_401),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_419),
.B(n_329),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_411),
.Y(n_493)
);

OAI21xp33_ASAP7_75t_SL g494 ( 
.A1(n_435),
.A2(n_284),
.B(n_353),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_405),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_417),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_417),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_443),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_422),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_406),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_443),
.B(n_452),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_434),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_399),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_437),
.A2(n_308),
.B1(n_189),
.B2(n_186),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_422),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_406),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_399),
.Y(n_507)
);

NOR2x1p5_ASAP7_75t_L g508 ( 
.A(n_461),
.B(n_169),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_413),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_452),
.B(n_262),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_461),
.B(n_359),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_424),
.B(n_353),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_438),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_438),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_413),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_461),
.B(n_346),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_396),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_400),
.B(n_381),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_438),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_462),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_424),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_462),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_462),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_416),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_410),
.B(n_332),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_416),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_396),
.Y(n_527)
);

OAI22xp33_ASAP7_75t_L g528 ( 
.A1(n_460),
.A2(n_213),
.B1(n_196),
.B2(n_333),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_462),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_462),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_436),
.B(n_447),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_424),
.Y(n_532)
);

INVx1_ASAP7_75t_SL g533 ( 
.A(n_464),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_414),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_462),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_418),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_465),
.A2(n_351),
.B1(n_254),
.B2(n_253),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_418),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_396),
.Y(n_539)
);

OR2x6_ASAP7_75t_L g540 ( 
.A(n_424),
.B(n_309),
.Y(n_540)
);

NAND3xp33_ASAP7_75t_L g541 ( 
.A(n_450),
.B(n_382),
.C(n_367),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_421),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_427),
.B(n_348),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_430),
.B(n_348),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_423),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_421),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_407),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_402),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_407),
.Y(n_549)
);

BUFx10_ASAP7_75t_L g550 ( 
.A(n_433),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_428),
.B(n_355),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_407),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_402),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_407),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_402),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_407),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_396),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_402),
.Y(n_558)
);

BUFx4f_ASAP7_75t_L g559 ( 
.A(n_458),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_403),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_458),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_458),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_403),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_403),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_403),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_432),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_428),
.B(n_355),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_408),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_458),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_432),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_429),
.B(n_358),
.Y(n_571)
);

INVx8_ASAP7_75t_L g572 ( 
.A(n_463),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_408),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_439),
.B(n_168),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_442),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_408),
.A2(n_420),
.B1(n_463),
.B2(n_423),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_408),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_420),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_420),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_420),
.Y(n_580)
);

AOI21x1_ASAP7_75t_L g581 ( 
.A1(n_429),
.A2(n_201),
.B(n_200),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_431),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_431),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_439),
.B(n_168),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_442),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_440),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_440),
.A2(n_265),
.B1(n_263),
.B2(n_276),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_449),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_441),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_449),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_441),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_454),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_445),
.Y(n_593)
);

NAND2x1p5_ASAP7_75t_L g594 ( 
.A(n_445),
.B(n_211),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_454),
.Y(n_595)
);

INVx5_ASAP7_75t_L g596 ( 
.A(n_398),
.Y(n_596)
);

NAND3xp33_ASAP7_75t_L g597 ( 
.A(n_446),
.B(n_358),
.C(n_360),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_446),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_448),
.B(n_241),
.Y(n_599)
);

BUFx6f_ASAP7_75t_SL g600 ( 
.A(n_463),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_448),
.B(n_360),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_456),
.Y(n_602)
);

AO21x2_ASAP7_75t_L g603 ( 
.A1(n_451),
.A2(n_222),
.B(n_313),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_456),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_451),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_457),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_453),
.Y(n_607)
);

OAI22xp33_ASAP7_75t_SL g608 ( 
.A1(n_453),
.A2(n_301),
.B1(n_291),
.B2(n_293),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_457),
.Y(n_609)
);

AO22x2_ASAP7_75t_L g610 ( 
.A1(n_490),
.A2(n_232),
.B1(n_235),
.B2(n_249),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_564),
.Y(n_611)
);

BUFx5_ASAP7_75t_L g612 ( 
.A(n_466),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_466),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_559),
.A2(n_426),
.B(n_425),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_498),
.A2(n_279),
.B1(n_268),
.B2(n_304),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_585),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_603),
.A2(n_463),
.B1(n_292),
.B2(n_246),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_498),
.B(n_492),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_545),
.B(n_463),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_585),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_545),
.B(n_463),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_564),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_501),
.B(n_426),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_564),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_469),
.Y(n_625)
);

OR2x6_ASAP7_75t_L g626 ( 
.A(n_540),
.B(n_361),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_469),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_534),
.B(n_160),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_482),
.B(n_162),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_488),
.B(n_216),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_585),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_588),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_478),
.B(n_361),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_468),
.B(n_455),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_481),
.B(n_162),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_510),
.B(n_171),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_478),
.B(n_455),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_528),
.B(n_171),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_588),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_588),
.Y(n_640)
);

A2O1A1Ixp33_ASAP7_75t_L g641 ( 
.A1(n_559),
.A2(n_217),
.B(n_312),
.C(n_258),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_517),
.B(n_227),
.Y(n_642)
);

INVxp67_ASAP7_75t_SL g643 ( 
.A(n_517),
.Y(n_643)
);

AO221x1_ASAP7_75t_L g644 ( 
.A1(n_587),
.A2(n_292),
.B1(n_246),
.B2(n_256),
.C(n_459),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_559),
.B(n_292),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_517),
.B(n_459),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_517),
.B(n_425),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_527),
.B(n_251),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_473),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_590),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_521),
.A2(n_264),
.B1(n_270),
.B2(n_299),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_473),
.B(n_288),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_527),
.B(n_257),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_590),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_543),
.B(n_288),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_589),
.B(n_178),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_468),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_489),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_468),
.A2(n_260),
.B1(n_178),
.B2(n_299),
.Y(n_659)
);

OAI221xp5_ASAP7_75t_L g660 ( 
.A1(n_494),
.A2(n_385),
.B1(n_392),
.B2(n_391),
.C(n_390),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_544),
.B(n_184),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_590),
.Y(n_662)
);

NOR2xp67_ASAP7_75t_SL g663 ( 
.A(n_596),
.B(n_292),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_592),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_527),
.B(n_292),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_589),
.B(n_184),
.Y(n_666)
);

BUFx6f_ASAP7_75t_SL g667 ( 
.A(n_550),
.Y(n_667)
);

NAND2xp33_ASAP7_75t_L g668 ( 
.A(n_521),
.B(n_193),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_592),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_SL g670 ( 
.A1(n_533),
.A2(n_241),
.B1(n_277),
.B2(n_276),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_477),
.B(n_193),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_527),
.B(n_539),
.Y(n_672)
);

BUFx6f_ASAP7_75t_SL g673 ( 
.A(n_550),
.Y(n_673)
);

OR2x6_ASAP7_75t_L g674 ( 
.A(n_540),
.B(n_385),
.Y(n_674)
);

NAND2xp33_ASAP7_75t_SL g675 ( 
.A(n_508),
.B(n_574),
.Y(n_675)
);

OAI22xp33_ASAP7_75t_L g676 ( 
.A1(n_504),
.A2(n_179),
.B1(n_194),
.B2(n_175),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_539),
.B(n_198),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_592),
.Y(n_678)
);

NAND2xp33_ASAP7_75t_L g679 ( 
.A(n_532),
.B(n_231),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_539),
.B(n_233),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_593),
.B(n_386),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_598),
.B(n_532),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_557),
.A2(n_386),
.B(n_392),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_471),
.B(n_233),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_598),
.B(n_468),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_540),
.A2(n_264),
.B1(n_270),
.B2(n_280),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_595),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_493),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_567),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_493),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_598),
.B(n_280),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_R g692 ( 
.A(n_550),
.B(n_281),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_466),
.B(n_282),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_603),
.A2(n_265),
.B1(n_174),
.B2(n_175),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_573),
.B(n_282),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_582),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_541),
.B(n_303),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_504),
.B(n_303),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_511),
.B(n_307),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_582),
.B(n_307),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_595),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_583),
.Y(n_702)
);

O2A1O1Ixp5_ASAP7_75t_L g703 ( 
.A1(n_561),
.A2(n_391),
.B(n_390),
.C(n_389),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_583),
.B(n_314),
.Y(n_704)
);

INVx8_ASAP7_75t_L g705 ( 
.A(n_540),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_573),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_567),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_573),
.B(n_314),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_595),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_512),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_602),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_551),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_586),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_512),
.B(n_550),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_602),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_508),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_591),
.B(n_203),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_602),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_605),
.B(n_398),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_607),
.Y(n_720)
);

NOR3xp33_ASAP7_75t_L g721 ( 
.A(n_537),
.B(n_389),
.C(n_387),
.Y(n_721)
);

HB1xp67_ASAP7_75t_L g722 ( 
.A(n_540),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_604),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_584),
.B(n_210),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_548),
.A2(n_398),
.B1(n_241),
.B2(n_277),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_548),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_571),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_573),
.B(n_398),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_578),
.B(n_398),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_604),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_578),
.B(n_277),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_578),
.B(n_215),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_494),
.B(n_220),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_553),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_495),
.B(n_230),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_495),
.B(n_234),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_553),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_500),
.B(n_506),
.Y(n_738)
);

AND2x6_ASAP7_75t_SL g739 ( 
.A(n_490),
.B(n_350),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_555),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_604),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_578),
.B(n_398),
.Y(n_742)
);

INVxp33_ASAP7_75t_L g743 ( 
.A(n_531),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_555),
.B(n_398),
.Y(n_744)
);

NOR2xp67_ASAP7_75t_L g745 ( 
.A(n_516),
.B(n_102),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_599),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_576),
.B(n_239),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_606),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_558),
.B(n_247),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_560),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_560),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_563),
.A2(n_248),
.B1(n_311),
.B2(n_310),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_563),
.B(n_352),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_565),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_565),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_606),
.Y(n_756)
);

OAI22xp33_ASAP7_75t_L g757 ( 
.A1(n_594),
.A2(n_287),
.B1(n_311),
.B2(n_310),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_568),
.B(n_263),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_568),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_577),
.B(n_352),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_577),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_579),
.B(n_580),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_579),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_580),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_606),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_500),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_566),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_506),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_509),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_509),
.B(n_305),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_657),
.Y(n_771)
);

INVx1_ASAP7_75t_SL g772 ( 
.A(n_649),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_613),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_657),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_635),
.A2(n_518),
.B1(n_515),
.B2(n_536),
.Y(n_775)
);

BUFx2_ASAP7_75t_L g776 ( 
.A(n_714),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_625),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_710),
.B(n_486),
.Y(n_778)
);

INVxp67_ASAP7_75t_L g779 ( 
.A(n_656),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_612),
.B(n_561),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_616),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_627),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_643),
.B(n_515),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_655),
.B(n_502),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_658),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_612),
.B(n_561),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_613),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_712),
.B(n_524),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_727),
.B(n_524),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_738),
.B(n_526),
.Y(n_790)
);

NAND2x1p5_ASAP7_75t_L g791 ( 
.A(n_613),
.B(n_706),
.Y(n_791)
);

CKINVDCx20_ASAP7_75t_R g792 ( 
.A(n_692),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_738),
.B(n_635),
.Y(n_793)
);

NAND2x2_ASAP7_75t_L g794 ( 
.A(n_746),
.B(n_486),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_689),
.B(n_707),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_613),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_767),
.Y(n_797)
);

BUFx2_ASAP7_75t_L g798 ( 
.A(n_674),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_629),
.B(n_526),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_688),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_706),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_767),
.Y(n_802)
);

OR2x2_ASAP7_75t_SL g803 ( 
.A(n_739),
.B(n_531),
.Y(n_803)
);

AOI211xp5_ASAP7_75t_L g804 ( 
.A1(n_676),
.A2(n_587),
.B(n_608),
.C(n_525),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_690),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_612),
.B(n_561),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_629),
.B(n_536),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_634),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_623),
.B(n_538),
.Y(n_809)
);

AND2x2_ASAP7_75t_SL g810 ( 
.A(n_617),
.B(n_538),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_612),
.B(n_562),
.Y(n_811)
);

INVxp67_ASAP7_75t_L g812 ( 
.A(n_656),
.Y(n_812)
);

AND2x4_ASAP7_75t_L g813 ( 
.A(n_634),
.B(n_597),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_705),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_726),
.Y(n_815)
);

A2O1A1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_733),
.A2(n_601),
.B(n_569),
.C(n_562),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_637),
.Y(n_817)
);

BUFx8_ASAP7_75t_L g818 ( 
.A(n_667),
.Y(n_818)
);

NOR3xp33_ASAP7_75t_L g819 ( 
.A(n_698),
.B(n_542),
.C(n_546),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_681),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_R g821 ( 
.A(n_675),
.B(n_600),
.Y(n_821)
);

BUFx12f_ASAP7_75t_L g822 ( 
.A(n_716),
.Y(n_822)
);

BUFx2_ASAP7_75t_L g823 ( 
.A(n_674),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_633),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_696),
.B(n_542),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_SL g826 ( 
.A1(n_610),
.A2(n_305),
.B1(n_172),
.B2(n_174),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_734),
.Y(n_827)
);

OAI21xp5_ASAP7_75t_L g828 ( 
.A1(n_645),
.A2(n_562),
.B(n_569),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_737),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_740),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_616),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_702),
.B(n_546),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_713),
.B(n_562),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_720),
.B(n_569),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_766),
.B(n_569),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_705),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_722),
.B(n_603),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_652),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_618),
.B(n_594),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_620),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_768),
.B(n_594),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_769),
.B(n_566),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_628),
.B(n_570),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_620),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_628),
.B(n_684),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_611),
.Y(n_846)
);

O2A1O1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_747),
.A2(n_609),
.B(n_575),
.C(n_505),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_671),
.B(n_575),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_694),
.A2(n_609),
.B1(n_497),
.B2(n_505),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_671),
.B(n_172),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_674),
.B(n_622),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_684),
.B(n_499),
.Y(n_852)
);

NAND2x2_ASAP7_75t_L g853 ( 
.A(n_770),
.B(n_581),
.Y(n_853)
);

OAI21x1_ASAP7_75t_L g854 ( 
.A1(n_614),
.A2(n_485),
.B(n_507),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_750),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_751),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_754),
.B(n_755),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_612),
.B(n_596),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_705),
.Y(n_859)
);

BUFx4f_ASAP7_75t_L g860 ( 
.A(n_626),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_612),
.B(n_596),
.Y(n_861)
);

BUFx12f_ASAP7_75t_L g862 ( 
.A(n_626),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_624),
.B(n_549),
.Y(n_863)
);

AND2x4_ASAP7_75t_SL g864 ( 
.A(n_759),
.B(n_761),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_694),
.A2(n_499),
.B1(n_484),
.B2(n_496),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_666),
.B(n_179),
.Y(n_866)
);

NAND2x1_ASAP7_75t_L g867 ( 
.A(n_631),
.B(n_480),
.Y(n_867)
);

INVxp67_ASAP7_75t_L g868 ( 
.A(n_758),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_763),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_764),
.B(n_549),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_685),
.B(n_596),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_672),
.B(n_480),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_762),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_753),
.Y(n_874)
);

INVx4_ASAP7_75t_L g875 ( 
.A(n_667),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_632),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_639),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_682),
.Y(n_878)
);

INVxp67_ASAP7_75t_SL g879 ( 
.A(n_646),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_639),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_717),
.B(n_735),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_SL g882 ( 
.A1(n_610),
.A2(n_194),
.B1(n_300),
.B2(n_295),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_765),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_717),
.B(n_480),
.Y(n_884)
);

NOR3xp33_ASAP7_75t_SL g885 ( 
.A(n_757),
.B(n_197),
.C(n_300),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_735),
.B(n_480),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_640),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_736),
.B(n_485),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_745),
.B(n_596),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_760),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_736),
.B(n_485),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_640),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_650),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_630),
.B(n_485),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_650),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_654),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_758),
.B(n_552),
.Y(n_897)
);

CKINVDCx20_ASAP7_75t_R g898 ( 
.A(n_661),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_749),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_654),
.Y(n_900)
);

OAI22xp5_ASAP7_75t_SL g901 ( 
.A1(n_743),
.A2(n_670),
.B1(n_724),
.B2(n_699),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_732),
.A2(n_731),
.B1(n_699),
.B2(n_708),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_636),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_700),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_619),
.B(n_596),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_644),
.A2(n_496),
.B1(n_491),
.B2(n_484),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_697),
.B(n_197),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_662),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_645),
.A2(n_680),
.B1(n_677),
.B2(n_642),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_721),
.B(n_552),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_733),
.A2(n_496),
.B1(n_491),
.B2(n_484),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_691),
.B(n_507),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_765),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_662),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_673),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_621),
.B(n_513),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_693),
.B(n_732),
.Y(n_917)
);

OAI22xp5_ASAP7_75t_L g918 ( 
.A1(n_648),
.A2(n_600),
.B1(n_487),
.B2(n_572),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_653),
.A2(n_600),
.B1(n_487),
.B2(n_572),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_731),
.A2(n_513),
.B1(n_535),
.B2(n_514),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_664),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_695),
.A2(n_535),
.B1(n_514),
.B2(n_519),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_728),
.B(n_514),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_695),
.A2(n_530),
.B1(n_519),
.B2(n_520),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_647),
.B(n_554),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_708),
.A2(n_530),
.B1(n_519),
.B2(n_520),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_664),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_704),
.B(n_554),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_669),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_669),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_678),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_678),
.B(n_556),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_687),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_687),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_747),
.A2(n_724),
.B1(n_668),
.B2(n_679),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_701),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_693),
.B(n_686),
.Y(n_937)
);

INVx4_ASAP7_75t_L g938 ( 
.A(n_673),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_638),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_729),
.B(n_520),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_697),
.B(n_285),
.Y(n_941)
);

INVxp67_ASAP7_75t_SL g942 ( 
.A(n_701),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_709),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_709),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_651),
.B(n_285),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_711),
.Y(n_946)
);

INVx4_ASAP7_75t_L g947 ( 
.A(n_814),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_779),
.B(n_752),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_793),
.B(n_683),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_845),
.B(n_756),
.Y(n_950)
);

A2O1A1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_845),
.A2(n_703),
.B(n_659),
.C(n_744),
.Y(n_951)
);

AOI21x1_ASAP7_75t_L g952 ( 
.A1(n_884),
.A2(n_665),
.B(n_748),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_879),
.A2(n_828),
.B(n_909),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_779),
.B(n_660),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_881),
.A2(n_615),
.B1(n_610),
.B2(n_617),
.Y(n_955)
);

A2O1A1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_902),
.A2(n_935),
.B(n_839),
.C(n_868),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_772),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_810),
.A2(n_790),
.B1(n_873),
.B2(n_937),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_809),
.B(n_711),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_930),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_812),
.B(n_878),
.Y(n_961)
);

O2A1O1Ixp33_ASAP7_75t_SL g962 ( 
.A1(n_816),
.A2(n_641),
.B(n_719),
.C(n_742),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_812),
.B(n_756),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_878),
.B(n_715),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_784),
.B(n_725),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_799),
.B(n_807),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_780),
.A2(n_487),
.B(n_572),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_817),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_810),
.A2(n_748),
.B1(n_741),
.B2(n_730),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_839),
.A2(n_741),
.B(n_730),
.C(n_723),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_777),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_824),
.B(n_715),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_818),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_L g974 ( 
.A1(n_937),
.A2(n_723),
.B1(n_718),
.B2(n_289),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_780),
.A2(n_806),
.B(n_786),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_868),
.A2(n_491),
.B(n_530),
.C(n_522),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_786),
.A2(n_487),
.B(n_572),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_843),
.B(n_556),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_782),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_811),
.A2(n_479),
.B(n_503),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_901),
.A2(n_600),
.B1(n_529),
.B2(n_522),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_930),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_816),
.A2(n_834),
.B(n_833),
.Y(n_983)
);

NOR3xp33_ASAP7_75t_L g984 ( 
.A(n_907),
.B(n_289),
.C(n_295),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_773),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_917),
.A2(n_522),
.B1(n_535),
.B2(n_529),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_835),
.A2(n_479),
.B(n_472),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_912),
.A2(n_479),
.B(n_472),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_917),
.A2(n_523),
.B1(n_529),
.B2(n_547),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_817),
.A2(n_581),
.B1(n_483),
.B2(n_467),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_814),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_942),
.A2(n_472),
.B(n_503),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_942),
.A2(n_472),
.B(n_503),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_945),
.A2(n_838),
.B(n_850),
.C(n_789),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_775),
.A2(n_523),
.B(n_547),
.C(n_476),
.Y(n_995)
);

AOI22xp33_ASAP7_75t_L g996 ( 
.A1(n_837),
.A2(n_941),
.B1(n_890),
.B2(n_874),
.Y(n_996)
);

AOI21x1_ASAP7_75t_L g997 ( 
.A1(n_886),
.A2(n_483),
.B(n_663),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_899),
.A2(n_503),
.B1(n_474),
.B2(n_472),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_788),
.B(n_476),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_934),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_785),
.Y(n_1001)
);

AOI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_837),
.A2(n_476),
.B1(n_475),
.B2(n_470),
.Y(n_1002)
);

INVx1_ASAP7_75t_SL g1003 ( 
.A(n_903),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_904),
.B(n_503),
.Y(n_1004)
);

INVxp67_ASAP7_75t_L g1005 ( 
.A(n_866),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_820),
.B(n_474),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_843),
.B(n_475),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_854),
.A2(n_475),
.B(n_470),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_776),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_SL g1010 ( 
.A(n_875),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_945),
.A2(n_467),
.B(n_470),
.C(n_4),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_800),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_820),
.A2(n_857),
.B1(n_827),
.B2(n_805),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_939),
.B(n_474),
.Y(n_1014)
);

OR2x6_ASAP7_75t_L g1015 ( 
.A(n_814),
.B(n_474),
.Y(n_1015)
);

O2A1O1Ixp33_ASAP7_75t_SL g1016 ( 
.A1(n_871),
.A2(n_467),
.B(n_72),
.C(n_156),
.Y(n_1016)
);

INVx6_ASAP7_75t_L g1017 ( 
.A(n_814),
.Y(n_1017)
);

BUFx8_ASAP7_75t_L g1018 ( 
.A(n_822),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_795),
.Y(n_1019)
);

O2A1O1Ixp5_ASAP7_75t_L g1020 ( 
.A1(n_852),
.A2(n_474),
.B(n_472),
.C(n_55),
.Y(n_1020)
);

OAI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_923),
.A2(n_155),
.B(n_146),
.Y(n_1021)
);

AOI21x1_ASAP7_75t_L g1022 ( 
.A1(n_888),
.A2(n_143),
.B(n_137),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_818),
.Y(n_1023)
);

NOR3xp33_ASAP7_75t_SL g1024 ( 
.A(n_915),
.B(n_0),
.C(n_3),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_898),
.B(n_4),
.Y(n_1025)
);

BUFx2_ASAP7_75t_L g1026 ( 
.A(n_798),
.Y(n_1026)
);

O2A1O1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_819),
.A2(n_7),
.B(n_13),
.C(n_18),
.Y(n_1027)
);

AO32x2_ASAP7_75t_L g1028 ( 
.A1(n_906),
.A2(n_7),
.A3(n_23),
.B1(n_26),
.B2(n_28),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_823),
.B(n_23),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_848),
.B(n_26),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_862),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_846),
.B(n_32),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_874),
.B(n_32),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_891),
.A2(n_84),
.B(n_130),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_934),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_826),
.B(n_35),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_890),
.B(n_35),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_792),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_819),
.A2(n_38),
.B(n_40),
.C(n_42),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_815),
.B(n_38),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_826),
.B(n_882),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_829),
.A2(n_40),
.B1(n_42),
.B2(n_44),
.Y(n_1042)
);

INVxp67_ASAP7_75t_L g1043 ( 
.A(n_778),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_SL g1044 ( 
.A1(n_871),
.A2(n_91),
.B(n_123),
.C(n_118),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_858),
.A2(n_80),
.B(n_113),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_830),
.B(n_44),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_855),
.B(n_45),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_869),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_858),
.A2(n_861),
.B(n_872),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_846),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_842),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_825),
.B(n_46),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_923),
.A2(n_94),
.B(n_107),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_773),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_841),
.A2(n_48),
.B(n_50),
.C(n_52),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_804),
.A2(n_52),
.B1(n_59),
.B2(n_88),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_876),
.Y(n_1057)
);

INVxp67_ASAP7_75t_L g1058 ( 
.A(n_778),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_783),
.A2(n_894),
.B(n_928),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_836),
.B(n_96),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_856),
.A2(n_98),
.B(n_132),
.C(n_864),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_877),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_875),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_832),
.B(n_856),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_808),
.B(n_813),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_887),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_925),
.A2(n_919),
.B(n_918),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_864),
.B(n_808),
.Y(n_1068)
);

OR2x6_ASAP7_75t_L g1069 ( 
.A(n_938),
.B(n_836),
.Y(n_1069)
);

NOR2xp67_ASAP7_75t_L g1070 ( 
.A(n_938),
.B(n_851),
.Y(n_1070)
);

NAND3xp33_ASAP7_75t_L g1071 ( 
.A(n_885),
.B(n_882),
.C(n_813),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_940),
.A2(n_911),
.B(n_906),
.Y(n_1072)
);

INVx4_ASAP7_75t_L g1073 ( 
.A(n_773),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_946),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_897),
.B(n_771),
.Y(n_1075)
);

O2A1O1Ixp5_ASAP7_75t_L g1076 ( 
.A1(n_889),
.A2(n_916),
.B(n_910),
.C(n_905),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_946),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_885),
.A2(n_910),
.B(n_897),
.C(n_847),
.Y(n_1078)
);

INVx1_ASAP7_75t_SL g1079 ( 
.A(n_803),
.Y(n_1079)
);

OR2x2_ASAP7_75t_L g1080 ( 
.A(n_851),
.B(n_859),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_771),
.B(n_774),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_774),
.A2(n_944),
.B(n_943),
.C(n_936),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_773),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_801),
.B(n_796),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_889),
.A2(n_932),
.B(n_801),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_796),
.B(n_797),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_953),
.A2(n_787),
.B(n_860),
.Y(n_1087)
);

AO31x2_ASAP7_75t_L g1088 ( 
.A1(n_990),
.A2(n_900),
.A3(n_929),
.B(n_927),
.Y(n_1088)
);

AO32x2_ASAP7_75t_L g1089 ( 
.A1(n_958),
.A2(n_853),
.A3(n_911),
.B1(n_865),
.B2(n_849),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1059),
.A2(n_787),
.B(n_860),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_971),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_965),
.B(n_859),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_980),
.A2(n_926),
.B(n_922),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_949),
.A2(n_787),
.B(n_791),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_948),
.A2(n_794),
.B1(n_853),
.B2(n_870),
.Y(n_1095)
);

OR2x6_ASAP7_75t_L g1096 ( 
.A(n_1069),
.B(n_787),
.Y(n_1096)
);

BUFx3_ASAP7_75t_L g1097 ( 
.A(n_957),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_956),
.A2(n_924),
.B(n_865),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_968),
.Y(n_1099)
);

NAND3xp33_ASAP7_75t_L g1100 ( 
.A(n_994),
.B(n_849),
.C(n_920),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1005),
.B(n_863),
.Y(n_1101)
);

OR2x2_ASAP7_75t_L g1102 ( 
.A(n_1003),
.B(n_802),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1067),
.A2(n_781),
.B(n_840),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_979),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_966),
.A2(n_867),
.B(n_933),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_1070),
.B(n_863),
.Y(n_1106)
);

AO21x2_ASAP7_75t_L g1107 ( 
.A1(n_952),
.A2(n_821),
.B(n_893),
.Y(n_1107)
);

BUFx8_ASAP7_75t_L g1108 ( 
.A(n_1010),
.Y(n_1108)
);

AOI21x1_ASAP7_75t_SL g1109 ( 
.A1(n_1030),
.A2(n_794),
.B(n_821),
.Y(n_1109)
);

OA21x2_ASAP7_75t_L g1110 ( 
.A1(n_983),
.A2(n_895),
.B(n_921),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1051),
.B(n_831),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_1069),
.B(n_844),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_954),
.A2(n_896),
.B(n_908),
.C(n_880),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_1038),
.Y(n_1114)
);

AOI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_984),
.A2(n_883),
.B1(n_892),
.B2(n_914),
.Y(n_1115)
);

AOI21x1_ASAP7_75t_L g1116 ( 
.A1(n_990),
.A2(n_931),
.B(n_913),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_955),
.A2(n_913),
.B1(n_933),
.B2(n_958),
.Y(n_1117)
);

CKINVDCx16_ASAP7_75t_R g1118 ( 
.A(n_1023),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_951),
.A2(n_913),
.B(n_933),
.Y(n_1119)
);

AOI21x1_ASAP7_75t_L g1120 ( 
.A1(n_997),
.A2(n_978),
.B(n_988),
.Y(n_1120)
);

OR2x2_ASAP7_75t_L g1121 ( 
.A(n_1009),
.B(n_961),
.Y(n_1121)
);

INVxp67_ASAP7_75t_L g1122 ( 
.A(n_1026),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1001),
.Y(n_1123)
);

BUFx4_ASAP7_75t_SL g1124 ( 
.A(n_973),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1007),
.A2(n_983),
.B(n_967),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_SL g1126 ( 
.A1(n_1041),
.A2(n_1036),
.B(n_1071),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_987),
.A2(n_975),
.B(n_993),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_991),
.Y(n_1128)
);

O2A1O1Ixp5_ASAP7_75t_SL g1129 ( 
.A1(n_1056),
.A2(n_1042),
.B(n_1048),
.C(n_1013),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_996),
.A2(n_950),
.B1(n_1072),
.B2(n_1056),
.Y(n_1130)
);

INVxp67_ASAP7_75t_L g1131 ( 
.A(n_1019),
.Y(n_1131)
);

NAND3xp33_ASAP7_75t_L g1132 ( 
.A(n_1027),
.B(n_1039),
.C(n_1037),
.Y(n_1132)
);

AO31x2_ASAP7_75t_L g1133 ( 
.A1(n_970),
.A2(n_969),
.A3(n_995),
.B(n_974),
.Y(n_1133)
);

AO21x2_ASAP7_75t_L g1134 ( 
.A1(n_1072),
.A2(n_978),
.B(n_992),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_SL g1135 ( 
.A1(n_1021),
.A2(n_1053),
.B(n_1078),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_977),
.A2(n_959),
.B(n_1064),
.Y(n_1136)
);

OA21x2_ASAP7_75t_L g1137 ( 
.A1(n_1020),
.A2(n_1076),
.B(n_1053),
.Y(n_1137)
);

INVx4_ASAP7_75t_SL g1138 ( 
.A(n_1017),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_959),
.A2(n_962),
.B(n_999),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1013),
.B(n_972),
.Y(n_1140)
);

NAND3xp33_ASAP7_75t_SL g1141 ( 
.A(n_1025),
.B(n_1079),
.C(n_1011),
.Y(n_1141)
);

O2A1O1Ixp5_ASAP7_75t_SL g1142 ( 
.A1(n_1042),
.A2(n_1048),
.B(n_974),
.C(n_1006),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_969),
.A2(n_976),
.B(n_1082),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1012),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1057),
.Y(n_1145)
);

O2A1O1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_1055),
.A2(n_1033),
.B(n_1046),
.C(n_1040),
.Y(n_1146)
);

AND2x6_ASAP7_75t_L g1147 ( 
.A(n_991),
.B(n_1060),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_1022),
.A2(n_1084),
.B(n_1086),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_963),
.B(n_964),
.Y(n_1149)
);

OA21x2_ASAP7_75t_L g1150 ( 
.A1(n_1021),
.A2(n_1034),
.B(n_1052),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1075),
.A2(n_989),
.B(n_986),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1004),
.A2(n_1081),
.B(n_1065),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_1068),
.B(n_1050),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_981),
.A2(n_1061),
.B(n_1047),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1045),
.A2(n_1066),
.B(n_1062),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1014),
.A2(n_1032),
.B(n_1043),
.C(n_1058),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_960),
.B(n_1035),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_982),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_1080),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1002),
.A2(n_1016),
.B(n_998),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1015),
.A2(n_1044),
.B(n_1000),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_985),
.A2(n_1077),
.B(n_1074),
.Y(n_1162)
);

BUFx10_ASAP7_75t_L g1163 ( 
.A(n_1010),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1060),
.A2(n_985),
.B(n_1015),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1054),
.B(n_1083),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1028),
.Y(n_1166)
);

AOI211x1_ASAP7_75t_L g1167 ( 
.A1(n_1028),
.A2(n_1024),
.B(n_1029),
.C(n_1054),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1028),
.Y(n_1168)
);

AO32x2_ASAP7_75t_L g1169 ( 
.A1(n_1073),
.A2(n_947),
.A3(n_1015),
.B1(n_1083),
.B2(n_1054),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1083),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_947),
.B(n_991),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1073),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1069),
.A2(n_1063),
.B(n_1031),
.Y(n_1173)
);

AO31x2_ASAP7_75t_L g1174 ( 
.A1(n_1017),
.A2(n_990),
.A3(n_953),
.B(n_956),
.Y(n_1174)
);

NAND2xp33_ASAP7_75t_R g1175 ( 
.A(n_1017),
.B(n_1018),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1018),
.B(n_966),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_948),
.B(n_534),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_953),
.A2(n_1059),
.B(n_909),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_971),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_966),
.A2(n_793),
.B1(n_881),
.B2(n_845),
.Y(n_1180)
);

AOI21xp33_ASAP7_75t_L g1181 ( 
.A1(n_994),
.A2(n_881),
.B(n_845),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_SL g1182 ( 
.A1(n_956),
.A2(n_881),
.B(n_793),
.C(n_845),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_953),
.A2(n_1059),
.B(n_909),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_966),
.B(n_845),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_953),
.A2(n_1059),
.B(n_909),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_957),
.Y(n_1186)
);

NOR2x1_ASAP7_75t_R g1187 ( 
.A(n_973),
.B(n_1023),
.Y(n_1187)
);

INVx2_ASAP7_75t_SL g1188 ( 
.A(n_957),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_957),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1008),
.A2(n_1085),
.B(n_1049),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_966),
.B(n_845),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_966),
.B(n_845),
.Y(n_1192)
);

NAND2x1_ASAP7_75t_L g1193 ( 
.A(n_1015),
.B(n_773),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_953),
.A2(n_1059),
.B(n_909),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1009),
.B(n_550),
.Y(n_1195)
);

OA21x2_ASAP7_75t_L g1196 ( 
.A1(n_953),
.A2(n_983),
.B(n_1067),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1008),
.A2(n_1085),
.B(n_1049),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_948),
.B(n_534),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_948),
.B(n_534),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_957),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_1038),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_966),
.B(n_793),
.Y(n_1202)
);

NAND2x1p5_ASAP7_75t_L g1203 ( 
.A(n_947),
.B(n_814),
.Y(n_1203)
);

NOR2x1_ASAP7_75t_L g1204 ( 
.A(n_947),
.B(n_434),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_971),
.Y(n_1205)
);

NAND2x1p5_ASAP7_75t_L g1206 ( 
.A(n_947),
.B(n_814),
.Y(n_1206)
);

OAI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_956),
.A2(n_953),
.B(n_845),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1041),
.A2(n_845),
.B1(n_901),
.B2(n_881),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_971),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1009),
.B(n_550),
.Y(n_1210)
);

AOI221xp5_ASAP7_75t_L g1211 ( 
.A1(n_1041),
.A2(n_528),
.B1(n_901),
.B2(n_676),
.C(n_845),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_SL g1212 ( 
.A1(n_1021),
.A2(n_1053),
.B(n_1078),
.Y(n_1212)
);

AO21x2_ASAP7_75t_L g1213 ( 
.A1(n_1067),
.A2(n_953),
.B(n_952),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_956),
.A2(n_845),
.B(n_881),
.C(n_793),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_971),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1008),
.A2(n_1085),
.B(n_1049),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1008),
.A2(n_1085),
.B(n_1049),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1008),
.A2(n_1085),
.B(n_1049),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_965),
.B(n_907),
.Y(n_1219)
);

O2A1O1Ixp5_ASAP7_75t_SL g1220 ( 
.A1(n_990),
.A2(n_1056),
.B(n_731),
.C(n_460),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_953),
.A2(n_1059),
.B(n_909),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_965),
.B(n_907),
.Y(n_1222)
);

NOR2x1_ASAP7_75t_L g1223 ( 
.A(n_947),
.B(n_434),
.Y(n_1223)
);

CKINVDCx14_ASAP7_75t_R g1224 ( 
.A(n_973),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_953),
.A2(n_1059),
.B(n_909),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_SL g1226 ( 
.A1(n_1021),
.A2(n_1053),
.B(n_1078),
.Y(n_1226)
);

AND2x6_ASAP7_75t_L g1227 ( 
.A(n_991),
.B(n_917),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_953),
.A2(n_1059),
.B(n_909),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1104),
.Y(n_1229)
);

OA21x2_ASAP7_75t_L g1230 ( 
.A1(n_1178),
.A2(n_1185),
.B(n_1183),
.Y(n_1230)
);

OA21x2_ASAP7_75t_L g1231 ( 
.A1(n_1194),
.A2(n_1225),
.B(n_1221),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1110),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1124),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_1174),
.Y(n_1234)
);

INVx4_ASAP7_75t_L g1235 ( 
.A(n_1138),
.Y(n_1235)
);

AO31x2_ASAP7_75t_L g1236 ( 
.A1(n_1228),
.A2(n_1125),
.A3(n_1130),
.B(n_1117),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1097),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1211),
.A2(n_1208),
.B1(n_1180),
.B2(n_1181),
.Y(n_1238)
);

INVxp33_ASAP7_75t_SL g1239 ( 
.A(n_1114),
.Y(n_1239)
);

AO31x2_ASAP7_75t_L g1240 ( 
.A1(n_1130),
.A2(n_1117),
.A3(n_1214),
.B(n_1136),
.Y(n_1240)
);

INVx4_ASAP7_75t_L g1241 ( 
.A(n_1138),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1123),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1207),
.A2(n_1180),
.B(n_1181),
.C(n_1098),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1207),
.A2(n_1098),
.B(n_1202),
.C(n_1198),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1182),
.A2(n_1139),
.B(n_1090),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1217),
.A2(n_1218),
.B(n_1127),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1205),
.Y(n_1247)
);

OAI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1202),
.A2(n_1126),
.B1(n_1177),
.B2(n_1199),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1116),
.A2(n_1120),
.B(n_1093),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1209),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1215),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1091),
.Y(n_1252)
);

INVx6_ASAP7_75t_SL g1253 ( 
.A(n_1096),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1219),
.B(n_1222),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1148),
.A2(n_1119),
.B(n_1087),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1094),
.A2(n_1119),
.B(n_1155),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1169),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1126),
.B(n_1141),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1146),
.A2(n_1129),
.B(n_1132),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1144),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1121),
.B(n_1149),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_1169),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1092),
.B(n_1101),
.Y(n_1263)
);

OAI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1154),
.A2(n_1220),
.B(n_1142),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1143),
.A2(n_1162),
.B(n_1161),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1151),
.A2(n_1152),
.B(n_1105),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1179),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1145),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1159),
.B(n_1102),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1157),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1157),
.Y(n_1271)
);

NAND3xp33_ASAP7_75t_L g1272 ( 
.A(n_1095),
.B(n_1156),
.C(n_1176),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_SL g1273 ( 
.A1(n_1164),
.A2(n_1140),
.B(n_1160),
.Y(n_1273)
);

BUFx2_ASAP7_75t_R g1274 ( 
.A(n_1201),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1088),
.Y(n_1275)
);

AOI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1100),
.A2(n_1137),
.B(n_1150),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_1112),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1160),
.A2(n_1196),
.B(n_1137),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1164),
.B(n_1112),
.Y(n_1279)
);

INVx1_ASAP7_75t_SL g1280 ( 
.A(n_1200),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_1186),
.Y(n_1281)
);

CKINVDCx11_ASAP7_75t_R g1282 ( 
.A(n_1163),
.Y(n_1282)
);

O2A1O1Ixp33_ASAP7_75t_SL g1283 ( 
.A1(n_1113),
.A2(n_1100),
.B(n_1168),
.C(n_1166),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1200),
.B(n_1099),
.Y(n_1284)
);

INVx6_ASAP7_75t_L g1285 ( 
.A(n_1138),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1196),
.A2(n_1150),
.B1(n_1153),
.B2(n_1204),
.Y(n_1286)
);

OA21x2_ASAP7_75t_L g1287 ( 
.A1(n_1111),
.A2(n_1115),
.B(n_1213),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1188),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1109),
.A2(n_1193),
.B(n_1173),
.Y(n_1289)
);

INVx3_ASAP7_75t_L g1290 ( 
.A(n_1106),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1108),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1173),
.A2(n_1165),
.B(n_1206),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1203),
.A2(n_1206),
.B(n_1165),
.Y(n_1293)
);

AOI22x1_ASAP7_75t_L g1294 ( 
.A1(n_1172),
.A2(n_1106),
.B1(n_1158),
.B2(n_1203),
.Y(n_1294)
);

NOR2xp67_ASAP7_75t_L g1295 ( 
.A(n_1189),
.B(n_1131),
.Y(n_1295)
);

NAND3xp33_ASAP7_75t_L g1296 ( 
.A(n_1167),
.B(n_1195),
.C(n_1210),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1223),
.A2(n_1170),
.B(n_1171),
.Y(n_1297)
);

CKINVDCx6p67_ASAP7_75t_R g1298 ( 
.A(n_1118),
.Y(n_1298)
);

OR2x6_ASAP7_75t_L g1299 ( 
.A(n_1096),
.B(n_1122),
.Y(n_1299)
);

OR2x2_ASAP7_75t_L g1300 ( 
.A(n_1096),
.B(n_1128),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1174),
.A2(n_1088),
.B(n_1107),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1224),
.A2(n_1147),
.B1(n_1169),
.B2(n_1227),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1088),
.A2(n_1107),
.B(n_1134),
.Y(n_1303)
);

CKINVDCx20_ASAP7_75t_R g1304 ( 
.A(n_1108),
.Y(n_1304)
);

OAI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1175),
.A2(n_1089),
.B1(n_1133),
.B2(n_1187),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1133),
.Y(n_1306)
);

AOI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1089),
.A2(n_901),
.B1(n_845),
.B2(n_327),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1208),
.A2(n_1184),
.B1(n_1192),
.B2(n_1191),
.Y(n_1308)
);

AO21x2_ASAP7_75t_L g1309 ( 
.A1(n_1178),
.A2(n_1225),
.B(n_1221),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1127),
.A2(n_1197),
.B(n_1190),
.Y(n_1310)
);

NAND3xp33_ASAP7_75t_L g1311 ( 
.A(n_1211),
.B(n_845),
.C(n_881),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1177),
.B(n_1198),
.Y(n_1312)
);

OAI22x1_ASAP7_75t_L g1313 ( 
.A1(n_1095),
.A2(n_1041),
.B1(n_1071),
.B2(n_1177),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1127),
.A2(n_1197),
.B(n_1190),
.Y(n_1314)
);

AOI22x1_ASAP7_75t_L g1315 ( 
.A1(n_1135),
.A2(n_1212),
.B1(n_1226),
.B2(n_1207),
.Y(n_1315)
);

OAI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1214),
.A2(n_845),
.B(n_881),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1127),
.A2(n_1197),
.B(n_1190),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1174),
.Y(n_1318)
);

O2A1O1Ixp33_ASAP7_75t_SL g1319 ( 
.A1(n_1214),
.A2(n_881),
.B(n_956),
.C(n_1056),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1177),
.B(n_1198),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_1124),
.Y(n_1321)
);

BUFx2_ASAP7_75t_R g1322 ( 
.A(n_1114),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1211),
.A2(n_1041),
.B1(n_845),
.B2(n_1208),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1097),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1219),
.B(n_1222),
.Y(n_1325)
);

NOR3xp33_ASAP7_75t_L g1326 ( 
.A(n_1211),
.B(n_881),
.C(n_845),
.Y(n_1326)
);

INVx1_ASAP7_75t_SL g1327 ( 
.A(n_1200),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_SL g1328 ( 
.A1(n_1208),
.A2(n_826),
.B1(n_882),
.B2(n_901),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1219),
.B(n_1222),
.Y(n_1329)
);

INVx1_ASAP7_75t_SL g1330 ( 
.A(n_1200),
.Y(n_1330)
);

NAND2x1p5_ASAP7_75t_L g1331 ( 
.A(n_1193),
.B(n_947),
.Y(n_1331)
);

OA21x2_ASAP7_75t_L g1332 ( 
.A1(n_1178),
.A2(n_1185),
.B(n_1183),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1127),
.A2(n_1197),
.B(n_1190),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_1097),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1112),
.Y(n_1335)
);

OA21x2_ASAP7_75t_L g1336 ( 
.A1(n_1178),
.A2(n_1185),
.B(n_1183),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1104),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1104),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_1169),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1110),
.Y(n_1340)
);

AND2x6_ASAP7_75t_SL g1341 ( 
.A(n_1176),
.B(n_1025),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1184),
.B(n_1191),
.Y(n_1342)
);

AOI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1177),
.A2(n_901),
.B1(n_845),
.B2(n_327),
.Y(n_1343)
);

O2A1O1Ixp5_ASAP7_75t_L g1344 ( 
.A1(n_1207),
.A2(n_845),
.B(n_881),
.C(n_1181),
.Y(n_1344)
);

OAI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1214),
.A2(n_845),
.B(n_881),
.Y(n_1345)
);

INVxp67_ASAP7_75t_L g1346 ( 
.A(n_1186),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1177),
.B(n_1198),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1177),
.B(n_1198),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1110),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1211),
.A2(n_1041),
.B1(n_845),
.B2(n_1208),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1178),
.A2(n_1225),
.B(n_1221),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1104),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1103),
.A2(n_1217),
.B(n_1216),
.Y(n_1353)
);

O2A1O1Ixp33_ASAP7_75t_L g1354 ( 
.A1(n_1214),
.A2(n_881),
.B(n_845),
.C(n_1181),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1312),
.A2(n_1320),
.B1(n_1348),
.B2(n_1347),
.Y(n_1355)
);

NOR2xp67_ASAP7_75t_L g1356 ( 
.A(n_1237),
.B(n_1272),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1263),
.B(n_1254),
.Y(n_1357)
);

OA21x2_ASAP7_75t_L g1358 ( 
.A1(n_1264),
.A2(n_1303),
.B(n_1245),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1261),
.B(n_1312),
.Y(n_1359)
);

O2A1O1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1320),
.A2(n_1347),
.B(n_1348),
.C(n_1326),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1279),
.B(n_1292),
.Y(n_1361)
);

O2A1O1Ixp5_ASAP7_75t_L g1362 ( 
.A1(n_1259),
.A2(n_1316),
.B(n_1345),
.C(n_1344),
.Y(n_1362)
);

O2A1O1Ixp33_ASAP7_75t_L g1363 ( 
.A1(n_1319),
.A2(n_1354),
.B(n_1248),
.C(n_1244),
.Y(n_1363)
);

OA21x2_ASAP7_75t_L g1364 ( 
.A1(n_1249),
.A2(n_1278),
.B(n_1301),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_1279),
.B(n_1292),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1267),
.Y(n_1366)
);

OA22x2_ASAP7_75t_L g1367 ( 
.A1(n_1328),
.A2(n_1343),
.B1(n_1307),
.B2(n_1313),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1252),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1325),
.B(n_1329),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1234),
.Y(n_1370)
);

AOI221xp5_ASAP7_75t_L g1371 ( 
.A1(n_1311),
.A2(n_1319),
.B1(n_1350),
.B2(n_1323),
.C(n_1238),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1342),
.B(n_1308),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1232),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1258),
.B(n_1269),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1279),
.B(n_1277),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1280),
.B(n_1327),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1244),
.B(n_1243),
.Y(n_1377)
);

INVxp67_ASAP7_75t_L g1378 ( 
.A(n_1284),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_SL g1379 ( 
.A1(n_1302),
.A2(n_1241),
.B(n_1235),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_1233),
.Y(n_1380)
);

OR2x2_ASAP7_75t_L g1381 ( 
.A(n_1330),
.B(n_1258),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1306),
.B(n_1257),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_SL g1383 ( 
.A1(n_1235),
.A2(n_1241),
.B(n_1339),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1335),
.B(n_1251),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1323),
.A2(n_1350),
.B1(n_1238),
.B2(n_1296),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1260),
.Y(n_1386)
);

CKINVDCx6p67_ASAP7_75t_R g1387 ( 
.A(n_1304),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1270),
.B(n_1271),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1299),
.A2(n_1295),
.B1(n_1346),
.B2(n_1281),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1251),
.B(n_1284),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1229),
.B(n_1242),
.Y(n_1391)
);

AO21x2_ASAP7_75t_L g1392 ( 
.A1(n_1351),
.A2(n_1276),
.B(n_1353),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1247),
.B(n_1250),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1268),
.B(n_1352),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_1289),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1309),
.A2(n_1230),
.B(n_1231),
.Y(n_1396)
);

O2A1O1Ixp5_ASAP7_75t_L g1397 ( 
.A1(n_1305),
.A2(n_1306),
.B(n_1275),
.C(n_1290),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1337),
.B(n_1338),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1290),
.B(n_1288),
.Y(n_1399)
);

CKINVDCx20_ASAP7_75t_R g1400 ( 
.A(n_1304),
.Y(n_1400)
);

NAND2x1_ASAP7_75t_L g1401 ( 
.A(n_1273),
.B(n_1285),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1324),
.B(n_1334),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1315),
.B(n_1305),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1285),
.A2(n_1253),
.B1(n_1286),
.B2(n_1300),
.Y(n_1404)
);

OA21x2_ASAP7_75t_L g1405 ( 
.A1(n_1265),
.A2(n_1256),
.B(n_1255),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1297),
.B(n_1289),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1298),
.B(n_1293),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1286),
.B(n_1331),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1285),
.A2(n_1253),
.B1(n_1294),
.B2(n_1239),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1309),
.A2(n_1230),
.B(n_1231),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1331),
.B(n_1322),
.Y(n_1411)
);

AOI21x1_ASAP7_75t_SL g1412 ( 
.A1(n_1318),
.A2(n_1341),
.B(n_1282),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1274),
.B(n_1262),
.Y(n_1413)
);

NAND2xp33_ASAP7_75t_SL g1414 ( 
.A(n_1257),
.B(n_1339),
.Y(n_1414)
);

O2A1O1Ixp5_ASAP7_75t_L g1415 ( 
.A1(n_1340),
.A2(n_1349),
.B(n_1240),
.C(n_1283),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1253),
.A2(n_1239),
.B1(n_1291),
.B2(n_1257),
.Y(n_1416)
);

OA22x2_ASAP7_75t_L g1417 ( 
.A1(n_1291),
.A2(n_1233),
.B1(n_1321),
.B2(n_1255),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1262),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1321),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1240),
.B(n_1287),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_1282),
.Y(n_1421)
);

OA21x2_ASAP7_75t_L g1422 ( 
.A1(n_1266),
.A2(n_1310),
.B(n_1333),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1240),
.B(n_1236),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1332),
.Y(n_1424)
);

OA21x2_ASAP7_75t_L g1425 ( 
.A1(n_1314),
.A2(n_1317),
.B(n_1333),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1336),
.A2(n_1317),
.B(n_1246),
.Y(n_1426)
);

INVx1_ASAP7_75t_SL g1427 ( 
.A(n_1280),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1234),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1263),
.B(n_1254),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1261),
.B(n_1269),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1261),
.B(n_1269),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1312),
.A2(n_1320),
.B1(n_1348),
.B2(n_1347),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1261),
.B(n_1269),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1312),
.A2(n_1320),
.B1(n_1348),
.B2(n_1347),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1261),
.B(n_1312),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_SL g1436 ( 
.A1(n_1244),
.A2(n_1056),
.B(n_1214),
.Y(n_1436)
);

A2O1A1Ixp33_ASAP7_75t_L g1437 ( 
.A1(n_1326),
.A2(n_845),
.B(n_881),
.C(n_1311),
.Y(n_1437)
);

INVx1_ASAP7_75t_SL g1438 ( 
.A(n_1280),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1261),
.B(n_1312),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1261),
.B(n_1312),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1312),
.A2(n_1320),
.B1(n_1348),
.B2(n_1347),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1261),
.B(n_1312),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1261),
.B(n_1312),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1312),
.A2(n_1320),
.B1(n_1348),
.B2(n_1347),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1423),
.B(n_1361),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1372),
.B(n_1377),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_SL g1447 ( 
.A1(n_1437),
.A2(n_1363),
.B(n_1371),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1361),
.B(n_1365),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1377),
.B(n_1359),
.Y(n_1449)
);

INVx2_ASAP7_75t_SL g1450 ( 
.A(n_1394),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1373),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1426),
.A2(n_1410),
.B(n_1396),
.Y(n_1452)
);

OA21x2_ASAP7_75t_L g1453 ( 
.A1(n_1397),
.A2(n_1362),
.B(n_1415),
.Y(n_1453)
);

NAND2xp33_ASAP7_75t_R g1454 ( 
.A(n_1421),
.B(n_1380),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1382),
.B(n_1361),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1365),
.B(n_1418),
.Y(n_1456)
);

AOI21xp5_ASAP7_75t_SL g1457 ( 
.A1(n_1437),
.A2(n_1385),
.B(n_1360),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1365),
.B(n_1406),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1367),
.A2(n_1355),
.B1(n_1441),
.B2(n_1434),
.Y(n_1459)
);

BUFx2_ASAP7_75t_L g1460 ( 
.A(n_1414),
.Y(n_1460)
);

NOR2x1_ASAP7_75t_R g1461 ( 
.A(n_1421),
.B(n_1380),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1435),
.B(n_1439),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1375),
.B(n_1420),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1366),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1368),
.Y(n_1465)
);

INVx2_ASAP7_75t_SL g1466 ( 
.A(n_1407),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1390),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1440),
.B(n_1442),
.Y(n_1468)
);

NOR3xp33_ASAP7_75t_L g1469 ( 
.A(n_1432),
.B(n_1444),
.C(n_1356),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1414),
.Y(n_1470)
);

OA21x2_ASAP7_75t_L g1471 ( 
.A1(n_1403),
.A2(n_1424),
.B(n_1386),
.Y(n_1471)
);

OR2x6_ASAP7_75t_L g1472 ( 
.A(n_1436),
.B(n_1383),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_1370),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1395),
.B(n_1408),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1370),
.B(n_1428),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1374),
.B(n_1384),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1425),
.Y(n_1477)
);

AO21x2_ASAP7_75t_L g1478 ( 
.A1(n_1392),
.A2(n_1436),
.B(n_1404),
.Y(n_1478)
);

OR2x6_ASAP7_75t_L g1479 ( 
.A(n_1383),
.B(n_1379),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1376),
.Y(n_1480)
);

OR2x6_ASAP7_75t_L g1481 ( 
.A(n_1379),
.B(n_1417),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1391),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1388),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1393),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1398),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1381),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1367),
.A2(n_1443),
.B1(n_1417),
.B2(n_1389),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1358),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1358),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1471),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1471),
.B(n_1364),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1465),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1477),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1471),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1477),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1471),
.Y(n_1496)
);

INVx2_ASAP7_75t_SL g1497 ( 
.A(n_1448),
.Y(n_1497)
);

OAI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1457),
.A2(n_1378),
.B(n_1401),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1448),
.B(n_1458),
.Y(n_1499)
);

INVxp67_ASAP7_75t_L g1500 ( 
.A(n_1486),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1448),
.B(n_1405),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1451),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1458),
.B(n_1405),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1483),
.B(n_1430),
.Y(n_1504)
);

AOI33xp33_ASAP7_75t_L g1505 ( 
.A1(n_1459),
.A2(n_1438),
.A3(n_1427),
.B1(n_1369),
.B2(n_1429),
.B3(n_1357),
.Y(n_1505)
);

AOI221xp5_ASAP7_75t_L g1506 ( 
.A1(n_1447),
.A2(n_1409),
.B1(n_1433),
.B2(n_1431),
.C(n_1416),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1458),
.B(n_1413),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1475),
.B(n_1422),
.Y(n_1508)
);

INVx5_ASAP7_75t_L g1509 ( 
.A(n_1472),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1483),
.B(n_1399),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1455),
.B(n_1422),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1473),
.Y(n_1512)
);

BUFx2_ASAP7_75t_SL g1513 ( 
.A(n_1460),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_SL g1514 ( 
.A1(n_1457),
.A2(n_1400),
.B1(n_1411),
.B2(n_1402),
.Y(n_1514)
);

OAI221xp5_ASAP7_75t_L g1515 ( 
.A1(n_1514),
.A2(n_1469),
.B1(n_1498),
.B2(n_1447),
.C(n_1487),
.Y(n_1515)
);

AND2x2_ASAP7_75t_SL g1516 ( 
.A(n_1505),
.B(n_1460),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1499),
.B(n_1474),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1499),
.B(n_1497),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1514),
.A2(n_1472),
.B1(n_1481),
.B2(n_1446),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_L g1520 ( 
.A(n_1512),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1493),
.Y(n_1521)
);

INVxp67_ASAP7_75t_L g1522 ( 
.A(n_1510),
.Y(n_1522)
);

OAI31xp33_ASAP7_75t_L g1523 ( 
.A1(n_1505),
.A2(n_1446),
.A3(n_1468),
.B(n_1462),
.Y(n_1523)
);

AOI222xp33_ASAP7_75t_L g1524 ( 
.A1(n_1506),
.A2(n_1449),
.B1(n_1480),
.B2(n_1461),
.C1(n_1400),
.C2(n_1482),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1506),
.A2(n_1472),
.B1(n_1481),
.B2(n_1479),
.Y(n_1525)
);

OAI33xp33_ASAP7_75t_L g1526 ( 
.A1(n_1500),
.A2(n_1449),
.A3(n_1482),
.B1(n_1485),
.B2(n_1484),
.B3(n_1464),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1508),
.B(n_1445),
.Y(n_1527)
);

INVxp67_ASAP7_75t_L g1528 ( 
.A(n_1510),
.Y(n_1528)
);

OAI221xp5_ASAP7_75t_L g1529 ( 
.A1(n_1498),
.A2(n_1481),
.B1(n_1472),
.B2(n_1466),
.C(n_1479),
.Y(n_1529)
);

OAI211xp5_ASAP7_75t_SL g1530 ( 
.A1(n_1500),
.A2(n_1485),
.B(n_1484),
.C(n_1466),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1509),
.A2(n_1472),
.B1(n_1481),
.B2(n_1479),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1502),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1504),
.B(n_1476),
.Y(n_1533)
);

BUFx12f_ASAP7_75t_L g1534 ( 
.A(n_1507),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1508),
.B(n_1445),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1509),
.A2(n_1481),
.B1(n_1474),
.B2(n_1478),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1511),
.B(n_1463),
.Y(n_1537)
);

AO21x2_ASAP7_75t_L g1538 ( 
.A1(n_1490),
.A2(n_1489),
.B(n_1488),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_SL g1539 ( 
.A1(n_1509),
.A2(n_1470),
.B1(n_1478),
.B2(n_1453),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1502),
.Y(n_1540)
);

OAI31xp33_ASAP7_75t_SL g1541 ( 
.A1(n_1507),
.A2(n_1412),
.A3(n_1463),
.B(n_1456),
.Y(n_1541)
);

INVx5_ASAP7_75t_L g1542 ( 
.A(n_1509),
.Y(n_1542)
);

OAI211xp5_ASAP7_75t_L g1543 ( 
.A1(n_1490),
.A2(n_1453),
.B(n_1470),
.C(n_1467),
.Y(n_1543)
);

INVxp67_ASAP7_75t_L g1544 ( 
.A(n_1504),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_SL g1545 ( 
.A(n_1509),
.B(n_1450),
.Y(n_1545)
);

INVx4_ASAP7_75t_L g1546 ( 
.A(n_1509),
.Y(n_1546)
);

OAI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1515),
.A2(n_1453),
.B(n_1509),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1538),
.Y(n_1548)
);

AOI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1543),
.A2(n_1496),
.B(n_1494),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1538),
.Y(n_1550)
);

OA21x2_ASAP7_75t_L g1551 ( 
.A1(n_1521),
.A2(n_1494),
.B(n_1496),
.Y(n_1551)
);

INVx4_ASAP7_75t_L g1552 ( 
.A(n_1542),
.Y(n_1552)
);

OAI21xp33_ASAP7_75t_L g1553 ( 
.A1(n_1524),
.A2(n_1516),
.B(n_1539),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1532),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1542),
.B(n_1495),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1542),
.Y(n_1556)
);

INVx2_ASAP7_75t_SL g1557 ( 
.A(n_1542),
.Y(n_1557)
);

OA21x2_ASAP7_75t_L g1558 ( 
.A1(n_1536),
.A2(n_1452),
.B(n_1491),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1523),
.B(n_1516),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1537),
.B(n_1501),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1542),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1522),
.B(n_1492),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1537),
.B(n_1501),
.Y(n_1563)
);

NAND3xp33_ASAP7_75t_SL g1564 ( 
.A(n_1523),
.B(n_1419),
.C(n_1461),
.Y(n_1564)
);

NAND3xp33_ASAP7_75t_SL g1565 ( 
.A(n_1524),
.B(n_1419),
.C(n_1512),
.Y(n_1565)
);

INVx4_ASAP7_75t_SL g1566 ( 
.A(n_1534),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1540),
.Y(n_1567)
);

OAI221xp5_ASAP7_75t_L g1568 ( 
.A1(n_1553),
.A2(n_1519),
.B1(n_1525),
.B2(n_1541),
.C(n_1529),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1567),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1556),
.Y(n_1570)
);

AND2x2_ASAP7_75t_SL g1571 ( 
.A(n_1552),
.B(n_1516),
.Y(n_1571)
);

AOI21xp33_ASAP7_75t_L g1572 ( 
.A1(n_1559),
.A2(n_1454),
.B(n_1541),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1560),
.B(n_1518),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1560),
.B(n_1518),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1559),
.B(n_1544),
.Y(n_1575)
);

NAND2xp33_ASAP7_75t_L g1576 ( 
.A(n_1553),
.B(n_1542),
.Y(n_1576)
);

NAND4xp25_ASAP7_75t_L g1577 ( 
.A(n_1559),
.B(n_1531),
.C(n_1546),
.D(n_1530),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1562),
.B(n_1528),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1562),
.B(n_1527),
.Y(n_1579)
);

NOR3xp33_ASAP7_75t_L g1580 ( 
.A(n_1564),
.B(n_1526),
.C(n_1546),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1562),
.B(n_1527),
.Y(n_1581)
);

CKINVDCx16_ASAP7_75t_R g1582 ( 
.A(n_1564),
.Y(n_1582)
);

NAND2xp33_ASAP7_75t_SL g1583 ( 
.A(n_1547),
.B(n_1545),
.Y(n_1583)
);

INVxp67_ASAP7_75t_SL g1584 ( 
.A(n_1548),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1553),
.B(n_1535),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1551),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1567),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1563),
.B(n_1517),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1552),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1563),
.B(n_1517),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1557),
.B(n_1546),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1551),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1557),
.B(n_1546),
.Y(n_1593)
);

AOI221xp5_ASAP7_75t_L g1594 ( 
.A1(n_1564),
.A2(n_1513),
.B1(n_1450),
.B2(n_1533),
.C(n_1520),
.Y(n_1594)
);

NAND3xp33_ASAP7_75t_L g1595 ( 
.A(n_1547),
.B(n_1453),
.C(n_1509),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1556),
.B(n_1503),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1556),
.B(n_1503),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1556),
.B(n_1503),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1554),
.B(n_1535),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1567),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1556),
.B(n_1501),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1551),
.Y(n_1602)
);

NOR2x1_ASAP7_75t_R g1603 ( 
.A(n_1575),
.B(n_1387),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1575),
.B(n_1547),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1570),
.B(n_1566),
.Y(n_1605)
);

INVxp67_ASAP7_75t_L g1606 ( 
.A(n_1571),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1582),
.B(n_1565),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1571),
.B(n_1588),
.Y(n_1608)
);

INVx2_ASAP7_75t_SL g1609 ( 
.A(n_1570),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1569),
.Y(n_1610)
);

INVx2_ASAP7_75t_SL g1611 ( 
.A(n_1570),
.Y(n_1611)
);

INVx1_ASAP7_75t_SL g1612 ( 
.A(n_1571),
.Y(n_1612)
);

AND2x4_ASAP7_75t_L g1613 ( 
.A(n_1588),
.B(n_1566),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1582),
.B(n_1580),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1569),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1573),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1580),
.B(n_1565),
.Y(n_1617)
);

NOR2x1_ASAP7_75t_L g1618 ( 
.A(n_1577),
.B(n_1561),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1588),
.B(n_1590),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1572),
.B(n_1387),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1573),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1587),
.Y(n_1622)
);

NOR2xp67_ASAP7_75t_L g1623 ( 
.A(n_1577),
.B(n_1552),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1585),
.B(n_1565),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1587),
.Y(n_1625)
);

AOI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1576),
.A2(n_1561),
.B(n_1558),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1590),
.B(n_1566),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1585),
.B(n_1578),
.Y(n_1628)
);

O2A1O1Ixp5_ASAP7_75t_L g1629 ( 
.A1(n_1572),
.A2(n_1549),
.B(n_1552),
.C(n_1555),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1590),
.B(n_1566),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1600),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1589),
.Y(n_1632)
);

NAND4xp25_ASAP7_75t_L g1633 ( 
.A(n_1594),
.B(n_1568),
.C(n_1595),
.D(n_1583),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1600),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1599),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1573),
.B(n_1566),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1574),
.B(n_1566),
.Y(n_1637)
);

NAND4xp25_ASAP7_75t_L g1638 ( 
.A(n_1594),
.B(n_1561),
.C(n_1552),
.D(n_1555),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1619),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1616),
.B(n_1578),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1619),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1614),
.B(n_1628),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1610),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1616),
.B(n_1579),
.Y(n_1644)
);

INVx1_ASAP7_75t_SL g1645 ( 
.A(n_1612),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1610),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1609),
.Y(n_1647)
);

AND2x2_ASAP7_75t_SL g1648 ( 
.A(n_1607),
.B(n_1552),
.Y(n_1648)
);

INVx3_ASAP7_75t_L g1649 ( 
.A(n_1613),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1624),
.B(n_1574),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1615),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1615),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1609),
.B(n_1574),
.Y(n_1653)
);

CKINVDCx16_ASAP7_75t_R g1654 ( 
.A(n_1620),
.Y(n_1654)
);

INVx4_ASAP7_75t_L g1655 ( 
.A(n_1605),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1621),
.B(n_1579),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1622),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1633),
.B(n_1568),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1622),
.Y(n_1659)
);

INVx1_ASAP7_75t_SL g1660 ( 
.A(n_1605),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1625),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1611),
.Y(n_1662)
);

OR2x6_ASAP7_75t_L g1663 ( 
.A(n_1611),
.B(n_1552),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1625),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1658),
.B(n_1606),
.Y(n_1665)
);

INVx2_ASAP7_75t_SL g1666 ( 
.A(n_1649),
.Y(n_1666)
);

OAI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1658),
.A2(n_1617),
.B1(n_1618),
.B2(n_1623),
.C(n_1604),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1649),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_SL g1669 ( 
.A1(n_1654),
.A2(n_1595),
.B1(n_1608),
.B2(n_1626),
.Y(n_1669)
);

INVx1_ASAP7_75t_SL g1670 ( 
.A(n_1660),
.Y(n_1670)
);

AOI221xp5_ASAP7_75t_L g1671 ( 
.A1(n_1642),
.A2(n_1629),
.B1(n_1638),
.B2(n_1635),
.C(n_1608),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1639),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1649),
.Y(n_1673)
);

AOI221xp5_ASAP7_75t_L g1674 ( 
.A1(n_1645),
.A2(n_1613),
.B1(n_1605),
.B2(n_1634),
.C(n_1631),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1639),
.Y(n_1675)
);

INVxp67_ASAP7_75t_L g1676 ( 
.A(n_1647),
.Y(n_1676)
);

AOI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1648),
.A2(n_1603),
.B(n_1631),
.Y(n_1677)
);

OAI21xp33_ASAP7_75t_L g1678 ( 
.A1(n_1650),
.A2(n_1637),
.B(n_1636),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1641),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1641),
.B(n_1621),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1643),
.Y(n_1681)
);

AOI221xp5_ASAP7_75t_L g1682 ( 
.A1(n_1662),
.A2(n_1613),
.B1(n_1634),
.B2(n_1636),
.C(n_1637),
.Y(n_1682)
);

AOI21xp33_ASAP7_75t_L g1683 ( 
.A1(n_1648),
.A2(n_1632),
.B(n_1630),
.Y(n_1683)
);

AOI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1662),
.A2(n_1630),
.B1(n_1627),
.B2(n_1558),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1663),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1676),
.B(n_1655),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1676),
.Y(n_1687)
);

INVx2_ASAP7_75t_SL g1688 ( 
.A(n_1666),
.Y(n_1688)
);

INVxp67_ASAP7_75t_L g1689 ( 
.A(n_1668),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1670),
.B(n_1655),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1674),
.B(n_1655),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1673),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1665),
.B(n_1640),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1669),
.A2(n_1627),
.B1(n_1653),
.B2(n_1656),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1678),
.B(n_1663),
.Y(n_1695)
);

INVx2_ASAP7_75t_SL g1696 ( 
.A(n_1680),
.Y(n_1696)
);

NAND5xp2_ASAP7_75t_L g1697 ( 
.A(n_1693),
.B(n_1694),
.C(n_1667),
.D(n_1671),
.E(n_1682),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1692),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1692),
.Y(n_1699)
);

NOR3xp33_ASAP7_75t_SL g1700 ( 
.A(n_1690),
.B(n_1677),
.C(n_1683),
.Y(n_1700)
);

NAND2x1p5_ASAP7_75t_L g1701 ( 
.A(n_1687),
.B(n_1696),
.Y(n_1701)
);

A2O1A1Ixp33_ASAP7_75t_L g1702 ( 
.A1(n_1691),
.A2(n_1669),
.B(n_1677),
.C(n_1684),
.Y(n_1702)
);

NOR4xp25_ASAP7_75t_L g1703 ( 
.A(n_1686),
.B(n_1681),
.C(n_1672),
.D(n_1675),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1689),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1688),
.B(n_1679),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1701),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1701),
.Y(n_1707)
);

AOI221xp5_ASAP7_75t_L g1708 ( 
.A1(n_1702),
.A2(n_1689),
.B1(n_1695),
.B2(n_1684),
.C(n_1685),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1705),
.B(n_1646),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1698),
.Y(n_1710)
);

OAI32xp33_ASAP7_75t_L g1711 ( 
.A1(n_1706),
.A2(n_1699),
.A3(n_1704),
.B1(n_1661),
.B2(n_1659),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1707),
.B(n_1703),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1708),
.B(n_1700),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1710),
.B(n_1651),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1709),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1706),
.B(n_1663),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1716),
.B(n_1663),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1712),
.B(n_1713),
.Y(n_1718)
);

XNOR2xp5_ASAP7_75t_L g1719 ( 
.A(n_1715),
.B(n_1714),
.Y(n_1719)
);

AOI322xp5_ASAP7_75t_L g1720 ( 
.A1(n_1711),
.A2(n_1697),
.A3(n_1664),
.B1(n_1657),
.B2(n_1652),
.C1(n_1584),
.C2(n_1632),
.Y(n_1720)
);

INVx1_ASAP7_75t_SL g1721 ( 
.A(n_1716),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1721),
.A2(n_1640),
.B1(n_1644),
.B2(n_1656),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1720),
.B(n_1717),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_R g1724 ( 
.A(n_1719),
.B(n_1589),
.Y(n_1724)
);

NAND4xp75_ASAP7_75t_L g1725 ( 
.A(n_1723),
.B(n_1718),
.C(n_1724),
.D(n_1722),
.Y(n_1725)
);

AOI322xp5_ASAP7_75t_L g1726 ( 
.A1(n_1725),
.A2(n_1584),
.A3(n_1602),
.B1(n_1592),
.B2(n_1586),
.C1(n_1589),
.C2(n_1550),
.Y(n_1726)
);

OAI31xp33_ASAP7_75t_SL g1727 ( 
.A1(n_1726),
.A2(n_1593),
.A3(n_1591),
.B(n_1592),
.Y(n_1727)
);

AOI221xp5_ASAP7_75t_L g1728 ( 
.A1(n_1726),
.A2(n_1589),
.B1(n_1644),
.B2(n_1591),
.C(n_1593),
.Y(n_1728)
);

OAI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1728),
.A2(n_1593),
.B(n_1591),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1727),
.B(n_1601),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1730),
.Y(n_1731)
);

AOI32xp33_ASAP7_75t_L g1732 ( 
.A1(n_1729),
.A2(n_1561),
.A3(n_1601),
.B1(n_1596),
.B2(n_1597),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1731),
.Y(n_1733)
);

O2A1O1Ixp33_ASAP7_75t_R g1734 ( 
.A1(n_1732),
.A2(n_1602),
.B(n_1586),
.C(n_1592),
.Y(n_1734)
);

OA21x2_ASAP7_75t_L g1735 ( 
.A1(n_1733),
.A2(n_1602),
.B(n_1586),
.Y(n_1735)
);

AOI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1735),
.A2(n_1734),
.B(n_1581),
.Y(n_1736)
);

HB1xp67_ASAP7_75t_L g1737 ( 
.A(n_1736),
.Y(n_1737)
);

AOI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1737),
.A2(n_1601),
.B1(n_1596),
.B2(n_1598),
.Y(n_1738)
);

AOI211xp5_ASAP7_75t_L g1739 ( 
.A1(n_1738),
.A2(n_1596),
.B(n_1598),
.C(n_1597),
.Y(n_1739)
);


endmodule