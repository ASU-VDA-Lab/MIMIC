module fake_jpeg_243_n_160 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_160);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_38),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_22),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_65),
.B(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_68),
.B(n_42),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_57),
.A2(n_47),
.B1(n_41),
.B2(n_53),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_72),
.A2(n_41),
.B1(n_55),
.B2(n_45),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_75),
.B(n_1),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_77),
.Y(n_95)
);

NOR2xp67_ASAP7_75t_SL g77 ( 
.A(n_74),
.B(n_53),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_74),
.A2(n_56),
.B1(n_43),
.B2(n_46),
.Y(n_78)
);

MAJx2_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_80),
.C(n_66),
.Y(n_94)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_49),
.B1(n_44),
.B2(n_52),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_41),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_84),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_64),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_86),
.B1(n_67),
.B2(n_3),
.Y(n_105)
);

OAI22x1_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_55),
.B1(n_45),
.B2(n_17),
.Y(n_86)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_88),
.B(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_70),
.Y(n_90)
);

INVxp33_ASAP7_75t_SL g93 ( 
.A(n_80),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_100),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_105),
.Y(n_111)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_87),
.Y(n_100)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_83),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_4),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_78),
.B(n_2),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_104),
.B(n_5),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_67),
.C(n_19),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_33),
.C(n_32),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_86),
.B1(n_16),
.B2(n_21),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_113),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_114),
.B(n_123),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_24),
.B1(n_39),
.B2(n_37),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_115),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_139)
);

AOI22x1_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_40),
.B1(n_35),
.B2(n_34),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_116),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_124),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_102),
.A2(n_5),
.B(n_6),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_118),
.A2(n_107),
.B(n_10),
.Y(n_128)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_121),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_6),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_7),
.B(n_9),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_122),
.A2(n_11),
.B(n_12),
.Y(n_134)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_92),
.Y(n_127)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_128),
.B(n_129),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_101),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_106),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_134),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_131),
.B(n_138),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_28),
.B(n_26),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_133),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_25),
.Y(n_138)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

AOI322xp5_ASAP7_75t_L g140 ( 
.A1(n_136),
.A2(n_118),
.A3(n_115),
.B1(n_116),
.B2(n_110),
.C1(n_122),
.C2(n_108),
.Y(n_140)
);

AOI321xp33_ASAP7_75t_L g148 ( 
.A1(n_140),
.A2(n_138),
.A3(n_126),
.B1(n_130),
.B2(n_132),
.C(n_129),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_137),
.B1(n_136),
.B2(n_135),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_149),
.B1(n_150),
.B2(n_146),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_148),
.B(n_144),
.C(n_143),
.Y(n_151)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_145),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

AOI211xp5_ASAP7_75t_SL g153 ( 
.A1(n_151),
.A2(n_152),
.B(n_148),
.C(n_146),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_119),
.B(n_141),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_13),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_157),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_124),
.C(n_14),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_15),
.Y(n_160)
);


endmodule