module fake_jpeg_5061_n_274 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_274);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx11_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_25),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_30),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

CKINVDCx12_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_42),
.B(n_54),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_44),
.Y(n_75)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_49),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_24),
.B1(n_15),
.B2(n_26),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_50),
.A2(n_24),
.B1(n_15),
.B2(n_26),
.Y(n_67)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_32),
.Y(n_52)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_33),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_23),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_21),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_56),
.B(n_18),
.Y(n_69)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_24),
.B1(n_19),
.B2(n_25),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_63),
.A2(n_64),
.B1(n_19),
.B2(n_23),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_24),
.B1(n_15),
.B2(n_31),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_67),
.A2(n_82),
.B1(n_85),
.B2(n_87),
.Y(n_99)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_69),
.Y(n_107)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_27),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_29),
.C(n_20),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_60),
.B(n_25),
.Y(n_72)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_23),
.Y(n_73)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_30),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_78),
.B1(n_87),
.B2(n_58),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_60),
.A2(n_19),
.B1(n_31),
.B2(n_16),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_50),
.A2(n_31),
.B1(n_16),
.B2(n_21),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_86),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_64),
.A2(n_16),
.B1(n_20),
.B2(n_40),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_88),
.B(n_89),
.Y(n_126)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_79),
.A2(n_20),
.B(n_51),
.C(n_58),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_90),
.A2(n_103),
.B1(n_28),
.B2(n_65),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_21),
.B(n_17),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_91),
.A2(n_93),
.B(n_84),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_98),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_71),
.A2(n_20),
.B(n_26),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_49),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_100),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_29),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_49),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_67),
.A2(n_51),
.B1(n_61),
.B2(n_53),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_102),
.A2(n_111),
.B1(n_86),
.B2(n_70),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_42),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_49),
.Y(n_104)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_29),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_105),
.B(n_68),
.Y(n_115)
);

MAJx2_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_41),
.C(n_40),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_106),
.A2(n_108),
.B(n_22),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_77),
.A2(n_46),
.B1(n_53),
.B2(n_20),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_113),
.A2(n_118),
.B1(n_122),
.B2(n_135),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_104),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_115),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_101),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_116),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_90),
.A2(n_46),
.B1(n_66),
.B2(n_83),
.Y(n_118)
);

O2A1O1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_66),
.B(n_22),
.C(n_28),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_119),
.A2(n_124),
.B(n_110),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_133),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_105),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_121),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_94),
.A2(n_22),
.B1(n_28),
.B2(n_59),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_128),
.Y(n_152)
);

HAxp5_ASAP7_75t_SL g125 ( 
.A(n_92),
.B(n_41),
.CON(n_125),
.SN(n_125)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_125),
.A2(n_109),
.B1(n_97),
.B2(n_99),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_41),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_127),
.A2(n_129),
.B(n_91),
.Y(n_148)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_93),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_100),
.A2(n_62),
.B1(n_59),
.B2(n_48),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_112),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_153),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_108),
.C(n_103),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_117),
.Y(n_164)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_140),
.B(n_144),
.Y(n_161)
);

INVxp67_ASAP7_75t_SL g141 ( 
.A(n_116),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_141),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_142),
.A2(n_148),
.B(n_149),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_115),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_143),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_135),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_150),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_110),
.B(n_107),
.Y(n_149)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_121),
.B(n_109),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_118),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_154),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_97),
.B1(n_88),
.B2(n_74),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_134),
.B1(n_124),
.B2(n_127),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_96),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_158),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_129),
.A2(n_62),
.B1(n_59),
.B2(n_48),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_159),
.A2(n_122),
.B1(n_119),
.B2(n_113),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_163),
.A2(n_159),
.B1(n_169),
.B2(n_145),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_172),
.Y(n_201)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_166),
.Y(n_200)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_173),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_120),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_182),
.Y(n_187)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_180),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_130),
.Y(n_176)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_136),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_178),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_154),
.A2(n_130),
.B1(n_127),
.B2(n_132),
.Y(n_179)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_136),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_181),
.A2(n_153),
.B(n_140),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_130),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_139),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_186),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_185),
.A2(n_167),
.B1(n_74),
.B2(n_65),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_148),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_142),
.C(n_150),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_189),
.C(n_161),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_149),
.C(n_157),
.Y(n_189)
);

FAx1_ASAP7_75t_SL g190 ( 
.A(n_176),
.B(n_157),
.CI(n_151),
.CON(n_190),
.SN(n_190)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_198),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_151),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_192),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_172),
.Y(n_192)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_194),
.Y(n_203)
);

AOI21x1_ASAP7_75t_SL g197 ( 
.A1(n_170),
.A2(n_132),
.B(n_138),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_177),
.Y(n_217)
);

AND2x6_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_138),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_174),
.Y(n_215)
);

AOI21x1_ASAP7_75t_L g202 ( 
.A1(n_173),
.A2(n_28),
.B(n_0),
.Y(n_202)
);

FAx1_ASAP7_75t_SL g214 ( 
.A(n_202),
.B(n_197),
.CI(n_191),
.CON(n_214),
.SN(n_214)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_200),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_204),
.B(n_207),
.Y(n_228)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_209),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_196),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_162),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_208),
.A2(n_211),
.B(n_212),
.Y(n_221)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_198),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_216),
.C(n_188),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_193),
.A2(n_177),
.B(n_160),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_192),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_217),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_187),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_180),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_189),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_223),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_210),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_183),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_214),
.C(n_217),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_187),
.C(n_199),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_2),
.C(n_3),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_186),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_232),
.Y(n_240)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_214),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_205),
.A2(n_96),
.B1(n_0),
.B2(n_2),
.Y(n_231)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_231),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_7),
.Y(n_232)
);

XNOR2x1_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_0),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_233),
.A2(n_226),
.B(n_232),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_224),
.A2(n_221),
.B(n_203),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_234),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_238),
.C(n_239),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_227),
.A2(n_211),
.B(n_208),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_241),
.B(n_6),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_242),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_233),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_1),
.C(n_2),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_245),
.C(n_240),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_254),
.Y(n_257)
);

NOR2xp67_ASAP7_75t_SL g247 ( 
.A(n_237),
.B(n_226),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_247),
.A2(n_235),
.B(n_9),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_236),
.A2(n_229),
.B1(n_4),
.B2(n_5),
.Y(n_248)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_248),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_253),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_9),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_8),
.Y(n_254)
);

NOR3xp33_ASAP7_75t_SL g255 ( 
.A(n_246),
.B(n_240),
.C(n_245),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_256),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_8),
.Y(n_258)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_258),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_254),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_251),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_10),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_248),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_264),
.A2(n_258),
.B(n_11),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_266),
.B(n_260),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_269),
.C(n_262),
.Y(n_271)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_268),
.Y(n_270)
);

AOI322xp5_ASAP7_75t_L g272 ( 
.A1(n_271),
.A2(n_10),
.A3(n_13),
.B1(n_14),
.B2(n_264),
.C1(n_265),
.C2(n_270),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_272),
.A2(n_13),
.B(n_14),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_14),
.Y(n_274)
);


endmodule