module fake_ariane_217_n_2082 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2082);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2082;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_851;
wire n_444;
wire n_355;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_1083;
wire n_967;
wire n_274;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_330;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_SL g217 ( 
.A(n_77),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_28),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_173),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g221 ( 
.A(n_89),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_75),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_39),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_215),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_66),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_29),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_183),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_209),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_80),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_94),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_133),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_129),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_40),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_162),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_163),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_193),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_41),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_45),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_63),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_78),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_8),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_154),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_169),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_196),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_17),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_14),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_138),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_188),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_167),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_24),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_132),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_126),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_13),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_55),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_56),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_69),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_176),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_46),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_185),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_78),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_187),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_145),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_84),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_204),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_125),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_192),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_112),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_110),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_165),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_120),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_127),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_135),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_85),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_123),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_208),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_121),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_38),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_113),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_40),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_106),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_51),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_1),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_157),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_118),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_102),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_137),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_142),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_92),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_8),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_195),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_26),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_213),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_31),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_26),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_19),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_97),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_49),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_203),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_148),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_105),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_13),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_115),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_41),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_45),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_70),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_172),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_131),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_214),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_72),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_122),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_156),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_11),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_15),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_87),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_206),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_60),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_216),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_47),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_75),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_7),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_55),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_91),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_66),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_202),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_34),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_60),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_7),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_63),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_68),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_117),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_152),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_80),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_17),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_199),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_99),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_1),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_61),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_168),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_134),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_68),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_151),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_210),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_205),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_10),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_130),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_73),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_171),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_82),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_181),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_70),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_101),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_48),
.Y(n_352)
);

INVxp33_ASAP7_75t_L g353 ( 
.A(n_170),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_109),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_24),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_27),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_150),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_95),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_149),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_0),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_124),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_43),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_31),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_54),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_155),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_107),
.Y(n_366)
);

BUFx5_ASAP7_75t_L g367 ( 
.A(n_56),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_175),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_161),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_212),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_49),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_19),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_178),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_25),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_39),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_81),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_62),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_0),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_180),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_86),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_194),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_57),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_27),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_81),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_20),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_12),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_116),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_108),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_90),
.Y(n_389)
);

CKINVDCx14_ASAP7_75t_R g390 ( 
.A(n_174),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_33),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_186),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_82),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_25),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_11),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_207),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_184),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_3),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_160),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_32),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_198),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_51),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_37),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_141),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_103),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_189),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_211),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_54),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_76),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_65),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_21),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_111),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_43),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_164),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_197),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_2),
.Y(n_416)
);

BUFx10_ASAP7_75t_L g417 ( 
.A(n_65),
.Y(n_417)
);

INVx2_ASAP7_75t_SL g418 ( 
.A(n_50),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_158),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_139),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_16),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_79),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_22),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_29),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_36),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_146),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_61),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_367),
.Y(n_428)
);

NOR2xp67_ASAP7_75t_L g429 ( 
.A(n_352),
.B(n_2),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_264),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_270),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_346),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_290),
.Y(n_433)
);

CKINVDCx14_ASAP7_75t_R g434 ( 
.A(n_390),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_381),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_367),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_367),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_389),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_367),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_367),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_397),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_426),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_367),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_346),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_333),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_416),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_333),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_416),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_280),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_367),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_225),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_294),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_294),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_222),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_293),
.B(n_3),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_237),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_380),
.B(n_4),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_233),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_238),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_367),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_239),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_367),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_240),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_291),
.Y(n_464)
);

NOR2xp67_ASAP7_75t_L g465 ( 
.A(n_352),
.B(n_4),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_219),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_332),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_380),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_241),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_219),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_220),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_411),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_280),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_220),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_231),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_231),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_234),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_246),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_269),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_234),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_236),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_236),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_243),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_269),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_250),
.Y(n_485)
);

INVxp67_ASAP7_75t_SL g486 ( 
.A(n_233),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_218),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_243),
.B(n_5),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_375),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_280),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_247),
.Y(n_491)
);

NOR2xp67_ASAP7_75t_L g492 ( 
.A(n_418),
.B(n_5),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_256),
.B(n_6),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_247),
.B(n_6),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_260),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_R g496 ( 
.A(n_227),
.B(n_83),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_233),
.B(n_9),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_281),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g499 ( 
.A(n_375),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_248),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_282),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_248),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_261),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_295),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_261),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_304),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_218),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_267),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_418),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_305),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_309),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_267),
.Y(n_512)
);

NOR2xp67_ASAP7_75t_L g513 ( 
.A(n_293),
.B(n_9),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_268),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_299),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_268),
.B(n_10),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_271),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_312),
.Y(n_518)
);

BUFx10_ASAP7_75t_L g519 ( 
.A(n_224),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_313),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_299),
.Y(n_521)
);

INVxp67_ASAP7_75t_SL g522 ( 
.A(n_223),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_299),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_271),
.B(n_12),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_272),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_272),
.B(n_14),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_275),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_316),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_275),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_284),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_318),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_284),
.Y(n_532)
);

INVxp67_ASAP7_75t_SL g533 ( 
.A(n_223),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_320),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_298),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_298),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_257),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_321),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_473),
.B(n_306),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_432),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_473),
.B(n_306),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_466),
.B(n_336),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_453),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_428),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_466),
.B(n_307),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_428),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_430),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_436),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_436),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_470),
.B(n_307),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_449),
.Y(n_551)
);

CKINVDCx8_ASAP7_75t_R g552 ( 
.A(n_431),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_437),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_458),
.B(n_486),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_437),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_439),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_439),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_440),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_440),
.Y(n_559)
);

CKINVDCx8_ASAP7_75t_R g560 ( 
.A(n_441),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_443),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_479),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_470),
.B(n_336),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_443),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_444),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_471),
.B(n_363),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_471),
.B(n_363),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_450),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_450),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_460),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_460),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_446),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_457),
.B(n_353),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_448),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_462),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_462),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_474),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_449),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_474),
.B(n_376),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_497),
.B(n_376),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_475),
.B(n_311),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_475),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_476),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_449),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_449),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_476),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_477),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_449),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_477),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_480),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_480),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_481),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_481),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_484),
.A2(n_245),
.B1(n_254),
.B2(n_217),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_482),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_482),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_445),
.Y(n_597)
);

BUFx8_ASAP7_75t_L g598 ( 
.A(n_509),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_454),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_483),
.B(n_257),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_483),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_497),
.B(n_257),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_491),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_491),
.Y(n_604)
);

OA21x2_ASAP7_75t_L g605 ( 
.A1(n_500),
.A2(n_314),
.B(n_311),
.Y(n_605)
);

AND2x6_ASAP7_75t_L g606 ( 
.A(n_500),
.B(n_252),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_502),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_502),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_503),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_503),
.B(n_314),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_505),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_505),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_508),
.Y(n_613)
);

AND2x6_ASAP7_75t_L g614 ( 
.A(n_508),
.B(n_252),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_512),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_512),
.B(n_322),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_514),
.B(n_257),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_514),
.Y(n_618)
);

NAND2x1p5_ASAP7_75t_L g619 ( 
.A(n_455),
.B(n_266),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_517),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_517),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_525),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_447),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_525),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_527),
.B(n_226),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_527),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_603),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_603),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_600),
.B(n_617),
.Y(n_629)
);

OAI22xp33_ASAP7_75t_L g630 ( 
.A1(n_619),
.A2(n_468),
.B1(n_455),
.B2(n_509),
.Y(n_630)
);

BUFx2_ASAP7_75t_L g631 ( 
.A(n_540),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_600),
.B(n_434),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_603),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_619),
.A2(n_468),
.B1(n_494),
.B2(n_488),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_573),
.B(n_456),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_603),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_551),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_603),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_600),
.B(n_617),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_599),
.B(n_459),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_606),
.Y(n_641)
);

CKINVDCx20_ASAP7_75t_R g642 ( 
.A(n_547),
.Y(n_642)
);

INVxp67_ASAP7_75t_SL g643 ( 
.A(n_596),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_544),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_603),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_603),
.Y(n_646)
);

INVx4_ASAP7_75t_L g647 ( 
.A(n_606),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_603),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_619),
.A2(n_524),
.B1(n_526),
.B2(n_516),
.Y(n_649)
);

HB1xp67_ASAP7_75t_L g650 ( 
.A(n_540),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_619),
.A2(n_515),
.B1(n_521),
.B2(n_490),
.Y(n_651)
);

INVx8_ASAP7_75t_L g652 ( 
.A(n_606),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_617),
.B(n_522),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_544),
.Y(n_654)
);

INVx4_ASAP7_75t_L g655 ( 
.A(n_606),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_606),
.Y(n_656)
);

INVxp67_ASAP7_75t_SL g657 ( 
.A(n_596),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_SL g658 ( 
.A1(n_598),
.A2(n_594),
.B1(n_537),
.B2(n_523),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_608),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_608),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g661 ( 
.A(n_599),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_608),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_608),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_619),
.A2(n_465),
.B1(n_492),
.B2(n_429),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_608),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_544),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_551),
.Y(n_667)
);

BUFx8_ASAP7_75t_SL g668 ( 
.A(n_547),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_556),
.Y(n_669)
);

BUFx2_ASAP7_75t_L g670 ( 
.A(n_598),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_554),
.B(n_519),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_551),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_573),
.B(n_461),
.Y(n_673)
);

INVx5_ASAP7_75t_L g674 ( 
.A(n_606),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_608),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_608),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_598),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_556),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g679 ( 
.A1(n_602),
.A2(n_327),
.B1(n_328),
.B2(n_326),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_608),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_556),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_599),
.B(n_463),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_577),
.Y(n_683)
);

AND2x6_ASAP7_75t_L g684 ( 
.A(n_580),
.B(n_322),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_556),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_558),
.Y(n_686)
);

NAND2x1p5_ASAP7_75t_L g687 ( 
.A(n_605),
.B(n_529),
.Y(n_687)
);

AND2x2_ASAP7_75t_SL g688 ( 
.A(n_605),
.B(n_263),
.Y(n_688)
);

INVx4_ASAP7_75t_L g689 ( 
.A(n_606),
.Y(n_689)
);

BUFx4f_ASAP7_75t_L g690 ( 
.A(n_605),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_558),
.Y(n_691)
);

INVx4_ASAP7_75t_L g692 ( 
.A(n_606),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_558),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_554),
.B(n_469),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_551),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_582),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_582),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_558),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_546),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_604),
.B(n_519),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_604),
.B(n_519),
.Y(n_701)
);

NAND2xp33_ASAP7_75t_L g702 ( 
.A(n_583),
.B(n_478),
.Y(n_702)
);

NOR3xp33_ASAP7_75t_L g703 ( 
.A(n_565),
.B(n_495),
.C(n_485),
.Y(n_703)
);

BUFx10_ASAP7_75t_L g704 ( 
.A(n_580),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_602),
.B(n_498),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_569),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_598),
.B(n_501),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_598),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_552),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_580),
.A2(n_529),
.B1(n_532),
.B2(n_530),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_569),
.Y(n_711)
);

CKINVDCx6p67_ASAP7_75t_R g712 ( 
.A(n_562),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_604),
.B(n_519),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_543),
.B(n_504),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_580),
.A2(n_530),
.B1(n_535),
.B2(n_532),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_604),
.B(n_535),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_552),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_569),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_546),
.Y(n_719)
);

BUFx10_ASAP7_75t_L g720 ( 
.A(n_580),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_580),
.B(n_536),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_569),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_571),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_597),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_583),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_583),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_606),
.A2(n_536),
.B1(n_513),
.B2(n_533),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_598),
.B(n_506),
.Y(n_728)
);

NAND2xp33_ASAP7_75t_L g729 ( 
.A(n_586),
.B(n_510),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_546),
.Y(n_730)
);

AND2x6_ASAP7_75t_L g731 ( 
.A(n_586),
.B(n_324),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_542),
.B(n_499),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_571),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_543),
.B(n_511),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_571),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_606),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_546),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_586),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_546),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_594),
.A2(n_337),
.B1(n_493),
.B2(n_344),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_597),
.B(n_442),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_623),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_591),
.Y(n_743)
);

INVxp67_ASAP7_75t_SL g744 ( 
.A(n_596),
.Y(n_744)
);

BUFx2_ASAP7_75t_L g745 ( 
.A(n_623),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_562),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_571),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_576),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_552),
.Y(n_749)
);

INVx4_ASAP7_75t_L g750 ( 
.A(n_606),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_546),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_565),
.B(n_518),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_591),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_572),
.B(n_520),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_587),
.B(n_528),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_560),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_625),
.B(n_452),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_548),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_591),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_572),
.B(n_531),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_576),
.Y(n_761)
);

INVx1_ASAP7_75t_SL g762 ( 
.A(n_574),
.Y(n_762)
);

AND2x6_ASAP7_75t_L g763 ( 
.A(n_593),
.B(n_324),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_576),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_587),
.B(n_534),
.Y(n_765)
);

AND3x2_ASAP7_75t_L g766 ( 
.A(n_574),
.B(n_452),
.C(n_489),
.Y(n_766)
);

OR2x6_ASAP7_75t_L g767 ( 
.A(n_625),
.B(n_487),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_605),
.Y(n_768)
);

HAxp5_ASAP7_75t_SL g769 ( 
.A(n_560),
.B(n_493),
.CON(n_769),
.SN(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_596),
.B(n_538),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_593),
.Y(n_771)
);

AND2x2_ASAP7_75t_SL g772 ( 
.A(n_605),
.B(n_263),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_593),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_595),
.Y(n_774)
);

INVx3_ASAP7_75t_L g775 ( 
.A(n_546),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_596),
.B(n_417),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_542),
.B(n_507),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_690),
.B(n_548),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_762),
.B(n_661),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_629),
.B(n_595),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_688),
.A2(n_605),
.B1(n_614),
.B2(n_590),
.Y(n_781)
);

INVxp67_ASAP7_75t_L g782 ( 
.A(n_631),
.Y(n_782)
);

NOR2xp67_ASAP7_75t_L g783 ( 
.A(n_714),
.B(n_545),
.Y(n_783)
);

INVx4_ASAP7_75t_L g784 ( 
.A(n_652),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_746),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_683),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_629),
.B(n_595),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_705),
.B(n_560),
.Y(n_788)
);

O2A1O1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_639),
.A2(n_548),
.B(n_553),
.C(n_549),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_694),
.B(n_601),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_755),
.B(n_601),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_635),
.A2(n_614),
.B1(n_589),
.B2(n_611),
.Y(n_792)
);

NAND2x1_ASAP7_75t_L g793 ( 
.A(n_641),
.B(n_601),
.Y(n_793)
);

OAI221xp5_ASAP7_75t_L g794 ( 
.A1(n_634),
.A2(n_289),
.B1(n_297),
.B2(n_279),
.C(n_301),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_765),
.B(n_611),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_673),
.B(n_539),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_653),
.B(n_611),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_653),
.B(n_612),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_630),
.B(n_612),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_666),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_666),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_653),
.B(n_612),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_653),
.B(n_615),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_684),
.A2(n_614),
.B1(n_589),
.B2(n_615),
.Y(n_804)
);

OAI22xp33_ASAP7_75t_L g805 ( 
.A1(n_767),
.A2(n_550),
.B1(n_581),
.B2(n_545),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_671),
.B(n_643),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_657),
.B(n_615),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_688),
.A2(n_614),
.B1(n_592),
.B2(n_607),
.Y(n_808)
);

BUFx6f_ASAP7_75t_SL g809 ( 
.A(n_757),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_770),
.B(n_632),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_744),
.B(n_732),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_767),
.B(n_539),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_732),
.B(n_621),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_710),
.B(n_621),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_715),
.B(n_664),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_649),
.B(n_621),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_721),
.B(n_624),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_631),
.Y(n_818)
);

INVx8_ASAP7_75t_L g819 ( 
.A(n_652),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_691),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_691),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_691),
.Y(n_822)
);

BUFx6f_ASAP7_75t_SL g823 ( 
.A(n_757),
.Y(n_823)
);

NAND2xp33_ASAP7_75t_L g824 ( 
.A(n_731),
.B(n_549),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_704),
.B(n_624),
.Y(n_825)
);

INVxp33_ASAP7_75t_L g826 ( 
.A(n_741),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_767),
.B(n_541),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_767),
.B(n_541),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_684),
.B(n_624),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_693),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_693),
.Y(n_831)
);

INVxp67_ASAP7_75t_L g832 ( 
.A(n_741),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_684),
.B(n_626),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_767),
.B(n_555),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_693),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_684),
.A2(n_614),
.B1(n_626),
.B2(n_625),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_684),
.B(n_626),
.Y(n_837)
);

BUFx6f_ASAP7_75t_SL g838 ( 
.A(n_757),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_668),
.Y(n_839)
);

BUFx6f_ASAP7_75t_SL g840 ( 
.A(n_757),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_684),
.B(n_555),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_696),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_688),
.A2(n_614),
.B1(n_592),
.B2(n_607),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_745),
.B(n_542),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_704),
.B(n_720),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_690),
.B(n_641),
.Y(n_846)
);

NAND3xp33_ASAP7_75t_L g847 ( 
.A(n_702),
.B(n_553),
.C(n_549),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_704),
.B(n_553),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_722),
.Y(n_849)
);

O2A1O1Ixp33_ASAP7_75t_L g850 ( 
.A1(n_716),
.A2(n_559),
.B(n_568),
.C(n_561),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_697),
.Y(n_851)
);

INVxp67_ASAP7_75t_L g852 ( 
.A(n_745),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_704),
.B(n_559),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_697),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_772),
.A2(n_614),
.B1(n_592),
.B2(n_607),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_772),
.A2(n_614),
.B1(n_592),
.B2(n_607),
.Y(n_856)
);

INVx8_ASAP7_75t_L g857 ( 
.A(n_652),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_684),
.B(n_559),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_777),
.B(n_561),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_777),
.B(n_561),
.Y(n_860)
);

AND2x4_ASAP7_75t_L g861 ( 
.A(n_670),
.B(n_563),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_690),
.B(n_568),
.Y(n_862)
);

BUFx5_ASAP7_75t_L g863 ( 
.A(n_758),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_720),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_725),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_758),
.B(n_568),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_720),
.B(n_776),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_772),
.A2(n_614),
.B1(n_609),
.B2(n_613),
.Y(n_868)
);

BUFx6f_ASAP7_75t_SL g869 ( 
.A(n_642),
.Y(n_869)
);

NOR2xp67_ASAP7_75t_L g870 ( 
.A(n_709),
.B(n_550),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_650),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_722),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_758),
.B(n_720),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_725),
.B(n_570),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_724),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_729),
.B(n_570),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_726),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_726),
.B(n_570),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_738),
.B(n_575),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_712),
.B(n_563),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_637),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_652),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_734),
.B(n_575),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_637),
.Y(n_884)
);

NOR3xp33_ASAP7_75t_L g885 ( 
.A(n_640),
.B(n_229),
.C(n_226),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_707),
.A2(n_614),
.B1(n_566),
.B2(n_567),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_738),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_731),
.A2(n_614),
.B1(n_590),
.B2(n_613),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_652),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_637),
.Y(n_890)
);

NAND3xp33_ASAP7_75t_L g891 ( 
.A(n_703),
.B(n_575),
.C(n_581),
.Y(n_891)
);

NOR3xp33_ASAP7_75t_L g892 ( 
.A(n_682),
.B(n_253),
.C(n_229),
.Y(n_892)
);

NAND2x1p5_ASAP7_75t_L g893 ( 
.A(n_670),
.B(n_590),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_722),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_667),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_641),
.B(n_576),
.Y(n_896)
);

INVxp67_ASAP7_75t_L g897 ( 
.A(n_742),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_667),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_747),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_743),
.B(n_590),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_743),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_731),
.A2(n_613),
.B1(n_618),
.B2(n_609),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_SL g903 ( 
.A(n_717),
.B(n_433),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_747),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_747),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_749),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_677),
.B(n_708),
.Y(n_907)
);

NOR2xp67_ASAP7_75t_L g908 ( 
.A(n_728),
.B(n_610),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_677),
.B(n_563),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_700),
.A2(n_610),
.B1(n_616),
.B2(n_613),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_753),
.B(n_609),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_701),
.B(n_713),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_753),
.B(n_609),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_667),
.Y(n_914)
);

INVx8_ASAP7_75t_L g915 ( 
.A(n_674),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_759),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_752),
.B(n_616),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_712),
.Y(n_918)
);

NAND2xp33_ASAP7_75t_SL g919 ( 
.A(n_708),
.B(n_618),
.Y(n_919)
);

INVxp33_ASAP7_75t_L g920 ( 
.A(n_754),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_760),
.B(n_618),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_641),
.B(n_546),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_759),
.A2(n_620),
.B(n_622),
.C(n_618),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_771),
.A2(n_622),
.B(n_620),
.C(n_253),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_771),
.B(n_620),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_748),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_672),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_647),
.B(n_557),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_773),
.Y(n_929)
);

INVx4_ASAP7_75t_L g930 ( 
.A(n_647),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_748),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_748),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_773),
.B(n_620),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_774),
.B(n_622),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_774),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_647),
.B(n_557),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_687),
.B(n_622),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_796),
.B(n_727),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_796),
.B(n_687),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_786),
.Y(n_940)
);

OAI21xp33_ASAP7_75t_L g941 ( 
.A1(n_790),
.A2(n_679),
.B(n_740),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_890),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_783),
.B(n_687),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_810),
.B(n_651),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_778),
.A2(n_768),
.B(n_739),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_810),
.A2(n_654),
.B(n_669),
.C(n_644),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_L g947 ( 
.A1(n_791),
.A2(n_768),
.B1(n_655),
.B2(n_656),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_917),
.B(n_812),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_778),
.A2(n_739),
.B(n_719),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_917),
.B(n_731),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_870),
.B(n_647),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_862),
.A2(n_912),
.B(n_876),
.Y(n_952)
);

NAND2x1p5_ASAP7_75t_L g953 ( 
.A(n_881),
.B(n_674),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_862),
.A2(n_739),
.B(n_719),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_912),
.A2(n_739),
.B(n_719),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_812),
.B(n_731),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_779),
.B(n_740),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_863),
.B(n_699),
.Y(n_958)
);

CKINVDCx20_ASAP7_75t_R g959 ( 
.A(n_839),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_937),
.A2(n_654),
.B(n_644),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_890),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_881),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_896),
.A2(n_678),
.B(n_669),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_844),
.B(n_658),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_805),
.A2(n_681),
.B(n_685),
.C(n_678),
.Y(n_965)
);

NOR2x1p5_ASAP7_75t_SL g966 ( 
.A(n_863),
.B(n_628),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_876),
.A2(n_775),
.B(n_719),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_795),
.A2(n_685),
.B(n_686),
.C(n_681),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_806),
.A2(n_775),
.B(n_698),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_818),
.Y(n_970)
);

AOI21x1_ASAP7_75t_L g971 ( 
.A1(n_874),
.A2(n_633),
.B(n_628),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_848),
.A2(n_656),
.B1(n_689),
.B2(n_655),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_827),
.B(n_731),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_827),
.B(n_731),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_828),
.B(n_763),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_914),
.Y(n_976)
);

OAI21xp5_ASAP7_75t_L g977 ( 
.A1(n_896),
.A2(n_698),
.B(n_686),
.Y(n_977)
);

BUFx3_ASAP7_75t_L g978 ( 
.A(n_785),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_811),
.B(n_756),
.Y(n_979)
);

AOI22xp5_ASAP7_75t_L g980 ( 
.A1(n_828),
.A2(n_763),
.B1(n_438),
.B2(n_435),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_859),
.B(n_763),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_860),
.B(n_763),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_832),
.B(n_775),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_883),
.A2(n_711),
.B(n_718),
.C(n_706),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_922),
.A2(n_775),
.B(n_711),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_922),
.A2(n_718),
.B(n_706),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_813),
.B(n_763),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_883),
.B(n_763),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_863),
.B(n_699),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_928),
.A2(n_733),
.B(n_723),
.Y(n_990)
);

CKINVDCx10_ASAP7_75t_R g991 ( 
.A(n_869),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_834),
.B(n_763),
.Y(n_992)
);

AOI33xp33_ASAP7_75t_L g993 ( 
.A1(n_871),
.A2(n_255),
.A3(n_427),
.B1(n_258),
.B2(n_277),
.B3(n_279),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_928),
.A2(n_733),
.B(n_723),
.Y(n_994)
);

AOI21xp33_ASAP7_75t_L g995 ( 
.A1(n_826),
.A2(n_761),
.B(n_735),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_936),
.A2(n_764),
.B(n_638),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_864),
.B(n_655),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_936),
.A2(n_638),
.B(n_633),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_853),
.A2(n_646),
.B(n_645),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_852),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_863),
.B(n_699),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_834),
.B(n_566),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_780),
.A2(n_255),
.B(n_277),
.C(n_258),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_797),
.B(n_566),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_861),
.B(n_909),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_853),
.A2(n_646),
.B(n_645),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_788),
.B(n_672),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_878),
.A2(n_659),
.B(n_648),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_879),
.A2(n_866),
.B(n_900),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_787),
.A2(n_289),
.B(n_301),
.C(n_297),
.Y(n_1010)
);

BUFx2_ASAP7_75t_SL g1011 ( 
.A(n_869),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_911),
.A2(n_925),
.B(n_913),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_809),
.A2(n_823),
.B1(n_840),
.B2(n_838),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_798),
.A2(n_303),
.B(n_323),
.C(n_319),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_890),
.Y(n_1015)
);

INVx4_ASAP7_75t_L g1016 ( 
.A(n_819),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_782),
.B(n_451),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_933),
.A2(n_659),
.B(n_648),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_934),
.A2(n_662),
.B(n_660),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_802),
.B(n_803),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_863),
.B(n_699),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_861),
.B(n_567),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_807),
.A2(n_662),
.B(n_660),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_793),
.A2(n_665),
.B(n_663),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_909),
.B(n_567),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_921),
.B(n_579),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_921),
.B(n_579),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_930),
.A2(n_665),
.B(n_663),
.Y(n_1028)
);

CKINVDCx8_ASAP7_75t_R g1029 ( 
.A(n_906),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_930),
.A2(n_675),
.B(n_656),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_842),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_867),
.A2(n_636),
.B(n_676),
.C(n_627),
.Y(n_1032)
);

INVx11_ASAP7_75t_L g1033 ( 
.A(n_903),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_873),
.A2(n_675),
.B(n_656),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_920),
.B(n_672),
.Y(n_1035)
);

OAI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_923),
.A2(n_636),
.B(n_627),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_891),
.B(n_695),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_824),
.A2(n_689),
.B(n_655),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_815),
.B(n_579),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_908),
.B(n_695),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_799),
.B(n_695),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_867),
.A2(n_636),
.B(n_676),
.C(n_627),
.Y(n_1042)
);

INVx4_ASAP7_75t_L g1043 ( 
.A(n_819),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_817),
.A2(n_303),
.B(n_323),
.C(n_319),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_910),
.A2(n_692),
.B(n_689),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_851),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_880),
.B(n_627),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_854),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_816),
.A2(n_676),
.B(n_636),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_825),
.A2(n_692),
.B(n_689),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_846),
.A2(n_736),
.B(n_692),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_846),
.A2(n_736),
.B(n_692),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_865),
.A2(n_750),
.B1(n_736),
.B2(n_680),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_800),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_918),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_877),
.B(n_676),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_800),
.A2(n_750),
.B(n_736),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_887),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_901),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_809),
.B(n_680),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_916),
.B(n_680),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_801),
.A2(n_750),
.B(n_680),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_823),
.A2(n_750),
.B1(n_699),
.B2(n_751),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_801),
.A2(n_737),
.B(n_730),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_820),
.A2(n_737),
.B(n_730),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_820),
.A2(n_737),
.B(n_730),
.Y(n_1066)
);

O2A1O1Ixp5_ASAP7_75t_L g1067 ( 
.A1(n_829),
.A2(n_585),
.B(n_588),
.C(n_578),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_821),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_838),
.B(n_766),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_850),
.A2(n_674),
.B(n_588),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_821),
.A2(n_737),
.B(n_730),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_929),
.B(n_730),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_935),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_822),
.A2(n_751),
.B(n_737),
.Y(n_1074)
);

NAND2x1p5_ASAP7_75t_L g1075 ( 
.A(n_914),
.B(n_927),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_864),
.B(n_751),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_863),
.B(n_674),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_875),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_822),
.A2(n_751),
.B(n_674),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_840),
.B(n_751),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_830),
.A2(n_674),
.B(n_564),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_897),
.B(n_464),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_794),
.B(n_557),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_882),
.B(n_557),
.Y(n_1084)
);

BUFx4f_ASAP7_75t_L g1085 ( 
.A(n_893),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_893),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_882),
.B(n_557),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_885),
.B(n_467),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_845),
.B(n_557),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_831),
.A2(n_564),
.B(n_557),
.Y(n_1090)
);

O2A1O1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_789),
.A2(n_383),
.B(n_350),
.C(n_378),
.Y(n_1091)
);

AO21x1_ASAP7_75t_L g1092 ( 
.A1(n_919),
.A2(n_338),
.B(n_331),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_831),
.A2(n_564),
.B(n_557),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_886),
.B(n_564),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_884),
.B(n_564),
.Y(n_1095)
);

INVx5_ASAP7_75t_L g1096 ( 
.A(n_819),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_814),
.B(n_585),
.Y(n_1097)
);

INVx4_ASAP7_75t_L g1098 ( 
.A(n_857),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_902),
.B(n_585),
.Y(n_1099)
);

NOR3xp33_ASAP7_75t_L g1100 ( 
.A(n_892),
.B(n_847),
.C(n_924),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_902),
.B(n_585),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_890),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_858),
.A2(n_588),
.B(n_585),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_932),
.B(n_472),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_835),
.B(n_588),
.Y(n_1105)
);

INVx4_ASAP7_75t_L g1106 ( 
.A(n_857),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_849),
.A2(n_894),
.B(n_872),
.Y(n_1107)
);

OAI21xp33_ASAP7_75t_L g1108 ( 
.A1(n_833),
.A2(n_348),
.B(n_340),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_849),
.A2(n_564),
.B(n_578),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_872),
.A2(n_564),
.B(n_578),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_837),
.A2(n_364),
.B1(n_356),
.B2(n_360),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_836),
.A2(n_841),
.B1(n_792),
.B2(n_907),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_952),
.A2(n_857),
.B(n_784),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_948),
.B(n_944),
.Y(n_1114)
);

INVx5_ASAP7_75t_L g1115 ( 
.A(n_1096),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_939),
.A2(n_784),
.B(n_915),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_979),
.B(n_1005),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_942),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1002),
.B(n_894),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1020),
.A2(n_808),
.B1(n_855),
.B2(n_843),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1012),
.A2(n_915),
.B(n_898),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_941),
.B(n_899),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_1000),
.A2(n_325),
.B(n_350),
.C(n_329),
.Y(n_1123)
);

INVxp33_ASAP7_75t_SL g1124 ( 
.A(n_1011),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_979),
.A2(n_769),
.B1(n_927),
.B2(n_804),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_1005),
.B(n_980),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_942),
.Y(n_1127)
);

NAND2x1p5_ASAP7_75t_L g1128 ( 
.A(n_1085),
.B(n_895),
.Y(n_1128)
);

AND2x2_ASAP7_75t_SL g1129 ( 
.A(n_1085),
.B(n_781),
.Y(n_1129)
);

INVx5_ASAP7_75t_L g1130 ( 
.A(n_1096),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_970),
.B(n_895),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_957),
.B(n_417),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_940),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_SL g1134 ( 
.A1(n_959),
.A2(n_769),
.B1(n_386),
.B2(n_372),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1067),
.A2(n_950),
.B(n_988),
.Y(n_1135)
);

INVx3_ASAP7_75t_SL g1136 ( 
.A(n_1055),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_1000),
.B(n_884),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1009),
.A2(n_915),
.B(n_898),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_964),
.B(n_970),
.Y(n_1139)
);

O2A1O1Ixp33_ASAP7_75t_SL g1140 ( 
.A1(n_1032),
.A2(n_932),
.B(n_931),
.C(n_926),
.Y(n_1140)
);

BUFx4f_ASAP7_75t_SL g1141 ( 
.A(n_1078),
.Y(n_1141)
);

INVx1_ASAP7_75t_SL g1142 ( 
.A(n_978),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_938),
.A2(n_888),
.B(n_855),
.C(n_808),
.Y(n_1143)
);

BUFx2_ASAP7_75t_L g1144 ( 
.A(n_1082),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_1022),
.A2(n_417),
.B1(n_781),
.B2(n_905),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1045),
.A2(n_889),
.B(n_882),
.Y(n_1146)
);

NOR2x1_ASAP7_75t_L g1147 ( 
.A(n_1080),
.B(n_895),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_942),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_SL g1149 ( 
.A1(n_1029),
.A2(n_362),
.B1(n_371),
.B2(n_393),
.Y(n_1149)
);

INVx8_ASAP7_75t_L g1150 ( 
.A(n_1096),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_960),
.A2(n_931),
.B(n_904),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1104),
.B(n_417),
.Y(n_1152)
);

INVxp67_ASAP7_75t_L g1153 ( 
.A(n_1022),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1025),
.B(n_899),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1091),
.A2(n_384),
.B(n_383),
.C(n_378),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1096),
.B(n_895),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_1086),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1004),
.B(n_904),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_983),
.B(n_905),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1107),
.A2(n_926),
.B(n_856),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_983),
.B(n_843),
.Y(n_1161)
);

NAND3xp33_ASAP7_75t_L g1162 ( 
.A(n_1100),
.B(n_868),
.C(n_856),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1035),
.B(n_868),
.Y(n_1163)
);

BUFx2_ASAP7_75t_L g1164 ( 
.A(n_1017),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_R g1165 ( 
.A(n_991),
.B(n_882),
.Y(n_1165)
);

OAI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_992),
.A2(n_889),
.B1(n_888),
.B2(n_395),
.Y(n_1166)
);

NAND2xp33_ASAP7_75t_SL g1167 ( 
.A(n_1016),
.B(n_889),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_981),
.A2(n_889),
.B1(n_325),
.B2(n_329),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1035),
.B(n_355),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1088),
.B(n_1013),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_R g1171 ( 
.A(n_1080),
.B(n_588),
.Y(n_1171)
);

INVxp67_ASAP7_75t_L g1172 ( 
.A(n_1047),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1026),
.B(n_374),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1031),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1083),
.A2(n_1039),
.B1(n_1048),
.B2(n_1046),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1016),
.B(n_377),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_SL g1177 ( 
.A1(n_1069),
.A2(n_403),
.B1(n_402),
.B2(n_425),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_972),
.A2(n_564),
.B(n_415),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1038),
.A2(n_414),
.B(n_578),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1027),
.B(n_1058),
.Y(n_1180)
);

O2A1O1Ixp33_ASAP7_75t_SL g1181 ( 
.A1(n_1042),
.A2(n_347),
.B(n_343),
.C(n_342),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_942),
.Y(n_1182)
);

OR2x2_ASAP7_75t_L g1183 ( 
.A(n_1059),
.B(n_384),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_1033),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_955),
.A2(n_584),
.B(n_224),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_1086),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_962),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_1043),
.B(n_1098),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_947),
.A2(n_584),
.B(n_351),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_943),
.A2(n_967),
.B(n_1062),
.Y(n_1190)
);

NOR3xp33_ASAP7_75t_SL g1191 ( 
.A(n_1003),
.B(n_385),
.C(n_382),
.Y(n_1191)
);

A2O1A1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1037),
.A2(n_392),
.B(n_388),
.C(n_366),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1069),
.B(n_391),
.Y(n_1193)
);

OR2x6_ASAP7_75t_SL g1194 ( 
.A(n_1111),
.B(n_394),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_SL g1195 ( 
.A1(n_1060),
.A2(n_398),
.B1(n_410),
.B2(n_413),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_958),
.A2(n_584),
.B(n_351),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1073),
.B(n_400),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_958),
.A2(n_584),
.B(n_370),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_962),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_993),
.B(n_409),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_1043),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1047),
.B(n_421),
.Y(n_1202)
);

O2A1O1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1010),
.A2(n_427),
.B(n_424),
.C(n_395),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1098),
.B(n_422),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_989),
.A2(n_370),
.B(n_296),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1106),
.B(n_408),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1106),
.B(n_423),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_1060),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_961),
.Y(n_1209)
);

AO32x2_ASAP7_75t_L g1210 ( 
.A1(n_1053),
.A2(n_408),
.A3(n_424),
.B1(n_18),
.B2(n_20),
.Y(n_1210)
);

O2A1O1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1044),
.A2(n_420),
.B(n_419),
.C(n_388),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1083),
.B(n_315),
.Y(n_1212)
);

A2O1A1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_1037),
.A2(n_338),
.B(n_420),
.C(n_419),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_956),
.B(n_335),
.Y(n_1214)
);

BUFx2_ASAP7_75t_L g1215 ( 
.A(n_976),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_989),
.A2(n_296),
.B(n_396),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1007),
.B(n_976),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1054),
.Y(n_1218)
);

AO21x1_ASAP7_75t_L g1219 ( 
.A1(n_973),
.A2(n_347),
.B(n_405),
.Y(n_1219)
);

CKINVDCx6p67_ASAP7_75t_R g1220 ( 
.A(n_961),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1001),
.A2(n_396),
.B(n_387),
.Y(n_1221)
);

CKINVDCx10_ASAP7_75t_R g1222 ( 
.A(n_995),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_974),
.B(n_496),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1001),
.A2(n_365),
.B(n_339),
.Y(n_1224)
);

INVx1_ASAP7_75t_SL g1225 ( 
.A(n_1075),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_975),
.A2(n_339),
.B(n_366),
.C(n_331),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1021),
.A2(n_343),
.B(n_392),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1112),
.B(n_412),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1014),
.B(n_404),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_SL g1230 ( 
.A1(n_1089),
.A2(n_404),
.B(n_405),
.C(n_18),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1075),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1094),
.A2(n_266),
.B(n_283),
.C(n_368),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_961),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1100),
.B(n_15),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1068),
.B(n_961),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_982),
.B(n_16),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1021),
.A2(n_407),
.B(n_406),
.Y(n_1237)
);

BUFx12f_ASAP7_75t_L g1238 ( 
.A(n_1015),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_969),
.A2(n_1095),
.B(n_987),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1015),
.B(n_228),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1041),
.B(n_21),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1072),
.A2(n_401),
.B1(n_399),
.B2(n_379),
.Y(n_1242)
);

INVx1_ASAP7_75t_SL g1243 ( 
.A(n_1015),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1094),
.A2(n_283),
.B(n_368),
.C(n_369),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1015),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1102),
.B(n_22),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1108),
.B(n_23),
.Y(n_1247)
);

NOR3xp33_ASAP7_75t_L g1248 ( 
.A(n_1067),
.B(n_373),
.C(n_361),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1105),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1056),
.B(n_30),
.Y(n_1250)
);

AOI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1092),
.A2(n_1063),
.B1(n_1089),
.B2(n_951),
.Y(n_1251)
);

INVx3_ASAP7_75t_SL g1252 ( 
.A(n_1102),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1102),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1095),
.A2(n_359),
.B(n_358),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1102),
.B(n_32),
.Y(n_1255)
);

INVx3_ASAP7_75t_L g1256 ( 
.A(n_953),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1040),
.B(n_357),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1099),
.A2(n_221),
.B1(n_349),
.B2(n_345),
.Y(n_1258)
);

O2A1O1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_946),
.A2(n_33),
.B(n_34),
.C(n_35),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1061),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1133),
.Y(n_1261)
);

AO31x2_ASAP7_75t_L g1262 ( 
.A1(n_1219),
.A2(n_984),
.A3(n_1097),
.B(n_1023),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1141),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1138),
.A2(n_1087),
.B(n_1084),
.Y(n_1264)
);

OA21x2_ASAP7_75t_L g1265 ( 
.A1(n_1239),
.A2(n_971),
.B(n_1049),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1132),
.B(n_35),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1190),
.A2(n_1019),
.B(n_1018),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1121),
.A2(n_1084),
.B(n_1087),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1247),
.A2(n_966),
.B(n_968),
.C(n_965),
.Y(n_1269)
);

BUFx2_ASAP7_75t_R g1270 ( 
.A(n_1184),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1151),
.A2(n_1008),
.B(n_1066),
.Y(n_1271)
);

O2A1O1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1234),
.A2(n_1070),
.B(n_1076),
.C(n_1036),
.Y(n_1272)
);

AO31x2_ASAP7_75t_L g1273 ( 
.A1(n_1122),
.A2(n_1006),
.A3(n_999),
.B(n_1071),
.Y(n_1273)
);

O2A1O1Ixp33_ASAP7_75t_SL g1274 ( 
.A1(n_1172),
.A2(n_997),
.B(n_1028),
.C(n_1077),
.Y(n_1274)
);

AO32x2_ASAP7_75t_L g1275 ( 
.A1(n_1120),
.A2(n_994),
.A3(n_977),
.B1(n_963),
.B2(n_1110),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1114),
.B(n_1101),
.Y(n_1276)
);

AO32x2_ASAP7_75t_L g1277 ( 
.A1(n_1168),
.A2(n_1109),
.A3(n_1103),
.B1(n_990),
.B2(n_986),
.Y(n_1277)
);

AO21x2_ASAP7_75t_L g1278 ( 
.A1(n_1248),
.A2(n_1064),
.B(n_1074),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1113),
.A2(n_945),
.B(n_1065),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1116),
.A2(n_1034),
.B(n_949),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1172),
.B(n_954),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1146),
.A2(n_996),
.B(n_998),
.Y(n_1282)
);

OR2x2_ASAP7_75t_L g1283 ( 
.A(n_1144),
.B(n_1090),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1141),
.Y(n_1284)
);

INVx3_ASAP7_75t_L g1285 ( 
.A(n_1150),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1136),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1117),
.B(n_230),
.Y(n_1287)
);

A2O1A1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1247),
.A2(n_1051),
.B(n_1052),
.C(n_1057),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1165),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1180),
.B(n_985),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1135),
.A2(n_1140),
.B(n_1159),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_SL g1292 ( 
.A(n_1129),
.B(n_953),
.Y(n_1292)
);

AOI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1139),
.A2(n_1050),
.B1(n_288),
.B2(n_232),
.Y(n_1293)
);

AO31x2_ASAP7_75t_L g1294 ( 
.A1(n_1232),
.A2(n_1244),
.A3(n_1143),
.B(n_1226),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1161),
.A2(n_1030),
.B(n_1093),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1165),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1158),
.A2(n_1079),
.B(n_1024),
.Y(n_1297)
);

A2O1A1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1214),
.A2(n_1081),
.B(n_354),
.C(n_341),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1139),
.B(n_36),
.Y(n_1299)
);

AOI221xp5_ASAP7_75t_L g1300 ( 
.A1(n_1123),
.A2(n_334),
.B1(n_330),
.B2(n_317),
.C(n_310),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1119),
.A2(n_308),
.B(n_302),
.Y(n_1301)
);

AOI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1134),
.A2(n_300),
.B1(n_292),
.B2(n_287),
.Y(n_1302)
);

NAND2x1_ASAP7_75t_L g1303 ( 
.A(n_1118),
.B(n_119),
.Y(n_1303)
);

HB1xp67_ASAP7_75t_L g1304 ( 
.A(n_1164),
.Y(n_1304)
);

A2O1A1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1214),
.A2(n_286),
.B(n_285),
.C(n_278),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1175),
.B(n_37),
.Y(n_1306)
);

AOI221xp5_ASAP7_75t_L g1307 ( 
.A1(n_1155),
.A2(n_276),
.B1(n_274),
.B2(n_273),
.C(n_265),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1208),
.B(n_262),
.Y(n_1308)
);

AOI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1185),
.A2(n_221),
.B(n_251),
.Y(n_1309)
);

O2A1O1Ixp33_ASAP7_75t_SL g1310 ( 
.A1(n_1230),
.A2(n_38),
.B(n_42),
.C(n_44),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1160),
.A2(n_221),
.B(n_98),
.Y(n_1311)
);

INVx1_ASAP7_75t_SL g1312 ( 
.A(n_1142),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1223),
.A2(n_259),
.B(n_249),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1196),
.A2(n_221),
.B(n_93),
.Y(n_1314)
);

AOI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1125),
.A2(n_244),
.B1(n_242),
.B2(n_235),
.Y(n_1315)
);

NAND2x1_ASAP7_75t_L g1316 ( 
.A(n_1118),
.B(n_147),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1198),
.A2(n_221),
.B(n_201),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1178),
.A2(n_144),
.B(n_200),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1189),
.A2(n_1216),
.B(n_1205),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1136),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1162),
.A2(n_143),
.B(n_191),
.Y(n_1321)
);

INVx2_ASAP7_75t_SL g1322 ( 
.A(n_1157),
.Y(n_1322)
);

O2A1O1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1228),
.A2(n_42),
.B(n_44),
.C(n_46),
.Y(n_1323)
);

O2A1O1Ixp33_ASAP7_75t_SL g1324 ( 
.A1(n_1188),
.A2(n_1255),
.B(n_1246),
.C(n_1260),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1152),
.B(n_47),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1175),
.A2(n_140),
.B(n_190),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1126),
.A2(n_1170),
.B1(n_1129),
.B2(n_1229),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1153),
.B(n_48),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1212),
.A2(n_1181),
.B(n_1163),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1179),
.A2(n_136),
.B(n_182),
.Y(n_1330)
);

AO31x2_ASAP7_75t_L g1331 ( 
.A1(n_1249),
.A2(n_221),
.A3(n_179),
.B(n_166),
.Y(n_1331)
);

A2O1A1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1241),
.A2(n_50),
.B(n_52),
.C(n_53),
.Y(n_1332)
);

A2O1A1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1241),
.A2(n_52),
.B(n_53),
.C(n_57),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1174),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1153),
.B(n_58),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1227),
.A2(n_221),
.B(n_159),
.Y(n_1336)
);

AO31x2_ASAP7_75t_L g1337 ( 
.A1(n_1192),
.A2(n_221),
.A3(n_153),
.B(n_128),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1217),
.A2(n_1147),
.B(n_1221),
.Y(n_1338)
);

O2A1O1Ixp33_ASAP7_75t_SL g1339 ( 
.A1(n_1202),
.A2(n_58),
.B(n_59),
.C(n_62),
.Y(n_1339)
);

AND2x4_ASAP7_75t_L g1340 ( 
.A(n_1231),
.B(n_114),
.Y(n_1340)
);

NOR4xp25_ASAP7_75t_L g1341 ( 
.A(n_1213),
.B(n_59),
.C(n_64),
.D(n_67),
.Y(n_1341)
);

NOR3xp33_ASAP7_75t_L g1342 ( 
.A(n_1149),
.B(n_64),
.C(n_67),
.Y(n_1342)
);

OR2x6_ASAP7_75t_L g1343 ( 
.A(n_1150),
.B(n_69),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1251),
.A2(n_221),
.B(n_104),
.Y(n_1344)
);

AOI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1193),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_1345)
);

AOI221x1_ASAP7_75t_L g1346 ( 
.A1(n_1248),
.A2(n_71),
.B1(n_74),
.B2(n_76),
.C(n_77),
.Y(n_1346)
);

BUFx12f_ASAP7_75t_L g1347 ( 
.A(n_1209),
.Y(n_1347)
);

OAI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1236),
.A2(n_74),
.B(n_79),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1157),
.B(n_88),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1250),
.A2(n_96),
.B(n_100),
.Y(n_1350)
);

A2O1A1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1211),
.A2(n_1203),
.B(n_1250),
.C(n_1191),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1256),
.A2(n_1224),
.B(n_1156),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1194),
.B(n_1137),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1167),
.A2(n_1166),
.B(n_1154),
.Y(n_1354)
);

A2O1A1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1191),
.A2(n_1259),
.B(n_1169),
.C(n_1145),
.Y(n_1355)
);

BUFx2_ASAP7_75t_L g1356 ( 
.A(n_1186),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1257),
.A2(n_1240),
.B(n_1137),
.Y(n_1357)
);

AOI221x1_ASAP7_75t_L g1358 ( 
.A1(n_1173),
.A2(n_1242),
.B1(n_1254),
.B2(n_1195),
.C(n_1218),
.Y(n_1358)
);

O2A1O1Ixp5_ASAP7_75t_SL g1359 ( 
.A1(n_1131),
.A2(n_1186),
.B(n_1245),
.C(n_1207),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1245),
.A2(n_1145),
.B(n_1243),
.Y(n_1360)
);

O2A1O1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1176),
.A2(n_1204),
.B(n_1197),
.C(n_1200),
.Y(n_1361)
);

O2A1O1Ixp33_ASAP7_75t_L g1362 ( 
.A1(n_1206),
.A2(n_1183),
.B(n_1215),
.C(n_1199),
.Y(n_1362)
);

CKINVDCx20_ASAP7_75t_R g1363 ( 
.A(n_1220),
.Y(n_1363)
);

A2O1A1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1258),
.A2(n_1206),
.B(n_1237),
.C(n_1225),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_1124),
.B(n_1177),
.Y(n_1365)
);

OAI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1258),
.A2(n_1235),
.B(n_1187),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1256),
.A2(n_1128),
.B(n_1201),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1238),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1118),
.A2(n_1182),
.B(n_1127),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1118),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1253),
.B(n_1182),
.Y(n_1371)
);

O2A1O1Ixp33_ASAP7_75t_SL g1372 ( 
.A1(n_1201),
.A2(n_1150),
.B(n_1210),
.C(n_1130),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1127),
.A2(n_1253),
.B(n_1233),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1127),
.A2(n_1253),
.B(n_1233),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1210),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1127),
.A2(n_1253),
.B(n_1233),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1252),
.B(n_1210),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1148),
.A2(n_1182),
.B(n_1233),
.Y(n_1378)
);

AO31x2_ASAP7_75t_L g1379 ( 
.A1(n_1210),
.A2(n_1222),
.A3(n_1148),
.B(n_1182),
.Y(n_1379)
);

OAI22x1_ASAP7_75t_L g1380 ( 
.A1(n_1252),
.A2(n_1115),
.B1(n_1130),
.B2(n_1171),
.Y(n_1380)
);

CKINVDCx6p67_ASAP7_75t_R g1381 ( 
.A(n_1115),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1148),
.A2(n_1115),
.B(n_1130),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1115),
.Y(n_1383)
);

AOI31xp67_ASAP7_75t_L g1384 ( 
.A1(n_1130),
.A2(n_1251),
.A3(n_989),
.B(n_1001),
.Y(n_1384)
);

BUFx6f_ASAP7_75t_L g1385 ( 
.A(n_1238),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1114),
.B(n_948),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1190),
.A2(n_1239),
.B(n_1151),
.Y(n_1387)
);

CKINVDCx11_ASAP7_75t_R g1388 ( 
.A(n_1136),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_1184),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_SL g1390 ( 
.A(n_1129),
.B(n_670),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1133),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1138),
.A2(n_952),
.B(n_939),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1138),
.A2(n_952),
.B(n_939),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1133),
.Y(n_1394)
);

AOI221x1_ASAP7_75t_L g1395 ( 
.A1(n_1234),
.A2(n_1247),
.B1(n_941),
.B2(n_1213),
.C(n_1192),
.Y(n_1395)
);

NAND3xp33_ASAP7_75t_SL g1396 ( 
.A(n_1234),
.B(n_547),
.C(n_642),
.Y(n_1396)
);

OAI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1135),
.A2(n_952),
.B(n_948),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1190),
.A2(n_1239),
.B(n_1151),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1190),
.A2(n_1239),
.B(n_1151),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1150),
.Y(n_1400)
);

O2A1O1Ixp33_ASAP7_75t_SL g1401 ( 
.A1(n_1172),
.A2(n_948),
.B(n_939),
.C(n_1234),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1190),
.A2(n_1239),
.B(n_1151),
.Y(n_1402)
);

OAI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1194),
.A2(n_944),
.B1(n_980),
.B2(n_740),
.Y(n_1403)
);

AOI221xp5_ASAP7_75t_L g1404 ( 
.A1(n_1123),
.A2(n_941),
.B1(n_673),
.B2(n_635),
.C(n_694),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1138),
.A2(n_952),
.B(n_939),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_1141),
.Y(n_1406)
);

OA21x2_ASAP7_75t_L g1407 ( 
.A1(n_1239),
.A2(n_1190),
.B(n_1135),
.Y(n_1407)
);

AO31x2_ASAP7_75t_L g1408 ( 
.A1(n_1219),
.A2(n_1122),
.A3(n_1239),
.B(n_1232),
.Y(n_1408)
);

AO31x2_ASAP7_75t_L g1409 ( 
.A1(n_1219),
.A2(n_1122),
.A3(n_1239),
.B(n_1232),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1141),
.Y(n_1410)
);

O2A1O1Ixp33_ASAP7_75t_SL g1411 ( 
.A1(n_1172),
.A2(n_948),
.B(n_939),
.C(n_1234),
.Y(n_1411)
);

INVx1_ASAP7_75t_SL g1412 ( 
.A(n_1142),
.Y(n_1412)
);

NAND3xp33_ASAP7_75t_L g1413 ( 
.A(n_1234),
.B(n_941),
.C(n_1247),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1138),
.A2(n_952),
.B(n_939),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1190),
.A2(n_1239),
.B(n_1151),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1138),
.A2(n_952),
.B(n_939),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1135),
.A2(n_952),
.B(n_948),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1190),
.A2(n_1239),
.B(n_1151),
.Y(n_1418)
);

AOI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1239),
.A2(n_1190),
.B(n_1219),
.Y(n_1419)
);

OAI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1135),
.A2(n_952),
.B(n_948),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1132),
.B(n_957),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1144),
.B(n_957),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1381),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1261),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1403),
.A2(n_1404),
.B1(n_1413),
.B2(n_1327),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1404),
.A2(n_1351),
.B1(n_1413),
.B2(n_1386),
.Y(n_1426)
);

BUFx8_ASAP7_75t_L g1427 ( 
.A(n_1289),
.Y(n_1427)
);

INVx8_ASAP7_75t_L g1428 ( 
.A(n_1347),
.Y(n_1428)
);

INVx6_ASAP7_75t_L g1429 ( 
.A(n_1385),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_SL g1430 ( 
.A(n_1286),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1386),
.A2(n_1355),
.B1(n_1345),
.B2(n_1348),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1263),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1348),
.A2(n_1353),
.B1(n_1306),
.B2(n_1315),
.Y(n_1433)
);

INVx8_ASAP7_75t_L g1434 ( 
.A(n_1363),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1421),
.A2(n_1342),
.B1(n_1306),
.B2(n_1422),
.Y(n_1435)
);

AOI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1396),
.A2(n_1390),
.B1(n_1300),
.B2(n_1365),
.Y(n_1436)
);

INVx4_ASAP7_75t_L g1437 ( 
.A(n_1389),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1299),
.A2(n_1266),
.B1(n_1300),
.B2(n_1390),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1350),
.A2(n_1325),
.B1(n_1307),
.B2(n_1375),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_SL g1440 ( 
.A1(n_1380),
.A2(n_1350),
.B(n_1395),
.Y(n_1440)
);

AOI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1308),
.A2(n_1292),
.B1(n_1335),
.B2(n_1287),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_SL g1442 ( 
.A1(n_1292),
.A2(n_1377),
.B1(n_1343),
.B2(n_1366),
.Y(n_1442)
);

BUFx2_ASAP7_75t_SL g1443 ( 
.A(n_1320),
.Y(n_1443)
);

BUFx2_ASAP7_75t_R g1444 ( 
.A(n_1296),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1334),
.Y(n_1445)
);

INVx2_ASAP7_75t_SL g1446 ( 
.A(n_1385),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1391),
.Y(n_1447)
);

OAI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1343),
.A2(n_1346),
.B1(n_1276),
.B2(n_1358),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1356),
.B(n_1322),
.Y(n_1449)
);

INVx6_ASAP7_75t_L g1450 ( 
.A(n_1385),
.Y(n_1450)
);

BUFx10_ASAP7_75t_L g1451 ( 
.A(n_1343),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_SL g1452 ( 
.A1(n_1366),
.A2(n_1349),
.B1(n_1328),
.B2(n_1276),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1388),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1307),
.A2(n_1394),
.B1(n_1329),
.B2(n_1304),
.Y(n_1454)
);

INVx4_ASAP7_75t_L g1455 ( 
.A(n_1284),
.Y(n_1455)
);

INVx6_ASAP7_75t_L g1456 ( 
.A(n_1340),
.Y(n_1456)
);

AOI21xp33_ASAP7_75t_L g1457 ( 
.A1(n_1361),
.A2(n_1323),
.B(n_1362),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1406),
.Y(n_1458)
);

CKINVDCx20_ASAP7_75t_R g1459 ( 
.A(n_1368),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1283),
.A2(n_1420),
.B1(n_1397),
.B2(n_1417),
.Y(n_1460)
);

INVx6_ASAP7_75t_L g1461 ( 
.A(n_1340),
.Y(n_1461)
);

CKINVDCx11_ASAP7_75t_R g1462 ( 
.A(n_1312),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1397),
.A2(n_1420),
.B1(n_1417),
.B2(n_1326),
.Y(n_1463)
);

INVx2_ASAP7_75t_SL g1464 ( 
.A(n_1412),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1293),
.A2(n_1281),
.B1(n_1302),
.B2(n_1290),
.Y(n_1465)
);

AOI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1332),
.A2(n_1333),
.B1(n_1305),
.B2(n_1341),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_1270),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1281),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_SL g1469 ( 
.A1(n_1341),
.A2(n_1379),
.B1(n_1344),
.B2(n_1372),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1401),
.B(n_1411),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1290),
.Y(n_1471)
);

INVx2_ASAP7_75t_SL g1472 ( 
.A(n_1285),
.Y(n_1472)
);

INVx1_ASAP7_75t_SL g1473 ( 
.A(n_1371),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1357),
.B(n_1379),
.Y(n_1474)
);

NAND2x1p5_ASAP7_75t_L g1475 ( 
.A(n_1367),
.B(n_1383),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1370),
.Y(n_1476)
);

BUFx12f_ASAP7_75t_L g1477 ( 
.A(n_1339),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1379),
.A2(n_1354),
.B1(n_1360),
.B2(n_1321),
.Y(n_1478)
);

BUFx8_ASAP7_75t_L g1479 ( 
.A(n_1275),
.Y(n_1479)
);

INVxp67_ASAP7_75t_SL g1480 ( 
.A(n_1407),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_1400),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1400),
.B(n_1371),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1291),
.A2(n_1318),
.B1(n_1301),
.B2(n_1330),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1324),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1265),
.A2(n_1295),
.B1(n_1416),
.B2(n_1278),
.Y(n_1485)
);

INVx4_ASAP7_75t_L g1486 ( 
.A(n_1407),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1364),
.A2(n_1272),
.B1(n_1269),
.B2(n_1298),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_1376),
.Y(n_1488)
);

BUFx2_ASAP7_75t_SL g1489 ( 
.A(n_1382),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1369),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1265),
.A2(n_1416),
.B1(n_1278),
.B2(n_1336),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1392),
.A2(n_1405),
.B1(n_1414),
.B2(n_1393),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1331),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1331),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1338),
.Y(n_1495)
);

OAI21xp33_ASAP7_75t_SL g1496 ( 
.A1(n_1359),
.A2(n_1352),
.B(n_1311),
.Y(n_1496)
);

OAI22xp33_ASAP7_75t_SL g1497 ( 
.A1(n_1303),
.A2(n_1316),
.B1(n_1313),
.B2(n_1310),
.Y(n_1497)
);

INVx3_ASAP7_75t_L g1498 ( 
.A(n_1294),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_SL g1499 ( 
.A1(n_1294),
.A2(n_1337),
.B1(n_1317),
.B2(n_1314),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_SL g1500 ( 
.A1(n_1294),
.A2(n_1337),
.B1(n_1384),
.B2(n_1268),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1337),
.Y(n_1501)
);

OAI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1297),
.A2(n_1264),
.B1(n_1374),
.B2(n_1378),
.Y(n_1502)
);

CKINVDCx8_ASAP7_75t_R g1503 ( 
.A(n_1373),
.Y(n_1503)
);

OAI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1288),
.A2(n_1274),
.B(n_1282),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1419),
.A2(n_1280),
.B1(n_1279),
.B2(n_1282),
.Y(n_1505)
);

AOI22xp5_ASAP7_75t_SL g1506 ( 
.A1(n_1279),
.A2(n_1280),
.B1(n_1409),
.B2(n_1408),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_SL g1507 ( 
.A1(n_1319),
.A2(n_1267),
.B1(n_1409),
.B2(n_1408),
.Y(n_1507)
);

CKINVDCx6p67_ASAP7_75t_R g1508 ( 
.A(n_1408),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1271),
.A2(n_1398),
.B1(n_1415),
.B2(n_1402),
.Y(n_1509)
);

INVx4_ASAP7_75t_L g1510 ( 
.A(n_1277),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1387),
.A2(n_1418),
.B1(n_1399),
.B2(n_1275),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1409),
.Y(n_1512)
);

BUFx2_ASAP7_75t_SL g1513 ( 
.A(n_1277),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1275),
.A2(n_1262),
.B1(n_1277),
.B2(n_1273),
.Y(n_1514)
);

OAI21xp5_ASAP7_75t_SL g1515 ( 
.A1(n_1309),
.A2(n_1404),
.B(n_1348),
.Y(n_1515)
);

CKINVDCx6p67_ASAP7_75t_R g1516 ( 
.A(n_1273),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1261),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1403),
.A2(n_1404),
.B1(n_964),
.B2(n_1413),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_SL g1519 ( 
.A1(n_1413),
.A2(n_964),
.B1(n_944),
.B2(n_598),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1403),
.A2(n_1404),
.B1(n_964),
.B2(n_1413),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1404),
.A2(n_1351),
.B1(n_1234),
.B2(n_948),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_1410),
.Y(n_1522)
);

BUFx10_ASAP7_75t_L g1523 ( 
.A(n_1389),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1404),
.A2(n_1403),
.B1(n_642),
.B2(n_941),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1381),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1261),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1261),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1261),
.Y(n_1528)
);

INVx3_ASAP7_75t_SL g1529 ( 
.A(n_1389),
.Y(n_1529)
);

CKINVDCx6p67_ASAP7_75t_R g1530 ( 
.A(n_1388),
.Y(n_1530)
);

INVx3_ASAP7_75t_SL g1531 ( 
.A(n_1389),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1261),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1403),
.A2(n_1404),
.B1(n_964),
.B2(n_1413),
.Y(n_1533)
);

CKINVDCx6p67_ASAP7_75t_R g1534 ( 
.A(n_1388),
.Y(n_1534)
);

CKINVDCx16_ASAP7_75t_R g1535 ( 
.A(n_1363),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1403),
.A2(n_1404),
.B1(n_964),
.B2(n_1413),
.Y(n_1536)
);

OAI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1348),
.A2(n_1234),
.B1(n_1306),
.B2(n_1413),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1410),
.Y(n_1538)
);

BUFx3_ASAP7_75t_L g1539 ( 
.A(n_1410),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_SL g1540 ( 
.A1(n_1413),
.A2(n_964),
.B1(n_944),
.B2(n_598),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1404),
.A2(n_1351),
.B1(n_1234),
.B2(n_948),
.Y(n_1541)
);

INVx8_ASAP7_75t_L g1542 ( 
.A(n_1347),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1404),
.A2(n_1351),
.B1(n_1234),
.B2(n_948),
.Y(n_1543)
);

CKINVDCx14_ASAP7_75t_R g1544 ( 
.A(n_1388),
.Y(n_1544)
);

OAI21xp5_ASAP7_75t_SL g1545 ( 
.A1(n_1404),
.A2(n_1348),
.B(n_1345),
.Y(n_1545)
);

CKINVDCx20_ASAP7_75t_R g1546 ( 
.A(n_1388),
.Y(n_1546)
);

INVx1_ASAP7_75t_SL g1547 ( 
.A(n_1312),
.Y(n_1547)
);

AOI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1404),
.A2(n_1403),
.B1(n_642),
.B2(n_941),
.Y(n_1548)
);

INVx1_ASAP7_75t_SL g1549 ( 
.A(n_1312),
.Y(n_1549)
);

OAI21xp33_ASAP7_75t_L g1550 ( 
.A1(n_1348),
.A2(n_1404),
.B(n_941),
.Y(n_1550)
);

BUFx3_ASAP7_75t_L g1551 ( 
.A(n_1410),
.Y(n_1551)
);

BUFx2_ASAP7_75t_R g1552 ( 
.A(n_1389),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_SL g1553 ( 
.A1(n_1413),
.A2(n_964),
.B1(n_944),
.B2(n_598),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1261),
.Y(n_1554)
);

BUFx2_ASAP7_75t_R g1555 ( 
.A(n_1389),
.Y(n_1555)
);

INVx4_ASAP7_75t_SL g1556 ( 
.A(n_1379),
.Y(n_1556)
);

INVx6_ASAP7_75t_L g1557 ( 
.A(n_1347),
.Y(n_1557)
);

BUFx2_ASAP7_75t_L g1558 ( 
.A(n_1304),
.Y(n_1558)
);

OAI21xp33_ASAP7_75t_L g1559 ( 
.A1(n_1348),
.A2(n_1404),
.B(n_941),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1403),
.A2(n_1404),
.B1(n_964),
.B2(n_1413),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_SL g1561 ( 
.A1(n_1413),
.A2(n_964),
.B1(n_944),
.B2(n_598),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1261),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1422),
.B(n_1356),
.Y(n_1563)
);

INVx3_ASAP7_75t_L g1564 ( 
.A(n_1381),
.Y(n_1564)
);

INVx6_ASAP7_75t_L g1565 ( 
.A(n_1347),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1468),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1471),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_1490),
.Y(n_1568)
);

OAI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1504),
.A2(n_1505),
.B(n_1485),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1474),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1424),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1563),
.B(n_1510),
.Y(n_1572)
);

BUFx2_ASAP7_75t_L g1573 ( 
.A(n_1488),
.Y(n_1573)
);

INVx3_ASAP7_75t_L g1574 ( 
.A(n_1486),
.Y(n_1574)
);

OA21x2_ASAP7_75t_L g1575 ( 
.A1(n_1485),
.A2(n_1492),
.B(n_1491),
.Y(n_1575)
);

OAI21x1_ASAP7_75t_L g1576 ( 
.A1(n_1509),
.A2(n_1491),
.B(n_1492),
.Y(n_1576)
);

INVx2_ASAP7_75t_SL g1577 ( 
.A(n_1475),
.Y(n_1577)
);

CKINVDCx20_ASAP7_75t_R g1578 ( 
.A(n_1546),
.Y(n_1578)
);

AO31x2_ASAP7_75t_L g1579 ( 
.A1(n_1510),
.A2(n_1501),
.A3(n_1487),
.B(n_1494),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1519),
.A2(n_1561),
.B1(n_1553),
.B2(n_1540),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1519),
.A2(n_1561),
.B1(n_1553),
.B2(n_1540),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1558),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_SL g1583 ( 
.A(n_1441),
.B(n_1537),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1445),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_SL g1585 ( 
.A1(n_1433),
.A2(n_1431),
.B1(n_1543),
.B2(n_1541),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1447),
.Y(n_1586)
);

BUFx3_ASAP7_75t_L g1587 ( 
.A(n_1503),
.Y(n_1587)
);

INVx3_ASAP7_75t_L g1588 ( 
.A(n_1486),
.Y(n_1588)
);

AOI21x1_ASAP7_75t_L g1589 ( 
.A1(n_1470),
.A2(n_1521),
.B(n_1484),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1550),
.A2(n_1559),
.B1(n_1442),
.B2(n_1533),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1517),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1460),
.B(n_1513),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1449),
.Y(n_1593)
);

INVx3_ASAP7_75t_L g1594 ( 
.A(n_1516),
.Y(n_1594)
);

INVxp67_ASAP7_75t_L g1595 ( 
.A(n_1464),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_1475),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1526),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1527),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1528),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1532),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1554),
.Y(n_1601)
);

OAI21x1_ASAP7_75t_L g1602 ( 
.A1(n_1509),
.A2(n_1511),
.B(n_1495),
.Y(n_1602)
);

INVx3_ASAP7_75t_L g1603 ( 
.A(n_1498),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1460),
.B(n_1562),
.Y(n_1604)
);

OAI21x1_ASAP7_75t_L g1605 ( 
.A1(n_1511),
.A2(n_1480),
.B(n_1493),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1556),
.B(n_1512),
.Y(n_1606)
);

OAI21x1_ASAP7_75t_L g1607 ( 
.A1(n_1480),
.A2(n_1463),
.B(n_1483),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1508),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1514),
.B(n_1482),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1479),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1476),
.Y(n_1611)
);

BUFx3_ASAP7_75t_L g1612 ( 
.A(n_1525),
.Y(n_1612)
);

INVx3_ASAP7_75t_L g1613 ( 
.A(n_1525),
.Y(n_1613)
);

OAI21x1_ASAP7_75t_L g1614 ( 
.A1(n_1463),
.A2(n_1483),
.B(n_1514),
.Y(n_1614)
);

AOI21x1_ASAP7_75t_L g1615 ( 
.A1(n_1426),
.A2(n_1472),
.B(n_1496),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1506),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_SL g1617 ( 
.A1(n_1477),
.A2(n_1461),
.B1(n_1456),
.B2(n_1545),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1473),
.Y(n_1618)
);

OAI21x1_ASAP7_75t_L g1619 ( 
.A1(n_1515),
.A2(n_1440),
.B(n_1465),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1547),
.Y(n_1620)
);

INVx3_ASAP7_75t_L g1621 ( 
.A(n_1525),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1549),
.B(n_1537),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1525),
.Y(n_1623)
);

BUFx2_ASAP7_75t_SL g1624 ( 
.A(n_1451),
.Y(n_1624)
);

INVxp67_ASAP7_75t_L g1625 ( 
.A(n_1443),
.Y(n_1625)
);

CKINVDCx20_ASAP7_75t_R g1626 ( 
.A(n_1544),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1432),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1489),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1451),
.Y(n_1629)
);

BUFx12f_ASAP7_75t_L g1630 ( 
.A(n_1462),
.Y(n_1630)
);

AOI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1524),
.A2(n_1548),
.B1(n_1560),
.B2(n_1520),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1436),
.A2(n_1438),
.B1(n_1439),
.B2(n_1533),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1462),
.B(n_1531),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1529),
.B(n_1531),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1518),
.B(n_1560),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1507),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1458),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1458),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1507),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1500),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1500),
.Y(n_1641)
);

BUFx3_ASAP7_75t_L g1642 ( 
.A(n_1423),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1502),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1455),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1466),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1423),
.Y(n_1646)
);

OAI21x1_ASAP7_75t_SL g1647 ( 
.A1(n_1439),
.A2(n_1454),
.B(n_1425),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1502),
.Y(n_1648)
);

INVx2_ASAP7_75t_SL g1649 ( 
.A(n_1557),
.Y(n_1649)
);

OAI21x1_ASAP7_75t_L g1650 ( 
.A1(n_1465),
.A2(n_1454),
.B(n_1425),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1564),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1469),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1469),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1518),
.B(n_1520),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1478),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1564),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1478),
.Y(n_1657)
);

AOI21x1_ASAP7_75t_L g1658 ( 
.A1(n_1499),
.A2(n_1448),
.B(n_1446),
.Y(n_1658)
);

OAI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1438),
.A2(n_1536),
.B1(n_1435),
.B2(n_1452),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1499),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1448),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1536),
.B(n_1442),
.Y(n_1662)
);

INVx3_ASAP7_75t_L g1663 ( 
.A(n_1429),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1452),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1497),
.Y(n_1665)
);

OAI21x1_ASAP7_75t_L g1666 ( 
.A1(n_1435),
.A2(n_1457),
.B(n_1481),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1430),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1430),
.Y(n_1668)
);

BUFx2_ASAP7_75t_L g1669 ( 
.A(n_1427),
.Y(n_1669)
);

BUFx3_ASAP7_75t_L g1670 ( 
.A(n_1427),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1450),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1529),
.B(n_1535),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1539),
.Y(n_1673)
);

OAI21x1_ASAP7_75t_L g1674 ( 
.A1(n_1444),
.A2(n_1565),
.B(n_1557),
.Y(n_1674)
);

AOI21x1_ASAP7_75t_L g1675 ( 
.A1(n_1539),
.A2(n_1434),
.B(n_1565),
.Y(n_1675)
);

INVx2_ASAP7_75t_SL g1676 ( 
.A(n_1557),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1437),
.B(n_1551),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1522),
.Y(n_1678)
);

BUFx2_ASAP7_75t_L g1679 ( 
.A(n_1459),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1538),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1585),
.A2(n_1544),
.B1(n_1565),
.B2(n_1467),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1627),
.B(n_1530),
.Y(n_1682)
);

OAI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1583),
.A2(n_1437),
.B(n_1453),
.Y(n_1683)
);

OAI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1619),
.A2(n_1434),
.B(n_1552),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1622),
.B(n_1534),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1638),
.B(n_1593),
.Y(n_1686)
);

AO21x2_ASAP7_75t_L g1687 ( 
.A1(n_1647),
.A2(n_1434),
.B(n_1428),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1575),
.A2(n_1428),
.B(n_1542),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_1578),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1571),
.Y(n_1690)
);

AOI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1632),
.A2(n_1428),
.B1(n_1542),
.B2(n_1523),
.Y(n_1691)
);

OAI21x1_ASAP7_75t_SL g1692 ( 
.A1(n_1647),
.A2(n_1542),
.B(n_1555),
.Y(n_1692)
);

AOI221xp5_ASAP7_75t_L g1693 ( 
.A1(n_1659),
.A2(n_1523),
.B1(n_1661),
.B2(n_1652),
.C(n_1653),
.Y(n_1693)
);

OAI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1619),
.A2(n_1650),
.B(n_1666),
.Y(n_1694)
);

AO21x1_ASAP7_75t_L g1695 ( 
.A1(n_1661),
.A2(n_1653),
.B(n_1652),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1572),
.B(n_1582),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1571),
.Y(n_1697)
);

OAI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1650),
.A2(n_1666),
.B(n_1589),
.Y(n_1698)
);

AO21x2_ASAP7_75t_L g1699 ( 
.A1(n_1658),
.A2(n_1657),
.B(n_1655),
.Y(n_1699)
);

OAI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1589),
.A2(n_1631),
.B(n_1645),
.Y(n_1700)
);

O2A1O1Ixp33_ASAP7_75t_SL g1701 ( 
.A1(n_1626),
.A2(n_1625),
.B(n_1644),
.C(n_1673),
.Y(n_1701)
);

AOI221xp5_ASAP7_75t_L g1702 ( 
.A1(n_1660),
.A2(n_1655),
.B1(n_1657),
.B2(n_1590),
.C(n_1664),
.Y(n_1702)
);

AO21x1_ASAP7_75t_L g1703 ( 
.A1(n_1658),
.A2(n_1645),
.B(n_1631),
.Y(n_1703)
);

NAND2xp33_ASAP7_75t_R g1704 ( 
.A(n_1662),
.B(n_1573),
.Y(n_1704)
);

AOI22xp33_ASAP7_75t_L g1705 ( 
.A1(n_1662),
.A2(n_1581),
.B1(n_1580),
.B2(n_1654),
.Y(n_1705)
);

AOI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1635),
.A2(n_1664),
.B1(n_1568),
.B2(n_1665),
.Y(n_1706)
);

INVxp67_ASAP7_75t_L g1707 ( 
.A(n_1616),
.Y(n_1707)
);

OAI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1665),
.A2(n_1616),
.B(n_1615),
.Y(n_1708)
);

O2A1O1Ixp33_ASAP7_75t_L g1709 ( 
.A1(n_1643),
.A2(n_1648),
.B(n_1620),
.C(n_1636),
.Y(n_1709)
);

AO32x2_ASAP7_75t_L g1710 ( 
.A1(n_1577),
.A2(n_1596),
.A3(n_1649),
.B1(n_1676),
.B2(n_1604),
.Y(n_1710)
);

O2A1O1Ixp33_ASAP7_75t_L g1711 ( 
.A1(n_1643),
.A2(n_1648),
.B(n_1636),
.C(n_1639),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1637),
.B(n_1609),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1568),
.B(n_1595),
.Y(n_1713)
);

A2O1A1Ixp33_ASAP7_75t_L g1714 ( 
.A1(n_1660),
.A2(n_1640),
.B(n_1641),
.C(n_1639),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1610),
.B(n_1608),
.Y(n_1715)
);

AOI221xp5_ASAP7_75t_L g1716 ( 
.A1(n_1640),
.A2(n_1570),
.B1(n_1641),
.B2(n_1592),
.C(n_1566),
.Y(n_1716)
);

AOI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1617),
.A2(n_1587),
.B1(n_1610),
.B2(n_1592),
.Y(n_1717)
);

AOI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1587),
.A2(n_1629),
.B1(n_1608),
.B2(n_1667),
.Y(n_1718)
);

BUFx3_ASAP7_75t_L g1719 ( 
.A(n_1642),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1606),
.B(n_1594),
.Y(n_1720)
);

A2O1A1Ixp33_ASAP7_75t_L g1721 ( 
.A1(n_1587),
.A2(n_1614),
.B(n_1674),
.C(n_1569),
.Y(n_1721)
);

A2O1A1Ixp33_ASAP7_75t_L g1722 ( 
.A1(n_1614),
.A2(n_1674),
.B(n_1569),
.C(n_1607),
.Y(n_1722)
);

INVxp67_ASAP7_75t_L g1723 ( 
.A(n_1570),
.Y(n_1723)
);

AO32x2_ASAP7_75t_L g1724 ( 
.A1(n_1577),
.A2(n_1596),
.A3(n_1676),
.B1(n_1649),
.B2(n_1618),
.Y(n_1724)
);

CKINVDCx5p33_ASAP7_75t_R g1725 ( 
.A(n_1630),
.Y(n_1725)
);

OA21x2_ASAP7_75t_L g1726 ( 
.A1(n_1576),
.A2(n_1607),
.B(n_1602),
.Y(n_1726)
);

OAI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1678),
.A2(n_1680),
.B1(n_1646),
.B2(n_1651),
.Y(n_1727)
);

NOR2x1_ASAP7_75t_L g1728 ( 
.A(n_1670),
.B(n_1667),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1606),
.B(n_1594),
.Y(n_1729)
);

O2A1O1Ixp33_ASAP7_75t_SL g1730 ( 
.A1(n_1634),
.A2(n_1633),
.B(n_1672),
.C(n_1668),
.Y(n_1730)
);

OAI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1615),
.A2(n_1576),
.B(n_1628),
.Y(n_1731)
);

A2O1A1Ixp33_ASAP7_75t_L g1732 ( 
.A1(n_1594),
.A2(n_1605),
.B(n_1624),
.C(n_1567),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_L g1733 ( 
.A(n_1675),
.B(n_1642),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1579),
.Y(n_1734)
);

OAI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1646),
.A2(n_1651),
.B1(n_1656),
.B2(n_1679),
.Y(n_1735)
);

INVx3_ASAP7_75t_L g1736 ( 
.A(n_1612),
.Y(n_1736)
);

NOR2x1_ASAP7_75t_SL g1737 ( 
.A(n_1630),
.B(n_1624),
.Y(n_1737)
);

A2O1A1Ixp33_ASAP7_75t_L g1738 ( 
.A1(n_1605),
.A2(n_1567),
.B(n_1566),
.C(n_1642),
.Y(n_1738)
);

OAI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1656),
.A2(n_1679),
.B1(n_1670),
.B2(n_1669),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1663),
.B(n_1623),
.Y(n_1740)
);

CKINVDCx20_ASAP7_75t_R g1741 ( 
.A(n_1669),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1663),
.B(n_1613),
.Y(n_1742)
);

O2A1O1Ixp33_ASAP7_75t_L g1743 ( 
.A1(n_1575),
.A2(n_1629),
.B(n_1671),
.C(n_1677),
.Y(n_1743)
);

OAI22xp5_ASAP7_75t_SL g1744 ( 
.A1(n_1613),
.A2(n_1621),
.B1(n_1623),
.B2(n_1575),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1712),
.B(n_1575),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1730),
.B(n_1621),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1690),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1726),
.B(n_1602),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1697),
.Y(n_1749)
);

OR2x2_ASAP7_75t_L g1750 ( 
.A(n_1696),
.B(n_1579),
.Y(n_1750)
);

AND2x4_ASAP7_75t_L g1751 ( 
.A(n_1720),
.B(n_1729),
.Y(n_1751)
);

BUFx6f_ASAP7_75t_L g1752 ( 
.A(n_1724),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1723),
.B(n_1600),
.Y(n_1753)
);

BUFx3_ASAP7_75t_L g1754 ( 
.A(n_1719),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1710),
.B(n_1588),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1723),
.Y(n_1756)
);

OAI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1705),
.A2(n_1600),
.B1(n_1599),
.B2(n_1598),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1710),
.B(n_1574),
.Y(n_1758)
);

INVx5_ASAP7_75t_L g1759 ( 
.A(n_1729),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1710),
.B(n_1574),
.Y(n_1760)
);

BUFx2_ASAP7_75t_L g1761 ( 
.A(n_1724),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1710),
.B(n_1574),
.Y(n_1762)
);

NAND3xp33_ASAP7_75t_L g1763 ( 
.A(n_1698),
.B(n_1597),
.C(n_1601),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1731),
.B(n_1686),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1707),
.B(n_1597),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1722),
.B(n_1584),
.Y(n_1766)
);

INVxp33_ASAP7_75t_SL g1767 ( 
.A(n_1689),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1722),
.B(n_1591),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1724),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1708),
.B(n_1586),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1724),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1738),
.B(n_1603),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1738),
.B(n_1603),
.Y(n_1773)
);

INVxp67_ASAP7_75t_L g1774 ( 
.A(n_1733),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1734),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1721),
.B(n_1611),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1727),
.Y(n_1777)
);

OAI31xp33_ASAP7_75t_L g1778 ( 
.A1(n_1757),
.A2(n_1714),
.A3(n_1681),
.B(n_1705),
.Y(n_1778)
);

INVxp67_ASAP7_75t_SL g1779 ( 
.A(n_1752),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1756),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1756),
.B(n_1743),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1766),
.B(n_1743),
.Y(n_1782)
);

INVx3_ASAP7_75t_L g1783 ( 
.A(n_1759),
.Y(n_1783)
);

INVx2_ASAP7_75t_SL g1784 ( 
.A(n_1759),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1753),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1775),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1766),
.B(n_1768),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1755),
.B(n_1732),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1775),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1750),
.B(n_1699),
.Y(n_1790)
);

AO21x2_ASAP7_75t_L g1791 ( 
.A1(n_1748),
.A2(n_1694),
.B(n_1700),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_SL g1792 ( 
.A1(n_1752),
.A2(n_1699),
.B1(n_1692),
.B2(n_1744),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1753),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1755),
.B(n_1732),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1747),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1755),
.B(n_1721),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1758),
.B(n_1736),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1750),
.B(n_1713),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1766),
.B(n_1733),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1775),
.Y(n_1800)
);

OAI221xp5_ASAP7_75t_L g1801 ( 
.A1(n_1757),
.A2(n_1693),
.B1(n_1706),
.B2(n_1702),
.C(n_1714),
.Y(n_1801)
);

INVx2_ASAP7_75t_SL g1802 ( 
.A(n_1759),
.Y(n_1802)
);

INVx2_ASAP7_75t_SL g1803 ( 
.A(n_1759),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1769),
.Y(n_1804)
);

OAI22xp5_ASAP7_75t_SL g1805 ( 
.A1(n_1752),
.A2(n_1741),
.B1(n_1685),
.B2(n_1725),
.Y(n_1805)
);

OAI22xp5_ASAP7_75t_L g1806 ( 
.A1(n_1761),
.A2(n_1717),
.B1(n_1691),
.B2(n_1716),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1747),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1749),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1758),
.B(n_1715),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1760),
.B(n_1715),
.Y(n_1810)
);

INVxp67_ASAP7_75t_SL g1811 ( 
.A(n_1752),
.Y(n_1811)
);

OAI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1763),
.A2(n_1709),
.B(n_1711),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1760),
.B(n_1740),
.Y(n_1813)
);

BUFx2_ASAP7_75t_L g1814 ( 
.A(n_1752),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1749),
.Y(n_1815)
);

HB1xp67_ASAP7_75t_L g1816 ( 
.A(n_1777),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1760),
.B(n_1740),
.Y(n_1817)
);

NAND2x1_ASAP7_75t_L g1818 ( 
.A(n_1751),
.B(n_1728),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1762),
.B(n_1745),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1768),
.B(n_1709),
.Y(n_1820)
);

INVxp67_ASAP7_75t_L g1821 ( 
.A(n_1777),
.Y(n_1821)
);

BUFx3_ASAP7_75t_L g1822 ( 
.A(n_1754),
.Y(n_1822)
);

OAI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1763),
.A2(n_1711),
.B(n_1688),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1768),
.B(n_1735),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1795),
.Y(n_1825)
);

HB1xp67_ASAP7_75t_L g1826 ( 
.A(n_1804),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1787),
.B(n_1761),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1814),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1795),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1821),
.B(n_1769),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1807),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1807),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1788),
.B(n_1752),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1788),
.B(n_1752),
.Y(n_1834)
);

HB1xp67_ASAP7_75t_L g1835 ( 
.A(n_1804),
.Y(n_1835)
);

INVx1_ASAP7_75t_SL g1836 ( 
.A(n_1822),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1814),
.Y(n_1837)
);

INVxp67_ASAP7_75t_L g1838 ( 
.A(n_1816),
.Y(n_1838)
);

NAND2x1p5_ASAP7_75t_L g1839 ( 
.A(n_1818),
.B(n_1759),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1788),
.B(n_1764),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_SL g1841 ( 
.A(n_1812),
.B(n_1746),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1821),
.Y(n_1842)
);

HB1xp67_ASAP7_75t_L g1843 ( 
.A(n_1785),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_SL g1844 ( 
.A(n_1812),
.B(n_1774),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1808),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1794),
.B(n_1764),
.Y(n_1846)
);

NOR2x1_ASAP7_75t_L g1847 ( 
.A(n_1818),
.B(n_1741),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1794),
.B(n_1764),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1794),
.B(n_1745),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1808),
.Y(n_1850)
);

INVx3_ASAP7_75t_L g1851 ( 
.A(n_1783),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1819),
.B(n_1745),
.Y(n_1852)
);

INVx3_ASAP7_75t_L g1853 ( 
.A(n_1783),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1819),
.B(n_1796),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1787),
.B(n_1771),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1819),
.B(n_1772),
.Y(n_1856)
);

HB1xp67_ASAP7_75t_L g1857 ( 
.A(n_1785),
.Y(n_1857)
);

INVxp67_ASAP7_75t_L g1858 ( 
.A(n_1781),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1815),
.Y(n_1859)
);

AOI211xp5_ASAP7_75t_L g1860 ( 
.A1(n_1778),
.A2(n_1684),
.B(n_1730),
.C(n_1685),
.Y(n_1860)
);

BUFx3_ASAP7_75t_L g1861 ( 
.A(n_1822),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1796),
.B(n_1809),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1796),
.B(n_1772),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1793),
.B(n_1771),
.Y(n_1864)
);

INVx1_ASAP7_75t_SL g1865 ( 
.A(n_1822),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1793),
.B(n_1780),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1809),
.B(n_1772),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1809),
.B(n_1773),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1815),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1781),
.B(n_1765),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1810),
.B(n_1797),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1780),
.B(n_1824),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1854),
.B(n_1810),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1828),
.Y(n_1874)
);

INVxp67_ASAP7_75t_L g1875 ( 
.A(n_1841),
.Y(n_1875)
);

NAND2x1p5_ASAP7_75t_L g1876 ( 
.A(n_1847),
.B(n_1783),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1854),
.B(n_1810),
.Y(n_1877)
);

OAI21xp33_ASAP7_75t_L g1878 ( 
.A1(n_1844),
.A2(n_1782),
.B(n_1820),
.Y(n_1878)
);

OAI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1841),
.A2(n_1778),
.B(n_1820),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1828),
.Y(n_1880)
);

INVxp33_ASAP7_75t_L g1881 ( 
.A(n_1847),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1870),
.B(n_1782),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1858),
.B(n_1824),
.Y(n_1883)
);

INVx2_ASAP7_75t_SL g1884 ( 
.A(n_1861),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1825),
.Y(n_1885)
);

AOI211xp5_ASAP7_75t_SL g1886 ( 
.A1(n_1860),
.A2(n_1805),
.B(n_1701),
.C(n_1806),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1858),
.B(n_1844),
.Y(n_1887)
);

NAND2xp33_ASAP7_75t_L g1888 ( 
.A(n_1842),
.B(n_1805),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1854),
.B(n_1813),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1838),
.B(n_1842),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1825),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1825),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1829),
.Y(n_1893)
);

AND2x4_ASAP7_75t_L g1894 ( 
.A(n_1862),
.B(n_1783),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1829),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1838),
.B(n_1799),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1862),
.B(n_1813),
.Y(n_1897)
);

NOR2xp33_ASAP7_75t_L g1898 ( 
.A(n_1836),
.B(n_1767),
.Y(n_1898)
);

BUFx3_ASAP7_75t_L g1899 ( 
.A(n_1861),
.Y(n_1899)
);

AOI211xp5_ASAP7_75t_L g1900 ( 
.A1(n_1860),
.A2(n_1806),
.B(n_1801),
.C(n_1823),
.Y(n_1900)
);

OAI21xp33_ASAP7_75t_L g1901 ( 
.A1(n_1833),
.A2(n_1811),
.B(n_1779),
.Y(n_1901)
);

OR2x2_ASAP7_75t_L g1902 ( 
.A(n_1870),
.B(n_1798),
.Y(n_1902)
);

OR2x2_ASAP7_75t_L g1903 ( 
.A(n_1870),
.B(n_1827),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1829),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1828),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1832),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1862),
.B(n_1813),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1832),
.Y(n_1908)
);

AND2x4_ASAP7_75t_L g1909 ( 
.A(n_1863),
.B(n_1784),
.Y(n_1909)
);

INVxp67_ASAP7_75t_L g1910 ( 
.A(n_1861),
.Y(n_1910)
);

OR2x2_ASAP7_75t_L g1911 ( 
.A(n_1827),
.B(n_1798),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1840),
.B(n_1817),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1840),
.B(n_1799),
.Y(n_1913)
);

INVx3_ASAP7_75t_L g1914 ( 
.A(n_1839),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1840),
.B(n_1791),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1846),
.B(n_1817),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1846),
.B(n_1791),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1832),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1846),
.B(n_1791),
.Y(n_1919)
);

INVx1_ASAP7_75t_SL g1920 ( 
.A(n_1899),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1885),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1873),
.B(n_1856),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1875),
.B(n_1836),
.Y(n_1923)
);

INVx1_ASAP7_75t_SL g1924 ( 
.A(n_1899),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1885),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1909),
.Y(n_1926)
);

INVxp67_ASAP7_75t_L g1927 ( 
.A(n_1898),
.Y(n_1927)
);

NAND2xp33_ASAP7_75t_L g1928 ( 
.A(n_1887),
.B(n_1865),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1882),
.B(n_1872),
.Y(n_1929)
);

NOR2x1p5_ASAP7_75t_L g1930 ( 
.A(n_1896),
.B(n_1861),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1891),
.Y(n_1931)
);

AND2x4_ASAP7_75t_L g1932 ( 
.A(n_1873),
.B(n_1863),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1879),
.B(n_1848),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1909),
.Y(n_1934)
);

OR2x6_ASAP7_75t_L g1935 ( 
.A(n_1884),
.B(n_1823),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1878),
.B(n_1848),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1877),
.B(n_1856),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1891),
.Y(n_1938)
);

OR2x2_ASAP7_75t_L g1939 ( 
.A(n_1882),
.B(n_1872),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1909),
.Y(n_1940)
);

OAI21xp33_ASAP7_75t_L g1941 ( 
.A1(n_1900),
.A2(n_1834),
.B(n_1833),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1883),
.B(n_1848),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1913),
.B(n_1863),
.Y(n_1943)
);

INVxp67_ASAP7_75t_SL g1944 ( 
.A(n_1888),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1877),
.B(n_1856),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1910),
.B(n_1865),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1890),
.B(n_1849),
.Y(n_1947)
);

INVx3_ASAP7_75t_L g1948 ( 
.A(n_1894),
.Y(n_1948)
);

INVx1_ASAP7_75t_SL g1949 ( 
.A(n_1903),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1906),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1912),
.B(n_1852),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1912),
.Y(n_1952)
);

INVx1_ASAP7_75t_SL g1953 ( 
.A(n_1903),
.Y(n_1953)
);

INVx2_ASAP7_75t_SL g1954 ( 
.A(n_1894),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1906),
.Y(n_1955)
);

OR2x2_ASAP7_75t_L g1956 ( 
.A(n_1902),
.B(n_1872),
.Y(n_1956)
);

OAI21xp33_ASAP7_75t_L g1957 ( 
.A1(n_1886),
.A2(n_1834),
.B(n_1833),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1908),
.Y(n_1958)
);

AOI33xp33_ASAP7_75t_L g1959 ( 
.A1(n_1949),
.A2(n_1953),
.A3(n_1924),
.B1(n_1920),
.B2(n_1931),
.B3(n_1958),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1931),
.Y(n_1960)
);

NAND2xp33_ASAP7_75t_R g1961 ( 
.A(n_1935),
.B(n_1914),
.Y(n_1961)
);

OAI222xp33_ASAP7_75t_L g1962 ( 
.A1(n_1933),
.A2(n_1801),
.B1(n_1919),
.B2(n_1917),
.C1(n_1915),
.C2(n_1792),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1923),
.B(n_1849),
.Y(n_1963)
);

AOI22xp5_ASAP7_75t_L g1964 ( 
.A1(n_1944),
.A2(n_1791),
.B1(n_1792),
.B2(n_1888),
.Y(n_1964)
);

AOI22xp5_ASAP7_75t_L g1965 ( 
.A1(n_1957),
.A2(n_1935),
.B1(n_1941),
.B2(n_1928),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1938),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1938),
.Y(n_1967)
);

AOI221xp5_ASAP7_75t_L g1968 ( 
.A1(n_1928),
.A2(n_1834),
.B1(n_1881),
.B2(n_1811),
.C(n_1779),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1958),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1921),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1925),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1950),
.Y(n_1972)
);

O2A1O1Ixp33_ASAP7_75t_L g1973 ( 
.A1(n_1935),
.A2(n_1835),
.B(n_1826),
.C(n_1901),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1932),
.B(n_1916),
.Y(n_1974)
);

AOI211xp5_ASAP7_75t_L g1975 ( 
.A1(n_1936),
.A2(n_1914),
.B(n_1827),
.C(n_1826),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1927),
.B(n_1884),
.Y(n_1976)
);

AOI222xp33_ASAP7_75t_L g1977 ( 
.A1(n_1942),
.A2(n_1849),
.B1(n_1830),
.B2(n_1776),
.C1(n_1835),
.C2(n_1748),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1955),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1956),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1932),
.B(n_1916),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1929),
.B(n_1897),
.Y(n_1981)
);

NAND2xp33_ASAP7_75t_SL g1982 ( 
.A(n_1930),
.B(n_1897),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1935),
.B(n_1902),
.Y(n_1983)
);

AOI22xp5_ASAP7_75t_L g1984 ( 
.A1(n_1932),
.A2(n_1703),
.B1(n_1695),
.B2(n_1687),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1922),
.B(n_1907),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1929),
.B(n_1907),
.Y(n_1986)
);

AO22x1_ASAP7_75t_L g1987 ( 
.A1(n_1946),
.A2(n_1894),
.B1(n_1914),
.B2(n_1889),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1974),
.B(n_1954),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1960),
.Y(n_1989)
);

HB1xp67_ASAP7_75t_L g1990 ( 
.A(n_1976),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1966),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1980),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1967),
.Y(n_1993)
);

AOI322xp5_ASAP7_75t_L g1994 ( 
.A1(n_1964),
.A2(n_1947),
.A3(n_1943),
.B1(n_1922),
.B2(n_1937),
.C1(n_1852),
.C2(n_1952),
.Y(n_1994)
);

OR2x2_ASAP7_75t_L g1995 ( 
.A(n_1981),
.B(n_1956),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1983),
.B(n_1939),
.Y(n_1996)
);

OAI311xp33_ASAP7_75t_L g1997 ( 
.A1(n_1965),
.A2(n_1939),
.A3(n_1948),
.B1(n_1937),
.C1(n_1911),
.Y(n_1997)
);

OAI22xp5_ASAP7_75t_L g1998 ( 
.A1(n_1975),
.A2(n_1876),
.B1(n_1945),
.B2(n_1952),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1985),
.B(n_1954),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1969),
.Y(n_2000)
);

AOI22xp5_ASAP7_75t_L g2001 ( 
.A1(n_1984),
.A2(n_1687),
.B1(n_1940),
.B2(n_1934),
.Y(n_2001)
);

AOI22xp33_ASAP7_75t_L g2002 ( 
.A1(n_1983),
.A2(n_1940),
.B1(n_1934),
.B2(n_1926),
.Y(n_2002)
);

OR2x2_ASAP7_75t_L g2003 ( 
.A(n_1986),
.B(n_1911),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1979),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1976),
.B(n_1945),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1970),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1959),
.B(n_1963),
.Y(n_2007)
);

OR2x2_ASAP7_75t_L g2008 ( 
.A(n_1971),
.B(n_1945),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1972),
.Y(n_2009)
);

AOI222xp33_ASAP7_75t_L g2010 ( 
.A1(n_1962),
.A2(n_1830),
.B1(n_1776),
.B2(n_1748),
.C1(n_1874),
.C2(n_1905),
.Y(n_2010)
);

OR2x2_ASAP7_75t_L g2011 ( 
.A(n_1995),
.B(n_1951),
.Y(n_2011)
);

INVx2_ASAP7_75t_SL g2012 ( 
.A(n_2005),
.Y(n_2012)
);

AOI21xp5_ASAP7_75t_L g2013 ( 
.A1(n_1997),
.A2(n_1973),
.B(n_1982),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_2003),
.Y(n_2014)
);

AOI21xp5_ASAP7_75t_L g2015 ( 
.A1(n_2007),
.A2(n_1990),
.B(n_1996),
.Y(n_2015)
);

AOI21xp33_ASAP7_75t_L g2016 ( 
.A1(n_2010),
.A2(n_1961),
.B(n_2002),
.Y(n_2016)
);

INVx1_ASAP7_75t_SL g2017 ( 
.A(n_2005),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1999),
.B(n_1959),
.Y(n_2018)
);

AOI222xp33_ASAP7_75t_L g2019 ( 
.A1(n_2004),
.A2(n_1968),
.B1(n_1978),
.B2(n_1987),
.C1(n_1961),
.C2(n_1880),
.Y(n_2019)
);

NOR2xp33_ASAP7_75t_R g2020 ( 
.A(n_1988),
.B(n_1948),
.Y(n_2020)
);

AOI21xp5_ASAP7_75t_L g2021 ( 
.A1(n_1998),
.A2(n_1926),
.B(n_1948),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_2003),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1995),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1999),
.B(n_1951),
.Y(n_2024)
);

O2A1O1Ixp5_ASAP7_75t_L g2025 ( 
.A1(n_1992),
.A2(n_1874),
.B(n_1880),
.C(n_1905),
.Y(n_2025)
);

OAI21xp5_ASAP7_75t_SL g2026 ( 
.A1(n_2002),
.A2(n_1977),
.B(n_1876),
.Y(n_2026)
);

NOR2xp67_ASAP7_75t_L g2027 ( 
.A(n_2012),
.B(n_1992),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_2011),
.Y(n_2028)
);

OAI21xp5_ASAP7_75t_L g2029 ( 
.A1(n_2013),
.A2(n_1994),
.B(n_1988),
.Y(n_2029)
);

NOR2xp33_ASAP7_75t_L g2030 ( 
.A(n_2017),
.B(n_2008),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_2024),
.Y(n_2031)
);

NOR3xp33_ASAP7_75t_L g2032 ( 
.A(n_2015),
.B(n_2009),
.C(n_2006),
.Y(n_2032)
);

NAND5xp2_ASAP7_75t_L g2033 ( 
.A(n_2019),
.B(n_1989),
.C(n_2000),
.D(n_1993),
.E(n_1991),
.Y(n_2033)
);

OAI21xp5_ASAP7_75t_L g2034 ( 
.A1(n_2016),
.A2(n_2001),
.B(n_2008),
.Y(n_2034)
);

AOI21xp33_ASAP7_75t_SL g2035 ( 
.A1(n_2018),
.A2(n_1876),
.B(n_1839),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2014),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_2022),
.B(n_2023),
.Y(n_2037)
);

NOR3xp33_ASAP7_75t_L g2038 ( 
.A(n_2026),
.B(n_2025),
.C(n_2021),
.Y(n_2038)
);

NOR3xp33_ASAP7_75t_L g2039 ( 
.A(n_2026),
.B(n_1683),
.C(n_1908),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_2020),
.B(n_1889),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_2024),
.B(n_1843),
.Y(n_2041)
);

OAI211xp5_ASAP7_75t_SL g2042 ( 
.A1(n_2013),
.A2(n_1853),
.B(n_1851),
.C(n_1918),
.Y(n_2042)
);

NOR2xp33_ASAP7_75t_L g2043 ( 
.A(n_2017),
.B(n_1851),
.Y(n_2043)
);

AOI221xp5_ASAP7_75t_L g2044 ( 
.A1(n_2033),
.A2(n_1918),
.B1(n_1904),
.B2(n_1895),
.C(n_1893),
.Y(n_2044)
);

AND4x1_ASAP7_75t_L g2045 ( 
.A(n_2030),
.B(n_1682),
.C(n_1868),
.D(n_1867),
.Y(n_2045)
);

AND5x1_ASAP7_75t_L g2046 ( 
.A(n_2038),
.B(n_1701),
.C(n_1718),
.D(n_1742),
.E(n_1737),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_2031),
.B(n_1852),
.Y(n_2047)
);

OAI21xp33_ASAP7_75t_SL g2048 ( 
.A1(n_2029),
.A2(n_1892),
.B(n_1853),
.Y(n_2048)
);

AOI211xp5_ASAP7_75t_L g2049 ( 
.A1(n_2038),
.A2(n_1739),
.B(n_1855),
.C(n_1828),
.Y(n_2049)
);

AOI221xp5_ASAP7_75t_L g2050 ( 
.A1(n_2034),
.A2(n_1864),
.B1(n_1855),
.B2(n_1843),
.C(n_1857),
.Y(n_2050)
);

OAI221xp5_ASAP7_75t_SL g2051 ( 
.A1(n_2039),
.A2(n_2032),
.B1(n_2037),
.B2(n_2036),
.C(n_2028),
.Y(n_2051)
);

OAI221xp5_ASAP7_75t_L g2052 ( 
.A1(n_2046),
.A2(n_2042),
.B1(n_2035),
.B2(n_2027),
.C(n_2040),
.Y(n_2052)
);

OAI211xp5_ASAP7_75t_SL g2053 ( 
.A1(n_2048),
.A2(n_2043),
.B(n_2041),
.C(n_1851),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_2047),
.B(n_1871),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_2045),
.B(n_1857),
.Y(n_2055)
);

HB1xp67_ASAP7_75t_L g2056 ( 
.A(n_2051),
.Y(n_2056)
);

AOI322xp5_ASAP7_75t_L g2057 ( 
.A1(n_2050),
.A2(n_1868),
.A3(n_1867),
.B1(n_1837),
.B2(n_1864),
.C1(n_1774),
.C2(n_1770),
.Y(n_2057)
);

AOI22xp5_ASAP7_75t_L g2058 ( 
.A1(n_2049),
.A2(n_1855),
.B1(n_1868),
.B2(n_1867),
.Y(n_2058)
);

OAI221xp5_ASAP7_75t_L g2059 ( 
.A1(n_2044),
.A2(n_1839),
.B1(n_1837),
.B2(n_1851),
.C(n_1853),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2054),
.Y(n_2060)
);

INVx1_ASAP7_75t_SL g2061 ( 
.A(n_2056),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_2055),
.B(n_1837),
.Y(n_2062)
);

AND2x4_ASAP7_75t_L g2063 ( 
.A(n_2058),
.B(n_1851),
.Y(n_2063)
);

NOR3xp33_ASAP7_75t_L g2064 ( 
.A(n_2052),
.B(n_2053),
.C(n_2059),
.Y(n_2064)
);

NAND2x1p5_ASAP7_75t_L g2065 ( 
.A(n_2057),
.B(n_1853),
.Y(n_2065)
);

NAND4xp75_ASAP7_75t_L g2066 ( 
.A(n_2055),
.B(n_1837),
.C(n_1784),
.D(n_1802),
.Y(n_2066)
);

OAI321xp33_ASAP7_75t_L g2067 ( 
.A1(n_2062),
.A2(n_1839),
.A3(n_1790),
.B1(n_1866),
.B2(n_1803),
.C(n_1784),
.Y(n_2067)
);

AOI22x1_ASAP7_75t_L g2068 ( 
.A1(n_2060),
.A2(n_1853),
.B1(n_1845),
.B2(n_1859),
.Y(n_2068)
);

AOI322xp5_ASAP7_75t_L g2069 ( 
.A1(n_2061),
.A2(n_1770),
.A3(n_1773),
.B1(n_1866),
.B2(n_1786),
.C1(n_1800),
.C2(n_1789),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_2069),
.B(n_2064),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2070),
.Y(n_2071)
);

OAI22xp5_ASAP7_75t_L g2072 ( 
.A1(n_2071),
.A2(n_2066),
.B1(n_2065),
.B2(n_2063),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_2071),
.Y(n_2073)
);

CKINVDCx20_ASAP7_75t_R g2074 ( 
.A(n_2073),
.Y(n_2074)
);

NOR2xp67_ASAP7_75t_L g2075 ( 
.A(n_2072),
.B(n_2067),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_2074),
.Y(n_2076)
);

AOI22xp5_ASAP7_75t_L g2077 ( 
.A1(n_2075),
.A2(n_2068),
.B1(n_1871),
.B2(n_1859),
.Y(n_2077)
);

OAI222xp33_ASAP7_75t_L g2078 ( 
.A1(n_2076),
.A2(n_1845),
.B1(n_1859),
.B2(n_1850),
.C1(n_1869),
.C2(n_1831),
.Y(n_2078)
);

AOI21xp33_ASAP7_75t_L g2079 ( 
.A1(n_2078),
.A2(n_2077),
.B(n_1790),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2079),
.Y(n_2080)
);

OAI221xp5_ASAP7_75t_R g2081 ( 
.A1(n_2080),
.A2(n_1704),
.B1(n_1850),
.B2(n_1845),
.C(n_1871),
.Y(n_2081)
);

AOI211xp5_ASAP7_75t_L g2082 ( 
.A1(n_2081),
.A2(n_1621),
.B(n_1623),
.C(n_1850),
.Y(n_2082)
);


endmodule