module fake_jpeg_29774_n_63 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_63);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_63;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_48;
wire n_35;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_7),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx12_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_9),
.A2(n_11),
.B1(n_16),
.B2(n_13),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_20),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_6),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_6),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_13),
.B(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_21),
.B(n_12),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_21),
.B(n_8),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_24),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_20),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_29),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_15),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_25),
.A2(n_17),
.B1(n_9),
.B2(n_11),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_14),
.B(n_12),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_23),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_SL g40 ( 
.A(n_34),
.B(n_12),
.C(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_16),
.C(n_11),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_14),
.C(n_10),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_14),
.B1(n_27),
.B2(n_3),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_48),
.B1(n_37),
.B2(n_2),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_45),
.B(n_47),
.Y(n_50)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_39),
.B1(n_42),
.B2(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_52),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_44),
.B(n_42),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_45),
.C(n_10),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_50),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_56),
.C(n_10),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_55),
.A2(n_51),
.B(n_53),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_1),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_61),
.B(n_60),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_5),
.Y(n_63)
);


endmodule