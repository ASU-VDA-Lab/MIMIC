module fake_jpeg_18277_n_161 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_161);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_161;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx8_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_31),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_0),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

INVx6_ASAP7_75t_SL g69 ( 
.A(n_30),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_34),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_5),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_52),
.B1(n_61),
.B2(n_75),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_0),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_77),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NAND2xp33_ASAP7_75t_SL g94 ( 
.A(n_83),
.B(n_84),
.Y(n_94)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_89),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_77),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_92),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_82),
.Y(n_89)
);

AND2x4_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_49),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_90),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_83),
.A2(n_55),
.B1(n_66),
.B2(n_62),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_101),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_60),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_103),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_70),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_90),
.B(n_74),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_104),
.B(n_107),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_80),
.B1(n_53),
.B2(n_73),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_106),
.A2(n_95),
.B1(n_51),
.B2(n_72),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_109),
.B(n_110),
.Y(n_111)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_114),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_72),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_67),
.C(n_76),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_3),
.C(n_4),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_101),
.A2(n_71),
.B(n_54),
.C(n_58),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_122),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_SL g117 ( 
.A1(n_98),
.A2(n_82),
.B(n_52),
.C(n_59),
.Y(n_117)
);

AO21x2_ASAP7_75t_L g129 ( 
.A1(n_117),
.A2(n_2),
.B(n_3),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_73),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_50),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_123),
.B(n_124),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_1),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_110),
.B(n_69),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_127),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_105),
.A2(n_68),
.B1(n_64),
.B2(n_28),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_126),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_1),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_129),
.A2(n_130),
.B1(n_139),
.B2(n_121),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_25),
.B1(n_46),
.B2(n_45),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_119),
.Y(n_141)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_135),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_6),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_113),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_140),
.A2(n_143),
.B1(n_137),
.B2(n_129),
.Y(n_147)
);

OA21x2_ASAP7_75t_SL g148 ( 
.A1(n_141),
.A2(n_142),
.B(n_116),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_128),
.B(n_138),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_130),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_146),
.A2(n_129),
.B(n_117),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_140),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_151),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_144),
.C(n_145),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_12),
.C(n_13),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_14),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_17),
.B(n_22),
.Y(n_156)
);

AOI21x1_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_24),
.B(n_29),
.Y(n_157)
);

AO21x1_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_32),
.B(n_33),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_35),
.B1(n_39),
.B2(n_41),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_159),
.B(n_42),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_43),
.Y(n_161)
);


endmodule