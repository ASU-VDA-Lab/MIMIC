module fake_jpeg_1352_n_58 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_58);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_0),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_1),
.Y(n_28)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_30),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_25),
.B1(n_18),
.B2(n_22),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_35),
.Y(n_38)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_24),
.B(n_16),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_1),
.B(n_2),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_18),
.B1(n_19),
.B2(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_26),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_7),
.C(n_13),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_34),
.B1(n_19),
.B2(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_43),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_40),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_44),
.B(n_5),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_6),
.Y(n_45)
);

XOR2x2_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_2),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_50),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_48),
.B(n_11),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_3),
.C(n_4),
.Y(n_51)
);

NAND2xp33_ASAP7_75t_R g50 ( 
.A(n_45),
.B(n_9),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_53),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_52),
.A2(n_46),
.B(n_50),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_54),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_15),
.Y(n_58)
);


endmodule