module fake_jpeg_6466_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_38),
.Y(n_49)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_45),
.Y(n_54)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_21),
.B1(n_20),
.B2(n_31),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_52),
.A2(n_19),
.B1(n_22),
.B2(n_23),
.Y(n_85)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_61),
.Y(n_80)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_29),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_27),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_37),
.B(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_64),
.Y(n_94)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_72),
.B1(n_30),
.B2(n_26),
.Y(n_83)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_38),
.Y(n_70)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_21),
.B1(n_30),
.B2(n_24),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_41),
.B(n_28),
.Y(n_73)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_78),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_77),
.B(n_27),
.Y(n_130)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_46),
.B1(n_43),
.B2(n_47),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_79),
.A2(n_83),
.B1(n_85),
.B2(n_96),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_50),
.A2(n_41),
.B1(n_46),
.B2(n_38),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_84),
.B(n_62),
.C(n_29),
.Y(n_127)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_88),
.Y(n_118)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_90),
.Y(n_120)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_92),
.Y(n_128)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_59),
.A2(n_41),
.B1(n_22),
.B2(n_31),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_100),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_77),
.B(n_60),
.Y(n_102)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_94),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_103),
.Y(n_143)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_106),
.Y(n_133)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_80),
.A2(n_100),
.B(n_84),
.C(n_76),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_110),
.A2(n_29),
.B(n_55),
.Y(n_148)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

INVxp67_ASAP7_75t_SL g140 ( 
.A(n_111),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_114),
.B(n_119),
.Y(n_157)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_68),
.B1(n_54),
.B2(n_49),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_116),
.A2(n_24),
.B1(n_26),
.B2(n_28),
.Y(n_135)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_121),
.B(n_122),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_99),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_82),
.Y(n_123)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_90),
.B(n_39),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_25),
.C(n_67),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_86),
.B(n_64),
.Y(n_125)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_25),
.B1(n_23),
.B2(n_26),
.Y(n_147)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_153),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_144),
.B1(n_130),
.B2(n_106),
.Y(n_165)
);

AOI22x1_ASAP7_75t_SL g136 ( 
.A1(n_124),
.A2(n_39),
.B1(n_55),
.B2(n_40),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

AND2x2_ASAP7_75t_SL g141 ( 
.A(n_108),
.B(n_74),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_141),
.A2(n_156),
.B(n_130),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_105),
.A2(n_116),
.B1(n_110),
.B2(n_127),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_150),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_148),
.A2(n_104),
.B1(n_111),
.B2(n_69),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_103),
.A2(n_42),
.B1(n_48),
.B2(n_40),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_149),
.A2(n_154),
.B1(n_117),
.B2(n_115),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_112),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_L g154 ( 
.A1(n_112),
.A2(n_42),
.B1(n_48),
.B2(n_40),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_155),
.B(n_158),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_123),
.A2(n_34),
.B(n_1),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_157),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_159),
.B(n_160),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_146),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_165),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_164),
.A2(n_187),
.B(n_145),
.Y(n_210)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_166),
.B(n_168),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_128),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_170),
.C(n_174),
.Y(n_192)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

INVx13_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_121),
.C(n_119),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_140),
.Y(n_171)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_131),
.Y(n_173)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_129),
.C(n_126),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_135),
.Y(n_175)
);

BUFx24_ASAP7_75t_SL g208 ( 
.A(n_175),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_176),
.A2(n_155),
.B1(n_152),
.B2(n_134),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_147),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_184),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_143),
.A2(n_109),
.B1(n_122),
.B2(n_114),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_179),
.A2(n_183),
.B1(n_145),
.B2(n_137),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_153),
.Y(n_180)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_180),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_137),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_181),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_182),
.Y(n_196)
);

OAI32xp33_ASAP7_75t_L g184 ( 
.A1(n_138),
.A2(n_113),
.A3(n_42),
.B1(n_48),
.B2(n_18),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_101),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_186),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_132),
.B(n_101),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_154),
.Y(n_189)
);

XOR2x2_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_190),
.Y(n_216)
);

AND2x2_ASAP7_75t_SL g190 ( 
.A(n_187),
.B(n_132),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_193),
.A2(n_204),
.B1(n_183),
.B2(n_173),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_164),
.A2(n_151),
.B(n_139),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_206),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_177),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_162),
.C(n_184),
.Y(n_221)
);

OAI32xp33_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_151),
.A3(n_134),
.B1(n_33),
.B2(n_35),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_210),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_186),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_213),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_172),
.A2(n_165),
.B1(n_174),
.B2(n_168),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_162),
.B(n_34),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_163),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_207),
.B(n_10),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_169),
.A2(n_58),
.B1(n_63),
.B2(n_51),
.Y(n_211)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_185),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_180),
.A2(n_142),
.B(n_101),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_35),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_201),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_217),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_197),
.B(n_204),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_218),
.B(n_221),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_208),
.B(n_178),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_219),
.B(n_228),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_212),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_220),
.B(n_229),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_225),
.A2(n_231),
.B1(n_238),
.B2(n_242),
.Y(n_261)
);

INVxp33_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_230),
.B(n_234),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_189),
.A2(n_107),
.B1(n_35),
.B2(n_33),
.Y(n_231)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_203),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_192),
.B(n_58),
.C(n_51),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_214),
.C(n_209),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_192),
.Y(n_245)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_200),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_239),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_189),
.A2(n_35),
.B1(n_33),
.B2(n_63),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_193),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_190),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_198),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_190),
.Y(n_241)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_241),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_191),
.A2(n_33),
.B1(n_1),
.B2(n_2),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_4),
.Y(n_275)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_246),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_223),
.A2(n_194),
.B1(n_210),
.B2(n_188),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_247),
.A2(n_249),
.B1(n_238),
.B2(n_226),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_250),
.C(n_0),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_216),
.A2(n_188),
.B1(n_214),
.B2(n_199),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_206),
.C(n_199),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_221),
.B(n_195),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_254),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_216),
.Y(n_257)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_257),
.Y(n_280)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_222),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_258),
.B(n_10),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_209),
.Y(n_260)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_225),
.A2(n_196),
.B1(n_1),
.B2(n_2),
.Y(n_262)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

AOI21xp33_ASAP7_75t_L g263 ( 
.A1(n_232),
.A2(n_8),
.B(n_15),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_263),
.B(n_5),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_0),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_242),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_244),
.A2(n_227),
.B1(n_224),
.B2(n_231),
.Y(n_266)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_266),
.Y(n_288)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_267),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_268),
.B(n_260),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_244),
.A2(n_226),
.B(n_235),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_269),
.A2(n_278),
.B(n_284),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_247),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_271)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_271),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_249),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_272)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_272),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_274),
.C(n_265),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_276),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_5),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_282),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_255),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_251),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_6),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_6),
.C(n_7),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_277),
.C(n_282),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_286),
.Y(n_312)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_287),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_245),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_268),
.Y(n_302)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_290),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_281),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_294),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_280),
.A2(n_253),
.B1(n_261),
.B2(n_252),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_292),
.A2(n_299),
.B1(n_293),
.B2(n_296),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_270),
.A2(n_264),
.B1(n_246),
.B2(n_243),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_298),
.A2(n_267),
.B1(n_283),
.B2(n_275),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_248),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_243),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_305),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_290),
.B(n_272),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_303),
.B(n_304),
.C(n_307),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_274),
.C(n_253),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_275),
.C(n_271),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_310),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_309),
.A2(n_7),
.B1(n_14),
.B2(n_15),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_259),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_6),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_313),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_7),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_303),
.B(n_288),
.Y(n_315)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_315),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_301),
.B(n_294),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_317),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_314),
.A2(n_295),
.B1(n_9),
.B2(n_11),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_304),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_321),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_308),
.A2(n_295),
.B1(n_13),
.B2(n_14),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_16),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_318),
.A2(n_306),
.B(n_305),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_328),
.A2(n_329),
.B(n_330),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_312),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_323),
.A2(n_311),
.B(n_14),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_315),
.Y(n_331)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_331),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_332),
.A2(n_322),
.B(n_319),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_334),
.B(n_336),
.Y(n_338)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_327),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_319),
.C(n_16),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_337),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_338),
.B(n_335),
.Y(n_340)
);

BUFx24_ASAP7_75t_SL g341 ( 
.A(n_340),
.Y(n_341)
);

BUFx24_ASAP7_75t_SL g342 ( 
.A(n_341),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_342),
.B(n_339),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_325),
.B(n_333),
.Y(n_344)
);


endmodule