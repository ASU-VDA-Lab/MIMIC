module fake_jpeg_30376_n_403 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_403);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_403;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_34),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_56),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_77),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_36),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_74),
.A2(n_30),
.B1(n_24),
.B2(n_23),
.Y(n_111)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_34),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_47),
.A2(n_44),
.B1(n_20),
.B2(n_21),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_86),
.A2(n_102),
.B1(n_44),
.B2(n_20),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_48),
.A2(n_44),
.B1(n_20),
.B2(n_21),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_60),
.A2(n_61),
.B1(n_58),
.B2(n_57),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_105),
.A2(n_111),
.B1(n_113),
.B2(n_30),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_31),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_31),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_22),
.C(n_40),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_32),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_73),
.A2(n_41),
.B1(n_25),
.B2(n_39),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_94),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_123),
.Y(n_159)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_122),
.Y(n_171)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_127),
.Y(n_164)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_126),
.Y(n_160)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

AOI22x1_ASAP7_75t_L g128 ( 
.A1(n_90),
.A2(n_67),
.B1(n_68),
.B2(n_51),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_128),
.A2(n_138),
.B1(n_120),
.B2(n_81),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

INVx3_ASAP7_75t_SL g183 ( 
.A(n_129),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_33),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_130),
.B(n_134),
.Y(n_173)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_139),
.B1(n_140),
.B2(n_155),
.Y(n_157)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_25),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_24),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_148),
.Y(n_158)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_86),
.A2(n_76),
.B1(n_62),
.B2(n_65),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_95),
.A2(n_63),
.B1(n_50),
.B2(n_52),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_83),
.A2(n_55),
.B1(n_49),
.B2(n_35),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_32),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_142),
.Y(n_174)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

INVx4_ASAP7_75t_SL g166 ( 
.A(n_146),
.Y(n_166)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_84),
.B(n_41),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_149),
.B(n_153),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_88),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_151),
.Y(n_163)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_154),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_39),
.Y(n_153)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

INVx11_ASAP7_75t_L g155 ( 
.A(n_112),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_161),
.A2(n_81),
.B1(n_120),
.B2(n_112),
.Y(n_204)
);

XNOR2x1_ASAP7_75t_SL g165 ( 
.A(n_146),
.B(n_72),
.Y(n_165)
);

XNOR2x1_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_128),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_118),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_175),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_118),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_131),
.B(n_114),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_181),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_114),
.Y(n_181)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_162),
.Y(n_187)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_173),
.B(n_164),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_188),
.B(n_189),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_163),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_172),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_192),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_175),
.B(n_130),
.Y(n_192)
);

OAI22x1_ASAP7_75t_SL g193 ( 
.A1(n_165),
.A2(n_128),
.B1(n_105),
.B2(n_144),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_166),
.B1(n_176),
.B2(n_157),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_181),
.A2(n_157),
.B1(n_166),
.B2(n_158),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_194),
.A2(n_204),
.B1(n_179),
.B2(n_170),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_195),
.B(n_206),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_196),
.Y(n_212)
);

FAx1_ASAP7_75t_SL g197 ( 
.A(n_158),
.B(n_135),
.CI(n_133),
.CON(n_197),
.SN(n_197)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_206),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_173),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_203),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_124),
.C(n_147),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_184),
.C(n_170),
.Y(n_214)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_163),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_205),
.A2(n_207),
.B1(n_162),
.B2(n_171),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_165),
.A2(n_122),
.B(n_152),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_210),
.A2(n_219),
.B1(n_221),
.B2(n_225),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_214),
.B(n_216),
.C(n_220),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_168),
.Y(n_216)
);

AOI322xp5_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_168),
.A3(n_174),
.B1(n_164),
.B2(n_161),
.C1(n_166),
.C2(n_157),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_233),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_202),
.A2(n_166),
.B(n_182),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_218),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_193),
.A2(n_82),
.B1(n_109),
.B2(n_155),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_184),
.C(n_182),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_208),
.A2(n_183),
.B1(n_143),
.B2(n_129),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_189),
.A2(n_178),
.B(n_160),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_222),
.A2(n_160),
.B(n_199),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_223),
.A2(n_69),
.B1(n_53),
.B2(n_78),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_224),
.B(n_228),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_208),
.A2(n_183),
.B1(n_179),
.B2(n_180),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_180),
.C(n_171),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_72),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_231),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_234),
.B(n_252),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_219),
.A2(n_194),
.B1(n_203),
.B2(n_205),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_236),
.A2(n_250),
.B1(n_254),
.B2(n_255),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_223),
.A2(n_207),
.B1(n_195),
.B2(n_197),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_237),
.A2(n_239),
.B1(n_240),
.B2(n_243),
.Y(n_278)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_238),
.Y(n_266)
);

OA22x2_ASAP7_75t_L g239 ( 
.A1(n_230),
.A2(n_197),
.B1(n_186),
.B2(n_185),
.Y(n_239)
);

OA22x2_ASAP7_75t_L g240 ( 
.A1(n_228),
.A2(n_186),
.B1(n_200),
.B2(n_171),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_241),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_242),
.A2(n_209),
.B(n_215),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_229),
.A2(n_198),
.B1(n_188),
.B2(n_183),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_244),
.Y(n_284)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_248),
.Y(n_267)
);

AND2x2_ASAP7_75t_SL g247 ( 
.A(n_224),
.B(n_201),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_247),
.Y(n_282)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_257),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_229),
.A2(n_183),
.B1(n_196),
.B2(n_187),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_216),
.B(n_213),
.Y(n_251)
);

NAND3xp33_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_29),
.C(n_40),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_167),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_231),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_253),
.B(n_259),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_227),
.A2(n_196),
.B1(n_160),
.B2(n_154),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_225),
.A2(n_160),
.B1(n_110),
.B2(n_104),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_221),
.A2(n_104),
.B1(n_137),
.B2(n_126),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_263),
.Y(n_279)
);

AOI22x1_ASAP7_75t_L g259 ( 
.A1(n_218),
.A2(n_148),
.B1(n_151),
.B2(n_144),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_261),
.A2(n_35),
.B1(n_29),
.B2(n_85),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_222),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_262),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_214),
.A2(n_212),
.B1(n_209),
.B2(n_232),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_232),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_264),
.B(n_275),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_215),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_286),
.C(n_287),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_248),
.B(n_33),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_271),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_256),
.A2(n_85),
.B(n_23),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_273),
.B(n_290),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_274),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_22),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_276),
.A2(n_236),
.B1(n_250),
.B2(n_255),
.Y(n_292)
);

NAND3xp33_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_12),
.C(n_18),
.Y(n_277)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_277),
.Y(n_295)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_259),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_281),
.Y(n_302)
);

XOR2x2_ASAP7_75t_L g283 ( 
.A(n_247),
.B(n_66),
.Y(n_283)
);

XNOR2x1_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_286),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_247),
.B(n_80),
.C(n_66),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_79),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_243),
.B(n_8),
.Y(n_289)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_289),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_256),
.A2(n_54),
.B(n_1),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_292),
.A2(n_303),
.B1(n_313),
.B2(n_283),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_281),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_293),
.B(n_304),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_294),
.B(n_268),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_280),
.A2(n_246),
.B1(n_271),
.B2(n_272),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_296),
.A2(n_306),
.B1(n_308),
.B2(n_310),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_263),
.C(n_242),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_311),
.C(n_268),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_278),
.A2(n_235),
.B1(n_288),
.B2(n_282),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_267),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_285),
.Y(n_305)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_305),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_280),
.A2(n_237),
.B1(n_254),
.B2(n_235),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_239),
.Y(n_307)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_307),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_279),
.A2(n_240),
.B1(n_239),
.B2(n_259),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_285),
.Y(n_309)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_309),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_266),
.A2(n_245),
.B1(n_244),
.B2(n_241),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_264),
.B(n_240),
.C(n_239),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_278),
.A2(n_265),
.B1(n_240),
.B2(n_290),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_275),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_314),
.B(n_321),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_315),
.B(n_323),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_316),
.A2(n_306),
.B1(n_308),
.B2(n_313),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_318),
.B(n_319),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_299),
.B(n_287),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_273),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_320),
.B(n_324),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_300),
.B(n_238),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_294),
.B(n_276),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_297),
.B(n_258),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_291),
.B(n_284),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_325),
.B(n_327),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_291),
.B(n_54),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_297),
.B(n_42),
.C(n_8),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_328),
.B(n_312),
.C(n_307),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_312),
.Y(n_329)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_329),
.Y(n_335)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_302),
.Y(n_330)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_330),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_301),
.B(n_8),
.Y(n_332)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_332),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_295),
.B(n_7),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_333),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_336),
.B(n_320),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_331),
.A2(n_312),
.B(n_302),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_337),
.A2(n_317),
.B(n_327),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_325),
.B(n_303),
.C(n_296),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_346),
.C(n_14),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_334),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_342),
.B(n_328),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_343),
.A2(n_13),
.B1(n_12),
.B2(n_9),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_322),
.A2(n_7),
.B1(n_18),
.B2(n_17),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_345),
.A2(n_348),
.B1(n_9),
.B2(n_1),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_318),
.B(n_42),
.C(n_17),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_324),
.A2(n_17),
.B1(n_14),
.B2(n_13),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_352),
.A2(n_355),
.B(n_357),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_353),
.B(n_354),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_340),
.B(n_326),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_347),
.B(n_319),
.Y(n_355)
);

OR2x2_ASAP7_75t_L g356 ( 
.A(n_335),
.B(n_323),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_356),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_347),
.B(n_315),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_358),
.A2(n_364),
.B(n_351),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_359),
.B(n_361),
.C(n_363),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_360),
.B(n_348),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_339),
.B(n_9),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_362),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_339),
.B(n_0),
.C(n_2),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_350),
.B(n_0),
.C(n_2),
.Y(n_364)
);

NOR2x1_ASAP7_75t_SL g365 ( 
.A(n_336),
.B(n_2),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_365),
.Y(n_373)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_367),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_355),
.B(n_338),
.Y(n_370)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_370),
.Y(n_384)
);

FAx1_ASAP7_75t_SL g371 ( 
.A(n_357),
.B(n_341),
.CI(n_350),
.CON(n_371),
.SN(n_371)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_371),
.B(n_341),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_375),
.B(n_3),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_356),
.A2(n_344),
.B1(n_359),
.B2(n_346),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_376),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_366),
.A2(n_363),
.B(n_364),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_377),
.B(n_379),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_378),
.B(n_381),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_370),
.A2(n_349),
.B(n_4),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_372),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_383),
.B(n_385),
.C(n_367),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_371),
.B(n_3),
.Y(n_385)
);

NOR2xp67_ASAP7_75t_SL g386 ( 
.A(n_369),
.B(n_3),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_386),
.B(n_369),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_384),
.B(n_373),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_387),
.A2(n_388),
.B(n_389),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_380),
.B(n_368),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_382),
.B(n_374),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_391),
.A2(n_393),
.B(n_5),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_387),
.A2(n_382),
.B(n_385),
.Y(n_395)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_395),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_390),
.A2(n_4),
.B(n_5),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_396),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_398),
.A2(n_394),
.B(n_397),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_400),
.A2(n_399),
.B(n_392),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_401),
.B(n_6),
.Y(n_402)
);

NAND2x1_ASAP7_75t_L g403 ( 
.A(n_402),
.B(n_6),
.Y(n_403)
);


endmodule