module fake_jpeg_31913_n_509 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_509);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_509;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_53),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_54),
.Y(n_152)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_55),
.Y(n_126)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_46),
.B(n_17),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_57),
.B(n_91),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_17),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_58),
.B(n_59),
.Y(n_104)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_61),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_22),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_63),
.Y(n_108)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_20),
.B(n_0),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_64),
.B(n_93),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_22),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_66),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_51),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_67),
.B(n_75),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_69),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_70),
.Y(n_158)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_72),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_73),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_41),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_76),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_78),
.B(n_80),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_79),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_26),
.B(n_16),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_81),
.B(n_83),
.Y(n_134)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_50),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_84),
.B(n_88),
.Y(n_137)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx11_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_87),
.Y(n_151)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

INVx6_ASAP7_75t_SL g91 ( 
.A(n_49),
.Y(n_91)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_29),
.Y(n_93)
);

OR2x2_ASAP7_75t_SL g94 ( 
.A(n_39),
.B(n_16),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_96),
.Y(n_138)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

INVx3_ASAP7_75t_SL g97 ( 
.A(n_33),
.Y(n_97)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_28),
.B(n_27),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_100),
.Y(n_148)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_28),
.B(n_15),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_21),
.Y(n_101)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_95),
.A2(n_49),
.B1(n_40),
.B2(n_44),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_107),
.A2(n_109),
.B1(n_112),
.B2(n_115),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_64),
.A2(n_49),
.B1(n_40),
.B2(n_33),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_91),
.A2(n_48),
.B1(n_44),
.B2(n_35),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_97),
.A2(n_48),
.B1(n_44),
.B2(n_35),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_58),
.B(n_36),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_116),
.B(n_132),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_48),
.B1(n_45),
.B2(n_26),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_117),
.A2(n_125),
.B1(n_131),
.B2(n_154),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_94),
.A2(n_27),
.B1(n_34),
.B2(n_36),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_119),
.B(n_142),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_80),
.B(n_45),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_121),
.B(n_128),
.Y(n_175)
);

BUFx4f_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_124),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_93),
.A2(n_43),
.B1(n_35),
.B2(n_38),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_71),
.B(n_42),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_89),
.A2(n_43),
.B1(n_35),
.B2(n_38),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_79),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_60),
.A2(n_30),
.B1(n_34),
.B2(n_42),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_55),
.B(n_30),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_156),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_82),
.A2(n_43),
.B1(n_86),
.B2(n_99),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_66),
.B(n_43),
.Y(n_156)
);

OA22x2_ASAP7_75t_L g157 ( 
.A1(n_92),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_157)
);

OA22x2_ASAP7_75t_L g173 ( 
.A1(n_157),
.A2(n_81),
.B1(n_2),
.B2(n_3),
.Y(n_173)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_160),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_67),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_161),
.B(n_162),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_104),
.B(n_56),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

INVx3_ASAP7_75t_SL g215 ( 
.A(n_164),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_70),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_165),
.B(n_167),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_117),
.A2(n_76),
.B1(n_90),
.B2(n_87),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_166),
.A2(n_173),
.B1(n_179),
.B2(n_202),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_70),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_122),
.B(n_73),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_168),
.Y(n_245)
);

NAND2xp33_ASAP7_75t_SL g169 ( 
.A(n_128),
.B(n_72),
.Y(n_169)
);

OAI21xp33_ASAP7_75t_L g238 ( 
.A1(n_169),
.A2(n_182),
.B(n_203),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_111),
.A2(n_106),
.B1(n_85),
.B2(n_96),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_170),
.A2(n_172),
.B1(n_135),
.B2(n_152),
.Y(n_225)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_111),
.Y(n_171)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_171),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_106),
.A2(n_96),
.B1(n_81),
.B2(n_72),
.Y(n_172)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_174),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_122),
.A2(n_69),
.B1(n_15),
.B2(n_74),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_179),
.B(n_184),
.Y(n_253)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_102),
.Y(n_180)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_180),
.Y(n_233)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_121),
.B(n_69),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_142),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_108),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_186),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_110),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_129),
.Y(n_187)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_187),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_141),
.Y(n_188)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_188),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_122),
.B(n_77),
.C(n_68),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_189),
.B(n_207),
.Y(n_235)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_134),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_192),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_127),
.B(n_54),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_105),
.B(n_53),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_195),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_138),
.B(n_109),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_194),
.B(n_202),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_119),
.B(n_0),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_129),
.Y(n_196)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_196),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_132),
.B(n_2),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_210),
.Y(n_229)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_118),
.Y(n_198)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_198),
.Y(n_232)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_102),
.Y(n_199)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_199),
.Y(n_256)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_118),
.Y(n_200)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_200),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_124),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_201),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_157),
.B(n_52),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_157),
.B(n_3),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_157),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_205),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_255)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_113),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_113),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_208),
.Y(n_250)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_114),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_209),
.B(n_158),
.Y(n_252)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_114),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_124),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_212),
.Y(n_240)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_133),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_184),
.A2(n_123),
.B1(n_103),
.B2(n_151),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_218),
.A2(n_230),
.B1(n_237),
.B2(n_239),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_224),
.A2(n_227),
.B1(n_231),
.B2(n_236),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_225),
.A2(n_144),
.B(n_188),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_194),
.A2(n_123),
.B1(n_103),
.B2(n_151),
.Y(n_227)
);

AO22x1_ASAP7_75t_SL g228 ( 
.A1(n_203),
.A2(n_163),
.B1(n_173),
.B2(n_169),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_228),
.B(n_248),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_204),
.A2(n_140),
.B1(n_120),
.B2(n_147),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_206),
.A2(n_139),
.B1(n_145),
.B2(n_140),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_206),
.A2(n_139),
.B1(n_145),
.B2(n_146),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_173),
.A2(n_147),
.B1(n_146),
.B2(n_133),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_173),
.A2(n_136),
.B1(n_149),
.B2(n_153),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_175),
.A2(n_126),
.B(n_152),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_241),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_189),
.A2(n_136),
.B1(n_149),
.B2(n_153),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_247),
.A2(n_144),
.B1(n_177),
.B2(n_183),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_198),
.B(n_126),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_200),
.B(n_171),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_181),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_255),
.A2(n_257),
.B1(n_168),
.B2(n_191),
.Y(n_275)
);

AO21x2_ASAP7_75t_L g257 ( 
.A1(n_203),
.A2(n_197),
.B(n_211),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_214),
.Y(n_259)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_259),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_244),
.B(n_249),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_260),
.B(n_263),
.Y(n_320)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_214),
.Y(n_262)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_262),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_244),
.B(n_175),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_232),
.Y(n_264)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_264),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_222),
.B(n_186),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_265),
.B(n_271),
.Y(n_328)
);

INVx8_ASAP7_75t_L g266 ( 
.A(n_213),
.Y(n_266)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_266),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_252),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_268),
.B(n_270),
.Y(n_317)
);

MAJx2_ASAP7_75t_L g269 ( 
.A(n_235),
.B(n_168),
.C(n_159),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_269),
.B(n_281),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_240),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_229),
.B(n_185),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_272),
.B(n_276),
.Y(n_319)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_232),
.Y(n_273)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_273),
.Y(n_332)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_233),
.Y(n_274)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_274),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_275),
.A2(n_294),
.B1(n_245),
.B2(n_224),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_176),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_242),
.B(n_196),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_277),
.B(n_285),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_251),
.Y(n_278)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_278),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_215),
.A2(n_178),
.B1(n_160),
.B2(n_135),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_279),
.Y(n_313)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_280),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_235),
.B(n_190),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_258),
.Y(n_282)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_282),
.Y(n_321)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_220),
.Y(n_284)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_284),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_248),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_216),
.B(n_209),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_286),
.Y(n_315)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_220),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_287),
.Y(n_325)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_221),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_289),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_223),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_290),
.A2(n_292),
.B(n_296),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_226),
.B(n_207),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_245),
.B(n_187),
.Y(n_293)
);

BUFx24_ASAP7_75t_SL g318 ( 
.A(n_293),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_227),
.A2(n_177),
.B1(n_212),
.B2(n_201),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_295),
.A2(n_298),
.B1(n_299),
.B2(n_243),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_241),
.B(n_210),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_297),
.A2(n_246),
.B1(n_243),
.B2(n_215),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_234),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_221),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_228),
.B(n_208),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_247),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_296),
.A2(n_253),
.B(n_225),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_302),
.A2(n_305),
.B(n_261),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_303),
.B(n_307),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_304),
.A2(n_335),
.B1(n_283),
.B2(n_284),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_267),
.A2(n_257),
.B(n_253),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_291),
.A2(n_253),
.B(n_257),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_310),
.A2(n_316),
.B(n_293),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_281),
.B(n_238),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_312),
.B(n_324),
.C(n_327),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_314),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_291),
.A2(n_267),
.B(n_300),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_269),
.B(n_228),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_269),
.B(n_228),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_263),
.B(n_231),
.C(n_236),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_331),
.B(n_333),
.C(n_270),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_260),
.B(n_250),
.C(n_246),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_275),
.A2(n_257),
.B1(n_255),
.B2(n_250),
.Y(n_335)
);

AO22x1_ASAP7_75t_L g336 ( 
.A1(n_285),
.A2(n_257),
.B1(n_215),
.B2(n_199),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_336),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_288),
.A2(n_257),
.B1(n_180),
.B2(n_217),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_337),
.B(n_283),
.Y(n_353)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_323),
.Y(n_339)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_339),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_340),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_334),
.B(n_271),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_343),
.B(n_351),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_328),
.B(n_290),
.Y(n_344)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_344),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_346),
.B(n_348),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_324),
.B(n_286),
.C(n_272),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_347),
.B(n_356),
.C(n_367),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_319),
.B(n_265),
.Y(n_349)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_349),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_315),
.B(n_292),
.Y(n_350)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_350),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_334),
.B(n_288),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_311),
.Y(n_352)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_352),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_353),
.A2(n_354),
.B1(n_355),
.B2(n_360),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_338),
.B(n_278),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_328),
.B(n_280),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_327),
.B(n_294),
.C(n_297),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_336),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_357),
.A2(n_302),
.B1(n_325),
.B2(n_329),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_311),
.Y(n_358)
);

INVxp33_ASAP7_75t_SL g386 ( 
.A(n_358),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_312),
.B(n_264),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_359),
.B(n_366),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_320),
.B(n_262),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_321),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g397 ( 
.A1(n_361),
.A2(n_254),
.B1(n_274),
.B2(n_256),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_320),
.B(n_282),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_362),
.A2(n_363),
.B1(n_365),
.B2(n_317),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_309),
.B(n_259),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_309),
.B(n_273),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_310),
.B(n_333),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_307),
.B(n_289),
.C(n_287),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_316),
.B(n_299),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_368),
.B(n_371),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_369),
.A2(n_337),
.B1(n_336),
.B2(n_303),
.Y(n_373)
);

XNOR2x1_ASAP7_75t_SL g370 ( 
.A(n_318),
.B(n_298),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_370),
.B(n_301),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_305),
.A2(n_266),
.B(n_251),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_373),
.A2(n_375),
.B1(n_391),
.B2(n_394),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_369),
.A2(n_304),
.B1(n_313),
.B2(n_335),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_376),
.B(n_372),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_353),
.A2(n_313),
.B1(n_331),
.B2(n_321),
.Y(n_378)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_378),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_383),
.B(n_398),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_345),
.A2(n_329),
.B1(n_325),
.B2(n_332),
.Y(n_384)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_384),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_341),
.B(n_326),
.C(n_322),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_385),
.B(n_393),
.C(n_396),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_345),
.A2(n_308),
.B1(n_330),
.B2(n_306),
.Y(n_387)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_387),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_389),
.B(n_6),
.Y(n_426)
);

BUFx5_ASAP7_75t_L g390 ( 
.A(n_364),
.Y(n_390)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_390),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_357),
.A2(n_330),
.B1(n_306),
.B2(n_301),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_341),
.B(n_219),
.C(n_213),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_363),
.A2(n_266),
.B1(n_217),
.B2(n_219),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_346),
.B(n_254),
.C(n_234),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_397),
.A2(n_342),
.B(n_360),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_340),
.A2(n_256),
.B1(n_233),
.B2(n_201),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_356),
.A2(n_164),
.B1(n_174),
.B2(n_183),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_401),
.A2(n_371),
.B1(n_364),
.B2(n_348),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_404),
.A2(n_413),
.B1(n_418),
.B2(n_401),
.Y(n_430)
);

BUFx24_ASAP7_75t_SL g405 ( 
.A(n_392),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_405),
.B(n_10),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_390),
.B(n_355),
.Y(n_408)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_408),
.Y(n_427)
);

NAND3xp33_ASAP7_75t_L g409 ( 
.A(n_388),
.B(n_365),
.C(n_370),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_409),
.B(n_420),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_377),
.B(n_351),
.C(n_366),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_410),
.B(n_422),
.C(n_425),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_381),
.B(n_347),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_414),
.B(n_417),
.Y(n_435)
);

CKINVDCx14_ASAP7_75t_R g436 ( 
.A(n_415),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_400),
.B(n_379),
.Y(n_416)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_416),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_381),
.B(n_343),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_399),
.A2(n_368),
.B1(n_342),
.B2(n_359),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_377),
.B(n_382),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_419),
.B(n_421),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_380),
.B(n_367),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_382),
.B(n_374),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_374),
.B(n_396),
.C(n_385),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_391),
.B(n_5),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_424),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_393),
.B(n_183),
.C(n_7),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_426),
.B(n_386),
.Y(n_440)
);

OA21x2_ASAP7_75t_L g428 ( 
.A1(n_402),
.A2(n_383),
.B(n_399),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_428),
.B(n_429),
.Y(n_447)
);

BUFx12_ASAP7_75t_L g429 ( 
.A(n_413),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_430),
.B(n_415),
.Y(n_449)
);

INVx13_ASAP7_75t_L g433 ( 
.A(n_423),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_433),
.B(n_440),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_417),
.B(n_395),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_434),
.B(n_439),
.Y(n_450)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_412),
.Y(n_437)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_437),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_414),
.B(n_395),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_406),
.A2(n_375),
.B1(n_389),
.B2(n_373),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_442),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_407),
.A2(n_398),
.B1(n_7),
.B2(n_8),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_443),
.A2(n_444),
.B1(n_408),
.B2(n_441),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_411),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_446),
.B(n_438),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_449),
.B(n_427),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_437),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_451),
.B(n_458),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_431),
.B(n_403),
.C(n_422),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_452),
.B(n_453),
.C(n_462),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_431),
.B(n_403),
.C(n_410),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_454),
.Y(n_469)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_455),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_445),
.B(n_419),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_456),
.B(n_457),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_429),
.A2(n_402),
.B(n_424),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_428),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_436),
.A2(n_418),
.B1(n_425),
.B2(n_421),
.Y(n_459)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_459),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_432),
.B(n_13),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_464),
.B(n_439),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_460),
.B(n_428),
.Y(n_465)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_465),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_457),
.B(n_455),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_468),
.B(n_476),
.Y(n_479)
);

OA21x2_ASAP7_75t_SL g470 ( 
.A1(n_447),
.A2(n_429),
.B(n_434),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_470),
.B(n_473),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_448),
.A2(n_461),
.B1(n_449),
.B2(n_459),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_471),
.A2(n_472),
.B1(n_475),
.B2(n_470),
.Y(n_488)
);

INVx11_ASAP7_75t_L g473 ( 
.A(n_448),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_452),
.B(n_432),
.C(n_435),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_474),
.A2(n_14),
.B(n_475),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_462),
.B(n_440),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_477),
.B(n_478),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_466),
.B(n_453),
.C(n_450),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_471),
.B(n_450),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_480),
.B(n_482),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_466),
.B(n_435),
.C(n_433),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_481),
.B(n_484),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_465),
.B(n_13),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_469),
.B(n_13),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_463),
.B(n_14),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_485),
.B(n_487),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_488),
.B(n_472),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_489),
.B(n_491),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_479),
.A2(n_463),
.B(n_467),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_490),
.B(n_464),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_483),
.B(n_469),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_480),
.A2(n_467),
.B(n_468),
.Y(n_494)
);

INVxp33_ASAP7_75t_L g500 ( 
.A(n_494),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_L g497 ( 
.A(n_493),
.B(n_486),
.Y(n_497)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_497),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_492),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_498),
.B(n_499),
.C(n_493),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_502),
.B(n_503),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_501),
.B(n_495),
.C(n_474),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_504),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_505),
.B(n_485),
.C(n_496),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_507),
.A2(n_506),
.B(n_482),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_508),
.A2(n_500),
.B1(n_473),
.B2(n_476),
.Y(n_509)
);


endmodule