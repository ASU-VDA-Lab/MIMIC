module fake_ariane_2901_n_1842 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1842);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1842;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_279;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_236;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_186),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_108),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_180),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_179),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_189),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_95),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_34),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_123),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_31),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_130),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_28),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_112),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_1),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_120),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_169),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_41),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_124),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_23),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_159),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_1),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_182),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_28),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_64),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_7),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

INVxp33_ASAP7_75t_L g221 ( 
.A(n_100),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_170),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_116),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_23),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_190),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_161),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_156),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_164),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_31),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_7),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_72),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_9),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_119),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_150),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_74),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_57),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_168),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_97),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_91),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_110),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_160),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_9),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_82),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_145),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_39),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_133),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_151),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_2),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_86),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_14),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_154),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_62),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_4),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_193),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_60),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_104),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_70),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_90),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_0),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_53),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_39),
.Y(n_261)
);

BUFx10_ASAP7_75t_L g262 ( 
.A(n_92),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_139),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_56),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_71),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_17),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_76),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_136),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_172),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_0),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_127),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_35),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_173),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_38),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_84),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_63),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_33),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_107),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_85),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_158),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_99),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_115),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_83),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_157),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_66),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_53),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_25),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_75),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_46),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_29),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_187),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_49),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_80),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_149),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_194),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_144),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_50),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_176),
.Y(n_298)
);

BUFx8_ASAP7_75t_SL g299 ( 
.A(n_12),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_137),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_153),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_45),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_143),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_27),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_25),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_135),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_51),
.Y(n_307)
);

BUFx10_ASAP7_75t_L g308 ( 
.A(n_175),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_117),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_32),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_47),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_49),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_192),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_101),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_129),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_32),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_81),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_191),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_26),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_114),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_106),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_94),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_141),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_68),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_47),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_87),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_122),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_79),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_184),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_118),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_17),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_163),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_14),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_2),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_181),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_67),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_174),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_88),
.Y(n_338)
);

BUFx5_ASAP7_75t_L g339 ( 
.A(n_6),
.Y(n_339)
);

INVxp33_ASAP7_75t_SL g340 ( 
.A(n_73),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_165),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_46),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_103),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_98),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_113),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_29),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_128),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_77),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_33),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_5),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_45),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_44),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_105),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_125),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_162),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_50),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_142),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_37),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_15),
.Y(n_359)
);

BUFx5_ASAP7_75t_L g360 ( 
.A(n_96),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_27),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_93),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_26),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_51),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_19),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_148),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_40),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_188),
.Y(n_368)
);

BUFx5_ASAP7_75t_L g369 ( 
.A(n_5),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_134),
.Y(n_370)
);

BUFx5_ASAP7_75t_L g371 ( 
.A(n_147),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_109),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_21),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_36),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_183),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_19),
.Y(n_376)
);

BUFx5_ASAP7_75t_L g377 ( 
.A(n_3),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_178),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_132),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_171),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_56),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_12),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_61),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_52),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_6),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_30),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_166),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_69),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_41),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_111),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_44),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_359),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_339),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_359),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_385),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_299),
.Y(n_396)
);

BUFx6f_ASAP7_75t_SL g397 ( 
.A(n_262),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_290),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_290),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_299),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_239),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_339),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_219),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_263),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_339),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_263),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_276),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_339),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_385),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_339),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_339),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_339),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_369),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_369),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_369),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_282),
.Y(n_416)
);

INVxp33_ASAP7_75t_SL g417 ( 
.A(n_391),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_282),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_369),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_369),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_306),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_369),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_369),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_306),
.Y(n_424)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_232),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_323),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_219),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_323),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_328),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_377),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_201),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_377),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_377),
.Y(n_433)
);

INVxp33_ASAP7_75t_L g434 ( 
.A(n_207),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g435 ( 
.A(n_232),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_377),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_377),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_377),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_210),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_215),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_328),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_245),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_262),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_248),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_253),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_270),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_262),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_272),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_274),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_269),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_287),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_297),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_305),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_242),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_307),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g456 ( 
.A(n_232),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_269),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_310),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_312),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_232),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_316),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_331),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_349),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g464 ( 
.A(n_242),
.Y(n_464)
);

CKINVDCx14_ASAP7_75t_R g465 ( 
.A(n_238),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_351),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_352),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_363),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_367),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_391),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_224),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_196),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_250),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_250),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_350),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_350),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_196),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_269),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_223),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_308),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_223),
.Y(n_481)
);

CKINVDCx14_ASAP7_75t_R g482 ( 
.A(n_308),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_233),
.Y(n_483)
);

INVxp67_ASAP7_75t_SL g484 ( 
.A(n_217),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_233),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_313),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_313),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_308),
.Y(n_488)
);

INVxp33_ASAP7_75t_SL g489 ( 
.A(n_203),
.Y(n_489)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_214),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_344),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_488),
.B(n_221),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_460),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_393),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_488),
.B(n_220),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_393),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_430),
.Y(n_497)
);

INVx6_ASAP7_75t_L g498 ( 
.A(n_477),
.Y(n_498)
);

AND2x2_ASAP7_75t_SL g499 ( 
.A(n_427),
.B(n_344),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_488),
.B(n_318),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_490),
.B(n_489),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_396),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_394),
.B(n_200),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_402),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_402),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_430),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_443),
.B(n_195),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_460),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_477),
.B(n_409),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_432),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_405),
.Y(n_511)
);

OAI21x1_ASAP7_75t_L g512 ( 
.A1(n_432),
.A2(n_321),
.B(n_213),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_427),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_405),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_433),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_408),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_472),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_472),
.B(n_220),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_436),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_408),
.Y(n_520)
);

NOR2x1_ASAP7_75t_L g521 ( 
.A(n_479),
.B(n_247),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_406),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_437),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_425),
.B(n_247),
.Y(n_524)
);

OR2x6_ASAP7_75t_L g525 ( 
.A(n_431),
.B(n_227),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_438),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_443),
.B(n_340),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_482),
.B(n_208),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_447),
.A2(n_389),
.B1(n_261),
.B2(n_342),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_435),
.B(n_227),
.Y(n_530)
);

OA21x2_ASAP7_75t_L g531 ( 
.A1(n_410),
.A2(n_241),
.B(n_235),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_465),
.B(n_249),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_410),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_411),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_411),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_412),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_412),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_401),
.A2(n_261),
.B1(n_389),
.B2(n_342),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_456),
.B(n_252),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_407),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_413),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_413),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_434),
.B(n_212),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_414),
.Y(n_544)
);

INVx5_ASAP7_75t_L g545 ( 
.A(n_414),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_415),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_447),
.B(n_254),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_415),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_419),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_419),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_420),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_450),
.B(n_256),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_420),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_422),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_407),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_422),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_423),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_396),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_392),
.B(n_304),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_416),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_423),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_479),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_481),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_416),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_481),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_483),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_401),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_450),
.B(n_258),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_397),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_454),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_464),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_517),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_497),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_497),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_517),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_519),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_519),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_534),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_506),
.Y(n_579)
);

OR2x6_ASAP7_75t_L g580 ( 
.A(n_525),
.B(n_395),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_492),
.B(n_457),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_499),
.B(n_340),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_495),
.B(n_457),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_523),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_523),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_506),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_510),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_495),
.B(n_509),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_545),
.Y(n_589)
);

INVxp33_ASAP7_75t_SL g590 ( 
.A(n_540),
.Y(n_590)
);

INVxp33_ASAP7_75t_SL g591 ( 
.A(n_540),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_543),
.Y(n_592)
);

BUFx10_ASAP7_75t_L g593 ( 
.A(n_501),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_534),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_495),
.B(n_478),
.Y(n_595)
);

INVx1_ASAP7_75t_SL g596 ( 
.A(n_571),
.Y(n_596)
);

INVx2_ASAP7_75t_SL g597 ( 
.A(n_543),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_509),
.B(n_478),
.Y(n_598)
);

NAND3xp33_ASAP7_75t_SL g599 ( 
.A(n_527),
.B(n_373),
.C(n_418),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_510),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_499),
.B(n_480),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_553),
.Y(n_602)
);

INVxp67_ASAP7_75t_SL g603 ( 
.A(n_509),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_553),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_533),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_533),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_553),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_499),
.A2(n_417),
.B1(n_397),
.B2(n_403),
.Y(n_608)
);

INVxp33_ASAP7_75t_L g609 ( 
.A(n_538),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_548),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_513),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_548),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_565),
.Y(n_613)
);

BUFx10_ASAP7_75t_L g614 ( 
.A(n_498),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_530),
.B(n_480),
.Y(n_615)
);

NAND2xp33_ASAP7_75t_L g616 ( 
.A(n_534),
.B(n_360),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_557),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_530),
.B(n_483),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_498),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_557),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_534),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_565),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_525),
.B(n_439),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_566),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_530),
.B(n_485),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_570),
.Y(n_626)
);

INVxp67_ASAP7_75t_SL g627 ( 
.A(n_534),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_561),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_535),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_561),
.Y(n_630)
);

NAND2xp33_ASAP7_75t_L g631 ( 
.A(n_535),
.B(n_360),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_535),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_535),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_535),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_498),
.Y(n_635)
);

INVx1_ASAP7_75t_SL g636 ( 
.A(n_522),
.Y(n_636)
);

BUFx10_ASAP7_75t_L g637 ( 
.A(n_498),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_500),
.B(n_485),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_525),
.A2(n_484),
.B1(n_397),
.B2(n_373),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_536),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_536),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_566),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_536),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_494),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_494),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_567),
.B(n_404),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_536),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_536),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_525),
.A2(n_470),
.B1(n_205),
.B2(n_230),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_537),
.Y(n_650)
);

INVx4_ASAP7_75t_L g651 ( 
.A(n_545),
.Y(n_651)
);

NAND2xp33_ASAP7_75t_L g652 ( 
.A(n_537),
.B(n_360),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_496),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_537),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_500),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_537),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_555),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_496),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_515),
.B(n_267),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_515),
.B(n_273),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_537),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_541),
.Y(n_662)
);

OAI22xp33_ASAP7_75t_L g663 ( 
.A1(n_529),
.A2(n_399),
.B1(n_398),
.B2(n_418),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_541),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_524),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_541),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_541),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_541),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_528),
.B(n_486),
.Y(n_669)
);

OR2x6_ASAP7_75t_L g670 ( 
.A(n_569),
.B(n_440),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_555),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_504),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_515),
.B(n_278),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_504),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_559),
.A2(n_487),
.B1(n_491),
.B2(n_486),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_505),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_505),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_511),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_511),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_544),
.Y(n_680)
);

BUFx10_ASAP7_75t_L g681 ( 
.A(n_524),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_547),
.B(n_487),
.Y(n_682)
);

INVx5_ASAP7_75t_L g683 ( 
.A(n_544),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_544),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_515),
.B(n_280),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_524),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_544),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_569),
.B(n_491),
.Y(n_688)
);

OAI22xp33_ASAP7_75t_L g689 ( 
.A1(n_552),
.A2(n_424),
.B1(n_426),
.B2(n_421),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_514),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_544),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_SL g692 ( 
.A(n_569),
.B(n_195),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_514),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_550),
.Y(n_694)
);

OAI22xp33_ASAP7_75t_SL g695 ( 
.A1(n_503),
.A2(n_424),
.B1(n_426),
.B2(n_421),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_516),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_515),
.B(n_293),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_550),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_559),
.A2(n_444),
.B1(n_445),
.B2(n_442),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_568),
.B(n_446),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_516),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_520),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_550),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_526),
.B(n_317),
.Y(n_704)
);

OA22x2_ASAP7_75t_L g705 ( 
.A1(n_562),
.A2(n_461),
.B1(n_448),
.B2(n_451),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_520),
.Y(n_706)
);

AND2x6_ASAP7_75t_L g707 ( 
.A(n_542),
.B(n_213),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_550),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_550),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_554),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_532),
.B(n_507),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_546),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_554),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_546),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_539),
.B(n_449),
.Y(n_715)
);

INVxp33_ASAP7_75t_L g716 ( 
.A(n_567),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_549),
.Y(n_717)
);

CKINVDCx6p67_ASAP7_75t_R g718 ( 
.A(n_502),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_644),
.Y(n_719)
);

OAI22xp33_ASAP7_75t_L g720 ( 
.A1(n_609),
.A2(n_429),
.B1(n_441),
.B2(n_428),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_711),
.B(n_554),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_681),
.Y(n_722)
);

NOR2x1p5_ASAP7_75t_L g723 ( 
.A(n_718),
.B(n_560),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_601),
.B(n_549),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_700),
.B(n_551),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_645),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_653),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_580),
.B(n_502),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_592),
.B(n_558),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_609),
.A2(n_531),
.B1(n_563),
.B2(n_562),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_596),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_603),
.B(n_551),
.Y(n_732)
);

NOR3xp33_ASAP7_75t_L g733 ( 
.A(n_599),
.B(n_560),
.C(n_564),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_573),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_623),
.B(n_554),
.Y(n_735)
);

BUFx2_ASAP7_75t_R g736 ( 
.A(n_657),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_597),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_669),
.B(n_518),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_582),
.A2(n_531),
.B1(n_563),
.B2(n_518),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_601),
.B(n_526),
.Y(n_740)
);

INVx8_ASAP7_75t_L g741 ( 
.A(n_670),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_682),
.B(n_518),
.Y(n_742)
);

INVxp67_ASAP7_75t_L g743 ( 
.A(n_611),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_629),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_573),
.Y(n_745)
);

NOR2xp67_ASAP7_75t_SL g746 ( 
.A(n_657),
.B(n_671),
.Y(n_746)
);

NAND2xp33_ASAP7_75t_SL g747 ( 
.A(n_581),
.B(n_564),
.Y(n_747)
);

BUFx3_ASAP7_75t_L g748 ( 
.A(n_614),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_574),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_597),
.Y(n_750)
);

OR2x2_ASAP7_75t_L g751 ( 
.A(n_636),
.B(n_428),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_574),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_623),
.B(n_554),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_658),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_582),
.B(n_526),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_579),
.Y(n_756)
);

INVxp67_ASAP7_75t_L g757 ( 
.A(n_646),
.Y(n_757)
);

INVx8_ASAP7_75t_L g758 ( 
.A(n_670),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_623),
.B(n_556),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_672),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_674),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_655),
.B(n_556),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_655),
.B(n_556),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_676),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_L g765 ( 
.A1(n_588),
.A2(n_333),
.B1(n_236),
.B2(n_259),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_715),
.B(n_556),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_646),
.B(n_429),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_579),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_586),
.Y(n_769)
);

NAND2xp33_ASAP7_75t_L g770 ( 
.A(n_707),
.B(n_556),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_677),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_578),
.B(n_526),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_665),
.B(n_526),
.Y(n_773)
);

O2A1O1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_638),
.A2(n_468),
.B(n_452),
.C(n_453),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_578),
.B(n_545),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_665),
.B(n_521),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_678),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_580),
.B(n_455),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_578),
.B(n_545),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_615),
.B(n_545),
.Y(n_780)
);

HB1xp67_ASAP7_75t_L g781 ( 
.A(n_626),
.Y(n_781)
);

O2A1O1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_613),
.A2(n_624),
.B(n_642),
.C(n_622),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_578),
.B(n_545),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_716),
.B(n_441),
.Y(n_784)
);

OR2x6_ASAP7_75t_L g785 ( 
.A(n_580),
.B(n_458),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_679),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_690),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_693),
.A2(n_512),
.B(n_459),
.C(n_466),
.Y(n_788)
);

INVxp67_ASAP7_75t_SL g789 ( 
.A(n_686),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_578),
.B(n_656),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_696),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_701),
.Y(n_792)
);

NOR3xp33_ASAP7_75t_L g793 ( 
.A(n_671),
.B(n_260),
.C(n_229),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_598),
.B(n_521),
.Y(n_794)
);

INVxp67_ASAP7_75t_L g795 ( 
.A(n_583),
.Y(n_795)
);

O2A1O1Ixp5_ASAP7_75t_L g796 ( 
.A1(n_594),
.A2(n_372),
.B(n_380),
.C(n_324),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_702),
.A2(n_531),
.B1(n_462),
.B2(n_463),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_629),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_686),
.B(n_618),
.Y(n_799)
);

NOR2xp67_ASAP7_75t_L g800 ( 
.A(n_595),
.B(n_639),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_625),
.B(n_531),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_706),
.A2(n_467),
.B1(n_469),
.B2(n_284),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_712),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_656),
.B(n_512),
.Y(n_804)
);

OAI21xp33_ASAP7_75t_L g805 ( 
.A1(n_714),
.A2(n_266),
.B(n_264),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_717),
.Y(n_806)
);

OAI221xp5_ASAP7_75t_L g807 ( 
.A1(n_608),
.A2(n_699),
.B1(n_675),
.B2(n_649),
.C(n_580),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_707),
.A2(n_246),
.B1(n_300),
.B2(n_284),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_656),
.B(n_216),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_572),
.B(n_225),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_656),
.B(n_216),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_587),
.Y(n_812)
);

NOR2xp67_ASAP7_75t_L g813 ( 
.A(n_688),
.B(n_471),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_656),
.B(n_218),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_707),
.A2(n_300),
.B1(n_246),
.B2(n_474),
.Y(n_815)
);

AND2x6_ASAP7_75t_SL g816 ( 
.A(n_590),
.B(n_400),
.Y(n_816)
);

OAI21xp5_ASAP7_75t_L g817 ( 
.A1(n_602),
.A2(n_315),
.B(n_283),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_593),
.B(n_277),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_716),
.B(n_473),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_575),
.B(n_234),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_681),
.B(n_237),
.Y(n_821)
);

NAND2x1p5_ASAP7_75t_L g822 ( 
.A(n_683),
.B(n_320),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_605),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_587),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_600),
.B(n_322),
.Y(n_825)
);

INVxp67_ASAP7_75t_SL g826 ( 
.A(n_694),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_606),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_600),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_593),
.B(n_286),
.Y(n_829)
);

NOR2xp67_ASAP7_75t_L g830 ( 
.A(n_619),
.B(n_475),
.Y(n_830)
);

NAND2x1_ASAP7_75t_L g831 ( 
.A(n_707),
.B(n_213),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_606),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_610),
.Y(n_833)
);

NAND2xp33_ASAP7_75t_L g834 ( 
.A(n_707),
.B(n_218),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_694),
.B(n_294),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_718),
.B(n_475),
.Y(n_836)
);

O2A1O1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_604),
.A2(n_476),
.B(n_388),
.C(n_343),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_694),
.B(n_294),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_692),
.A2(n_390),
.B1(n_355),
.B2(n_336),
.Y(n_839)
);

OR2x2_ASAP7_75t_SL g840 ( 
.A(n_590),
.B(n_591),
.Y(n_840)
);

NOR2xp67_ASAP7_75t_L g841 ( 
.A(n_619),
.B(n_476),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_607),
.B(n_387),
.Y(n_842)
);

INVx8_ASAP7_75t_L g843 ( 
.A(n_670),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_576),
.B(n_355),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_694),
.B(n_390),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_707),
.A2(n_366),
.B1(n_493),
.B2(n_508),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_577),
.B(n_289),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_610),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_612),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_612),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_584),
.B(n_292),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_617),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_617),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_694),
.B(n_337),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_591),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_705),
.B(n_302),
.Y(n_856)
);

BUFx6f_ASAP7_75t_SL g857 ( 
.A(n_670),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_585),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_614),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_594),
.B(n_311),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_594),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_705),
.Y(n_862)
);

INVx8_ASAP7_75t_L g863 ( 
.A(n_683),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_692),
.A2(n_341),
.B1(n_288),
.B2(n_285),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_689),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_621),
.B(n_319),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_620),
.B(n_325),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_629),
.B(n_360),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_628),
.B(n_334),
.Y(n_869)
);

NAND2xp33_ASAP7_75t_L g870 ( 
.A(n_629),
.B(n_346),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_641),
.B(n_360),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_628),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_630),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_641),
.B(n_360),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_659),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_756),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_785),
.B(n_635),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_719),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_722),
.B(n_695),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_725),
.B(n_630),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_724),
.B(n_621),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_724),
.B(n_621),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_731),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_722),
.B(n_637),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_726),
.B(n_633),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_865),
.A2(n_663),
.B1(n_633),
.B2(n_709),
.Y(n_886)
);

INVx4_ASAP7_75t_L g887 ( 
.A(n_741),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_727),
.B(n_654),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_863),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_754),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_863),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_863),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_SL g893 ( 
.A1(n_855),
.A2(n_356),
.B1(n_358),
.B2(n_386),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_760),
.B(n_654),
.Y(n_894)
);

NOR3xp33_ASAP7_75t_SL g895 ( 
.A(n_747),
.B(n_829),
.C(n_818),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_728),
.Y(n_896)
);

INVx5_ASAP7_75t_L g897 ( 
.A(n_741),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_744),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_761),
.B(n_654),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_785),
.B(n_635),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_799),
.B(n_666),
.Y(n_901)
);

OR2x2_ASAP7_75t_SL g902 ( 
.A(n_767),
.B(n_366),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_764),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_738),
.B(n_666),
.Y(n_904)
);

AND2x6_ASAP7_75t_SL g905 ( 
.A(n_784),
.B(n_361),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_742),
.B(n_666),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_744),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_729),
.B(n_364),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_728),
.B(n_641),
.Y(n_909)
);

AOI22xp33_ASAP7_75t_SL g910 ( 
.A1(n_807),
.A2(n_382),
.B1(n_365),
.B2(n_374),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_771),
.Y(n_911)
);

AND3x1_ASAP7_75t_L g912 ( 
.A(n_733),
.B(n_668),
.C(n_667),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_777),
.B(n_667),
.Y(n_913)
);

INVx4_ASAP7_75t_L g914 ( 
.A(n_741),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_786),
.B(n_667),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_787),
.B(n_668),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_791),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_862),
.A2(n_659),
.B1(n_660),
.B2(n_673),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_720),
.B(n_668),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_792),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_744),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_795),
.B(n_680),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_803),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_778),
.B(n_708),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_798),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_798),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_806),
.B(n_680),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_732),
.B(n_680),
.Y(n_928)
);

AOI22xp33_ASAP7_75t_L g929 ( 
.A1(n_856),
.A2(n_660),
.B1(n_673),
.B2(n_685),
.Y(n_929)
);

BUFx2_ASAP7_75t_L g930 ( 
.A(n_781),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_SL g931 ( 
.A1(n_857),
.A2(n_376),
.B1(n_381),
.B2(n_384),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_766),
.B(n_684),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_720),
.A2(n_685),
.B1(n_697),
.B2(n_704),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_798),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_794),
.B(n_684),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_757),
.B(n_704),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_778),
.B(n_708),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_751),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_794),
.B(n_684),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_782),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_832),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_839),
.A2(n_703),
.B1(n_709),
.B2(n_710),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_743),
.B(n_703),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_800),
.A2(n_703),
.B1(n_709),
.B2(n_627),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_818),
.B(n_632),
.Y(n_945)
);

OR2x2_ASAP7_75t_L g946 ( 
.A(n_840),
.B(n_632),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_833),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_833),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_858),
.Y(n_949)
);

BUFx12f_ASAP7_75t_L g950 ( 
.A(n_816),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_836),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_798),
.Y(n_952)
);

AND2x6_ASAP7_75t_SL g953 ( 
.A(n_829),
.B(n_3),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_748),
.B(n_708),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_734),
.Y(n_955)
);

INVxp67_ASAP7_75t_L g956 ( 
.A(n_819),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_755),
.B(n_634),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_745),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_788),
.A2(n_713),
.B(n_710),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_780),
.A2(n_713),
.B(n_634),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_749),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_812),
.Y(n_962)
);

AND2x6_ASAP7_75t_SL g963 ( 
.A(n_736),
.B(n_4),
.Y(n_963)
);

INVx5_ASAP7_75t_L g964 ( 
.A(n_758),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_789),
.B(n_640),
.Y(n_965)
);

NAND2x1p5_ASAP7_75t_L g966 ( 
.A(n_735),
.B(n_683),
.Y(n_966)
);

INVx4_ASAP7_75t_L g967 ( 
.A(n_758),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_755),
.B(n_698),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_752),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_824),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_801),
.B(n_691),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_828),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_768),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_785),
.B(n_640),
.Y(n_974)
);

NAND3xp33_ASAP7_75t_SL g975 ( 
.A(n_793),
.B(n_240),
.C(n_383),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_730),
.B(n_687),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_769),
.Y(n_977)
);

OAI21xp33_ASAP7_75t_SL g978 ( 
.A1(n_817),
.A2(n_664),
.B(n_662),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_730),
.B(n_643),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_758),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_873),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_821),
.B(n_643),
.Y(n_982)
);

BUFx8_ASAP7_75t_L g983 ( 
.A(n_857),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_753),
.B(n_647),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_740),
.B(n_664),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_740),
.B(n_647),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_797),
.B(n_662),
.Y(n_987)
);

BUFx4f_ASAP7_75t_L g988 ( 
.A(n_843),
.Y(n_988)
);

AND2x6_ASAP7_75t_L g989 ( 
.A(n_859),
.B(n_648),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_823),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_827),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_848),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_797),
.B(n_721),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_759),
.B(n_650),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_721),
.B(n_661),
.Y(n_995)
);

INVx2_ASAP7_75t_SL g996 ( 
.A(n_723),
.Y(n_996)
);

AOI22xp5_ASAP7_75t_L g997 ( 
.A1(n_759),
.A2(n_652),
.B1(n_631),
.B2(n_616),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_849),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_843),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_859),
.Y(n_1000)
);

AOI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_737),
.A2(n_652),
.B1(n_631),
.B2(n_616),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_850),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_750),
.B(n_589),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_861),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_864),
.B(n_651),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_852),
.Y(n_1006)
);

INVx1_ASAP7_75t_SL g1007 ( 
.A(n_773),
.Y(n_1007)
);

NAND3xp33_ASAP7_75t_SL g1008 ( 
.A(n_765),
.B(n_206),
.C(n_379),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_853),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_861),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_872),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_810),
.B(n_820),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_SL g1013 ( 
.A1(n_808),
.A2(n_204),
.B1(n_378),
.B2(n_375),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_875),
.B(n_776),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_762),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_762),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_763),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_808),
.A2(n_508),
.B1(n_493),
.B2(n_321),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_763),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_822),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_830),
.Y(n_1021)
);

NOR2x1p5_ASAP7_75t_L g1022 ( 
.A(n_746),
.B(n_321),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_802),
.A2(n_508),
.B1(n_493),
.B2(n_651),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_860),
.A2(n_199),
.B1(n_370),
.B2(n_368),
.Y(n_1024)
);

OAI21xp33_ASAP7_75t_L g1025 ( 
.A1(n_860),
.A2(n_197),
.B(n_362),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_739),
.B(n_508),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_772),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_867),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_869),
.Y(n_1029)
);

XNOR2xp5_ASAP7_75t_L g1030 ( 
.A(n_822),
.B(n_198),
.Y(n_1030)
);

INVx5_ASAP7_75t_L g1031 ( 
.A(n_770),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_805),
.B(n_202),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_847),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_739),
.B(n_508),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_842),
.B(n_209),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_841),
.Y(n_1036)
);

NOR3xp33_ASAP7_75t_L g1037 ( 
.A(n_774),
.B(n_345),
.C(n_296),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_851),
.Y(n_1038)
);

CKINVDCx20_ASAP7_75t_R g1039 ( 
.A(n_809),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_825),
.B(n_211),
.Y(n_1040)
);

NAND3xp33_ASAP7_75t_SL g1041 ( 
.A(n_837),
.B(n_815),
.C(n_844),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_813),
.B(n_222),
.Y(n_1042)
);

AOI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_866),
.A2(n_301),
.B1(n_228),
.B2(n_357),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_831),
.Y(n_1044)
);

NOR2x2_ASAP7_75t_L g1045 ( 
.A(n_866),
.B(n_8),
.Y(n_1045)
);

INVx5_ASAP7_75t_L g1046 ( 
.A(n_846),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_SL g1047 ( 
.A(n_988),
.B(n_826),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_876),
.Y(n_1048)
);

OAI21xp33_ASAP7_75t_L g1049 ( 
.A1(n_1024),
.A2(n_838),
.B(n_811),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_1033),
.B(n_815),
.Y(n_1050)
);

BUFx2_ASAP7_75t_L g1051 ( 
.A(n_930),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_878),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_1046),
.A2(n_780),
.B1(n_845),
.B2(n_838),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_889),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_881),
.A2(n_804),
.B(n_834),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_956),
.B(n_1012),
.Y(n_1056)
);

CKINVDCx11_ASAP7_75t_R g1057 ( 
.A(n_963),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_951),
.B(n_809),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_1046),
.A2(n_814),
.B1(n_835),
.B2(n_845),
.Y(n_1059)
);

NAND2xp33_ASAP7_75t_R g1060 ( 
.A(n_895),
.B(n_226),
.Y(n_1060)
);

INVx1_ASAP7_75t_SL g1061 ( 
.A(n_883),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_908),
.B(n_811),
.Y(n_1062)
);

INVx4_ASAP7_75t_L g1063 ( 
.A(n_897),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_896),
.B(n_846),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_881),
.A2(n_804),
.B(n_790),
.Y(n_1065)
);

NOR3xp33_ASAP7_75t_SL g1066 ( 
.A(n_975),
.B(n_835),
.C(n_788),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_1046),
.A2(n_790),
.B1(n_772),
.B2(n_854),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_936),
.B(n_919),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_882),
.A2(n_880),
.B(n_935),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_889),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_941),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1007),
.B(n_870),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_910),
.A2(n_854),
.B1(n_871),
.B2(n_868),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_947),
.Y(n_1074)
);

AO21x1_ASAP7_75t_L g1075 ( 
.A1(n_945),
.A2(n_874),
.B(n_783),
.Y(n_1075)
);

BUFx2_ASAP7_75t_SL g1076 ( 
.A(n_897),
.Y(n_1076)
);

AOI221xp5_ASAP7_75t_L g1077 ( 
.A1(n_893),
.A2(n_796),
.B1(n_309),
.B2(n_303),
.C(n_243),
.Y(n_1077)
);

INVx2_ASAP7_75t_SL g1078 ( 
.A(n_983),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_938),
.B(n_943),
.Y(n_1079)
);

HB1xp67_ASAP7_75t_L g1080 ( 
.A(n_877),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_1038),
.B(n_775),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_983),
.Y(n_1082)
);

INVx5_ASAP7_75t_L g1083 ( 
.A(n_1046),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_948),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_882),
.A2(n_783),
.B(n_779),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_940),
.A2(n_779),
.B1(n_775),
.B2(n_314),
.Y(n_1086)
);

OAI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_890),
.A2(n_295),
.B1(n_354),
.B2(n_353),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_903),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_980),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_877),
.B(n_231),
.Y(n_1090)
);

INVxp67_ASAP7_75t_L g1091 ( 
.A(n_946),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_955),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_897),
.B(n_493),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_1028),
.B(n_244),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_1039),
.A2(n_298),
.B1(n_348),
.B2(n_347),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_SL g1096 ( 
.A1(n_902),
.A2(n_251),
.B1(n_255),
.B2(n_257),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_959),
.A2(n_371),
.B(n_89),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_980),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_911),
.A2(n_920),
.B1(n_923),
.B2(n_917),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_1013),
.A2(n_326),
.B1(n_338),
.B2(n_335),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_1029),
.A2(n_281),
.B1(n_332),
.B2(n_330),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1007),
.B(n_8),
.Y(n_1102)
);

NOR2xp67_ASAP7_75t_L g1103 ( 
.A(n_897),
.B(n_265),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_880),
.A2(n_279),
.B(n_329),
.Y(n_1104)
);

CKINVDCx16_ASAP7_75t_R g1105 ( 
.A(n_950),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_935),
.A2(n_327),
.B(n_291),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_949),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_R g1108 ( 
.A(n_988),
.B(n_275),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_980),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_885),
.A2(n_271),
.B1(n_268),
.B2(n_13),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_939),
.A2(n_371),
.B(n_11),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_939),
.A2(n_371),
.B(n_11),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1035),
.B(n_10),
.Y(n_1113)
);

INVx1_ASAP7_75t_SL g1114 ( 
.A(n_1045),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_932),
.A2(n_371),
.B(n_13),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_1014),
.B(n_10),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_900),
.Y(n_1117)
);

INVx1_ASAP7_75t_SL g1118 ( 
.A(n_900),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_879),
.B(n_15),
.Y(n_1119)
);

CKINVDCx20_ASAP7_75t_R g1120 ( 
.A(n_1030),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_958),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_887),
.B(n_16),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1040),
.B(n_16),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_932),
.A2(n_371),
.B(n_20),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_886),
.B(n_18),
.Y(n_1125)
);

O2A1O1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_1008),
.A2(n_18),
.B(n_20),
.C(n_21),
.Y(n_1126)
);

OA22x2_ASAP7_75t_L g1127 ( 
.A1(n_909),
.A2(n_22),
.B1(n_24),
.B2(n_30),
.Y(n_1127)
);

O2A1O1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_922),
.A2(n_22),
.B(n_24),
.C(n_34),
.Y(n_1128)
);

NOR3xp33_ASAP7_75t_SL g1129 ( 
.A(n_1022),
.B(n_35),
.C(n_36),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_931),
.B(n_37),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_964),
.B(n_38),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_999),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_999),
.B(n_40),
.Y(n_1133)
);

NAND3xp33_ASAP7_75t_L g1134 ( 
.A(n_1032),
.B(n_1043),
.C(n_1037),
.Y(n_1134)
);

O2A1O1Ixp5_ASAP7_75t_L g1135 ( 
.A1(n_1005),
.A2(n_42),
.B(n_43),
.C(n_48),
.Y(n_1135)
);

INVx4_ASAP7_75t_L g1136 ( 
.A(n_964),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_887),
.B(n_42),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_R g1138 ( 
.A(n_999),
.B(n_126),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_962),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_928),
.A2(n_971),
.B(n_906),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_974),
.B(n_43),
.Y(n_1141)
);

NOR2x1_ASAP7_75t_SL g1142 ( 
.A(n_1031),
.B(n_371),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_914),
.B(n_48),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_928),
.A2(n_52),
.B(n_54),
.Y(n_1144)
);

AOI221xp5_ASAP7_75t_L g1145 ( 
.A1(n_1041),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.C(n_58),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_SL g1146 ( 
.A(n_914),
.B(n_55),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1025),
.A2(n_1019),
.B(n_1016),
.C(n_1017),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_1000),
.B(n_58),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_971),
.A2(n_59),
.B(n_65),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_970),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_972),
.Y(n_1151)
);

O2A1O1Ixp5_ASAP7_75t_L g1152 ( 
.A1(n_954),
.A2(n_78),
.B(n_102),
.C(n_121),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_885),
.A2(n_131),
.B1(n_138),
.B2(n_140),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_967),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_SL g1155 ( 
.A1(n_884),
.A2(n_146),
.B(n_152),
.C(n_155),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_981),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_1000),
.B(n_167),
.Y(n_1157)
);

BUFx8_ASAP7_75t_L g1158 ( 
.A(n_996),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_R g1159 ( 
.A(n_905),
.B(n_967),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_1031),
.B(n_974),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_953),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_1004),
.Y(n_1162)
);

A2O1A1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_1015),
.A2(n_978),
.B(n_933),
.C(n_993),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_SL g1164 ( 
.A1(n_1044),
.A2(n_926),
.B(n_934),
.C(n_888),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_961),
.A2(n_969),
.B1(n_973),
.B2(n_1011),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_984),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_904),
.A2(n_960),
.B(n_985),
.Y(n_1167)
);

NOR3xp33_ASAP7_75t_L g1168 ( 
.A(n_1042),
.B(n_924),
.C(n_937),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1010),
.B(n_1021),
.Y(n_1169)
);

NAND3xp33_ASAP7_75t_L g1170 ( 
.A(n_912),
.B(n_944),
.C(n_1001),
.Y(n_1170)
);

AO221x2_ASAP7_75t_L g1171 ( 
.A1(n_942),
.A2(n_927),
.B1(n_913),
.B2(n_888),
.C(n_899),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_985),
.A2(n_986),
.B(n_901),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_986),
.A2(n_968),
.B(n_957),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1003),
.B(n_1020),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_957),
.A2(n_968),
.B(n_915),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_984),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1020),
.B(n_1036),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1003),
.B(n_982),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_977),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1031),
.B(n_892),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_993),
.B(n_918),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_994),
.A2(n_989),
.B1(n_942),
.B2(n_916),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_SL g1183 ( 
.A(n_989),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_929),
.B(n_994),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_894),
.A2(n_916),
.B(n_927),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_998),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_894),
.A2(n_913),
.B(n_915),
.C(n_899),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_926),
.B(n_934),
.Y(n_1188)
);

INVx1_ASAP7_75t_SL g1189 ( 
.A(n_989),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_989),
.B(n_992),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1031),
.A2(n_997),
.B1(n_965),
.B2(n_921),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_995),
.A2(n_1034),
.B(n_1026),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1006),
.A2(n_1009),
.B1(n_990),
.B2(n_991),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1002),
.B(n_1027),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_987),
.B(n_976),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_995),
.A2(n_1034),
.B(n_1026),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_891),
.B(n_892),
.Y(n_1197)
);

AO31x2_ASAP7_75t_L g1198 ( 
.A1(n_1075),
.A2(n_976),
.A3(n_979),
.B(n_987),
.Y(n_1198)
);

INVx5_ASAP7_75t_SL g1199 ( 
.A(n_1154),
.Y(n_1199)
);

NOR2xp67_ASAP7_75t_L g1200 ( 
.A(n_1056),
.B(n_891),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1079),
.B(n_952),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_SL g1202 ( 
.A1(n_1183),
.A2(n_979),
.B(n_925),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1068),
.B(n_952),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1114),
.B(n_898),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1083),
.B(n_907),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1083),
.B(n_907),
.Y(n_1206)
);

INVx4_ASAP7_75t_L g1207 ( 
.A(n_1154),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1083),
.B(n_921),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1123),
.A2(n_1083),
.B1(n_1125),
.B2(n_1134),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1052),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1131),
.B(n_966),
.Y(n_1211)
);

BUFx4f_ASAP7_75t_SL g1212 ( 
.A(n_1158),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1069),
.A2(n_1018),
.B(n_1023),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1088),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_1131),
.B(n_1047),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_SL g1216 ( 
.A(n_1178),
.B(n_1072),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1192),
.A2(n_1196),
.B(n_1065),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1051),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1140),
.A2(n_1175),
.B(n_1185),
.Y(n_1219)
);

INVx3_ASAP7_75t_SL g1220 ( 
.A(n_1162),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1145),
.A2(n_1119),
.B1(n_1116),
.B2(n_1182),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1196),
.A2(n_1065),
.B(n_1055),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1049),
.A2(n_1081),
.B(n_1126),
.C(n_1170),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1107),
.Y(n_1224)
);

NAND2x1p5_ASAP7_75t_L g1225 ( 
.A(n_1160),
.B(n_1063),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1154),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1145),
.A2(n_1181),
.B1(n_1099),
.B2(n_1100),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1139),
.Y(n_1228)
);

NOR2xp67_ASAP7_75t_L g1229 ( 
.A(n_1136),
.B(n_1169),
.Y(n_1229)
);

NAND3x1_ASAP7_75t_L g1230 ( 
.A(n_1130),
.B(n_1062),
.C(n_1133),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_SL g1231 ( 
.A1(n_1164),
.A2(n_1157),
.B(n_1148),
.C(n_1187),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1122),
.A2(n_1137),
.B1(n_1163),
.B2(n_1102),
.Y(n_1232)
);

AO31x2_ASAP7_75t_L g1233 ( 
.A1(n_1173),
.A2(n_1140),
.A3(n_1172),
.B(n_1175),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1172),
.A2(n_1185),
.B(n_1191),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1091),
.B(n_1061),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1118),
.B(n_1050),
.Y(n_1236)
);

OAI21xp5_ASAP7_75t_SL g1237 ( 
.A1(n_1126),
.A2(n_1128),
.B(n_1077),
.Y(n_1237)
);

AO31x2_ASAP7_75t_L g1238 ( 
.A1(n_1195),
.A2(n_1053),
.A3(n_1059),
.B(n_1147),
.Y(n_1238)
);

AO31x2_ASAP7_75t_L g1239 ( 
.A1(n_1067),
.A2(n_1194),
.A3(n_1111),
.B(n_1112),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1094),
.B(n_1080),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1171),
.A2(n_1149),
.B(n_1085),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1117),
.B(n_1150),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1171),
.A2(n_1149),
.B(n_1106),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1111),
.A2(n_1112),
.B(n_1124),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_1158),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1184),
.B(n_1151),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1106),
.A2(n_1104),
.B(n_1153),
.Y(n_1247)
);

AO21x2_ASAP7_75t_L g1248 ( 
.A1(n_1190),
.A2(n_1115),
.B(n_1066),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1098),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1146),
.B(n_1174),
.Y(n_1250)
);

OR2x6_ASAP7_75t_L g1251 ( 
.A(n_1076),
.B(n_1078),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1104),
.A2(n_1086),
.B(n_1180),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1156),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1135),
.A2(n_1144),
.B(n_1152),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1095),
.B(n_1143),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1188),
.A2(n_1155),
.B(n_1189),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1166),
.B(n_1176),
.Y(n_1257)
);

INVx1_ASAP7_75t_SL g1258 ( 
.A(n_1141),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1144),
.A2(n_1073),
.B(n_1077),
.Y(n_1259)
);

NOR3xp33_ASAP7_75t_L g1260 ( 
.A(n_1090),
.B(n_1096),
.C(n_1110),
.Y(n_1260)
);

AO31x2_ASAP7_75t_L g1261 ( 
.A1(n_1142),
.A2(n_1084),
.A3(n_1074),
.B(n_1071),
.Y(n_1261)
);

AOI21xp33_ASAP7_75t_L g1262 ( 
.A1(n_1127),
.A2(n_1060),
.B(n_1064),
.Y(n_1262)
);

INVx1_ASAP7_75t_SL g1263 ( 
.A(n_1132),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1058),
.B(n_1177),
.Y(n_1264)
);

AOI221x1_ASAP7_75t_L g1265 ( 
.A1(n_1168),
.A2(n_1087),
.B1(n_1186),
.B2(n_1092),
.C(n_1179),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1120),
.B(n_1089),
.Y(n_1266)
);

INVx2_ASAP7_75t_SL g1267 ( 
.A(n_1089),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1054),
.A2(n_1070),
.B(n_1193),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1121),
.B(n_1108),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1089),
.B(n_1109),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1109),
.B(n_1136),
.Y(n_1271)
);

CKINVDCx20_ASAP7_75t_R g1272 ( 
.A(n_1105),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1127),
.A2(n_1129),
.B1(n_1183),
.B2(n_1101),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1109),
.B(n_1197),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_1159),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1165),
.Y(n_1276)
);

AO21x1_ASAP7_75t_L g1277 ( 
.A1(n_1093),
.A2(n_1197),
.B(n_1103),
.Y(n_1277)
);

NAND2x1p5_ASAP7_75t_L g1278 ( 
.A(n_1093),
.B(n_1070),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1138),
.A2(n_1082),
.B(n_1161),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1057),
.A2(n_1097),
.B(n_1167),
.Y(n_1280)
);

NOR2x1_ASAP7_75t_SL g1281 ( 
.A(n_1083),
.B(n_1076),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1097),
.A2(n_1167),
.B(n_1192),
.Y(n_1282)
);

NOR2x1_ASAP7_75t_SL g1283 ( 
.A(n_1083),
.B(n_1076),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1097),
.A2(n_1167),
.B(n_1192),
.Y(n_1284)
);

AND2x4_ASAP7_75t_L g1285 ( 
.A(n_1083),
.B(n_887),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1052),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1097),
.A2(n_1167),
.B(n_1192),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1056),
.B(n_1068),
.Y(n_1288)
);

NAND3x1_ASAP7_75t_L g1289 ( 
.A(n_1130),
.B(n_1119),
.C(n_639),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1052),
.Y(n_1290)
);

AOI21xp33_ASAP7_75t_L g1291 ( 
.A1(n_1125),
.A2(n_1113),
.B(n_1123),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1069),
.A2(n_1140),
.B(n_1175),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1069),
.A2(n_1140),
.B(n_1175),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1051),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1069),
.A2(n_1140),
.B(n_1175),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1069),
.A2(n_1140),
.B(n_1175),
.Y(n_1296)
);

AOI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1119),
.A2(n_591),
.B1(n_590),
.B2(n_657),
.Y(n_1297)
);

OAI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1113),
.A2(n_609),
.B1(n_416),
.B2(n_418),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_1051),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1069),
.A2(n_1140),
.B(n_1175),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1052),
.Y(n_1301)
);

BUFx10_ASAP7_75t_L g1302 ( 
.A(n_1122),
.Y(n_1302)
);

INVx3_ASAP7_75t_L g1303 ( 
.A(n_1063),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1105),
.Y(n_1304)
);

AOI21x1_ASAP7_75t_SL g1305 ( 
.A1(n_1113),
.A2(n_1123),
.B(n_581),
.Y(n_1305)
);

BUFx10_ASAP7_75t_L g1306 ( 
.A(n_1122),
.Y(n_1306)
);

OAI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1069),
.A2(n_1065),
.B(n_1173),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1097),
.A2(n_1167),
.B(n_1192),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1048),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1097),
.A2(n_1167),
.B(n_1192),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1051),
.B(n_590),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1056),
.B(n_1068),
.Y(n_1312)
);

BUFx4f_ASAP7_75t_SL g1313 ( 
.A(n_1158),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1056),
.B(n_1068),
.Y(n_1314)
);

INVx5_ASAP7_75t_L g1315 ( 
.A(n_1083),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1051),
.B(n_590),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1083),
.B(n_1134),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1069),
.A2(n_1065),
.B(n_1173),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1069),
.A2(n_1065),
.B(n_1173),
.Y(n_1319)
);

OA21x2_ASAP7_75t_L g1320 ( 
.A1(n_1192),
.A2(n_1196),
.B(n_1167),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_SL g1321 ( 
.A1(n_1183),
.A2(n_1187),
.B(n_857),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1069),
.A2(n_1065),
.B(n_1173),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1097),
.A2(n_1167),
.B(n_1192),
.Y(n_1323)
);

AO31x2_ASAP7_75t_L g1324 ( 
.A1(n_1075),
.A2(n_1173),
.A3(n_1196),
.B(n_1192),
.Y(n_1324)
);

INVx3_ASAP7_75t_L g1325 ( 
.A(n_1063),
.Y(n_1325)
);

A2O1A1Ixp33_ASAP7_75t_L g1326 ( 
.A1(n_1113),
.A2(n_1123),
.B(n_1134),
.C(n_1119),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1048),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1052),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1056),
.B(n_1068),
.Y(n_1329)
);

A2O1A1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1113),
.A2(n_1123),
.B(n_1134),
.C(n_1119),
.Y(n_1330)
);

AOI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1119),
.A2(n_591),
.B1(n_590),
.B2(n_657),
.Y(n_1331)
);

AO31x2_ASAP7_75t_L g1332 ( 
.A1(n_1075),
.A2(n_1173),
.A3(n_1196),
.B(n_1192),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1069),
.A2(n_1065),
.B(n_1173),
.Y(n_1333)
);

O2A1O1Ixp33_ASAP7_75t_SL g1334 ( 
.A1(n_1113),
.A2(n_1123),
.B(n_1164),
.C(n_1134),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_SL g1335 ( 
.A1(n_1085),
.A2(n_1187),
.B(n_1068),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1079),
.B(n_609),
.Y(n_1336)
);

AOI221xp5_ASAP7_75t_SL g1337 ( 
.A1(n_1145),
.A2(n_1126),
.B1(n_1144),
.B2(n_1128),
.C(n_1113),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1210),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1221),
.B(n_1232),
.Y(n_1339)
);

OAI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1221),
.A2(n_1227),
.B1(n_1237),
.B2(n_1232),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1214),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1282),
.A2(n_1287),
.B(n_1284),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1336),
.B(n_1201),
.Y(n_1343)
);

INVxp67_ASAP7_75t_SL g1344 ( 
.A(n_1217),
.Y(n_1344)
);

OA21x2_ASAP7_75t_L g1345 ( 
.A1(n_1295),
.A2(n_1300),
.B(n_1296),
.Y(n_1345)
);

OAI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1326),
.A2(n_1330),
.B(n_1223),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1262),
.A2(n_1291),
.B1(n_1260),
.B2(n_1255),
.Y(n_1347)
);

AOI22x1_ASAP7_75t_L g1348 ( 
.A1(n_1243),
.A2(n_1244),
.B1(n_1247),
.B2(n_1241),
.Y(n_1348)
);

CKINVDCx20_ASAP7_75t_R g1349 ( 
.A(n_1272),
.Y(n_1349)
);

BUFx12f_ASAP7_75t_L g1350 ( 
.A(n_1304),
.Y(n_1350)
);

NOR2x1_ASAP7_75t_SL g1351 ( 
.A(n_1315),
.B(n_1251),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1218),
.Y(n_1352)
);

OAI31xp33_ASAP7_75t_L g1353 ( 
.A1(n_1298),
.A2(n_1273),
.A3(n_1209),
.B(n_1262),
.Y(n_1353)
);

AO31x2_ASAP7_75t_L g1354 ( 
.A1(n_1265),
.A2(n_1213),
.A3(n_1252),
.B(n_1246),
.Y(n_1354)
);

AO21x1_ASAP7_75t_L g1355 ( 
.A1(n_1291),
.A2(n_1317),
.B(n_1273),
.Y(n_1355)
);

OA21x2_ASAP7_75t_L g1356 ( 
.A1(n_1307),
.A2(n_1333),
.B(n_1322),
.Y(n_1356)
);

AOI221xp5_ASAP7_75t_L g1357 ( 
.A1(n_1337),
.A2(n_1334),
.B1(n_1297),
.B2(n_1331),
.C(n_1329),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1224),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1228),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1233),
.Y(n_1360)
);

INVx2_ASAP7_75t_SL g1361 ( 
.A(n_1220),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1318),
.A2(n_1319),
.B(n_1333),
.Y(n_1362)
);

OAI221xp5_ASAP7_75t_L g1363 ( 
.A1(n_1337),
.A2(n_1240),
.B1(n_1314),
.B2(n_1312),
.C(n_1288),
.Y(n_1363)
);

OA21x2_ASAP7_75t_L g1364 ( 
.A1(n_1319),
.A2(n_1322),
.B(n_1222),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1308),
.A2(n_1323),
.B(n_1310),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1264),
.B(n_1216),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1242),
.B(n_1294),
.Y(n_1367)
);

A2O1A1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1254),
.A2(n_1280),
.B(n_1234),
.C(n_1203),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1233),
.Y(n_1369)
);

INVx2_ASAP7_75t_SL g1370 ( 
.A(n_1245),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_SL g1371 ( 
.A1(n_1281),
.A2(n_1283),
.B(n_1277),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1258),
.B(n_1299),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1266),
.B(n_1204),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1253),
.Y(n_1374)
);

INVx2_ASAP7_75t_SL g1375 ( 
.A(n_1212),
.Y(n_1375)
);

AO31x2_ASAP7_75t_L g1376 ( 
.A1(n_1276),
.A2(n_1301),
.A3(n_1286),
.B(n_1328),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1290),
.Y(n_1377)
);

O2A1O1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1254),
.A2(n_1231),
.B(n_1250),
.C(n_1311),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1320),
.A2(n_1256),
.B(n_1268),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1320),
.A2(n_1305),
.B(n_1321),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1233),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1206),
.A2(n_1208),
.B(n_1225),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1324),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1313),
.Y(n_1384)
);

AOI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1215),
.A2(n_1229),
.B(n_1211),
.Y(n_1385)
);

A2O1A1Ixp33_ASAP7_75t_L g1386 ( 
.A1(n_1200),
.A2(n_1258),
.B(n_1279),
.C(n_1236),
.Y(n_1386)
);

OAI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1251),
.A2(n_1289),
.B1(n_1257),
.B2(n_1235),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1324),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_1249),
.Y(n_1389)
);

AO31x2_ASAP7_75t_L g1390 ( 
.A1(n_1309),
.A2(n_1327),
.A3(n_1238),
.B(n_1324),
.Y(n_1390)
);

AOI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1316),
.A2(n_1230),
.B1(n_1306),
.B2(n_1302),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1270),
.Y(n_1392)
);

OA21x2_ASAP7_75t_L g1393 ( 
.A1(n_1332),
.A2(n_1239),
.B(n_1238),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1332),
.Y(n_1394)
);

OAI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1251),
.A2(n_1274),
.B1(n_1275),
.B2(n_1269),
.Y(n_1395)
);

O2A1O1Ixp33_ASAP7_75t_SL g1396 ( 
.A1(n_1303),
.A2(n_1325),
.B(n_1267),
.C(n_1302),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1278),
.A2(n_1248),
.B(n_1239),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1306),
.B(n_1263),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1205),
.A2(n_1285),
.B(n_1239),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1261),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1199),
.B(n_1226),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1207),
.B(n_1285),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1271),
.Y(n_1403)
);

INVx2_ASAP7_75t_SL g1404 ( 
.A(n_1199),
.Y(n_1404)
);

BUFx6f_ASAP7_75t_L g1405 ( 
.A(n_1238),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1221),
.A2(n_609),
.B1(n_538),
.B2(n_1227),
.Y(n_1406)
);

AO31x2_ASAP7_75t_L g1407 ( 
.A1(n_1292),
.A2(n_1295),
.A3(n_1296),
.B(n_1293),
.Y(n_1407)
);

CKINVDCx11_ASAP7_75t_R g1408 ( 
.A(n_1272),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1315),
.B(n_1083),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1336),
.B(n_1201),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1210),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1221),
.B(n_1232),
.Y(n_1412)
);

A2O1A1Ixp33_ASAP7_75t_L g1413 ( 
.A1(n_1221),
.A2(n_1259),
.B(n_1330),
.C(n_1326),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1198),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1297),
.A2(n_1331),
.B1(n_1113),
.B2(n_1221),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1210),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1282),
.A2(n_1287),
.B(n_1284),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1221),
.B(n_1232),
.Y(n_1418)
);

INVx3_ASAP7_75t_SL g1419 ( 
.A(n_1304),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1212),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1221),
.B(n_1232),
.Y(n_1421)
);

NAND2x1_ASAP7_75t_L g1422 ( 
.A(n_1321),
.B(n_1335),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1210),
.Y(n_1423)
);

OAI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1232),
.A2(n_1330),
.B(n_1326),
.Y(n_1424)
);

INVx3_ASAP7_75t_SL g1425 ( 
.A(n_1304),
.Y(n_1425)
);

OA21x2_ASAP7_75t_L g1426 ( 
.A1(n_1219),
.A2(n_1293),
.B(n_1292),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1198),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_1212),
.Y(n_1428)
);

O2A1O1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1326),
.A2(n_1330),
.B(n_1232),
.C(n_1221),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1210),
.Y(n_1430)
);

OA21x2_ASAP7_75t_L g1431 ( 
.A1(n_1219),
.A2(n_1293),
.B(n_1292),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1210),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_1212),
.Y(n_1433)
);

OAI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1221),
.A2(n_609),
.B1(n_1068),
.B2(n_1125),
.Y(n_1434)
);

OA21x2_ASAP7_75t_L g1435 ( 
.A1(n_1219),
.A2(n_1293),
.B(n_1292),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1210),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1198),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1210),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1221),
.A2(n_609),
.B1(n_538),
.B2(n_1227),
.Y(n_1439)
);

AND2x4_ASAP7_75t_L g1440 ( 
.A(n_1315),
.B(n_1083),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1297),
.A2(n_1331),
.B1(n_1113),
.B2(n_1221),
.Y(n_1441)
);

OA21x2_ASAP7_75t_L g1442 ( 
.A1(n_1219),
.A2(n_1293),
.B(n_1292),
.Y(n_1442)
);

BUFx2_ASAP7_75t_L g1443 ( 
.A(n_1218),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1198),
.Y(n_1444)
);

NAND2x1p5_ASAP7_75t_L g1445 ( 
.A(n_1315),
.B(n_1083),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_SL g1446 ( 
.A1(n_1221),
.A2(n_1259),
.B(n_1335),
.Y(n_1446)
);

OR2x6_ASAP7_75t_L g1447 ( 
.A(n_1321),
.B(n_1202),
.Y(n_1447)
);

OAI211xp5_ASAP7_75t_L g1448 ( 
.A1(n_1326),
.A2(n_1330),
.B(n_1291),
.C(n_1297),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_SL g1449 ( 
.A1(n_1413),
.A2(n_1429),
.B(n_1346),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1339),
.A2(n_1421),
.B1(n_1412),
.B2(n_1418),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1340),
.A2(n_1412),
.B(n_1339),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1340),
.A2(n_1421),
.B(n_1418),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1367),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1413),
.A2(n_1362),
.B(n_1424),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1372),
.B(n_1352),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1443),
.B(n_1338),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1389),
.B(n_1403),
.Y(n_1457)
);

OA22x2_ASAP7_75t_L g1458 ( 
.A1(n_1391),
.A2(n_1415),
.B1(n_1441),
.B2(n_1446),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1366),
.B(n_1392),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1376),
.B(n_1363),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1373),
.B(n_1389),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1347),
.B(n_1398),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1347),
.B(n_1398),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1341),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1358),
.B(n_1359),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1408),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1374),
.B(n_1377),
.Y(n_1467)
);

O2A1O1Ixp33_ASAP7_75t_L g1468 ( 
.A1(n_1448),
.A2(n_1406),
.B(n_1439),
.C(n_1434),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1411),
.B(n_1416),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1423),
.Y(n_1470)
);

OA21x2_ASAP7_75t_L g1471 ( 
.A1(n_1417),
.A2(n_1342),
.B(n_1365),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1430),
.B(n_1432),
.Y(n_1472)
);

O2A1O1Ixp5_ASAP7_75t_L g1473 ( 
.A1(n_1422),
.A2(n_1355),
.B(n_1434),
.C(n_1399),
.Y(n_1473)
);

A2O1A1Ixp33_ASAP7_75t_L g1474 ( 
.A1(n_1406),
.A2(n_1439),
.B(n_1353),
.C(n_1378),
.Y(n_1474)
);

OAI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1357),
.A2(n_1387),
.B1(n_1348),
.B2(n_1356),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1436),
.B(n_1438),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_1408),
.Y(n_1477)
);

INVx2_ASAP7_75t_SL g1478 ( 
.A(n_1361),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1387),
.B(n_1390),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1402),
.B(n_1404),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1402),
.B(n_1401),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1349),
.A2(n_1395),
.B1(n_1370),
.B2(n_1368),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1447),
.B(n_1351),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1400),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1419),
.B(n_1425),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1349),
.A2(n_1395),
.B1(n_1368),
.B2(n_1388),
.Y(n_1486)
);

BUFx8_ASAP7_75t_L g1487 ( 
.A(n_1350),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1397),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_1384),
.Y(n_1489)
);

INVxp67_ASAP7_75t_L g1490 ( 
.A(n_1382),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1364),
.A2(n_1386),
.B1(n_1405),
.B2(n_1375),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1409),
.B(n_1440),
.Y(n_1492)
);

O2A1O1Ixp33_ASAP7_75t_L g1493 ( 
.A1(n_1396),
.A2(n_1394),
.B(n_1383),
.C(n_1360),
.Y(n_1493)
);

O2A1O1Ixp33_ASAP7_75t_L g1494 ( 
.A1(n_1396),
.A2(n_1394),
.B(n_1383),
.C(n_1360),
.Y(n_1494)
);

O2A1O1Ixp5_ASAP7_75t_L g1495 ( 
.A1(n_1385),
.A2(n_1381),
.B(n_1369),
.C(n_1344),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1364),
.A2(n_1405),
.B1(n_1445),
.B2(n_1393),
.Y(n_1496)
);

O2A1O1Ixp33_ASAP7_75t_L g1497 ( 
.A1(n_1369),
.A2(n_1381),
.B(n_1344),
.C(n_1371),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1350),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1354),
.B(n_1393),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1380),
.B(n_1354),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1445),
.A2(n_1420),
.B1(n_1384),
.B2(n_1428),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_1433),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1433),
.A2(n_1345),
.B1(n_1442),
.B2(n_1435),
.Y(n_1503)
);

OAI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1345),
.A2(n_1431),
.B1(n_1435),
.B2(n_1426),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1345),
.A2(n_1431),
.B1(n_1435),
.B2(n_1426),
.Y(n_1505)
);

AOI211xp5_ASAP7_75t_L g1506 ( 
.A1(n_1379),
.A2(n_1444),
.B(n_1437),
.C(n_1427),
.Y(n_1506)
);

AOI221x1_ASAP7_75t_SL g1507 ( 
.A1(n_1414),
.A2(n_1427),
.B1(n_1437),
.B2(n_1407),
.C(n_1442),
.Y(n_1507)
);

OA22x2_ASAP7_75t_L g1508 ( 
.A1(n_1424),
.A2(n_1346),
.B1(n_1221),
.B2(n_1391),
.Y(n_1508)
);

AOI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1340),
.A2(n_1412),
.B(n_1339),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1339),
.B(n_1412),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1339),
.B(n_1412),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1367),
.Y(n_1512)
);

AOI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1340),
.A2(n_1412),
.B(n_1339),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1339),
.B(n_1412),
.Y(n_1514)
);

BUFx12f_ASAP7_75t_L g1515 ( 
.A(n_1408),
.Y(n_1515)
);

A2O1A1Ixp33_ASAP7_75t_L g1516 ( 
.A1(n_1339),
.A2(n_1412),
.B(n_1421),
.C(n_1418),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1340),
.A2(n_1412),
.B(n_1339),
.Y(n_1517)
);

OAI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1339),
.A2(n_1412),
.B1(n_1421),
.B2(n_1418),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1339),
.B(n_1412),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1339),
.A2(n_1412),
.B1(n_1421),
.B2(n_1418),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1343),
.B(n_1410),
.Y(n_1521)
);

NOR2xp67_ASAP7_75t_L g1522 ( 
.A(n_1391),
.B(n_1398),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1453),
.B(n_1512),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1464),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1500),
.B(n_1467),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1470),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1469),
.B(n_1472),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1476),
.B(n_1461),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1484),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1465),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1510),
.B(n_1511),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1510),
.B(n_1511),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1460),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1519),
.B(n_1450),
.Y(n_1534)
);

INVx4_ASAP7_75t_SL g1535 ( 
.A(n_1483),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1460),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1455),
.B(n_1456),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_L g1538 ( 
.A(n_1514),
.B(n_1450),
.Y(n_1538)
);

INVx3_ASAP7_75t_L g1539 ( 
.A(n_1471),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1518),
.B(n_1520),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1490),
.Y(n_1541)
);

OR2x6_ASAP7_75t_L g1542 ( 
.A(n_1491),
.B(n_1479),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1499),
.Y(n_1543)
);

OAI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1474),
.A2(n_1513),
.B(n_1451),
.Y(n_1544)
);

AO21x2_ASAP7_75t_L g1545 ( 
.A1(n_1504),
.A2(n_1505),
.B(n_1479),
.Y(n_1545)
);

AO21x2_ASAP7_75t_L g1546 ( 
.A1(n_1504),
.A2(n_1505),
.B(n_1503),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1503),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1521),
.B(n_1516),
.Y(n_1548)
);

AO21x2_ASAP7_75t_L g1549 ( 
.A1(n_1496),
.A2(n_1486),
.B(n_1491),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1495),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1493),
.Y(n_1551)
);

NOR2xp67_ASAP7_75t_L g1552 ( 
.A(n_1454),
.B(n_1488),
.Y(n_1552)
);

BUFx2_ASAP7_75t_L g1553 ( 
.A(n_1457),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1494),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1497),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1518),
.B(n_1520),
.Y(n_1556)
);

OAI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1508),
.A2(n_1458),
.B1(n_1509),
.B2(n_1517),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_1489),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1462),
.B(n_1463),
.Y(n_1559)
);

OR2x6_ASAP7_75t_L g1560 ( 
.A(n_1486),
.B(n_1482),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1452),
.B(n_1481),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1459),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1533),
.B(n_1507),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1529),
.Y(n_1564)
);

BUFx6f_ASAP7_75t_L g1565 ( 
.A(n_1546),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1539),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1529),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1539),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1525),
.B(n_1527),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1543),
.Y(n_1570)
);

OAI21xp33_ASAP7_75t_SL g1571 ( 
.A1(n_1538),
.A2(n_1449),
.B(n_1458),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1535),
.B(n_1539),
.Y(n_1572)
);

NOR2x1_ASAP7_75t_L g1573 ( 
.A(n_1552),
.B(n_1482),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1541),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1524),
.Y(n_1575)
);

INVxp67_ASAP7_75t_L g1576 ( 
.A(n_1536),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1536),
.B(n_1507),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1547),
.B(n_1475),
.Y(n_1578)
);

BUFx3_ASAP7_75t_L g1579 ( 
.A(n_1553),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1547),
.B(n_1508),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1545),
.B(n_1506),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1545),
.B(n_1457),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1545),
.B(n_1473),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1526),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1535),
.B(n_1492),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1545),
.B(n_1480),
.Y(n_1586)
);

NAND4xp25_ASAP7_75t_SL g1587 ( 
.A(n_1540),
.B(n_1468),
.C(n_1485),
.D(n_1515),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1546),
.B(n_1522),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1564),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1571),
.B(n_1544),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1564),
.Y(n_1591)
);

AO21x2_ASAP7_75t_L g1592 ( 
.A1(n_1581),
.A2(n_1550),
.B(n_1546),
.Y(n_1592)
);

OAI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1565),
.A2(n_1560),
.B1(n_1544),
.B2(n_1557),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1564),
.Y(n_1594)
);

INVxp67_ASAP7_75t_SL g1595 ( 
.A(n_1588),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1567),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1567),
.Y(n_1597)
);

NAND3xp33_ASAP7_75t_L g1598 ( 
.A(n_1588),
.B(n_1540),
.C(n_1556),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1567),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1574),
.Y(n_1600)
);

INVxp67_ASAP7_75t_L g1601 ( 
.A(n_1588),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1575),
.Y(n_1602)
);

AOI31xp33_ASAP7_75t_L g1603 ( 
.A1(n_1571),
.A2(n_1534),
.A3(n_1548),
.B(n_1501),
.Y(n_1603)
);

AOI33xp33_ASAP7_75t_L g1604 ( 
.A1(n_1588),
.A2(n_1578),
.A3(n_1583),
.B1(n_1580),
.B2(n_1581),
.B3(n_1532),
.Y(n_1604)
);

INVx1_ASAP7_75t_SL g1605 ( 
.A(n_1586),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1575),
.Y(n_1606)
);

OAI33xp33_ASAP7_75t_L g1607 ( 
.A1(n_1563),
.A2(n_1534),
.A3(n_1523),
.B1(n_1530),
.B2(n_1562),
.B3(n_1537),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1569),
.B(n_1528),
.Y(n_1608)
);

INVx3_ASAP7_75t_L g1609 ( 
.A(n_1572),
.Y(n_1609)
);

OAI221xp5_ASAP7_75t_SL g1610 ( 
.A1(n_1571),
.A2(n_1583),
.B1(n_1560),
.B2(n_1581),
.C(n_1578),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1584),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1580),
.B(n_1531),
.Y(n_1612)
);

AOI31xp33_ASAP7_75t_L g1613 ( 
.A1(n_1573),
.A2(n_1501),
.A3(n_1561),
.B(n_1466),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1580),
.A2(n_1560),
.B1(n_1549),
.B2(n_1559),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1569),
.B(n_1528),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1580),
.B(n_1531),
.Y(n_1616)
);

BUFx2_ASAP7_75t_L g1617 ( 
.A(n_1585),
.Y(n_1617)
);

BUFx2_ASAP7_75t_L g1618 ( 
.A(n_1582),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_1579),
.Y(n_1619)
);

OAI31xp33_ASAP7_75t_L g1620 ( 
.A1(n_1587),
.A2(n_1555),
.A3(n_1551),
.B(n_1554),
.Y(n_1620)
);

AOI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1587),
.A2(n_1549),
.B1(n_1542),
.B2(n_1555),
.Y(n_1621)
);

BUFx4f_ASAP7_75t_SL g1622 ( 
.A(n_1579),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1573),
.A2(n_1549),
.B(n_1542),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1574),
.Y(n_1624)
);

OAI211xp5_ASAP7_75t_SL g1625 ( 
.A1(n_1563),
.A2(n_1478),
.B(n_1537),
.C(n_1523),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1589),
.Y(n_1626)
);

CKINVDCx16_ASAP7_75t_R g1627 ( 
.A(n_1590),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1591),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1594),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1596),
.Y(n_1630)
);

NAND3xp33_ASAP7_75t_SL g1631 ( 
.A(n_1604),
.B(n_1583),
.C(n_1578),
.Y(n_1631)
);

INVxp67_ASAP7_75t_SL g1632 ( 
.A(n_1595),
.Y(n_1632)
);

BUFx4f_ASAP7_75t_L g1633 ( 
.A(n_1618),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1600),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1624),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1618),
.B(n_1601),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1604),
.B(n_1576),
.Y(n_1637)
);

OA21x2_ASAP7_75t_L g1638 ( 
.A1(n_1623),
.A2(n_1583),
.B(n_1568),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1598),
.B(n_1576),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1597),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1592),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1599),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1602),
.Y(n_1643)
);

NOR3xp33_ASAP7_75t_L g1644 ( 
.A(n_1590),
.B(n_1577),
.C(n_1563),
.Y(n_1644)
);

INVx4_ASAP7_75t_SL g1645 ( 
.A(n_1622),
.Y(n_1645)
);

OA21x2_ASAP7_75t_L g1646 ( 
.A1(n_1621),
.A2(n_1568),
.B(n_1566),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1606),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1592),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1592),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1619),
.Y(n_1650)
);

INVxp67_ASAP7_75t_L g1651 ( 
.A(n_1603),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1613),
.B(n_1477),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1617),
.B(n_1586),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1609),
.B(n_1582),
.Y(n_1654)
);

BUFx2_ASAP7_75t_L g1655 ( 
.A(n_1619),
.Y(n_1655)
);

HB1xp67_ASAP7_75t_L g1656 ( 
.A(n_1611),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1633),
.B(n_1608),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1633),
.B(n_1605),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1633),
.B(n_1608),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1656),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1631),
.A2(n_1620),
.B(n_1610),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1656),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1631),
.B(n_1612),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1626),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1626),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1628),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1634),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1638),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1634),
.Y(n_1669)
);

INVx2_ASAP7_75t_SL g1670 ( 
.A(n_1633),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1653),
.B(n_1615),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1650),
.B(n_1609),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1628),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1644),
.B(n_1616),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1644),
.B(n_1627),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1629),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_1650),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1655),
.B(n_1609),
.Y(n_1678)
);

BUFx2_ASAP7_75t_L g1679 ( 
.A(n_1645),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1655),
.B(n_1654),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1637),
.B(n_1577),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1627),
.B(n_1586),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1629),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1637),
.B(n_1577),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1630),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1635),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1639),
.B(n_1651),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1630),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1638),
.Y(n_1689)
);

INVx3_ASAP7_75t_L g1690 ( 
.A(n_1638),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1638),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1639),
.B(n_1586),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1640),
.Y(n_1693)
);

AND2x2_ASAP7_75t_SL g1694 ( 
.A(n_1638),
.B(n_1565),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1635),
.B(n_1570),
.Y(n_1695)
);

BUFx6f_ASAP7_75t_L g1696 ( 
.A(n_1646),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1640),
.Y(n_1697)
);

NAND2x1_ASAP7_75t_L g1698 ( 
.A(n_1657),
.B(n_1659),
.Y(n_1698)
);

NAND2x1p5_ASAP7_75t_L g1699 ( 
.A(n_1679),
.B(n_1585),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1660),
.Y(n_1700)
);

INVxp67_ASAP7_75t_L g1701 ( 
.A(n_1675),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1660),
.Y(n_1702)
);

NOR2x1_ASAP7_75t_L g1703 ( 
.A(n_1679),
.B(n_1652),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1696),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1657),
.B(n_1645),
.Y(n_1705)
);

AOI21xp33_ASAP7_75t_L g1706 ( 
.A1(n_1675),
.A2(n_1651),
.B(n_1565),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1662),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1662),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1659),
.B(n_1645),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1680),
.B(n_1645),
.Y(n_1710)
);

OAI21xp33_ASAP7_75t_L g1711 ( 
.A1(n_1661),
.A2(n_1636),
.B(n_1625),
.Y(n_1711)
);

AOI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_1687),
.A2(n_1607),
.B1(n_1565),
.B2(n_1593),
.C(n_1614),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1674),
.B(n_1681),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1674),
.B(n_1642),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1680),
.B(n_1645),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1667),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1672),
.B(n_1654),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1681),
.B(n_1642),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1684),
.B(n_1643),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1667),
.Y(n_1720)
);

OA21x2_ASAP7_75t_L g1721 ( 
.A1(n_1661),
.A2(n_1648),
.B(n_1641),
.Y(n_1721)
);

NAND2x1_ASAP7_75t_L g1722 ( 
.A(n_1658),
.B(n_1636),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1684),
.B(n_1643),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1669),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1669),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1686),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1686),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1664),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1664),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1687),
.B(n_1632),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1672),
.B(n_1636),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1663),
.B(n_1647),
.Y(n_1732)
);

INVxp67_ASAP7_75t_SL g1733 ( 
.A(n_1696),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1696),
.A2(n_1565),
.B1(n_1549),
.B2(n_1614),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1713),
.B(n_1677),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1718),
.B(n_1663),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1718),
.B(n_1692),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1720),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1720),
.Y(n_1739)
);

BUFx3_ASAP7_75t_L g1740 ( 
.A(n_1716),
.Y(n_1740)
);

BUFx3_ASAP7_75t_L g1741 ( 
.A(n_1724),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1728),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1719),
.B(n_1692),
.Y(n_1743)
);

NOR2xp33_ASAP7_75t_L g1744 ( 
.A(n_1710),
.B(n_1487),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1729),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1721),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1721),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1719),
.Y(n_1748)
);

INVxp67_ASAP7_75t_L g1749 ( 
.A(n_1710),
.Y(n_1749)
);

INVxp67_ASAP7_75t_L g1750 ( 
.A(n_1715),
.Y(n_1750)
);

INVx1_ASAP7_75t_SL g1751 ( 
.A(n_1715),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1723),
.Y(n_1752)
);

BUFx2_ASAP7_75t_L g1753 ( 
.A(n_1705),
.Y(n_1753)
);

INVx1_ASAP7_75t_SL g1754 ( 
.A(n_1705),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1725),
.Y(n_1755)
);

OAI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1711),
.A2(n_1682),
.B(n_1694),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_SL g1757 ( 
.A(n_1709),
.B(n_1696),
.Y(n_1757)
);

CKINVDCx16_ASAP7_75t_R g1758 ( 
.A(n_1709),
.Y(n_1758)
);

INVx2_ASAP7_75t_SL g1759 ( 
.A(n_1698),
.Y(n_1759)
);

AOI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1712),
.A2(n_1694),
.B(n_1682),
.Y(n_1760)
);

NOR2xp67_ASAP7_75t_L g1761 ( 
.A(n_1731),
.B(n_1670),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1753),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1752),
.B(n_1726),
.Y(n_1763)
);

AOI32xp33_ASAP7_75t_L g1764 ( 
.A1(n_1736),
.A2(n_1690),
.A3(n_1734),
.B1(n_1730),
.B2(n_1703),
.Y(n_1764)
);

INVxp67_ASAP7_75t_L g1765 ( 
.A(n_1753),
.Y(n_1765)
);

NOR3xp33_ASAP7_75t_L g1766 ( 
.A(n_1758),
.B(n_1701),
.C(n_1706),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1751),
.B(n_1731),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1754),
.B(n_1717),
.Y(n_1768)
);

INVxp67_ASAP7_75t_L g1769 ( 
.A(n_1744),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1752),
.B(n_1727),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1736),
.B(n_1714),
.Y(n_1771)
);

AOI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1746),
.A2(n_1721),
.B1(n_1734),
.B2(n_1696),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1755),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1748),
.B(n_1700),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1740),
.B(n_1702),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1740),
.B(n_1741),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1741),
.B(n_1707),
.Y(n_1777)
);

AOI211xp5_ASAP7_75t_SL g1778 ( 
.A1(n_1749),
.A2(n_1733),
.B(n_1708),
.C(n_1704),
.Y(n_1778)
);

AOI21xp5_ASAP7_75t_SL g1779 ( 
.A1(n_1757),
.A2(n_1704),
.B(n_1670),
.Y(n_1779)
);

NAND3xp33_ASAP7_75t_L g1780 ( 
.A(n_1756),
.B(n_1696),
.C(n_1565),
.Y(n_1780)
);

O2A1O1Ixp33_ASAP7_75t_L g1781 ( 
.A1(n_1746),
.A2(n_1690),
.B(n_1732),
.C(n_1668),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1759),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1767),
.Y(n_1783)
);

HB1xp67_ASAP7_75t_L g1784 ( 
.A(n_1765),
.Y(n_1784)
);

INVx2_ASAP7_75t_SL g1785 ( 
.A(n_1768),
.Y(n_1785)
);

NAND2x1_ASAP7_75t_L g1786 ( 
.A(n_1779),
.B(n_1759),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1762),
.B(n_1750),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1771),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1778),
.B(n_1735),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1782),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1776),
.B(n_1757),
.Y(n_1791)
);

AOI222xp33_ASAP7_75t_L g1792 ( 
.A1(n_1763),
.A2(n_1747),
.B1(n_1739),
.B2(n_1738),
.C1(n_1745),
.C2(n_1742),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1778),
.B(n_1761),
.Y(n_1793)
);

NAND2x1_ASAP7_75t_L g1794 ( 
.A(n_1773),
.B(n_1678),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_SL g1795 ( 
.A(n_1785),
.B(n_1764),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1783),
.Y(n_1796)
);

AOI221x1_ASAP7_75t_L g1797 ( 
.A1(n_1789),
.A2(n_1766),
.B1(n_1775),
.B2(n_1777),
.C(n_1747),
.Y(n_1797)
);

AOI211xp5_ASAP7_75t_L g1798 ( 
.A1(n_1793),
.A2(n_1781),
.B(n_1780),
.C(n_1769),
.Y(n_1798)
);

AOI211xp5_ASAP7_75t_L g1799 ( 
.A1(n_1791),
.A2(n_1788),
.B(n_1790),
.C(n_1787),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1786),
.A2(n_1763),
.B(n_1772),
.Y(n_1800)
);

NOR2xp33_ASAP7_75t_L g1801 ( 
.A(n_1794),
.B(n_1770),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1784),
.B(n_1774),
.Y(n_1802)
);

AOI211xp5_ASAP7_75t_L g1803 ( 
.A1(n_1792),
.A2(n_1760),
.B(n_1743),
.C(n_1737),
.Y(n_1803)
);

OAI221xp5_ASAP7_75t_L g1804 ( 
.A1(n_1792),
.A2(n_1690),
.B1(n_1691),
.B2(n_1668),
.C(n_1689),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1783),
.B(n_1737),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1786),
.A2(n_1722),
.B(n_1670),
.Y(n_1806)
);

O2A1O1Ixp33_ASAP7_75t_L g1807 ( 
.A1(n_1795),
.A2(n_1800),
.B(n_1802),
.C(n_1803),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1805),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1796),
.Y(n_1809)
);

NAND2xp33_ASAP7_75t_R g1810 ( 
.A(n_1801),
.B(n_1502),
.Y(n_1810)
);

NOR3xp33_ASAP7_75t_L g1811 ( 
.A(n_1798),
.B(n_1743),
.C(n_1690),
.Y(n_1811)
);

HB1xp67_ASAP7_75t_L g1812 ( 
.A(n_1799),
.Y(n_1812)
);

OAI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1797),
.A2(n_1699),
.B(n_1694),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1808),
.B(n_1806),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1812),
.Y(n_1815)
);

XOR2x2_ASAP7_75t_L g1816 ( 
.A(n_1811),
.B(n_1487),
.Y(n_1816)
);

AOI32xp33_ASAP7_75t_L g1817 ( 
.A1(n_1809),
.A2(n_1804),
.A3(n_1668),
.B1(n_1689),
.B2(n_1691),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1807),
.Y(n_1818)
);

INVxp67_ASAP7_75t_SL g1819 ( 
.A(n_1810),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1813),
.B(n_1665),
.Y(n_1820)
);

HB1xp67_ASAP7_75t_L g1821 ( 
.A(n_1814),
.Y(n_1821)
);

AO22x1_ASAP7_75t_L g1822 ( 
.A1(n_1819),
.A2(n_1810),
.B1(n_1498),
.B2(n_1558),
.Y(n_1822)
);

OAI221xp5_ASAP7_75t_L g1823 ( 
.A1(n_1817),
.A2(n_1689),
.B1(n_1691),
.B2(n_1699),
.C(n_1646),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_L g1824 ( 
.A(n_1818),
.B(n_1665),
.Y(n_1824)
);

NAND4xp75_ASAP7_75t_L g1825 ( 
.A(n_1815),
.B(n_1717),
.C(n_1658),
.D(n_1646),
.Y(n_1825)
);

AOI211xp5_ASAP7_75t_L g1826 ( 
.A1(n_1822),
.A2(n_1820),
.B(n_1816),
.C(n_1658),
.Y(n_1826)
);

CKINVDCx20_ASAP7_75t_R g1827 ( 
.A(n_1821),
.Y(n_1827)
);

NOR3xp33_ASAP7_75t_L g1828 ( 
.A(n_1824),
.B(n_1820),
.C(n_1648),
.Y(n_1828)
);

AND2x4_ASAP7_75t_L g1829 ( 
.A(n_1827),
.B(n_1678),
.Y(n_1829)
);

AOI322xp5_ASAP7_75t_L g1830 ( 
.A1(n_1829),
.A2(n_1828),
.A3(n_1825),
.B1(n_1823),
.B2(n_1826),
.C1(n_1641),
.C2(n_1648),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1830),
.Y(n_1831)
);

BUFx2_ASAP7_75t_L g1832 ( 
.A(n_1830),
.Y(n_1832)
);

OAI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1831),
.A2(n_1649),
.B(n_1641),
.Y(n_1833)
);

OAI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1832),
.A2(n_1695),
.B1(n_1697),
.B2(n_1693),
.Y(n_1834)
);

BUFx2_ASAP7_75t_L g1835 ( 
.A(n_1833),
.Y(n_1835)
);

OAI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1834),
.A2(n_1832),
.B1(n_1695),
.B2(n_1697),
.Y(n_1836)
);

XOR2xp5_ASAP7_75t_L g1837 ( 
.A(n_1836),
.B(n_1671),
.Y(n_1837)
);

AO221x2_ASAP7_75t_L g1838 ( 
.A1(n_1837),
.A2(n_1835),
.B1(n_1693),
.B2(n_1666),
.C(n_1673),
.Y(n_1838)
);

OAI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1838),
.A2(n_1649),
.B(n_1666),
.Y(n_1839)
);

AOI22xp33_ASAP7_75t_SL g1840 ( 
.A1(n_1839),
.A2(n_1649),
.B1(n_1673),
.B2(n_1676),
.Y(n_1840)
);

AOI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1840),
.A2(n_1676),
.B1(n_1683),
.B2(n_1685),
.Y(n_1841)
);

AOI211xp5_ASAP7_75t_L g1842 ( 
.A1(n_1841),
.A2(n_1685),
.B(n_1683),
.C(n_1688),
.Y(n_1842)
);


endmodule