module fake_jpeg_26614_n_314 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_314);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx2_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_26),
.B(n_35),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_25),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_46),
.Y(n_51)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_41),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_29),
.A2(n_18),
.B1(n_25),
.B2(n_24),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_45),
.A2(n_29),
.B1(n_33),
.B2(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_52),
.Y(n_79)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_69),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_54),
.B(n_61),
.Y(n_72)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_20),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_62),
.Y(n_73)
);

CKINVDCx9p33_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

BUFx2_ASAP7_75t_R g58 ( 
.A(n_44),
.Y(n_58)
);

AOI22x1_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_68),
.B1(n_44),
.B2(n_31),
.Y(n_75)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_32),
.B1(n_30),
.B2(n_26),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_65),
.B1(n_33),
.B2(n_26),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_31),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_24),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_41),
.A2(n_26),
.B1(n_30),
.B2(n_32),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_67),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_47),
.A2(n_24),
.B1(n_20),
.B2(n_22),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_61),
.B(n_58),
.Y(n_95)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_86),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_54),
.A2(n_20),
.B(n_22),
.C(n_24),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_19),
.B(n_61),
.Y(n_90)
);

MAJx2_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_43),
.C(n_29),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_37),
.C(n_43),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_66),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_37),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_37),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_60),
.A2(n_35),
.B1(n_69),
.B2(n_59),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_66),
.B1(n_64),
.B2(n_46),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_14),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_63),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_90),
.A2(n_95),
.B(n_96),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_93),
.Y(n_119)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_71),
.A2(n_52),
.B1(n_55),
.B2(n_53),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_97),
.B1(n_99),
.B2(n_102),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_72),
.A2(n_58),
.B(n_19),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_71),
.A2(n_52),
.B1(n_53),
.B2(n_64),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_85),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_98),
.B(n_100),
.Y(n_131)
);

AND2x6_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_81),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_104),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_105),
.Y(n_130)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_57),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_48),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_63),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_66),
.C(n_1),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_48),
.Y(n_108)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_83),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_112),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_48),
.C(n_39),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_89),
.C(n_80),
.Y(n_116)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_116),
.B(n_132),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_38),
.C(n_48),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_117),
.B(n_118),
.C(n_136),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_38),
.C(n_88),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_76),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_135),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_126),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_133),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_98),
.A2(n_79),
.B1(n_77),
.B2(n_70),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_128),
.A2(n_129),
.B1(n_34),
.B2(n_28),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_99),
.A2(n_79),
.B1(n_77),
.B2(n_70),
.Y(n_129)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_138),
.Y(n_166)
);

O2A1O1Ixp5_ASAP7_75t_L g135 ( 
.A1(n_100),
.A2(n_14),
.B(n_21),
.C(n_28),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_67),
.C(n_34),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_139),
.B(n_140),
.Y(n_151)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_31),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_104),
.A2(n_82),
.B1(n_67),
.B2(n_19),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_113),
.B1(n_93),
.B2(n_101),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_90),
.B(n_82),
.Y(n_143)
);

XNOR2x1_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_14),
.Y(n_169)
);

AO22x1_ASAP7_75t_SL g144 ( 
.A1(n_91),
.A2(n_87),
.B1(n_12),
.B2(n_17),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_23),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_87),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_145),
.A2(n_154),
.B(n_164),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_20),
.B(n_25),
.C(n_22),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_158),
.Y(n_185)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_153),
.Y(n_195)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_34),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_155),
.B(n_156),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_0),
.B(n_1),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_157),
.A2(n_165),
.B(n_172),
.Y(n_184)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_163),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_126),
.Y(n_160)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_160),
.Y(n_200)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_131),
.A2(n_19),
.B(n_22),
.Y(n_164)
);

AND2x6_ASAP7_75t_L g165 ( 
.A(n_115),
.B(n_0),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_167),
.A2(n_117),
.B1(n_125),
.B2(n_116),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_170),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_169),
.B(n_12),
.Y(n_197)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_142),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_115),
.A2(n_0),
.B(n_1),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_31),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_31),
.B(n_27),
.C(n_12),
.Y(n_199)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_114),
.Y(n_174)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

OA21x2_ASAP7_75t_L g188 ( 
.A1(n_175),
.A2(n_161),
.B(n_167),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_118),
.B(n_21),
.Y(n_176)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_122),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_132),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_180),
.B(n_207),
.Y(n_226)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_178),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_191),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_187),
.A2(n_206),
.B1(n_168),
.B2(n_159),
.Y(n_214)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_190),
.Y(n_231)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_146),
.A2(n_1),
.B(n_2),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_171),
.C(n_176),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_148),
.C(n_169),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_147),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_196),
.B(n_205),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_197),
.B(n_13),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_2),
.B(n_3),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_SL g212 ( 
.A(n_198),
.B(n_184),
.C(n_157),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_175),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_154),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_145),
.A2(n_23),
.B1(n_17),
.B2(n_15),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_162),
.B(n_21),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_148),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_208),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_216),
.C(n_218),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_211),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_212),
.B(n_215),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_214),
.A2(n_220),
.B1(n_229),
.B2(n_179),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_183),
.A2(n_145),
.B1(n_150),
.B2(n_165),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_173),
.C(n_164),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_197),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_180),
.B(n_23),
.C(n_17),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_202),
.A2(n_23),
.B1(n_17),
.B2(n_15),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_186),
.C(n_187),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_225),
.C(n_227),
.Y(n_235)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_223),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_23),
.C(n_17),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_23),
.C(n_17),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_184),
.A2(n_15),
.B1(n_21),
.B2(n_14),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_190),
.B(n_201),
.Y(n_230)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_230),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_234),
.A2(n_236),
.B1(n_239),
.B2(n_248),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_221),
.A2(n_203),
.B1(n_188),
.B2(n_189),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_244),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_209),
.A2(n_188),
.B1(n_179),
.B2(n_181),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_231),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_245),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_181),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_208),
.A2(n_200),
.B1(n_182),
.B2(n_185),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_218),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_224),
.A2(n_185),
.B1(n_206),
.B2(n_191),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_250),
.B(n_199),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_247),
.A2(n_219),
.B1(n_222),
.B2(n_211),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_251),
.A2(n_255),
.B1(n_4),
.B2(n_5),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_239),
.A2(n_198),
.B(n_216),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_253),
.A2(n_235),
.B(n_232),
.Y(n_270)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_233),
.A2(n_210),
.B1(n_226),
.B2(n_217),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_248),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_257),
.Y(n_266)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_236),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_262),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_261),
.B(n_264),
.Y(n_267)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_246),
.A2(n_2),
.B(n_3),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_263),
.A2(n_265),
.B(n_3),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_15),
.C(n_16),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_21),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_244),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_272),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_253),
.A2(n_241),
.B1(n_238),
.B2(n_235),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_269),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_13),
.B(n_6),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_237),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_276),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_274),
.A2(n_264),
.B1(n_252),
.B2(n_6),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_259),
.A2(n_16),
.B(n_14),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_275),
.A2(n_13),
.B(n_16),
.Y(n_284)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_15),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_5),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_289),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_4),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_280),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_4),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_285),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_284),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_267),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_287),
.C(n_288),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_16),
.C(n_13),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_16),
.C(n_13),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_7),
.Y(n_298)
);

NAND2xp33_ASAP7_75t_SL g291 ( 
.A(n_286),
.B(n_269),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_295),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_282),
.A2(n_283),
.B(n_288),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_268),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_298),
.Y(n_301)
);

NAND3xp33_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_276),
.C(n_8),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_9),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_8),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_302),
.A2(n_303),
.B(n_304),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_9),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_16),
.C(n_13),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_306),
.A2(n_293),
.B(n_297),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_301),
.C(n_292),
.Y(n_309)
);

A2O1A1Ixp33_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_305),
.B(n_301),
.C(n_294),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_310),
.A2(n_307),
.B(n_11),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_10),
.C(n_11),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_10),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_10),
.B(n_13),
.Y(n_314)
);


endmodule