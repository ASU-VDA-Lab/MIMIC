module fake_jpeg_13150_n_476 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_476);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_476;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_352;
wire n_350;
wire n_150;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_46),
.Y(n_111)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_48),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_50),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_12),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_51),
.B(n_65),
.Y(n_125)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_53),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_61),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_41),
.B(n_12),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_14),
.Y(n_69)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_70),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_27),
.B(n_11),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_71),
.B(n_96),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_72),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_74),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_75),
.Y(n_154)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_77),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_14),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_83),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_80),
.Y(n_146)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_13),
.Y(n_82)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx6_ASAP7_75t_SL g83 ( 
.A(n_14),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g148 ( 
.A(n_85),
.Y(n_148)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_13),
.Y(n_86)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_87),
.Y(n_153)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_13),
.Y(n_88)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_13),
.Y(n_90)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_14),
.Y(n_91)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_93),
.B(n_95),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_97),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_14),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_100),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_31),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_99),
.A2(n_27),
.B1(n_29),
.B2(n_36),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_15),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_15),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_101),
.B(n_15),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_29),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_108),
.B(n_42),
.Y(n_195)
);

AOI21xp33_ASAP7_75t_SL g113 ( 
.A1(n_51),
.A2(n_14),
.B(n_16),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_L g199 ( 
.A1(n_113),
.A2(n_24),
.B(n_23),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_69),
.A2(n_41),
.B1(n_26),
.B2(n_16),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_130),
.A2(n_132),
.B1(n_136),
.B2(n_143),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_58),
.A2(n_41),
.B1(n_16),
.B2(n_45),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_91),
.A2(n_16),
.B1(n_97),
.B2(n_39),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_76),
.A2(n_16),
.B1(n_39),
.B2(n_15),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_149),
.A2(n_42),
.B1(n_40),
.B2(n_23),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_65),
.B(n_36),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_156),
.B(n_157),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_75),
.B(n_45),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_125),
.B(n_33),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_160),
.B(n_184),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_158),
.A2(n_85),
.B1(n_92),
.B2(n_87),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_162),
.A2(n_163),
.B1(n_186),
.B2(n_40),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_119),
.A2(n_28),
.B1(n_22),
.B2(n_25),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_166),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_105),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_167),
.B(n_190),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_119),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_176),
.Y(n_210)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_169),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_132),
.A2(n_93),
.B1(n_96),
.B2(n_95),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_170),
.A2(n_183),
.B1(n_191),
.B2(n_196),
.Y(n_223)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_171),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

INVxp67_ASAP7_75t_SL g214 ( 
.A(n_172),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_173),
.Y(n_234)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_174),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_60),
.B1(n_84),
.B2(n_80),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_175),
.A2(n_148),
.B1(n_124),
.B2(n_140),
.Y(n_229)
);

AND2x4_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_16),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_112),
.Y(n_178)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_178),
.Y(n_228)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_138),
.Y(n_179)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_118),
.B(n_121),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_180),
.B(n_145),
.C(n_116),
.Y(n_226)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_182),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_143),
.A2(n_136),
.B1(n_130),
.B2(n_108),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_103),
.B(n_24),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_185),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_159),
.A2(n_49),
.B1(n_79),
.B2(n_73),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_188),
.Y(n_225)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_109),
.Y(n_189)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_189),
.Y(n_238)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_126),
.A2(n_66),
.B1(n_54),
.B2(n_98),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_126),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_195),
.Y(n_227)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_115),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_193),
.Y(n_217)
);

INVx11_ASAP7_75t_L g194 ( 
.A(n_104),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_194),
.A2(n_201),
.B1(n_202),
.B2(n_204),
.Y(n_218)
);

AO22x1_ASAP7_75t_SL g197 ( 
.A1(n_104),
.A2(n_38),
.B1(n_28),
.B2(n_25),
.Y(n_197)
);

AO22x1_ASAP7_75t_SL g212 ( 
.A1(n_197),
.A2(n_169),
.B1(n_194),
.B2(n_179),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_145),
.B(n_15),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_198),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_128),
.Y(n_208)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_107),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_127),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_131),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_111),
.A2(n_38),
.B1(n_22),
.B2(n_33),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_107),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_203),
.Y(n_236)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_129),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_208),
.Y(n_261)
);

NOR2x1p5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_32),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_209),
.B(n_212),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_161),
.B(n_120),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_211),
.B(n_180),
.C(n_171),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_222),
.A2(n_230),
.B1(n_170),
.B2(n_191),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_223),
.A2(n_163),
.B1(n_176),
.B2(n_114),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_226),
.B(n_176),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_229),
.A2(n_133),
.B1(n_117),
.B2(n_146),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_175),
.A2(n_114),
.B1(n_148),
.B2(n_146),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_233),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_161),
.B(n_129),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_235),
.B(n_197),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_239),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_231),
.A2(n_183),
.B1(n_187),
.B2(n_168),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_240),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_242),
.A2(n_246),
.B1(n_251),
.B2(n_262),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_243),
.A2(n_254),
.B1(n_258),
.B2(n_173),
.Y(n_277)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_237),
.Y(n_244)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_244),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_211),
.B(n_160),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_248),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_223),
.A2(n_192),
.B1(n_185),
.B2(n_180),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_210),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_247),
.B(n_253),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_219),
.B(n_167),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_232),
.B(n_164),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_265),
.Y(n_276)
);

AOI32xp33_ASAP7_75t_L g250 ( 
.A1(n_208),
.A2(n_200),
.A3(n_188),
.B1(n_181),
.B2(n_94),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_250),
.A2(n_217),
.B(n_216),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_233),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_231),
.A2(n_133),
.B1(n_117),
.B2(n_109),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_237),
.Y(n_255)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_260),
.C(n_226),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_212),
.A2(n_140),
.B1(n_124),
.B2(n_127),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_225),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_263),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_174),
.C(n_203),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_229),
.A2(n_197),
.B1(n_190),
.B2(n_165),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_210),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_227),
.B(n_225),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_264),
.B(n_259),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_210),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_224),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_241),
.B(n_235),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_267),
.B(n_280),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_252),
.A2(n_218),
.B(n_209),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_269),
.A2(n_290),
.B(n_293),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_248),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_271),
.B(n_275),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_252),
.Y(n_273)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_273),
.Y(n_307)
);

NAND2xp33_ASAP7_75t_SL g274 ( 
.A(n_247),
.B(n_209),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_274),
.A2(n_220),
.B(n_207),
.Y(n_311)
);

OA21x2_ASAP7_75t_L g275 ( 
.A1(n_265),
.A2(n_212),
.B(n_230),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_277),
.A2(n_256),
.B1(n_234),
.B2(n_205),
.Y(n_320)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_244),
.Y(n_281)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_281),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_255),
.Y(n_282)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_282),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_257),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_288),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_246),
.A2(n_206),
.B1(n_217),
.B2(n_238),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_289),
.A2(n_292),
.B1(n_258),
.B2(n_254),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_264),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_291),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_240),
.A2(n_206),
.B1(n_220),
.B2(n_207),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_239),
.A2(n_253),
.B(n_261),
.Y(n_293)
);

INVxp33_ASAP7_75t_L g295 ( 
.A(n_288),
.Y(n_295)
);

INVx11_ASAP7_75t_L g344 ( 
.A(n_295),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_296),
.B(n_304),
.C(n_312),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_267),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_297),
.B(n_302),
.Y(n_326)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_298),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_277),
.A2(n_242),
.B1(n_241),
.B2(n_262),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_299),
.A2(n_320),
.B1(n_279),
.B2(n_275),
.Y(n_343)
);

OA21x2_ASAP7_75t_L g300 ( 
.A1(n_273),
.A2(n_251),
.B(n_243),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_300),
.A2(n_275),
.B(n_277),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_275),
.A2(n_257),
.B1(n_266),
.B2(n_250),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_245),
.C(n_260),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_271),
.B(n_249),
.Y(n_305)
);

AOI21xp33_ASAP7_75t_L g336 ( 
.A1(n_305),
.A2(n_276),
.B(n_270),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_275),
.A2(n_260),
.B1(n_251),
.B2(n_256),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_306),
.B(n_310),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_289),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_311),
.A2(n_274),
.B(n_286),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_284),
.B(n_216),
.C(n_236),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_268),
.Y(n_313)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_313),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_283),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_314),
.B(n_315),
.Y(n_337)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_268),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_281),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_317),
.Y(n_322)
);

NAND3xp33_ASAP7_75t_L g319 ( 
.A(n_280),
.B(n_276),
.C(n_286),
.Y(n_319)
);

NOR3xp33_ASAP7_75t_SL g338 ( 
.A(n_319),
.B(n_291),
.C(n_283),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_296),
.B(n_278),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_321),
.B(n_330),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_318),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_323),
.B(n_333),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_324),
.A2(n_327),
.B(n_329),
.Y(n_369)
);

OAI31xp33_ASAP7_75t_L g361 ( 
.A1(n_325),
.A2(n_300),
.A3(n_298),
.B(n_309),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_308),
.A2(n_285),
.B(n_293),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_304),
.B(n_270),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_328),
.B(n_316),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_308),
.A2(n_290),
.B(n_293),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_312),
.B(n_302),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_318),
.A2(n_273),
.B(n_269),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_294),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_334),
.B(n_335),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_294),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_336),
.Y(n_355)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_338),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_311),
.B(n_292),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_342),
.C(n_345),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_314),
.B(n_292),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_343),
.A2(n_346),
.B1(n_282),
.B2(n_272),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_297),
.B(n_269),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_299),
.A2(n_279),
.B1(n_282),
.B2(n_272),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_320),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_347),
.B(n_316),
.Y(n_349)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_349),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_343),
.A2(n_306),
.B1(n_310),
.B2(n_307),
.Y(n_350)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_350),
.Y(n_376)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_337),
.Y(n_352)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_352),
.Y(n_381)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_337),
.Y(n_353)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_353),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_354),
.B(n_324),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_321),
.B(n_330),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_356),
.B(n_357),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_328),
.B(n_340),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_340),
.B(n_301),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_359),
.B(n_341),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_345),
.B(n_307),
.C(n_315),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_360),
.B(n_362),
.C(n_364),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_361),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_329),
.B(n_317),
.C(n_313),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_322),
.Y(n_363)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_363),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_326),
.B(n_342),
.C(n_327),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_331),
.A2(n_300),
.B1(n_303),
.B2(n_309),
.Y(n_365)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_365),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_326),
.B(n_303),
.C(n_300),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_366),
.B(n_341),
.C(n_287),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_367),
.B(n_325),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_331),
.A2(n_287),
.B1(n_205),
.B2(n_234),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_368),
.B(n_370),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_344),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_351),
.A2(n_346),
.B1(n_332),
.B2(n_338),
.Y(n_373)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_373),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_348),
.B(n_344),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_375),
.B(n_384),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_377),
.A2(n_362),
.B1(n_369),
.B2(n_360),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_382),
.B(n_388),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_355),
.B(n_213),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_366),
.A2(n_332),
.B1(n_333),
.B2(n_339),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_385),
.A2(n_393),
.B1(n_178),
.B2(n_177),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_359),
.B(n_213),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_386),
.B(n_392),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_389),
.B(n_221),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_371),
.B(n_214),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_391),
.B(n_368),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_372),
.A2(n_287),
.B1(n_228),
.B2(n_189),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_364),
.A2(n_228),
.B1(n_201),
.B2(n_193),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_378),
.B(n_357),
.C(n_371),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_395),
.B(n_399),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_374),
.Y(n_396)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_396),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_397),
.B(n_406),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_378),
.A2(n_358),
.B(n_369),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_388),
.B(n_356),
.C(n_358),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_400),
.B(n_407),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_382),
.A2(n_361),
.B(n_354),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g414 ( 
.A(n_401),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_379),
.A2(n_350),
.B(n_365),
.Y(n_403)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_403),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_389),
.B(n_221),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_408),
.B(n_413),
.Y(n_420)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_394),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_409),
.B(n_387),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_410),
.B(n_411),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_376),
.A2(n_215),
.B1(n_111),
.B2(n_150),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_385),
.B(n_215),
.C(n_204),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_412),
.B(n_394),
.C(n_390),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_376),
.A2(n_150),
.B1(n_131),
.B2(n_154),
.Y(n_413)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_415),
.Y(n_436)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_418),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_408),
.B(n_377),
.C(n_390),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_421),
.B(n_422),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_402),
.B(n_383),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_SL g423 ( 
.A1(n_405),
.A2(n_379),
.B1(n_381),
.B2(n_393),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_423),
.A2(n_412),
.B1(n_413),
.B2(n_406),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_396),
.B(n_383),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_424),
.B(n_10),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_395),
.B(n_380),
.C(n_391),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_425),
.B(n_397),
.Y(n_431)
);

FAx1_ASAP7_75t_SL g426 ( 
.A(n_400),
.B(n_380),
.CI(n_10),
.CON(n_426),
.SN(n_426)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_426),
.B(n_414),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_403),
.A2(n_110),
.B(n_142),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_428),
.A2(n_0),
.B(n_2),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_431),
.B(n_437),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_429),
.B(n_404),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_432),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_419),
.A2(n_410),
.B1(n_398),
.B2(n_411),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_433),
.B(n_435),
.Y(n_446)
);

MAJx2_ASAP7_75t_L g450 ( 
.A(n_434),
.B(n_418),
.C(n_420),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_417),
.B(n_404),
.Y(n_435)
);

NAND3xp33_ASAP7_75t_L g439 ( 
.A(n_427),
.B(n_9),
.C(n_8),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_439),
.B(n_440),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_416),
.B(n_0),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_429),
.B(n_32),
.C(n_1),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_442),
.B(n_444),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_443),
.B(n_3),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_441),
.B(n_421),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_448),
.B(n_451),
.Y(n_456)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_450),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_432),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_436),
.B(n_439),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_452),
.B(n_453),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_438),
.B(n_423),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_454),
.B(n_3),
.Y(n_461)
);

NAND2xp33_ASAP7_75t_L g457 ( 
.A(n_446),
.B(n_426),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_457),
.A2(n_458),
.B(n_460),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_451),
.A2(n_425),
.B(n_442),
.Y(n_458)
);

OR2x6_ASAP7_75t_SL g460 ( 
.A(n_445),
.B(n_430),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_461),
.B(n_3),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_449),
.Y(n_463)
);

OA21x2_ASAP7_75t_L g468 ( 
.A1(n_463),
.A2(n_420),
.B(n_4),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_456),
.A2(n_455),
.B(n_447),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_464),
.B(n_465),
.C(n_468),
.Y(n_469)
);

O2A1O1Ixp33_ASAP7_75t_SL g467 ( 
.A1(n_462),
.A2(n_434),
.B(n_450),
.C(n_430),
.Y(n_467)
);

AOI321xp33_ASAP7_75t_L g471 ( 
.A1(n_467),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_466),
.B(n_459),
.C(n_460),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_470),
.B(n_471),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_469),
.B(n_7),
.C(n_3),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_472),
.B(n_4),
.C(n_7),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_474),
.B(n_473),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_475),
.Y(n_476)
);


endmodule