module fake_jpeg_19633_n_188 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_188);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_SL g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_2),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_44),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_2),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_33),
.B(n_40),
.Y(n_64)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_21),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_25),
.B(n_2),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_25),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_49),
.B(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_26),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_40),
.B(n_32),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_32),
.Y(n_67)
);

OR2x2_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_20),
.Y(n_57)
);

OR2x2_ASAP7_75t_SL g81 ( 
.A(n_57),
.B(n_20),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_61),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_19),
.Y(n_60)
);

AO21x1_ASAP7_75t_L g89 ( 
.A1(n_60),
.A2(n_62),
.B(n_35),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_31),
.B(n_26),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_57),
.A2(n_41),
.B1(n_29),
.B2(n_44),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_65),
.A2(n_69),
.B1(n_72),
.B2(n_76),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_67),
.B(n_80),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_36),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_68),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_50),
.A2(n_23),
.B1(n_29),
.B2(n_27),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_34),
.B1(n_41),
.B2(n_43),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_71),
.A2(n_75),
.B1(n_63),
.B2(n_52),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_43),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_77),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_58),
.A2(n_34),
.B1(n_43),
.B2(n_38),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_23),
.B1(n_16),
.B2(n_24),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_24),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_78),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_20),
.B(n_15),
.C(n_19),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_85),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_15),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_3),
.B(n_4),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_47),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_82),
.B(n_84),
.Y(n_115)
);

INVx5_ASAP7_75t_SL g83 ( 
.A(n_47),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_86),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_19),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_60),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_19),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_90),
.Y(n_113)
);

NAND2x1_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_35),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_18),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_97),
.B1(n_100),
.B2(n_114),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_71),
.A2(n_63),
.B1(n_52),
.B2(n_56),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_67),
.A2(n_35),
.B1(n_37),
.B2(n_24),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_79),
.Y(n_124)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_108),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_73),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_74),
.A2(n_90),
.B1(n_85),
.B2(n_77),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_124),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_70),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_120),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_96),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_66),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_121),
.B(n_132),
.Y(n_135)
);

AND2x6_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_81),
.Y(n_123)
);

A2O1A1O1Ixp25_ASAP7_75t_L g133 ( 
.A1(n_123),
.A2(n_125),
.B(n_110),
.C(n_102),
.D(n_114),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_109),
.A2(n_68),
.B(n_89),
.C(n_20),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_75),
.B(n_92),
.C(n_87),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_127),
.A2(n_115),
.B(n_111),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_128),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_68),
.B1(n_83),
.B2(n_23),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_129),
.A2(n_130),
.B1(n_94),
.B2(n_106),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_102),
.A2(n_91),
.B1(n_88),
.B2(n_35),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_101),
.B(n_13),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_133),
.A2(n_138),
.B(n_141),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_122),
.A2(n_113),
.B(n_99),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_132),
.B(n_120),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_122),
.A2(n_99),
.B(n_96),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_100),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_146),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_144),
.A2(n_127),
.B1(n_130),
.B2(n_116),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_118),
.Y(n_145)
);

NOR3xp33_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_131),
.C(n_117),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_124),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_144),
.B1(n_140),
.B2(n_142),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_148),
.B(n_135),
.Y(n_167)
);

AOI21xp33_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_129),
.B(n_126),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_150),
.B(n_153),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_151),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_116),
.C(n_95),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_133),
.C(n_18),
.Y(n_164)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_154),
.Y(n_165)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_155),
.A2(n_107),
.B1(n_95),
.B2(n_137),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_93),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_136),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_162),
.B(n_152),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_164),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_147),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_166),
.A2(n_157),
.B(n_148),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_174),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_159),
.B(n_158),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_170),
.B(n_165),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_171),
.A2(n_162),
.B1(n_163),
.B2(n_165),
.Y(n_175)
);

AOI31xp67_ASAP7_75t_L g172 ( 
.A1(n_167),
.A2(n_157),
.A3(n_158),
.B(n_156),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_172),
.A2(n_28),
.B(n_11),
.C(n_37),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_175),
.A2(n_176),
.B(n_178),
.Y(n_180)
);

OAI221xp5_ASAP7_75t_L g181 ( 
.A1(n_177),
.A2(n_11),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_173),
.A2(n_168),
.B(n_169),
.Y(n_178)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_181),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_179),
.A2(n_28),
.B1(n_5),
.B2(n_7),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_3),
.B1(n_5),
.B2(n_8),
.Y(n_183)
);

OAI21x1_ASAP7_75t_L g185 ( 
.A1(n_183),
.A2(n_180),
.B(n_8),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_185),
.A2(n_184),
.B1(n_8),
.B2(n_9),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_9),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_9),
.Y(n_188)
);


endmodule