module fake_netlist_6_149_n_2340 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_507, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_396, n_495, n_350, n_78, n_84, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_522, n_466, n_506, n_56, n_360, n_119, n_235, n_536, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_521, n_363, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_513, n_321, n_331, n_105, n_227, n_132, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_33, n_477, n_533, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_537, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_487, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2340);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_507;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_536;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_33;
input n_477;
input n_533;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_537;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2340;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2291;
wire n_830;
wire n_2299;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2129;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_572;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2207;
wire n_1970;
wire n_608;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_2073;
wire n_2273;
wire n_792;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2193;
wire n_1655;
wire n_928;
wire n_1214;
wire n_835;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_2178;
wire n_950;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_2069;
wire n_2307;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_2231;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_811;
wire n_683;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2204;
wire n_1520;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2289;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_1905;
wire n_2016;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_2278;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_2302;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_1997;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_654;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_806;
wire n_959;
wire n_879;
wire n_2310;
wire n_584;
wire n_2141;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_1045;
wire n_706;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_646;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_1283;
wire n_918;
wire n_748;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_2287;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_1028;
wire n_576;
wire n_2106;
wire n_2265;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_709;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_924;
wire n_1582;
wire n_2318;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_570;
wire n_2033;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_1218;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_985;
wire n_2233;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1996;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_1025;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_364),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_153),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_36),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_326),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_496),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_421),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_45),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_319),
.Y(n_551)
);

BUFx10_ASAP7_75t_L g552 ( 
.A(n_370),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_343),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_348),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_129),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_415),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_440),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_63),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_154),
.Y(n_559)
);

BUFx2_ASAP7_75t_L g560 ( 
.A(n_487),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_371),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_494),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_9),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_533),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_477),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_384),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_2),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_102),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_8),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_132),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_301),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_423),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_50),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_501),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_332),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_383),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_377),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_512),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_472),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_276),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_136),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_135),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_377),
.Y(n_583)
);

CKINVDCx16_ASAP7_75t_R g584 ( 
.A(n_242),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_316),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_410),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_300),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_204),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_137),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_373),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_462),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_231),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_95),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_446),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_205),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_212),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_354),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_468),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_543),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_190),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_91),
.Y(n_601)
);

BUFx10_ASAP7_75t_L g602 ( 
.A(n_203),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_397),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_19),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_90),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_195),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_109),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_11),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_482),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_529),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_288),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_82),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_382),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_444),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_91),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_153),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_145),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_233),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_226),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_471),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_126),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_264),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_499),
.Y(n_623)
);

BUFx2_ASAP7_75t_L g624 ( 
.A(n_73),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_461),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_283),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_78),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_68),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_380),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_378),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_264),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_328),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_233),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_226),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_204),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_355),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_414),
.Y(n_637)
);

INVx1_ASAP7_75t_SL g638 ( 
.A(n_320),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_261),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_344),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_162),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_520),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_346),
.Y(n_643)
);

BUFx10_ASAP7_75t_L g644 ( 
.A(n_287),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_164),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_95),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_244),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_347),
.Y(n_648)
);

CKINVDCx16_ASAP7_75t_R g649 ( 
.A(n_2),
.Y(n_649)
);

INVx1_ASAP7_75t_SL g650 ( 
.A(n_515),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_144),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_522),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_465),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_441),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_279),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_418),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_509),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_232),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_390),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_183),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_230),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_261),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_56),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_30),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_365),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_98),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_191),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_53),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_189),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_167),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_73),
.Y(n_671)
);

INVx1_ASAP7_75t_SL g672 ( 
.A(n_80),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_257),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_202),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_117),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_521),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_511),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_184),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_83),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_513),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_106),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_416),
.Y(n_682)
);

BUFx3_ASAP7_75t_L g683 ( 
.A(n_448),
.Y(n_683)
);

BUFx8_ASAP7_75t_SL g684 ( 
.A(n_319),
.Y(n_684)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_532),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_54),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_45),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_60),
.Y(n_688)
);

BUFx5_ASAP7_75t_L g689 ( 
.A(n_154),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_117),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_265),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_324),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_334),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_313),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_445),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_484),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_139),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_430),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_454),
.Y(n_699)
);

CKINVDCx20_ASAP7_75t_R g700 ( 
.A(n_271),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_35),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_54),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_387),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_523),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_188),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_466),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_127),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_15),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_330),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_74),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_493),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_248),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_283),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_220),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_194),
.Y(n_715)
);

BUFx10_ASAP7_75t_L g716 ( 
.A(n_436),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_166),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_381),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_61),
.Y(n_719)
);

HB1xp67_ASAP7_75t_L g720 ( 
.A(n_85),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_122),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_38),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_216),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_528),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_27),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_64),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_167),
.Y(n_727)
);

BUFx10_ASAP7_75t_L g728 ( 
.A(n_417),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_309),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_51),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_292),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_428),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_196),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_476),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_278),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_375),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_442),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_5),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_87),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_185),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_327),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_61),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_134),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_198),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_170),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_303),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_178),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_14),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_481),
.Y(n_749)
);

BUFx10_ASAP7_75t_L g750 ( 
.A(n_366),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_307),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_470),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_301),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_374),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_222),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_309),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_459),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_224),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_230),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_83),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_684),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_689),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_689),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_689),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_689),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_680),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_689),
.Y(n_767)
);

CKINVDCx16_ASAP7_75t_R g768 ( 
.A(n_584),
.Y(n_768)
);

INVxp33_ASAP7_75t_L g769 ( 
.A(n_720),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_689),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_689),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_660),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_680),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_684),
.Y(n_774)
);

HB1xp67_ASAP7_75t_L g775 ( 
.A(n_649),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_683),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_660),
.Y(n_777)
);

INVxp67_ASAP7_75t_SL g778 ( 
.A(n_560),
.Y(n_778)
);

CKINVDCx20_ASAP7_75t_R g779 ( 
.A(n_554),
.Y(n_779)
);

BUFx10_ASAP7_75t_L g780 ( 
.A(n_561),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_561),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_561),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_561),
.Y(n_783)
);

INVxp33_ASAP7_75t_SL g784 ( 
.A(n_559),
.Y(n_784)
);

NOR2xp67_ASAP7_75t_L g785 ( 
.A(n_567),
.B(n_0),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_612),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_544),
.Y(n_787)
);

INVxp33_ASAP7_75t_L g788 ( 
.A(n_573),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_624),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_612),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_691),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_691),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_712),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_712),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_612),
.Y(n_795)
);

INVxp33_ASAP7_75t_L g796 ( 
.A(n_645),
.Y(n_796)
);

INVxp33_ASAP7_75t_L g797 ( 
.A(n_713),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_667),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_667),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_546),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_667),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_667),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_683),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_555),
.Y(n_804)
);

NOR2xp67_ASAP7_75t_L g805 ( 
.A(n_621),
.B(n_0),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_571),
.Y(n_806)
);

INVxp67_ASAP7_75t_SL g807 ( 
.A(n_565),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_575),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_559),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_577),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_581),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_563),
.Y(n_812)
);

CKINVDCx14_ASAP7_75t_R g813 ( 
.A(n_552),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_590),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_605),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_606),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_611),
.Y(n_817)
);

INVxp33_ASAP7_75t_SL g818 ( 
.A(n_563),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_613),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_616),
.Y(n_820)
);

CKINVDCx14_ASAP7_75t_R g821 ( 
.A(n_552),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_545),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_547),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_627),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_628),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_631),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_633),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_545),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_639),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_655),
.Y(n_830)
);

INVxp67_ASAP7_75t_SL g831 ( 
.A(n_572),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_550),
.Y(n_832)
);

CKINVDCx16_ASAP7_75t_R g833 ( 
.A(n_574),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_669),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_675),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_551),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_549),
.B(n_3),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_626),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_708),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_710),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_714),
.Y(n_841)
);

INVxp33_ASAP7_75t_L g842 ( 
.A(n_626),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_715),
.Y(n_843)
);

INVx1_ASAP7_75t_SL g844 ( 
.A(n_552),
.Y(n_844)
);

NOR2xp67_ASAP7_75t_L g845 ( 
.A(n_621),
.B(n_1),
.Y(n_845)
);

OR2x2_ASAP7_75t_L g846 ( 
.A(n_718),
.B(n_1),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_549),
.Y(n_847)
);

INVxp33_ASAP7_75t_SL g848 ( 
.A(n_566),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_719),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_730),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_739),
.Y(n_851)
);

INVx1_ASAP7_75t_SL g852 ( 
.A(n_602),
.Y(n_852)
);

INVxp33_ASAP7_75t_L g853 ( 
.A(n_646),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_566),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_646),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_663),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_553),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_742),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_847),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_781),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_847),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_847),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_766),
.B(n_707),
.Y(n_863)
);

AND2x2_ASAP7_75t_SL g864 ( 
.A(n_837),
.B(n_591),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_847),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_781),
.Y(n_866)
);

OR2x2_ASAP7_75t_L g867 ( 
.A(n_844),
.B(n_707),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_782),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_782),
.Y(n_869)
);

OAI21x1_ASAP7_75t_L g870 ( 
.A1(n_763),
.A2(n_652),
.B(n_591),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_807),
.B(n_652),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_847),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_775),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_783),
.Y(n_874)
);

CKINVDCx16_ASAP7_75t_R g875 ( 
.A(n_768),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_831),
.B(n_704),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_786),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_764),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_776),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_786),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_780),
.Y(n_881)
);

BUFx2_ASAP7_75t_L g882 ( 
.A(n_787),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_778),
.B(n_650),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_790),
.Y(n_884)
);

AOI22x1_ASAP7_75t_SL g885 ( 
.A1(n_779),
.A2(n_758),
.B1(n_554),
.B2(n_582),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_765),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_780),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_790),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_795),
.Y(n_889)
);

OA21x2_ASAP7_75t_L g890 ( 
.A1(n_762),
.A2(n_770),
.B(n_767),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_771),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_809),
.Y(n_892)
);

BUFx12f_ASAP7_75t_L g893 ( 
.A(n_774),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_787),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_762),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_776),
.B(n_704),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_800),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_798),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_800),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_823),
.Y(n_900)
);

NOR2x1_ASAP7_75t_L g901 ( 
.A(n_799),
.B(n_578),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_801),
.Y(n_902)
);

INVx4_ASAP7_75t_L g903 ( 
.A(n_776),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_776),
.B(n_586),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_776),
.Y(n_905)
);

BUFx2_ASAP7_75t_L g906 ( 
.A(n_823),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_803),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_802),
.Y(n_908)
);

INVx4_ASAP7_75t_L g909 ( 
.A(n_803),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_803),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_803),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_803),
.Y(n_912)
);

INVx5_ASAP7_75t_L g913 ( 
.A(n_780),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_832),
.B(n_557),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_822),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_822),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_828),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_766),
.B(n_594),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_773),
.B(n_663),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_828),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_838),
.Y(n_921)
);

INVx4_ASAP7_75t_L g922 ( 
.A(n_838),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_916),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_875),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_891),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_891),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_878),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_863),
.B(n_773),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_916),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_878),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_918),
.B(n_804),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_878),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_862),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_878),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_SL g935 ( 
.A1(n_875),
.A2(n_558),
.B1(n_593),
.B2(n_582),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_916),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_878),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_862),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_900),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_882),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_886),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_893),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_864),
.B(n_832),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_882),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_SL g945 ( 
.A1(n_883),
.A2(n_558),
.B1(n_608),
.B2(n_593),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_893),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_899),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_899),
.Y(n_948)
);

BUFx8_ASAP7_75t_L g949 ( 
.A(n_906),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_886),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_906),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_885),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_886),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_886),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_916),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_886),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_916),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_916),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_886),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_905),
.Y(n_960)
);

BUFx10_ASAP7_75t_L g961 ( 
.A(n_914),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_895),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_895),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_885),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_905),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_920),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_894),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_867),
.Y(n_968)
);

NOR2xp67_ASAP7_75t_L g969 ( 
.A(n_913),
.B(n_857),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_905),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_895),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_895),
.Y(n_972)
);

INVxp67_ASAP7_75t_L g973 ( 
.A(n_873),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_920),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_SL g975 ( 
.A1(n_864),
.A2(n_821),
.B1(n_813),
.B2(n_608),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_897),
.Y(n_976)
);

BUFx2_ASAP7_75t_L g977 ( 
.A(n_892),
.Y(n_977)
);

OAI21x1_ASAP7_75t_L g978 ( 
.A1(n_870),
.A2(n_599),
.B(n_598),
.Y(n_978)
);

CKINVDCx20_ASAP7_75t_R g979 ( 
.A(n_881),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_881),
.B(n_784),
.Y(n_980)
);

INVxp67_ASAP7_75t_L g981 ( 
.A(n_919),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_887),
.B(n_784),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_864),
.B(n_836),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_887),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_918),
.B(n_806),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_918),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_895),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_918),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_R g989 ( 
.A(n_876),
.B(n_836),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_895),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_896),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_871),
.B(n_857),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_863),
.B(n_919),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_896),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_920),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_871),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_871),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_871),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_889),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_896),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_913),
.B(n_818),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_889),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_896),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_904),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_904),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_904),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_904),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_862),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_991),
.Y(n_1009)
);

OR2x6_ASAP7_75t_L g1010 ( 
.A(n_948),
.B(n_846),
.Y(n_1010)
);

BUFx12f_ASAP7_75t_L g1011 ( 
.A(n_924),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_939),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_994),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_939),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_1000),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_SL g1016 ( 
.A(n_961),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_1003),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_999),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_931),
.Y(n_1019)
);

AO21x2_ASAP7_75t_L g1020 ( 
.A1(n_943),
.A2(n_637),
.B(n_625),
.Y(n_1020)
);

NAND3xp33_ASAP7_75t_L g1021 ( 
.A(n_983),
.B(n_854),
.C(n_812),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1002),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1004),
.Y(n_1023)
);

INVx4_ASAP7_75t_L g1024 ( 
.A(n_996),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_1005),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_996),
.B(n_890),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_1006),
.Y(n_1027)
);

BUFx4f_ASAP7_75t_L g1028 ( 
.A(n_984),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1007),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_997),
.B(n_998),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_993),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_931),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_985),
.Y(n_1033)
);

INVxp67_ASAP7_75t_SL g1034 ( 
.A(n_981),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_928),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_925),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_985),
.Y(n_1037)
);

NAND2xp33_ASAP7_75t_L g1038 ( 
.A(n_997),
.B(n_548),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_SL g1039 ( 
.A(n_961),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_926),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_989),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_998),
.B(n_992),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_968),
.B(n_788),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_924),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_1008),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_942),
.Y(n_1046)
);

INVx2_ASAP7_75t_SL g1047 ( 
.A(n_928),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_1008),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_985),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_980),
.B(n_818),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_986),
.B(n_808),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_933),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_969),
.B(n_962),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_963),
.B(n_890),
.Y(n_1054)
);

CKINVDCx6p67_ASAP7_75t_R g1055 ( 
.A(n_940),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_982),
.B(n_848),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_923),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_923),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_971),
.B(n_890),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_988),
.B(n_848),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_929),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_972),
.B(n_890),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_961),
.B(n_973),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_929),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_936),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_933),
.Y(n_1066)
);

OR2x6_ASAP7_75t_L g1067 ( 
.A(n_935),
.B(n_846),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_936),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_977),
.B(n_788),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_978),
.Y(n_1070)
);

NAND2xp33_ASAP7_75t_L g1071 ( 
.A(n_1001),
.B(n_556),
.Y(n_1071)
);

BUFx10_ASAP7_75t_L g1072 ( 
.A(n_942),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_978),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_955),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_975),
.B(n_796),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_947),
.A2(n_685),
.B1(n_737),
.B2(n_574),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_955),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_979),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_957),
.B(n_903),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_987),
.A2(n_737),
.B1(n_685),
.B2(n_990),
.Y(n_1080)
);

CKINVDCx20_ASAP7_75t_R g1081 ( 
.A(n_946),
.Y(n_1081)
);

OAI21xp33_ASAP7_75t_SL g1082 ( 
.A1(n_927),
.A2(n_845),
.B(n_805),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_957),
.Y(n_1083)
);

NAND2xp33_ASAP7_75t_SL g1084 ( 
.A(n_979),
.B(n_774),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_958),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_958),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_967),
.Y(n_1087)
);

INVxp33_ASAP7_75t_SL g1088 ( 
.A(n_946),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_966),
.B(n_903),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_967),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_940),
.Y(n_1091)
);

BUFx4f_ASAP7_75t_L g1092 ( 
.A(n_930),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_976),
.Y(n_1093)
);

CKINVDCx6p67_ASAP7_75t_R g1094 ( 
.A(n_944),
.Y(n_1094)
);

INVx6_ASAP7_75t_L g1095 ( 
.A(n_949),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_974),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_SL g1097 ( 
.A(n_949),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_995),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_995),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_933),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_938),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_938),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_1008),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_932),
.B(n_903),
.Y(n_1104)
);

BUFx8_ASAP7_75t_SL g1105 ( 
.A(n_944),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_934),
.B(n_950),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_945),
.A2(n_738),
.B1(n_741),
.B2(n_665),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_976),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_1008),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_1008),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_947),
.Y(n_1111)
);

OR2x6_ASAP7_75t_L g1112 ( 
.A(n_949),
.B(n_772),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_960),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_937),
.B(n_796),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_960),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_941),
.B(n_903),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_953),
.B(n_954),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_956),
.B(n_909),
.Y(n_1118)
);

INVx2_ASAP7_75t_SL g1119 ( 
.A(n_951),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_959),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_960),
.B(n_909),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_960),
.B(n_879),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_951),
.B(n_797),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_965),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_965),
.Y(n_1125)
);

AND2x6_ASAP7_75t_L g1126 ( 
.A(n_965),
.B(n_654),
.Y(n_1126)
);

BUFx4f_ASAP7_75t_L g1127 ( 
.A(n_965),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_970),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_SL g1129 ( 
.A1(n_952),
.A2(n_833),
.B1(n_779),
.B2(n_761),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_970),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_970),
.Y(n_1131)
);

NAND3xp33_ASAP7_75t_L g1132 ( 
.A(n_952),
.B(n_789),
.C(n_785),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_964),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_964),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_1050),
.B(n_1056),
.Y(n_1135)
);

OR2x2_ASAP7_75t_L g1136 ( 
.A(n_1076),
.B(n_852),
.Y(n_1136)
);

INVxp33_ASAP7_75t_L g1137 ( 
.A(n_1069),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1009),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1009),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1015),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_1042),
.B(n_913),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1034),
.B(n_922),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_1014),
.Y(n_1143)
);

NAND2xp33_ASAP7_75t_L g1144 ( 
.A(n_1026),
.B(n_579),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1017),
.Y(n_1145)
);

CKINVDCx20_ASAP7_75t_R g1146 ( 
.A(n_1081),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1054),
.A2(n_901),
.B(n_861),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_1049),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_1011),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_1042),
.B(n_913),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1031),
.B(n_922),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_1019),
.B(n_913),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1017),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_1050),
.B(n_797),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1043),
.B(n_769),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1025),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1025),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1013),
.B(n_922),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1023),
.B(n_879),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1029),
.B(n_1056),
.Y(n_1160)
);

NOR2xp67_ASAP7_75t_L g1161 ( 
.A(n_1041),
.B(n_777),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1027),
.B(n_909),
.Y(n_1162)
);

INVxp67_ASAP7_75t_L g1163 ( 
.A(n_1114),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_1123),
.B(n_761),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_1019),
.B(n_913),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_1060),
.B(n_769),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1060),
.B(n_671),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1035),
.B(n_671),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_1049),
.B(n_1035),
.Y(n_1169)
);

NOR3xp33_ASAP7_75t_L g1170 ( 
.A(n_1030),
.B(n_638),
.C(n_604),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1027),
.B(n_909),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1028),
.B(n_562),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_1091),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1047),
.B(n_859),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1036),
.Y(n_1175)
);

NAND2x1p5_ASAP7_75t_L g1176 ( 
.A(n_1045),
.B(n_905),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1057),
.Y(n_1177)
);

BUFx5_ASAP7_75t_L g1178 ( 
.A(n_1070),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1036),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_SL g1180 ( 
.A(n_1088),
.B(n_690),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1114),
.B(n_859),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_1063),
.B(n_690),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1040),
.B(n_861),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_1028),
.B(n_564),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1040),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1032),
.B(n_1033),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1024),
.B(n_564),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_SL g1188 ( 
.A(n_1072),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1058),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1037),
.B(n_865),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_SL g1191 ( 
.A(n_1046),
.B(n_700),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1020),
.B(n_865),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1020),
.B(n_872),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1059),
.B(n_872),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1120),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1063),
.B(n_700),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1030),
.A2(n_676),
.B1(n_677),
.B2(n_659),
.Y(n_1197)
);

INVxp67_ASAP7_75t_L g1198 ( 
.A(n_1051),
.Y(n_1198)
);

NOR2xp67_ASAP7_75t_L g1199 ( 
.A(n_1087),
.B(n_791),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1061),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1062),
.B(n_682),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1051),
.B(n_810),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1064),
.B(n_699),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1064),
.B(n_732),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_1018),
.B(n_1022),
.Y(n_1205)
);

NOR3xp33_ASAP7_75t_L g1206 ( 
.A(n_1021),
.B(n_722),
.C(n_672),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1065),
.B(n_734),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1080),
.B(n_758),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1065),
.B(n_749),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1068),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1068),
.B(n_752),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1075),
.B(n_842),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1074),
.B(n_757),
.Y(n_1213)
);

INVxp67_ASAP7_75t_L g1214 ( 
.A(n_1010),
.Y(n_1214)
);

NOR2xp67_ASAP7_75t_L g1215 ( 
.A(n_1093),
.B(n_792),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1119),
.B(n_842),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1010),
.B(n_853),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_1127),
.B(n_1090),
.Y(n_1218)
);

INVx2_ASAP7_75t_SL g1219 ( 
.A(n_1010),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1083),
.B(n_1085),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1067),
.B(n_853),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_1127),
.B(n_603),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1079),
.A2(n_862),
.B(n_912),
.Y(n_1223)
);

NOR3xp33_ASAP7_75t_L g1224 ( 
.A(n_1132),
.B(n_794),
.C(n_793),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1083),
.Y(n_1225)
);

NOR3xp33_ASAP7_75t_L g1226 ( 
.A(n_1111),
.B(n_1133),
.C(n_1129),
.Y(n_1226)
);

NAND2xp33_ASAP7_75t_L g1227 ( 
.A(n_1045),
.B(n_609),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_SL g1228 ( 
.A(n_1072),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1086),
.B(n_860),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1086),
.B(n_860),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1096),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1108),
.B(n_576),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_1044),
.B(n_580),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1096),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1098),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1100),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1077),
.B(n_866),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1099),
.B(n_866),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1100),
.Y(n_1239)
);

OAI21xp33_ASAP7_75t_L g1240 ( 
.A1(n_1107),
.A2(n_569),
.B(n_568),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_1082),
.B(n_610),
.Y(n_1241)
);

NAND2xp33_ASAP7_75t_SL g1242 ( 
.A(n_1016),
.B(n_614),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1092),
.B(n_620),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1067),
.B(n_583),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1102),
.B(n_868),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1102),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1113),
.B(n_868),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1012),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1106),
.Y(n_1249)
);

AND2x4_ASAP7_75t_L g1250 ( 
.A(n_1112),
.B(n_811),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1113),
.B(n_869),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1124),
.B(n_869),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1124),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1078),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1052),
.Y(n_1255)
);

OR2x2_ASAP7_75t_L g1256 ( 
.A(n_1067),
.B(n_814),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1115),
.B(n_623),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1101),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1107),
.B(n_602),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1038),
.B(n_585),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1066),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1125),
.B(n_874),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1016),
.B(n_587),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1117),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1110),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1117),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1115),
.B(n_642),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1110),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1128),
.B(n_877),
.Y(n_1269)
);

NAND3xp33_ASAP7_75t_L g1270 ( 
.A(n_1071),
.B(n_589),
.C(n_588),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1130),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1131),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1045),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1122),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1079),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1115),
.B(n_1048),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1048),
.B(n_1103),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1048),
.B(n_877),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1048),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1103),
.B(n_880),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1103),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1103),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_1105),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1109),
.B(n_1115),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1039),
.B(n_592),
.Y(n_1285)
);

BUFx8_ASAP7_75t_L g1286 ( 
.A(n_1097),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1089),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1109),
.B(n_880),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1109),
.B(n_888),
.Y(n_1289)
);

INVxp67_ASAP7_75t_L g1290 ( 
.A(n_1078),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1104),
.Y(n_1291)
);

NOR3xp33_ASAP7_75t_L g1292 ( 
.A(n_1084),
.B(n_1134),
.C(n_816),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1073),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1104),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1053),
.B(n_888),
.Y(n_1295)
);

OR2x2_ASAP7_75t_L g1296 ( 
.A(n_1055),
.B(n_815),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1116),
.B(n_920),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1116),
.B(n_653),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1118),
.B(n_920),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1118),
.B(n_920),
.Y(n_1300)
);

INVxp67_ASAP7_75t_L g1301 ( 
.A(n_1126),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1121),
.B(n_905),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1121),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1126),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1126),
.B(n_905),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1112),
.B(n_656),
.Y(n_1306)
);

INVx2_ASAP7_75t_SL g1307 ( 
.A(n_1094),
.Y(n_1307)
);

OR2x2_ASAP7_75t_SL g1308 ( 
.A(n_1136),
.B(n_1095),
.Y(n_1308)
);

NAND3xp33_ASAP7_75t_SL g1309 ( 
.A(n_1135),
.B(n_569),
.C(n_568),
.Y(n_1309)
);

OAI221xp5_ASAP7_75t_L g1310 ( 
.A1(n_1135),
.A2(n_1112),
.B1(n_736),
.B2(n_740),
.C(n_651),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1140),
.Y(n_1311)
);

INVx4_ASAP7_75t_L g1312 ( 
.A(n_1148),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1138),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1139),
.Y(n_1314)
);

OAI221xp5_ASAP7_75t_L g1315 ( 
.A1(n_1154),
.A2(n_736),
.B1(n_740),
.B2(n_651),
.C(n_570),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1200),
.Y(n_1316)
);

NAND2x1p5_ASAP7_75t_L g1317 ( 
.A(n_1148),
.B(n_907),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1145),
.Y(n_1318)
);

INVxp67_ASAP7_75t_L g1319 ( 
.A(n_1155),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1154),
.A2(n_695),
.B1(n_696),
.B2(n_657),
.Y(n_1320)
);

NAND2x1p5_ASAP7_75t_L g1321 ( 
.A(n_1148),
.B(n_1169),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1156),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1212),
.B(n_1095),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1169),
.B(n_817),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_SL g1325 ( 
.A(n_1160),
.B(n_698),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1157),
.Y(n_1326)
);

OAI221xp5_ASAP7_75t_L g1327 ( 
.A1(n_1167),
.A2(n_744),
.B1(n_745),
.B2(n_743),
.C(n_570),
.Y(n_1327)
);

OR2x2_ASAP7_75t_SL g1328 ( 
.A(n_1256),
.B(n_1095),
.Y(n_1328)
);

AOI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1212),
.A2(n_706),
.B1(n_711),
.B2(n_703),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1153),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_1283),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1175),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1198),
.B(n_819),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1179),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1185),
.Y(n_1335)
);

NAND2x1p5_ASAP7_75t_L g1336 ( 
.A(n_1273),
.B(n_907),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_1254),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1166),
.B(n_1216),
.Y(n_1338)
);

NAND2x1_ASAP7_75t_L g1339 ( 
.A(n_1273),
.B(n_1126),
.Y(n_1339)
);

OR2x6_ASAP7_75t_L g1340 ( 
.A(n_1248),
.B(n_1097),
.Y(n_1340)
);

AO22x2_ASAP7_75t_L g1341 ( 
.A1(n_1259),
.A2(n_1170),
.B1(n_1226),
.B2(n_1206),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1166),
.B(n_602),
.Y(n_1342)
);

CKINVDCx14_ASAP7_75t_R g1343 ( 
.A(n_1146),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1186),
.Y(n_1344)
);

OAI221xp5_ASAP7_75t_L g1345 ( 
.A1(n_1167),
.A2(n_745),
.B1(n_759),
.B2(n_744),
.C(n_743),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1210),
.Y(n_1346)
);

OAI221xp5_ASAP7_75t_L g1347 ( 
.A1(n_1208),
.A2(n_759),
.B1(n_597),
.B2(n_600),
.C(n_596),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1177),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1163),
.B(n_1249),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1225),
.Y(n_1350)
);

AO22x2_ASAP7_75t_L g1351 ( 
.A1(n_1170),
.A2(n_1226),
.B1(n_1206),
.B2(n_1163),
.Y(n_1351)
);

INVxp67_ASAP7_75t_L g1352 ( 
.A(n_1205),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1231),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1234),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1189),
.Y(n_1355)
);

AO22x2_ASAP7_75t_L g1356 ( 
.A1(n_1214),
.A2(n_741),
.B1(n_751),
.B2(n_746),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1219),
.B(n_820),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1202),
.B(n_824),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1182),
.B(n_595),
.Y(n_1359)
);

AND2x6_ASAP7_75t_L g1360 ( 
.A(n_1304),
.B(n_754),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1195),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1237),
.Y(n_1362)
);

INVx3_ASAP7_75t_L g1363 ( 
.A(n_1273),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_1143),
.Y(n_1364)
);

BUFx8_ASAP7_75t_L g1365 ( 
.A(n_1188),
.Y(n_1365)
);

INVxp67_ASAP7_75t_L g1366 ( 
.A(n_1205),
.Y(n_1366)
);

OR2x2_ASAP7_75t_SL g1367 ( 
.A(n_1296),
.B(n_755),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1142),
.B(n_1126),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1238),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1202),
.B(n_825),
.Y(n_1370)
);

AO22x2_ASAP7_75t_L g1371 ( 
.A1(n_1214),
.A2(n_756),
.B1(n_827),
.B2(n_826),
.Y(n_1371)
);

BUFx3_ASAP7_75t_L g1372 ( 
.A(n_1173),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_1254),
.Y(n_1373)
);

INVxp67_ASAP7_75t_L g1374 ( 
.A(n_1217),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1239),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1246),
.Y(n_1376)
);

OR2x6_ASAP7_75t_L g1377 ( 
.A(n_1149),
.B(n_829),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1235),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1245),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1262),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_1188),
.Y(n_1381)
);

NAND2x1p5_ASAP7_75t_L g1382 ( 
.A(n_1218),
.B(n_907),
.Y(n_1382)
);

AO22x2_ASAP7_75t_L g1383 ( 
.A1(n_1208),
.A2(n_834),
.B1(n_835),
.B2(n_830),
.Y(n_1383)
);

OAI221xp5_ASAP7_75t_L g1384 ( 
.A1(n_1196),
.A2(n_615),
.B1(n_617),
.B2(n_607),
.C(n_601),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1228),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1269),
.Y(n_1386)
);

NAND2x1p5_ASAP7_75t_L g1387 ( 
.A(n_1307),
.B(n_907),
.Y(n_1387)
);

AOI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1260),
.A2(n_724),
.B1(n_728),
.B2(n_716),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1229),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1230),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1247),
.Y(n_1391)
);

INVx3_ASAP7_75t_L g1392 ( 
.A(n_1253),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1251),
.Y(n_1393)
);

OAI221xp5_ASAP7_75t_L g1394 ( 
.A1(n_1196),
.A2(n_622),
.B1(n_629),
.B2(n_619),
.C(n_618),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1274),
.B(n_915),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1228),
.Y(n_1396)
);

XOR2xp5_ASAP7_75t_L g1397 ( 
.A(n_1137),
.B(n_385),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1252),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1236),
.Y(n_1399)
);

AO22x2_ASAP7_75t_L g1400 ( 
.A1(n_1290),
.A2(n_840),
.B1(n_841),
.B2(n_839),
.Y(n_1400)
);

AO22x2_ASAP7_75t_L g1401 ( 
.A1(n_1306),
.A2(n_849),
.B1(n_850),
.B2(n_843),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1174),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1190),
.Y(n_1403)
);

OAI221xp5_ASAP7_75t_L g1404 ( 
.A1(n_1168),
.A2(n_634),
.B1(n_635),
.B2(n_632),
.C(n_630),
.Y(n_1404)
);

INVx2_ASAP7_75t_SL g1405 ( 
.A(n_1250),
.Y(n_1405)
);

AOI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1260),
.A2(n_728),
.B1(n_716),
.B2(n_898),
.Y(n_1406)
);

CKINVDCx20_ASAP7_75t_R g1407 ( 
.A(n_1286),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1258),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1293),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_1286),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1271),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1272),
.Y(n_1412)
);

OAI221xp5_ASAP7_75t_L g1413 ( 
.A1(n_1168),
.A2(n_641),
.B1(n_643),
.B2(n_640),
.C(n_636),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1264),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1266),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1261),
.Y(n_1416)
);

AO22x2_ASAP7_75t_L g1417 ( 
.A1(n_1303),
.A2(n_858),
.B1(n_851),
.B2(n_750),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1183),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1220),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1221),
.B(n_644),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1250),
.B(n_855),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_SL g1422 ( 
.A(n_1191),
.Y(n_1422)
);

BUFx8_ASAP7_75t_L g1423 ( 
.A(n_1255),
.Y(n_1423)
);

AO22x2_ASAP7_75t_L g1424 ( 
.A1(n_1291),
.A2(n_750),
.B1(n_644),
.B2(n_855),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1203),
.Y(n_1425)
);

INVxp67_ASAP7_75t_L g1426 ( 
.A(n_1217),
.Y(n_1426)
);

BUFx2_ASAP7_75t_L g1427 ( 
.A(n_1279),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1204),
.Y(n_1428)
);

NAND2x1p5_ASAP7_75t_L g1429 ( 
.A(n_1281),
.B(n_907),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1207),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1265),
.Y(n_1431)
);

INVxp67_ASAP7_75t_L g1432 ( 
.A(n_1232),
.Y(n_1432)
);

INVxp67_ASAP7_75t_L g1433 ( 
.A(n_1233),
.Y(n_1433)
);

XOR2xp5_ASAP7_75t_L g1434 ( 
.A(n_1270),
.B(n_386),
.Y(n_1434)
);

OAI221xp5_ASAP7_75t_L g1435 ( 
.A1(n_1244),
.A2(n_648),
.B1(n_661),
.B2(n_658),
.C(n_647),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1268),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1209),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_1164),
.B(n_662),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1211),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1221),
.B(n_856),
.Y(n_1440)
);

NAND3xp33_ASAP7_75t_SL g1441 ( 
.A(n_1180),
.B(n_666),
.C(n_664),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1213),
.Y(n_1442)
);

AO22x2_ASAP7_75t_L g1443 ( 
.A1(n_1294),
.A2(n_644),
.B1(n_750),
.B2(n_856),
.Y(n_1443)
);

NAND2xp33_ASAP7_75t_L g1444 ( 
.A(n_1178),
.B(n_760),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1181),
.B(n_915),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1159),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1151),
.B(n_917),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1278),
.Y(n_1448)
);

AO22x2_ASAP7_75t_L g1449 ( 
.A1(n_1275),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_1449)
);

OAI221xp5_ASAP7_75t_L g1450 ( 
.A1(n_1244),
.A2(n_673),
.B1(n_674),
.B2(n_670),
.C(n_668),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1280),
.Y(n_1451)
);

OAI221xp5_ASAP7_75t_L g1452 ( 
.A1(n_1240),
.A2(n_681),
.B1(n_686),
.B2(n_679),
.C(n_678),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1288),
.Y(n_1453)
);

NAND2x1p5_ASAP7_75t_L g1454 ( 
.A(n_1282),
.B(n_910),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1287),
.Y(n_1455)
);

AO22x2_ASAP7_75t_L g1456 ( 
.A1(n_1241),
.A2(n_7),
.B1(n_4),
.B2(n_6),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1289),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1295),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1158),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1276),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_SL g1461 ( 
.A(n_1292),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1199),
.B(n_921),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1178),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1178),
.Y(n_1464)
);

AND2x4_ASAP7_75t_L g1465 ( 
.A(n_1215),
.B(n_1161),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1172),
.B(n_687),
.Y(n_1466)
);

OAI22xp33_ASAP7_75t_SL g1467 ( 
.A1(n_1187),
.A2(n_692),
.B1(n_693),
.B2(n_688),
.Y(n_1467)
);

AND2x4_ASAP7_75t_L g1468 ( 
.A(n_1301),
.B(n_921),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_SL g1469 ( 
.A(n_1197),
.B(n_716),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1194),
.B(n_898),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1162),
.Y(n_1471)
);

CKINVDCx16_ASAP7_75t_R g1472 ( 
.A(n_1242),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1201),
.B(n_902),
.Y(n_1473)
);

OAI221xp5_ASAP7_75t_L g1474 ( 
.A1(n_1224),
.A2(n_701),
.B1(n_702),
.B2(n_697),
.C(n_694),
.Y(n_1474)
);

CKINVDCx20_ASAP7_75t_R g1475 ( 
.A(n_1184),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1178),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1144),
.B(n_908),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_1284),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1192),
.Y(n_1479)
);

AO22x2_ASAP7_75t_L g1480 ( 
.A1(n_1141),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_1480)
);

OAI221xp5_ASAP7_75t_L g1481 ( 
.A1(n_1224),
.A2(n_717),
.B1(n_721),
.B2(n_709),
.C(n_705),
.Y(n_1481)
);

AO22x2_ASAP7_75t_L g1482 ( 
.A1(n_1150),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1193),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1277),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1178),
.Y(n_1485)
);

OR2x6_ASAP7_75t_L g1486 ( 
.A(n_1263),
.B(n_910),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1298),
.A2(n_728),
.B1(n_884),
.B2(n_725),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1171),
.A2(n_726),
.B1(n_727),
.B2(n_723),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1459),
.A2(n_1147),
.B(n_1297),
.Y(n_1489)
);

O2A1O1Ixp33_ASAP7_75t_L g1490 ( 
.A1(n_1359),
.A2(n_1292),
.B(n_1263),
.C(n_1285),
.Y(n_1490)
);

O2A1O1Ixp5_ASAP7_75t_L g1491 ( 
.A1(n_1438),
.A2(n_1222),
.B(n_1267),
.C(n_1257),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1458),
.B(n_1243),
.Y(n_1492)
);

AOI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1444),
.A2(n_1300),
.B(n_1299),
.Y(n_1493)
);

AOI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1338),
.A2(n_1227),
.B1(n_1165),
.B2(n_1152),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1368),
.A2(n_1302),
.B(n_1223),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1344),
.A2(n_1352),
.B1(n_1366),
.B2(n_1349),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1316),
.Y(n_1497)
);

INVxp67_ASAP7_75t_L g1498 ( 
.A(n_1337),
.Y(n_1498)
);

CKINVDCx20_ASAP7_75t_R g1499 ( 
.A(n_1364),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1342),
.B(n_729),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_SL g1501 ( 
.A(n_1432),
.B(n_1305),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1362),
.A2(n_1176),
.B1(n_733),
.B2(n_735),
.Y(n_1502)
);

NOR3xp33_ASAP7_75t_L g1503 ( 
.A(n_1347),
.B(n_747),
.C(n_731),
.Y(n_1503)
);

INVx1_ASAP7_75t_SL g1504 ( 
.A(n_1372),
.Y(n_1504)
);

AOI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1471),
.A2(n_1447),
.B(n_1473),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1369),
.A2(n_753),
.B1(n_748),
.B2(n_910),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1433),
.B(n_1374),
.Y(n_1507)
);

O2A1O1Ixp33_ASAP7_75t_L g1508 ( 
.A1(n_1327),
.A2(n_884),
.B(n_13),
.C(n_10),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1380),
.A2(n_910),
.B1(n_912),
.B2(n_911),
.Y(n_1509)
);

AO21x1_ASAP7_75t_L g1510 ( 
.A1(n_1479),
.A2(n_12),
.B(n_13),
.Y(n_1510)
);

AOI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1483),
.A2(n_912),
.B(n_911),
.Y(n_1511)
);

O2A1O1Ixp5_ASAP7_75t_L g1512 ( 
.A1(n_1325),
.A2(n_15),
.B(n_12),
.C(n_14),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1386),
.B(n_911),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1426),
.B(n_16),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1402),
.B(n_911),
.Y(n_1515)
);

AOI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1323),
.A2(n_912),
.B1(n_862),
.B2(n_18),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1420),
.B(n_16),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1405),
.B(n_542),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1361),
.Y(n_1519)
);

OA22x2_ASAP7_75t_L g1520 ( 
.A1(n_1388),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1389),
.B(n_17),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1471),
.A2(n_389),
.B(n_388),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_SL g1523 ( 
.A(n_1465),
.B(n_20),
.Y(n_1523)
);

O2A1O1Ixp33_ASAP7_75t_L g1524 ( 
.A1(n_1345),
.A2(n_22),
.B(n_20),
.C(n_21),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_1465),
.B(n_21),
.Y(n_1525)
);

AOI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1425),
.A2(n_392),
.B(n_391),
.Y(n_1526)
);

AOI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1428),
.A2(n_394),
.B(n_393),
.Y(n_1527)
);

BUFx12f_ASAP7_75t_L g1528 ( 
.A(n_1410),
.Y(n_1528)
);

AOI21x1_ASAP7_75t_L g1529 ( 
.A1(n_1470),
.A2(n_541),
.B(n_396),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1319),
.B(n_22),
.Y(n_1530)
);

AOI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1430),
.A2(n_398),
.B(n_395),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_L g1532 ( 
.A(n_1312),
.Y(n_1532)
);

OAI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1437),
.A2(n_400),
.B(n_399),
.Y(n_1533)
);

O2A1O1Ixp33_ASAP7_75t_L g1534 ( 
.A1(n_1309),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_1534)
);

AOI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1341),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_1535)
);

OAI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1439),
.A2(n_540),
.B(n_402),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1390),
.B(n_26),
.Y(n_1537)
);

OAI22x1_ASAP7_75t_L g1538 ( 
.A1(n_1406),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_SL g1539 ( 
.A(n_1422),
.B(n_28),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1441),
.B(n_29),
.Y(n_1540)
);

AO21x1_ASAP7_75t_L g1541 ( 
.A1(n_1445),
.A2(n_29),
.B(n_30),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1379),
.B(n_31),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1442),
.A2(n_403),
.B(n_401),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1419),
.B(n_31),
.Y(n_1544)
);

OAI21xp5_ASAP7_75t_L g1545 ( 
.A1(n_1446),
.A2(n_539),
.B(n_405),
.Y(n_1545)
);

OAI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1448),
.A2(n_406),
.B(n_404),
.Y(n_1546)
);

AOI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1477),
.A2(n_408),
.B(n_407),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1391),
.B(n_32),
.Y(n_1548)
);

INVx11_ASAP7_75t_L g1549 ( 
.A(n_1423),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1393),
.B(n_32),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1398),
.B(n_33),
.Y(n_1551)
);

INVx3_ASAP7_75t_L g1552 ( 
.A(n_1312),
.Y(n_1552)
);

OAI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1418),
.A2(n_411),
.B(n_409),
.Y(n_1553)
);

INVxp67_ASAP7_75t_L g1554 ( 
.A(n_1373),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1451),
.B(n_33),
.Y(n_1555)
);

OAI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1453),
.A2(n_413),
.B(n_412),
.Y(n_1556)
);

NOR2x1p5_ASAP7_75t_SL g1557 ( 
.A(n_1463),
.B(n_419),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1457),
.A2(n_422),
.B(n_420),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1403),
.B(n_34),
.Y(n_1559)
);

AO21x1_ASAP7_75t_L g1560 ( 
.A1(n_1484),
.A2(n_34),
.B(n_36),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1341),
.B(n_37),
.Y(n_1561)
);

AOI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1475),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_1562)
);

BUFx3_ASAP7_75t_L g1563 ( 
.A(n_1423),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1409),
.Y(n_1564)
);

OAI21xp33_ASAP7_75t_L g1565 ( 
.A1(n_1466),
.A2(n_39),
.B(n_40),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1414),
.B(n_40),
.Y(n_1566)
);

BUFx2_ASAP7_75t_L g1567 ( 
.A(n_1324),
.Y(n_1567)
);

OAI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1395),
.A2(n_538),
.B(n_425),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1464),
.A2(n_426),
.B(n_424),
.Y(n_1569)
);

A2O1A1Ixp33_ASAP7_75t_L g1570 ( 
.A1(n_1384),
.A2(n_1394),
.B(n_1310),
.C(n_1415),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1351),
.B(n_41),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1351),
.B(n_41),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1411),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1440),
.B(n_1478),
.Y(n_1574)
);

INVx1_ASAP7_75t_SL g1575 ( 
.A(n_1324),
.Y(n_1575)
);

AOI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1476),
.A2(n_429),
.B(n_427),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1455),
.B(n_42),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1346),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_L g1579 ( 
.A(n_1321),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1383),
.B(n_43),
.Y(n_1580)
);

OAI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1460),
.A2(n_432),
.B(n_431),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1422),
.B(n_44),
.Y(n_1582)
);

NOR2xp67_ASAP7_75t_L g1583 ( 
.A(n_1331),
.B(n_537),
.Y(n_1583)
);

AOI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1485),
.A2(n_434),
.B(n_433),
.Y(n_1584)
);

AOI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1486),
.A2(n_437),
.B(n_435),
.Y(n_1585)
);

BUFx12f_ASAP7_75t_L g1586 ( 
.A(n_1365),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1350),
.Y(n_1587)
);

AOI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1486),
.A2(n_439),
.B(n_438),
.Y(n_1588)
);

AOI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1461),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1353),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1412),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1435),
.B(n_49),
.Y(n_1592)
);

NOR2xp67_ASAP7_75t_L g1593 ( 
.A(n_1416),
.B(n_443),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_L g1594 ( 
.A(n_1450),
.B(n_50),
.Y(n_1594)
);

INVx3_ASAP7_75t_L g1595 ( 
.A(n_1339),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1333),
.B(n_51),
.Y(n_1596)
);

AO21x1_ASAP7_75t_L g1597 ( 
.A1(n_1469),
.A2(n_52),
.B(n_53),
.Y(n_1597)
);

INVx1_ASAP7_75t_SL g1598 ( 
.A(n_1427),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1333),
.B(n_52),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1308),
.B(n_55),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1358),
.Y(n_1601)
);

O2A1O1Ixp5_ASAP7_75t_L g1602 ( 
.A1(n_1313),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_1602)
);

INVxp67_ASAP7_75t_L g1603 ( 
.A(n_1358),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1408),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_1604)
);

AOI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1314),
.A2(n_1322),
.B(n_1318),
.Y(n_1605)
);

NOR2x1_ASAP7_75t_L g1606 ( 
.A(n_1363),
.B(n_447),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1326),
.A2(n_450),
.B(n_449),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1328),
.Y(n_1608)
);

A2O1A1Ixp33_ASAP7_75t_L g1609 ( 
.A1(n_1315),
.A2(n_62),
.B(n_58),
.C(n_60),
.Y(n_1609)
);

A2O1A1Ixp33_ASAP7_75t_L g1610 ( 
.A1(n_1320),
.A2(n_64),
.B(n_62),
.C(n_63),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1383),
.B(n_65),
.Y(n_1611)
);

O2A1O1Ixp5_ASAP7_75t_L g1612 ( 
.A1(n_1332),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_1612)
);

INVxp67_ASAP7_75t_L g1613 ( 
.A(n_1370),
.Y(n_1613)
);

OAI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1334),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_1614)
);

INVx11_ASAP7_75t_L g1615 ( 
.A(n_1365),
.Y(n_1615)
);

AOI21x1_ASAP7_75t_L g1616 ( 
.A1(n_1375),
.A2(n_536),
.B(n_452),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_SL g1617 ( 
.A(n_1467),
.B(n_1472),
.Y(n_1617)
);

NAND3xp33_ASAP7_75t_L g1618 ( 
.A(n_1404),
.B(n_69),
.C(n_70),
.Y(n_1618)
);

AOI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1335),
.A2(n_453),
.B(n_451),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1413),
.B(n_69),
.Y(n_1620)
);

BUFx4f_ASAP7_75t_L g1621 ( 
.A(n_1340),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1354),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1376),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1401),
.B(n_71),
.Y(n_1624)
);

AOI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1461),
.A2(n_75),
.B1(n_72),
.B2(n_74),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1367),
.B(n_76),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1462),
.B(n_76),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1462),
.B(n_77),
.Y(n_1628)
);

OAI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1330),
.A2(n_456),
.B(n_455),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1370),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1311),
.B(n_77),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1378),
.A2(n_1392),
.B1(n_1431),
.B2(n_1329),
.Y(n_1632)
);

OAI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1468),
.A2(n_458),
.B(n_457),
.Y(n_1633)
);

NOR2xp67_ASAP7_75t_L g1634 ( 
.A(n_1436),
.B(n_535),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1357),
.B(n_78),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1348),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1468),
.B(n_79),
.Y(n_1637)
);

AOI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1397),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_1638)
);

INVx1_ASAP7_75t_SL g1639 ( 
.A(n_1421),
.Y(n_1639)
);

INVx1_ASAP7_75t_SL g1640 ( 
.A(n_1421),
.Y(n_1640)
);

OAI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1436),
.A2(n_84),
.B1(n_81),
.B2(n_82),
.Y(n_1641)
);

AOI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1343),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1642)
);

AOI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1434),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1474),
.B(n_1481),
.Y(n_1644)
);

NAND2x1_ASAP7_75t_L g1645 ( 
.A(n_1363),
.B(n_460),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1355),
.B(n_88),
.Y(n_1646)
);

OAI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1399),
.A2(n_464),
.B(n_463),
.Y(n_1647)
);

A2O1A1Ixp33_ASAP7_75t_L g1648 ( 
.A1(n_1487),
.A2(n_92),
.B(n_89),
.C(n_90),
.Y(n_1648)
);

AOI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1317),
.A2(n_469),
.B(n_467),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1400),
.B(n_1488),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1452),
.B(n_1382),
.Y(n_1651)
);

INVx3_ASAP7_75t_L g1652 ( 
.A(n_1336),
.Y(n_1652)
);

O2A1O1Ixp33_ASAP7_75t_L g1653 ( 
.A1(n_1490),
.A2(n_1377),
.B(n_1340),
.C(n_1387),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1519),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_SL g1655 ( 
.A(n_1496),
.B(n_1381),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1574),
.B(n_1400),
.Y(n_1656)
);

AOI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1644),
.A2(n_1377),
.B1(n_1396),
.B2(n_1385),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1507),
.B(n_1407),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1505),
.A2(n_1449),
.B(n_1480),
.Y(n_1659)
);

BUFx3_ASAP7_75t_L g1660 ( 
.A(n_1499),
.Y(n_1660)
);

INVx4_ASAP7_75t_L g1661 ( 
.A(n_1532),
.Y(n_1661)
);

O2A1O1Ixp5_ASAP7_75t_L g1662 ( 
.A1(n_1651),
.A2(n_1482),
.B(n_1480),
.C(n_1456),
.Y(n_1662)
);

OAI21xp33_ASAP7_75t_L g1663 ( 
.A1(n_1592),
.A2(n_1443),
.B(n_1424),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1492),
.B(n_1417),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1639),
.B(n_1417),
.Y(n_1665)
);

INVxp67_ASAP7_75t_L g1666 ( 
.A(n_1601),
.Y(n_1666)
);

AND2x4_ASAP7_75t_SL g1667 ( 
.A(n_1579),
.B(n_1360),
.Y(n_1667)
);

CKINVDCx11_ASAP7_75t_R g1668 ( 
.A(n_1586),
.Y(n_1668)
);

INVx5_ASAP7_75t_L g1669 ( 
.A(n_1532),
.Y(n_1669)
);

INVx3_ASAP7_75t_L g1670 ( 
.A(n_1532),
.Y(n_1670)
);

BUFx8_ASAP7_75t_L g1671 ( 
.A(n_1528),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1489),
.A2(n_1449),
.B(n_1482),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1640),
.B(n_1371),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1640),
.B(n_1356),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1500),
.B(n_1356),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1575),
.B(n_1424),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1575),
.B(n_1443),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1530),
.B(n_1360),
.Y(n_1678)
);

O2A1O1Ixp33_ASAP7_75t_L g1679 ( 
.A1(n_1594),
.A2(n_1429),
.B(n_1454),
.C(n_1360),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_SL g1680 ( 
.A(n_1621),
.B(n_473),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1497),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1630),
.B(n_92),
.Y(n_1682)
);

OAI21xp33_ASAP7_75t_L g1683 ( 
.A1(n_1620),
.A2(n_93),
.B(n_94),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1564),
.Y(n_1684)
);

AOI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1493),
.A2(n_534),
.B(n_475),
.Y(n_1685)
);

INVx4_ASAP7_75t_L g1686 ( 
.A(n_1549),
.Y(n_1686)
);

BUFx12f_ASAP7_75t_L g1687 ( 
.A(n_1567),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1495),
.A2(n_478),
.B(n_474),
.Y(n_1688)
);

O2A1O1Ixp33_ASAP7_75t_L g1689 ( 
.A1(n_1570),
.A2(n_97),
.B(n_94),
.C(n_96),
.Y(n_1689)
);

BUFx8_ASAP7_75t_L g1690 ( 
.A(n_1608),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1603),
.B(n_96),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1503),
.B(n_97),
.Y(n_1692)
);

BUFx4f_ASAP7_75t_L g1693 ( 
.A(n_1579),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_R g1694 ( 
.A(n_1621),
.B(n_479),
.Y(n_1694)
);

BUFx6f_ASAP7_75t_L g1695 ( 
.A(n_1579),
.Y(n_1695)
);

CKINVDCx10_ASAP7_75t_R g1696 ( 
.A(n_1615),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1578),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_SL g1698 ( 
.A(n_1517),
.B(n_98),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1565),
.A2(n_1540),
.B1(n_1618),
.B2(n_1520),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1587),
.Y(n_1700)
);

AOI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1617),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_1701)
);

BUFx12f_ASAP7_75t_L g1702 ( 
.A(n_1600),
.Y(n_1702)
);

INVxp67_ASAP7_75t_L g1703 ( 
.A(n_1504),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1590),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1623),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1613),
.B(n_99),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1521),
.B(n_100),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1598),
.B(n_101),
.Y(n_1708)
);

BUFx6f_ASAP7_75t_L g1709 ( 
.A(n_1563),
.Y(n_1709)
);

BUFx6f_ASAP7_75t_L g1710 ( 
.A(n_1552),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1537),
.B(n_102),
.Y(n_1711)
);

AOI21xp5_ASAP7_75t_L g1712 ( 
.A1(n_1491),
.A2(n_531),
.B(n_483),
.Y(n_1712)
);

AOI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1568),
.A2(n_530),
.B(n_485),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_SL g1714 ( 
.A1(n_1539),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_SL g1715 ( 
.A(n_1598),
.B(n_103),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1504),
.B(n_480),
.Y(n_1716)
);

AOI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1546),
.A2(n_1556),
.B(n_1647),
.Y(n_1717)
);

AOI21x1_ASAP7_75t_L g1718 ( 
.A1(n_1511),
.A2(n_488),
.B(n_486),
.Y(n_1718)
);

OAI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1554),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1542),
.B(n_107),
.Y(n_1720)
);

BUFx6f_ASAP7_75t_L g1721 ( 
.A(n_1552),
.Y(n_1721)
);

O2A1O1Ixp33_ASAP7_75t_L g1722 ( 
.A1(n_1609),
.A2(n_109),
.B(n_107),
.C(n_108),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1636),
.Y(n_1723)
);

OAI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1650),
.A2(n_111),
.B1(n_108),
.B2(n_110),
.Y(n_1724)
);

O2A1O1Ixp33_ASAP7_75t_SL g1725 ( 
.A1(n_1610),
.A2(n_112),
.B(n_110),
.C(n_111),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1548),
.B(n_112),
.Y(n_1726)
);

OAI21x1_ASAP7_75t_L g1727 ( 
.A1(n_1529),
.A2(n_490),
.B(n_489),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1523),
.B(n_491),
.Y(n_1728)
);

O2A1O1Ixp5_ASAP7_75t_SL g1729 ( 
.A1(n_1501),
.A2(n_115),
.B(n_113),
.C(n_114),
.Y(n_1729)
);

BUFx2_ASAP7_75t_L g1730 ( 
.A(n_1498),
.Y(n_1730)
);

AO21x1_ASAP7_75t_L g1731 ( 
.A1(n_1561),
.A2(n_113),
.B(n_114),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1525),
.B(n_492),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1631),
.Y(n_1733)
);

AOI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1629),
.A2(n_497),
.B(n_495),
.Y(n_1734)
);

AND2x2_ASAP7_75t_SL g1735 ( 
.A(n_1539),
.B(n_115),
.Y(n_1735)
);

AOI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1581),
.A2(n_527),
.B(n_500),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1550),
.B(n_116),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1646),
.Y(n_1738)
);

BUFx6f_ASAP7_75t_L g1739 ( 
.A(n_1518),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1533),
.A2(n_526),
.B(n_502),
.Y(n_1740)
);

AOI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1533),
.A2(n_525),
.B(n_503),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1643),
.A2(n_119),
.B1(n_116),
.B2(n_118),
.Y(n_1742)
);

A2O1A1Ixp33_ASAP7_75t_L g1743 ( 
.A1(n_1508),
.A2(n_1524),
.B(n_1633),
.C(n_1536),
.Y(n_1743)
);

NOR2xp33_ASAP7_75t_L g1744 ( 
.A(n_1627),
.B(n_498),
.Y(n_1744)
);

BUFx6f_ASAP7_75t_L g1745 ( 
.A(n_1518),
.Y(n_1745)
);

AOI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1536),
.A2(n_505),
.B(n_504),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1551),
.B(n_118),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1515),
.Y(n_1748)
);

INVx1_ASAP7_75t_SL g1749 ( 
.A(n_1596),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_SL g1750 ( 
.A(n_1544),
.B(n_120),
.Y(n_1750)
);

INVx6_ASAP7_75t_L g1751 ( 
.A(n_1580),
.Y(n_1751)
);

AOI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1553),
.A2(n_1545),
.B(n_1513),
.Y(n_1752)
);

OAI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1494),
.A2(n_120),
.B(n_121),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1577),
.Y(n_1754)
);

OAI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1516),
.A2(n_121),
.B(n_122),
.Y(n_1755)
);

INVx3_ASAP7_75t_L g1756 ( 
.A(n_1595),
.Y(n_1756)
);

AOI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1553),
.A2(n_507),
.B(n_506),
.Y(n_1757)
);

OAI21x1_ASAP7_75t_L g1758 ( 
.A1(n_1616),
.A2(n_510),
.B(n_508),
.Y(n_1758)
);

BUFx4f_ASAP7_75t_L g1759 ( 
.A(n_1652),
.Y(n_1759)
);

AOI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1545),
.A2(n_516),
.B(n_514),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1566),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1520),
.A2(n_1572),
.B1(n_1571),
.B2(n_1538),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1555),
.B(n_123),
.Y(n_1763)
);

INVx5_ASAP7_75t_L g1764 ( 
.A(n_1595),
.Y(n_1764)
);

OAI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1559),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1605),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1637),
.B(n_124),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1652),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1632),
.Y(n_1769)
);

O2A1O1Ixp33_ASAP7_75t_L g1770 ( 
.A1(n_1648),
.A2(n_127),
.B(n_125),
.C(n_126),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_L g1771 ( 
.A(n_1628),
.B(n_517),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1514),
.B(n_128),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1645),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1510),
.Y(n_1774)
);

AOI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1626),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1599),
.B(n_130),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1522),
.A2(n_524),
.B(n_519),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1635),
.B(n_518),
.Y(n_1778)
);

OAI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1535),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.Y(n_1779)
);

OAI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1638),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_SL g1781 ( 
.A(n_1582),
.B(n_1593),
.Y(n_1781)
);

AOI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1589),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1512),
.Y(n_1783)
);

BUFx6f_ASAP7_75t_L g1784 ( 
.A(n_1624),
.Y(n_1784)
);

O2A1O1Ixp33_ASAP7_75t_L g1785 ( 
.A1(n_1611),
.A2(n_140),
.B(n_138),
.C(n_139),
.Y(n_1785)
);

A2O1A1Ixp33_ASAP7_75t_L g1786 ( 
.A1(n_1534),
.A2(n_142),
.B(n_140),
.C(n_141),
.Y(n_1786)
);

INVx4_ASAP7_75t_L g1787 ( 
.A(n_1557),
.Y(n_1787)
);

OAI22xp33_ASAP7_75t_L g1788 ( 
.A1(n_1625),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.Y(n_1788)
);

BUFx2_ASAP7_75t_L g1789 ( 
.A(n_1606),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1502),
.B(n_143),
.Y(n_1790)
);

O2A1O1Ixp33_ASAP7_75t_L g1791 ( 
.A1(n_1573),
.A2(n_147),
.B(n_145),
.C(n_146),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_L g1792 ( 
.A(n_1642),
.B(n_146),
.Y(n_1792)
);

AOI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1547),
.A2(n_384),
.B(n_147),
.Y(n_1793)
);

OAI221xp5_ASAP7_75t_L g1794 ( 
.A1(n_1562),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.C(n_151),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1506),
.B(n_148),
.Y(n_1795)
);

AOI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1558),
.A2(n_149),
.B(n_150),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_1591),
.Y(n_1797)
);

AOI21x1_ASAP7_75t_L g1798 ( 
.A1(n_1718),
.A2(n_1541),
.B(n_1509),
.Y(n_1798)
);

BUFx2_ASAP7_75t_L g1799 ( 
.A(n_1687),
.Y(n_1799)
);

BUFx6f_ASAP7_75t_L g1800 ( 
.A(n_1669),
.Y(n_1800)
);

BUFx3_ASAP7_75t_L g1801 ( 
.A(n_1660),
.Y(n_1801)
);

BUFx12f_ASAP7_75t_L g1802 ( 
.A(n_1668),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1769),
.B(n_1560),
.Y(n_1803)
);

OAI21x1_ASAP7_75t_L g1804 ( 
.A1(n_1688),
.A2(n_1576),
.B(n_1569),
.Y(n_1804)
);

OA21x2_ASAP7_75t_L g1805 ( 
.A1(n_1752),
.A2(n_1612),
.B(n_1602),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1717),
.A2(n_1588),
.B(n_1585),
.Y(n_1806)
);

OAI21x1_ASAP7_75t_L g1807 ( 
.A1(n_1758),
.A2(n_1584),
.B(n_1527),
.Y(n_1807)
);

CKINVDCx14_ASAP7_75t_R g1808 ( 
.A(n_1686),
.Y(n_1808)
);

OAI21x1_ASAP7_75t_L g1809 ( 
.A1(n_1712),
.A2(n_1727),
.B(n_1685),
.Y(n_1809)
);

NOR2x1_ASAP7_75t_L g1810 ( 
.A(n_1781),
.B(n_1583),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1749),
.B(n_1597),
.Y(n_1811)
);

AND2x4_ASAP7_75t_L g1812 ( 
.A(n_1739),
.B(n_1634),
.Y(n_1812)
);

INVx2_ASAP7_75t_SL g1813 ( 
.A(n_1693),
.Y(n_1813)
);

OAI21x1_ASAP7_75t_L g1814 ( 
.A1(n_1766),
.A2(n_1531),
.B(n_1526),
.Y(n_1814)
);

AO31x2_ASAP7_75t_L g1815 ( 
.A1(n_1672),
.A2(n_1607),
.A3(n_1619),
.B(n_1543),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1654),
.Y(n_1816)
);

AO22x2_ASAP7_75t_L g1817 ( 
.A1(n_1659),
.A2(n_1604),
.B1(n_1622),
.B2(n_1614),
.Y(n_1817)
);

OAI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1743),
.A2(n_1649),
.B(n_1641),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1684),
.Y(n_1819)
);

OAI21x1_ASAP7_75t_SL g1820 ( 
.A1(n_1731),
.A2(n_1653),
.B(n_1753),
.Y(n_1820)
);

OAI21xp5_ASAP7_75t_L g1821 ( 
.A1(n_1713),
.A2(n_151),
.B(n_152),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1784),
.B(n_152),
.Y(n_1822)
);

AOI221xp5_ASAP7_75t_SL g1823 ( 
.A1(n_1788),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.C(n_158),
.Y(n_1823)
);

NOR4xp25_ASAP7_75t_L g1824 ( 
.A(n_1689),
.B(n_157),
.C(n_155),
.D(n_156),
.Y(n_1824)
);

OAI21x1_ASAP7_75t_L g1825 ( 
.A1(n_1777),
.A2(n_158),
.B(n_159),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_SL g1826 ( 
.A(n_1738),
.B(n_160),
.Y(n_1826)
);

AOI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1734),
.A2(n_161),
.B(n_162),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1784),
.B(n_161),
.Y(n_1828)
);

AOI21x1_ASAP7_75t_L g1829 ( 
.A1(n_1740),
.A2(n_163),
.B(n_165),
.Y(n_1829)
);

AOI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1736),
.A2(n_165),
.B(n_166),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1784),
.B(n_168),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1739),
.B(n_168),
.Y(n_1832)
);

BUFx3_ASAP7_75t_L g1833 ( 
.A(n_1730),
.Y(n_1833)
);

AOI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1741),
.A2(n_169),
.B(n_171),
.Y(n_1834)
);

AOI21xp5_ASAP7_75t_L g1835 ( 
.A1(n_1746),
.A2(n_171),
.B(n_172),
.Y(n_1835)
);

AOI21x1_ASAP7_75t_L g1836 ( 
.A1(n_1757),
.A2(n_1760),
.B(n_1774),
.Y(n_1836)
);

INVx1_ASAP7_75t_SL g1837 ( 
.A(n_1673),
.Y(n_1837)
);

AOI221x1_ASAP7_75t_L g1838 ( 
.A1(n_1663),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.C(n_176),
.Y(n_1838)
);

NAND3x1_ASAP7_75t_L g1839 ( 
.A(n_1792),
.B(n_176),
.C(n_177),
.Y(n_1839)
);

OA21x2_ASAP7_75t_L g1840 ( 
.A1(n_1662),
.A2(n_1796),
.B(n_1793),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1761),
.B(n_177),
.Y(n_1841)
);

OAI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1782),
.A2(n_180),
.B1(n_178),
.B2(n_179),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1723),
.Y(n_1843)
);

BUFx6f_ASAP7_75t_L g1844 ( 
.A(n_1669),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1697),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1700),
.Y(n_1846)
);

NOR2x1_ASAP7_75t_SL g1847 ( 
.A(n_1764),
.B(n_181),
.Y(n_1847)
);

OAI21x1_ASAP7_75t_SL g1848 ( 
.A1(n_1722),
.A2(n_181),
.B(n_182),
.Y(n_1848)
);

BUFx2_ASAP7_75t_L g1849 ( 
.A(n_1703),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1674),
.Y(n_1850)
);

NAND3x1_ASAP7_75t_L g1851 ( 
.A(n_1657),
.B(n_182),
.C(n_183),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1678),
.B(n_184),
.Y(n_1852)
);

A2O1A1Ixp33_ASAP7_75t_L g1853 ( 
.A1(n_1755),
.A2(n_187),
.B(n_185),
.C(n_186),
.Y(n_1853)
);

AND2x4_ASAP7_75t_L g1854 ( 
.A(n_1739),
.B(n_186),
.Y(n_1854)
);

O2A1O1Ixp5_ASAP7_75t_L g1855 ( 
.A1(n_1692),
.A2(n_187),
.B(n_188),
.C(n_189),
.Y(n_1855)
);

OA21x2_ASAP7_75t_L g1856 ( 
.A1(n_1783),
.A2(n_190),
.B(n_191),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_1789),
.B(n_192),
.Y(n_1857)
);

AOI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1764),
.A2(n_192),
.B(n_193),
.Y(n_1858)
);

CKINVDCx11_ASAP7_75t_R g1859 ( 
.A(n_1686),
.Y(n_1859)
);

INVx4_ASAP7_75t_L g1860 ( 
.A(n_1669),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1764),
.A2(n_193),
.B(n_194),
.Y(n_1861)
);

NOR2xp33_ASAP7_75t_R g1862 ( 
.A(n_1696),
.B(n_195),
.Y(n_1862)
);

AOI221x1_ASAP7_75t_L g1863 ( 
.A1(n_1683),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.C(n_199),
.Y(n_1863)
);

AOI21xp5_ASAP7_75t_L g1864 ( 
.A1(n_1679),
.A2(n_197),
.B(n_199),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1699),
.B(n_200),
.Y(n_1865)
);

AOI21xp5_ASAP7_75t_L g1866 ( 
.A1(n_1680),
.A2(n_1748),
.B(n_1725),
.Y(n_1866)
);

OAI21x1_ASAP7_75t_L g1867 ( 
.A1(n_1756),
.A2(n_200),
.B(n_201),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1754),
.B(n_201),
.Y(n_1868)
);

AOI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1742),
.A2(n_202),
.B1(n_203),
.B2(n_205),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1704),
.Y(n_1870)
);

OAI21x1_ASAP7_75t_L g1871 ( 
.A1(n_1756),
.A2(n_206),
.B(n_207),
.Y(n_1871)
);

A2O1A1Ixp33_ASAP7_75t_L g1872 ( 
.A1(n_1770),
.A2(n_206),
.B(n_207),
.C(n_208),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1705),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1733),
.B(n_1762),
.Y(n_1874)
);

OAI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1735),
.A2(n_1794),
.B1(n_1797),
.B2(n_1714),
.Y(n_1875)
);

OAI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1786),
.A2(n_208),
.B(n_209),
.Y(n_1876)
);

NAND2x1p5_ASAP7_75t_L g1877 ( 
.A(n_1787),
.B(n_209),
.Y(n_1877)
);

AOI21xp5_ASAP7_75t_L g1878 ( 
.A1(n_1773),
.A2(n_210),
.B(n_211),
.Y(n_1878)
);

OA21x2_ASAP7_75t_L g1879 ( 
.A1(n_1664),
.A2(n_210),
.B(n_211),
.Y(n_1879)
);

OAI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1795),
.A2(n_212),
.B(n_213),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1656),
.B(n_213),
.Y(n_1881)
);

OAI22xp33_ASAP7_75t_L g1882 ( 
.A1(n_1775),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1681),
.B(n_214),
.Y(n_1883)
);

AOI21x1_ASAP7_75t_L g1884 ( 
.A1(n_1665),
.A2(n_215),
.B(n_217),
.Y(n_1884)
);

OAI21x1_ASAP7_75t_L g1885 ( 
.A1(n_1729),
.A2(n_217),
.B(n_218),
.Y(n_1885)
);

O2A1O1Ixp33_ASAP7_75t_SL g1886 ( 
.A1(n_1790),
.A2(n_218),
.B(n_219),
.C(n_220),
.Y(n_1886)
);

AOI221x1_ASAP7_75t_L g1887 ( 
.A1(n_1724),
.A2(n_219),
.B1(n_221),
.B2(n_222),
.C(n_223),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_1859),
.Y(n_1888)
);

AO21x2_ASAP7_75t_L g1889 ( 
.A1(n_1806),
.A2(n_1836),
.B(n_1821),
.Y(n_1889)
);

BUFx3_ASAP7_75t_L g1890 ( 
.A(n_1800),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1837),
.B(n_1676),
.Y(n_1891)
);

CKINVDCx6p67_ASAP7_75t_R g1892 ( 
.A(n_1802),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1816),
.Y(n_1893)
);

OA21x2_ASAP7_75t_L g1894 ( 
.A1(n_1809),
.A2(n_1677),
.B(n_1675),
.Y(n_1894)
);

OA21x2_ASAP7_75t_L g1895 ( 
.A1(n_1814),
.A2(n_1711),
.B(n_1707),
.Y(n_1895)
);

HB1xp67_ASAP7_75t_L g1896 ( 
.A(n_1850),
.Y(n_1896)
);

AOI21x1_ASAP7_75t_L g1897 ( 
.A1(n_1798),
.A2(n_1655),
.B(n_1750),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1845),
.Y(n_1898)
);

OAI21x1_ASAP7_75t_L g1899 ( 
.A1(n_1807),
.A2(n_1785),
.B(n_1791),
.Y(n_1899)
);

OA21x2_ASAP7_75t_L g1900 ( 
.A1(n_1803),
.A2(n_1726),
.B(n_1720),
.Y(n_1900)
);

OAI21x1_ASAP7_75t_L g1901 ( 
.A1(n_1804),
.A2(n_1747),
.B(n_1737),
.Y(n_1901)
);

HB1xp67_ASAP7_75t_L g1902 ( 
.A(n_1837),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1801),
.B(n_1658),
.Y(n_1903)
);

NAND2x1p5_ASAP7_75t_L g1904 ( 
.A(n_1856),
.B(n_1787),
.Y(n_1904)
);

OAI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1834),
.A2(n_1744),
.B(n_1779),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1846),
.B(n_1751),
.Y(n_1906)
);

AOI21x1_ASAP7_75t_L g1907 ( 
.A1(n_1829),
.A2(n_1763),
.B(n_1765),
.Y(n_1907)
);

A2O1A1Ixp33_ASAP7_75t_L g1908 ( 
.A1(n_1821),
.A2(n_1701),
.B(n_1732),
.C(n_1728),
.Y(n_1908)
);

OAI21xp5_ASAP7_75t_L g1909 ( 
.A1(n_1835),
.A2(n_1778),
.B(n_1771),
.Y(n_1909)
);

OR2x2_ASAP7_75t_L g1910 ( 
.A(n_1870),
.B(n_1776),
.Y(n_1910)
);

NAND2x1_ASAP7_75t_L g1911 ( 
.A(n_1856),
.B(n_1710),
.Y(n_1911)
);

OAI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1827),
.A2(n_1780),
.B(n_1772),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1873),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1803),
.Y(n_1914)
);

AOI22xp33_ASAP7_75t_L g1915 ( 
.A1(n_1875),
.A2(n_1751),
.B1(n_1702),
.B2(n_1698),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1811),
.B(n_1831),
.Y(n_1916)
);

OAI21x1_ASAP7_75t_L g1917 ( 
.A1(n_1825),
.A2(n_1768),
.B(n_1767),
.Y(n_1917)
);

OAI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1875),
.A2(n_1745),
.B1(n_1716),
.B2(n_1759),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1874),
.B(n_1666),
.Y(n_1919)
);

NAND2x1p5_ASAP7_75t_L g1920 ( 
.A(n_1840),
.B(n_1745),
.Y(n_1920)
);

O2A1O1Ixp33_ASAP7_75t_L g1921 ( 
.A1(n_1853),
.A2(n_1719),
.B(n_1708),
.C(n_1715),
.Y(n_1921)
);

AND2x4_ASAP7_75t_L g1922 ( 
.A(n_1819),
.B(n_1695),
.Y(n_1922)
);

BUFx2_ASAP7_75t_L g1923 ( 
.A(n_1833),
.Y(n_1923)
);

OAI22xp33_ASAP7_75t_L g1924 ( 
.A1(n_1869),
.A2(n_1745),
.B1(n_1682),
.B2(n_1691),
.Y(n_1924)
);

BUFx3_ASAP7_75t_L g1925 ( 
.A(n_1800),
.Y(n_1925)
);

OAI21x1_ASAP7_75t_L g1926 ( 
.A1(n_1805),
.A2(n_1670),
.B(n_1706),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1849),
.B(n_1716),
.Y(n_1927)
);

NAND2x1p5_ASAP7_75t_L g1928 ( 
.A(n_1840),
.B(n_1661),
.Y(n_1928)
);

HB1xp67_ASAP7_75t_L g1929 ( 
.A(n_1843),
.Y(n_1929)
);

AOI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1818),
.A2(n_1667),
.B(n_1710),
.Y(n_1930)
);

BUFx12f_ASAP7_75t_L g1931 ( 
.A(n_1813),
.Y(n_1931)
);

AO21x2_ASAP7_75t_L g1932 ( 
.A1(n_1820),
.A2(n_1694),
.B(n_1710),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1881),
.B(n_1695),
.Y(n_1933)
);

INVx4_ASAP7_75t_L g1934 ( 
.A(n_1800),
.Y(n_1934)
);

BUFx3_ASAP7_75t_L g1935 ( 
.A(n_1844),
.Y(n_1935)
);

AO21x2_ASAP7_75t_L g1936 ( 
.A1(n_1818),
.A2(n_1721),
.B(n_1695),
.Y(n_1936)
);

OA21x2_ASAP7_75t_L g1937 ( 
.A1(n_1864),
.A2(n_221),
.B(n_223),
.Y(n_1937)
);

HB1xp67_ASAP7_75t_L g1938 ( 
.A(n_1902),
.Y(n_1938)
);

AOI21x1_ASAP7_75t_L g1939 ( 
.A1(n_1897),
.A2(n_1911),
.B(n_1884),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_1888),
.Y(n_1940)
);

AOI22xp33_ASAP7_75t_SL g1941 ( 
.A1(n_1909),
.A2(n_1876),
.B1(n_1880),
.B2(n_1865),
.Y(n_1941)
);

INVx8_ASAP7_75t_L g1942 ( 
.A(n_1931),
.Y(n_1942)
);

HB1xp67_ASAP7_75t_L g1943 ( 
.A(n_1896),
.Y(n_1943)
);

INVx1_ASAP7_75t_SL g1944 ( 
.A(n_1923),
.Y(n_1944)
);

AO21x1_ASAP7_75t_SL g1945 ( 
.A1(n_1914),
.A2(n_1876),
.B(n_1880),
.Y(n_1945)
);

BUFx6f_ASAP7_75t_L g1946 ( 
.A(n_1890),
.Y(n_1946)
);

CKINVDCx16_ASAP7_75t_R g1947 ( 
.A(n_1916),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1891),
.B(n_1881),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1893),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_1888),
.Y(n_1950)
);

AND2x4_ASAP7_75t_L g1951 ( 
.A(n_1893),
.B(n_1815),
.Y(n_1951)
);

BUFx10_ASAP7_75t_L g1952 ( 
.A(n_1922),
.Y(n_1952)
);

BUFx6f_ASAP7_75t_L g1953 ( 
.A(n_1890),
.Y(n_1953)
);

HB1xp67_ASAP7_75t_L g1954 ( 
.A(n_1929),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1913),
.Y(n_1955)
);

BUFx2_ASAP7_75t_L g1956 ( 
.A(n_1894),
.Y(n_1956)
);

HB1xp67_ASAP7_75t_L g1957 ( 
.A(n_1894),
.Y(n_1957)
);

AOI22xp5_ASAP7_75t_SL g1958 ( 
.A1(n_1900),
.A2(n_1879),
.B1(n_1865),
.B2(n_1839),
.Y(n_1958)
);

INVx6_ASAP7_75t_L g1959 ( 
.A(n_1934),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1898),
.Y(n_1960)
);

HB1xp67_ASAP7_75t_L g1961 ( 
.A(n_1894),
.Y(n_1961)
);

NAND2x1p5_ASAP7_75t_L g1962 ( 
.A(n_1911),
.B(n_1879),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1900),
.B(n_1822),
.Y(n_1963)
);

HB1xp67_ASAP7_75t_L g1964 ( 
.A(n_1936),
.Y(n_1964)
);

AOI22xp33_ASAP7_75t_L g1965 ( 
.A1(n_1905),
.A2(n_1882),
.B1(n_1842),
.B2(n_1830),
.Y(n_1965)
);

INVx11_ASAP7_75t_L g1966 ( 
.A(n_1931),
.Y(n_1966)
);

AOI22xp33_ASAP7_75t_SL g1967 ( 
.A1(n_1912),
.A2(n_1848),
.B1(n_1817),
.B2(n_1847),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1900),
.B(n_1822),
.Y(n_1968)
);

INVx1_ASAP7_75t_SL g1969 ( 
.A(n_1923),
.Y(n_1969)
);

OAI22xp5_ASAP7_75t_L g1970 ( 
.A1(n_1941),
.A2(n_1908),
.B1(n_1851),
.B2(n_1869),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1949),
.Y(n_1971)
);

AOI22xp33_ASAP7_75t_SL g1972 ( 
.A1(n_1958),
.A2(n_1918),
.B1(n_1937),
.B2(n_1889),
.Y(n_1972)
);

BUFx3_ASAP7_75t_L g1973 ( 
.A(n_1946),
.Y(n_1973)
);

AOI22xp33_ASAP7_75t_SL g1974 ( 
.A1(n_1958),
.A2(n_1937),
.B1(n_1889),
.B2(n_1817),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1938),
.B(n_1914),
.Y(n_1975)
);

AOI22xp33_ASAP7_75t_L g1976 ( 
.A1(n_1945),
.A2(n_1924),
.B1(n_1889),
.B2(n_1895),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1949),
.Y(n_1977)
);

OR2x2_ASAP7_75t_L g1978 ( 
.A(n_1963),
.B(n_1910),
.Y(n_1978)
);

AOI22xp33_ASAP7_75t_SL g1979 ( 
.A1(n_1947),
.A2(n_1937),
.B1(n_1932),
.B2(n_1877),
.Y(n_1979)
);

CKINVDCx11_ASAP7_75t_R g1980 ( 
.A(n_1942),
.Y(n_1980)
);

OAI22xp33_ASAP7_75t_L g1981 ( 
.A1(n_1947),
.A2(n_1887),
.B1(n_1838),
.B2(n_1863),
.Y(n_1981)
);

AOI22xp33_ASAP7_75t_L g1982 ( 
.A1(n_1945),
.A2(n_1895),
.B1(n_1932),
.B2(n_1915),
.Y(n_1982)
);

INVx3_ASAP7_75t_L g1983 ( 
.A(n_1952),
.Y(n_1983)
);

OAI22xp5_ASAP7_75t_L g1984 ( 
.A1(n_1965),
.A2(n_1872),
.B1(n_1810),
.B2(n_1877),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1944),
.B(n_1916),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1955),
.Y(n_1986)
);

CKINVDCx5p33_ASAP7_75t_R g1987 ( 
.A(n_1940),
.Y(n_1987)
);

AOI22xp33_ASAP7_75t_SL g1988 ( 
.A1(n_1942),
.A2(n_1932),
.B1(n_1899),
.B2(n_1895),
.Y(n_1988)
);

OAI21xp5_ASAP7_75t_SL g1989 ( 
.A1(n_1967),
.A2(n_1921),
.B(n_1878),
.Y(n_1989)
);

BUFx12f_ASAP7_75t_L g1990 ( 
.A(n_1940),
.Y(n_1990)
);

NOR2xp33_ASAP7_75t_L g1991 ( 
.A(n_1990),
.B(n_1950),
.Y(n_1991)
);

INVxp67_ASAP7_75t_L g1992 ( 
.A(n_1985),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1971),
.Y(n_1993)
);

NOR2xp33_ASAP7_75t_R g1994 ( 
.A(n_1987),
.B(n_1950),
.Y(n_1994)
);

NAND2xp33_ASAP7_75t_R g1995 ( 
.A(n_1987),
.B(n_1862),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_1990),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1986),
.Y(n_1997)
);

AND2x4_ASAP7_75t_L g1998 ( 
.A(n_1973),
.B(n_1951),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1985),
.B(n_1969),
.Y(n_1999)
);

AND2x4_ASAP7_75t_L g2000 ( 
.A(n_1973),
.B(n_1951),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1993),
.Y(n_2001)
);

HB1xp67_ASAP7_75t_L g2002 ( 
.A(n_1997),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1992),
.Y(n_2003)
);

OR2x2_ASAP7_75t_L g2004 ( 
.A(n_1999),
.B(n_1978),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1997),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1999),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_2002),
.Y(n_2007)
);

HB1xp67_ASAP7_75t_L g2008 ( 
.A(n_2002),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_2006),
.B(n_1998),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_2001),
.Y(n_2010)
);

OR2x2_ASAP7_75t_L g2011 ( 
.A(n_2004),
.B(n_1978),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_2005),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_2003),
.B(n_1998),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_2001),
.Y(n_2014)
);

HB1xp67_ASAP7_75t_L g2015 ( 
.A(n_2002),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_SL g2016 ( 
.A(n_2003),
.B(n_1994),
.Y(n_2016)
);

AND2x4_ASAP7_75t_L g2017 ( 
.A(n_2016),
.B(n_1996),
.Y(n_2017)
);

AND2x4_ASAP7_75t_L g2018 ( 
.A(n_2016),
.B(n_1996),
.Y(n_2018)
);

NOR2xp67_ASAP7_75t_L g2019 ( 
.A(n_2008),
.B(n_1991),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_2008),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_2013),
.B(n_1892),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_2010),
.B(n_1943),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_2014),
.B(n_2007),
.Y(n_2023)
);

INVxp67_ASAP7_75t_L g2024 ( 
.A(n_2015),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_2015),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_2009),
.B(n_1892),
.Y(n_2026)
);

OR2x2_ASAP7_75t_L g2027 ( 
.A(n_2011),
.B(n_1968),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_2026),
.Y(n_2028)
);

NAND3xp33_ASAP7_75t_SL g2029 ( 
.A(n_2024),
.B(n_1989),
.C(n_1970),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_2021),
.B(n_2007),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_2020),
.B(n_2012),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_2025),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_2017),
.B(n_2000),
.Y(n_2033)
);

AND2x4_ASAP7_75t_L g2034 ( 
.A(n_2019),
.B(n_1998),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_2023),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_2023),
.B(n_1977),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_2032),
.B(n_2017),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_2034),
.Y(n_2038)
);

NOR2x1_ASAP7_75t_SL g2039 ( 
.A(n_2029),
.B(n_2022),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_2033),
.B(n_2018),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_2040),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_2037),
.Y(n_2042)
);

OAI21xp5_ASAP7_75t_L g2043 ( 
.A1(n_2037),
.A2(n_2018),
.B(n_2035),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_2038),
.B(n_2030),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_2044),
.Y(n_2045)
);

AOI22xp33_ASAP7_75t_L g2046 ( 
.A1(n_2041),
.A2(n_2028),
.B1(n_2034),
.B2(n_2031),
.Y(n_2046)
);

OAI21xp5_ASAP7_75t_SL g2047 ( 
.A1(n_2043),
.A2(n_2031),
.B(n_2039),
.Y(n_2047)
);

INVxp67_ASAP7_75t_SL g2048 ( 
.A(n_2043),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_2042),
.Y(n_2049)
);

AOI21xp5_ASAP7_75t_L g2050 ( 
.A1(n_2043),
.A2(n_2036),
.B(n_2022),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_2045),
.B(n_2036),
.Y(n_2051)
);

OR2x2_ASAP7_75t_L g2052 ( 
.A(n_2048),
.B(n_2027),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_2049),
.Y(n_2053)
);

OAI32xp33_ASAP7_75t_L g2054 ( 
.A1(n_2046),
.A2(n_1995),
.A3(n_1984),
.B1(n_1857),
.B2(n_1903),
.Y(n_2054)
);

AOI21xp5_ASAP7_75t_L g2055 ( 
.A1(n_2048),
.A2(n_1808),
.B(n_1942),
.Y(n_2055)
);

OR2x2_ASAP7_75t_L g2056 ( 
.A(n_2047),
.B(n_1975),
.Y(n_2056)
);

NAND3xp33_ASAP7_75t_L g2057 ( 
.A(n_2050),
.B(n_1671),
.C(n_1823),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_2045),
.B(n_1709),
.Y(n_2058)
);

NAND3xp33_ASAP7_75t_SL g2059 ( 
.A(n_2047),
.B(n_1799),
.C(n_1972),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_2048),
.B(n_2000),
.Y(n_2060)
);

OAI22xp5_ASAP7_75t_L g2061 ( 
.A1(n_2052),
.A2(n_1966),
.B1(n_1979),
.B2(n_1974),
.Y(n_2061)
);

OR2x2_ASAP7_75t_L g2062 ( 
.A(n_2060),
.B(n_1948),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2051),
.Y(n_2063)
);

INVxp67_ASAP7_75t_L g2064 ( 
.A(n_2058),
.Y(n_2064)
);

OAI22xp5_ASAP7_75t_L g2065 ( 
.A1(n_2056),
.A2(n_1966),
.B1(n_1982),
.B2(n_1942),
.Y(n_2065)
);

AOI21xp5_ASAP7_75t_L g2066 ( 
.A1(n_2055),
.A2(n_1942),
.B(n_1886),
.Y(n_2066)
);

NOR2xp33_ASAP7_75t_L g2067 ( 
.A(n_2053),
.B(n_1671),
.Y(n_2067)
);

OAI22xp33_ASAP7_75t_L g2068 ( 
.A1(n_2057),
.A2(n_1709),
.B1(n_1953),
.B2(n_1946),
.Y(n_2068)
);

NOR2xp33_ASAP7_75t_L g2069 ( 
.A(n_2054),
.B(n_1709),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2059),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2060),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_2058),
.B(n_2000),
.Y(n_2072)
);

AOI22xp5_ASAP7_75t_L g2073 ( 
.A1(n_2059),
.A2(n_1980),
.B1(n_1690),
.B2(n_1823),
.Y(n_2073)
);

NOR3xp33_ASAP7_75t_L g2074 ( 
.A(n_2067),
.B(n_1980),
.C(n_1841),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2063),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_2071),
.B(n_1690),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_2064),
.B(n_1983),
.Y(n_2077)
);

NOR2xp33_ASAP7_75t_L g2078 ( 
.A(n_2070),
.B(n_1841),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2069),
.B(n_1906),
.Y(n_2079)
);

AOI211xp5_ASAP7_75t_L g2080 ( 
.A1(n_2068),
.A2(n_1824),
.B(n_1861),
.C(n_1858),
.Y(n_2080)
);

NOR2xp33_ASAP7_75t_L g2081 ( 
.A(n_2062),
.B(n_1868),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2072),
.Y(n_2082)
);

AOI21xp33_ASAP7_75t_L g2083 ( 
.A1(n_2065),
.A2(n_1828),
.B(n_1868),
.Y(n_2083)
);

AOI221xp5_ASAP7_75t_L g2084 ( 
.A1(n_2061),
.A2(n_1824),
.B1(n_1981),
.B2(n_1976),
.C(n_1855),
.Y(n_2084)
);

NOR2xp33_ASAP7_75t_L g2085 ( 
.A(n_2066),
.B(n_1828),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_SL g2086 ( 
.A(n_2073),
.B(n_1844),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_2063),
.B(n_1906),
.Y(n_2087)
);

AOI21xp5_ASAP7_75t_L g2088 ( 
.A1(n_2067),
.A2(n_1826),
.B(n_1852),
.Y(n_2088)
);

OAI211xp5_ASAP7_75t_SL g2089 ( 
.A1(n_2082),
.A2(n_1883),
.B(n_1919),
.C(n_1988),
.Y(n_2089)
);

OAI221xp5_ASAP7_75t_SL g2090 ( 
.A1(n_2075),
.A2(n_2076),
.B1(n_2077),
.B2(n_2074),
.C(n_2079),
.Y(n_2090)
);

O2A1O1Ixp33_ASAP7_75t_L g2091 ( 
.A1(n_2078),
.A2(n_1883),
.B(n_227),
.C(n_224),
.Y(n_2091)
);

O2A1O1Ixp33_ASAP7_75t_L g2092 ( 
.A1(n_2086),
.A2(n_228),
.B(n_225),
.C(n_227),
.Y(n_2092)
);

AOI211xp5_ASAP7_75t_L g2093 ( 
.A1(n_2085),
.A2(n_1854),
.B(n_1832),
.C(n_1844),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_2081),
.B(n_1910),
.Y(n_2094)
);

NOR2xp33_ASAP7_75t_L g2095 ( 
.A(n_2087),
.B(n_225),
.Y(n_2095)
);

NAND2xp33_ASAP7_75t_SL g2096 ( 
.A(n_2083),
.B(n_1661),
.Y(n_2096)
);

NAND3xp33_ASAP7_75t_L g2097 ( 
.A(n_2080),
.B(n_1854),
.C(n_1832),
.Y(n_2097)
);

OAI22xp5_ASAP7_75t_L g2098 ( 
.A1(n_2084),
.A2(n_1959),
.B1(n_1983),
.B2(n_1953),
.Y(n_2098)
);

OAI21xp5_ASAP7_75t_L g2099 ( 
.A1(n_2088),
.A2(n_1901),
.B(n_1871),
.Y(n_2099)
);

A2O1A1Ixp33_ASAP7_75t_L g2100 ( 
.A1(n_2078),
.A2(n_1901),
.B(n_1867),
.C(n_1983),
.Y(n_2100)
);

AND5x1_ASAP7_75t_L g2101 ( 
.A(n_2078),
.B(n_1930),
.C(n_1866),
.D(n_231),
.E(n_232),
.Y(n_2101)
);

AOI22xp5_ASAP7_75t_L g2102 ( 
.A1(n_2074),
.A2(n_1959),
.B1(n_1953),
.B2(n_1946),
.Y(n_2102)
);

NAND3xp33_ASAP7_75t_L g2103 ( 
.A(n_2092),
.B(n_1860),
.C(n_228),
.Y(n_2103)
);

AOI211xp5_ASAP7_75t_L g2104 ( 
.A1(n_2090),
.A2(n_235),
.B(n_229),
.C(n_234),
.Y(n_2104)
);

AOI221x1_ASAP7_75t_SL g2105 ( 
.A1(n_2095),
.A2(n_1933),
.B1(n_1927),
.B2(n_235),
.C(n_236),
.Y(n_2105)
);

OAI21xp33_ASAP7_75t_SL g2106 ( 
.A1(n_2102),
.A2(n_1934),
.B(n_1860),
.Y(n_2106)
);

OAI21xp5_ASAP7_75t_SL g2107 ( 
.A1(n_2091),
.A2(n_1962),
.B(n_1907),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_2094),
.B(n_229),
.Y(n_2108)
);

NOR2xp67_ASAP7_75t_L g2109 ( 
.A(n_2097),
.B(n_234),
.Y(n_2109)
);

AOI21xp5_ASAP7_75t_L g2110 ( 
.A1(n_2096),
.A2(n_1917),
.B(n_236),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_2093),
.B(n_237),
.Y(n_2111)
);

NAND4xp75_ASAP7_75t_L g2112 ( 
.A(n_2099),
.B(n_239),
.C(n_237),
.D(n_238),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2098),
.Y(n_2113)
);

NAND4xp25_ASAP7_75t_L g2114 ( 
.A(n_2089),
.B(n_1935),
.C(n_1925),
.D(n_1934),
.Y(n_2114)
);

AOI211xp5_ASAP7_75t_L g2115 ( 
.A1(n_2100),
.A2(n_238),
.B(n_239),
.C(n_240),
.Y(n_2115)
);

OAI211xp5_ASAP7_75t_L g2116 ( 
.A1(n_2101),
.A2(n_240),
.B(n_241),
.C(n_242),
.Y(n_2116)
);

OA21x2_ASAP7_75t_L g2117 ( 
.A1(n_2095),
.A2(n_1885),
.B(n_241),
.Y(n_2117)
);

OAI21xp33_ASAP7_75t_L g2118 ( 
.A1(n_2102),
.A2(n_1935),
.B(n_1925),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_2095),
.B(n_243),
.Y(n_2119)
);

NOR2xp33_ASAP7_75t_L g2120 ( 
.A(n_2090),
.B(n_243),
.Y(n_2120)
);

OAI221xp5_ASAP7_75t_L g2121 ( 
.A1(n_2090),
.A2(n_1962),
.B1(n_1959),
.B2(n_1907),
.C(n_1953),
.Y(n_2121)
);

O2A1O1Ixp33_ASAP7_75t_L g2122 ( 
.A1(n_2092),
.A2(n_244),
.B(n_245),
.C(n_246),
.Y(n_2122)
);

OAI21xp5_ASAP7_75t_L g2123 ( 
.A1(n_2092),
.A2(n_1917),
.B(n_1926),
.Y(n_2123)
);

AOI221xp5_ASAP7_75t_L g2124 ( 
.A1(n_2120),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.C(n_248),
.Y(n_2124)
);

AOI221xp5_ASAP7_75t_L g2125 ( 
.A1(n_2122),
.A2(n_247),
.B1(n_249),
.B2(n_250),
.C(n_251),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_2112),
.Y(n_2126)
);

AOI21xp5_ASAP7_75t_L g2127 ( 
.A1(n_2119),
.A2(n_249),
.B(n_250),
.Y(n_2127)
);

AOI211xp5_ASAP7_75t_L g2128 ( 
.A1(n_2103),
.A2(n_251),
.B(n_252),
.C(n_253),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_SL g2129 ( 
.A(n_2104),
.B(n_1946),
.Y(n_2129)
);

NAND2xp33_ASAP7_75t_SL g2130 ( 
.A(n_2108),
.B(n_1721),
.Y(n_2130)
);

INVx2_ASAP7_75t_SL g2131 ( 
.A(n_2113),
.Y(n_2131)
);

OAI211xp5_ASAP7_75t_L g2132 ( 
.A1(n_2109),
.A2(n_252),
.B(n_253),
.C(n_254),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2111),
.Y(n_2133)
);

AOI322xp5_ASAP7_75t_L g2134 ( 
.A1(n_2106),
.A2(n_1956),
.A3(n_1961),
.B1(n_1957),
.B2(n_1964),
.C1(n_1954),
.C2(n_1953),
.Y(n_2134)
);

AOI221xp5_ASAP7_75t_L g2135 ( 
.A1(n_2116),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.C(n_257),
.Y(n_2135)
);

AOI211xp5_ASAP7_75t_L g2136 ( 
.A1(n_2115),
.A2(n_255),
.B(n_256),
.C(n_258),
.Y(n_2136)
);

AOI211x1_ASAP7_75t_L g2137 ( 
.A1(n_2110),
.A2(n_1939),
.B(n_1897),
.C(n_260),
.Y(n_2137)
);

AOI221xp5_ASAP7_75t_L g2138 ( 
.A1(n_2121),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.C(n_262),
.Y(n_2138)
);

NAND4xp25_ASAP7_75t_L g2139 ( 
.A(n_2105),
.B(n_259),
.C(n_262),
.D(n_263),
.Y(n_2139)
);

NAND4xp25_ASAP7_75t_L g2140 ( 
.A(n_2114),
.B(n_263),
.C(n_265),
.D(n_266),
.Y(n_2140)
);

AOI221xp5_ASAP7_75t_L g2141 ( 
.A1(n_2107),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.C(n_269),
.Y(n_2141)
);

OAI221xp5_ASAP7_75t_L g2142 ( 
.A1(n_2118),
.A2(n_1962),
.B1(n_1959),
.B2(n_1904),
.C(n_1946),
.Y(n_2142)
);

AND4x1_ASAP7_75t_L g2143 ( 
.A(n_2123),
.B(n_267),
.C(n_268),
.D(n_269),
.Y(n_2143)
);

AOI221x1_ASAP7_75t_L g2144 ( 
.A1(n_2117),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.C(n_273),
.Y(n_2144)
);

AOI311xp33_ASAP7_75t_L g2145 ( 
.A1(n_2117),
.A2(n_270),
.A3(n_272),
.B(n_273),
.C(n_274),
.Y(n_2145)
);

O2A1O1Ixp33_ASAP7_75t_L g2146 ( 
.A1(n_2120),
.A2(n_274),
.B(n_275),
.C(n_276),
.Y(n_2146)
);

OAI221xp5_ASAP7_75t_L g2147 ( 
.A1(n_2105),
.A2(n_1904),
.B1(n_1956),
.B2(n_1939),
.C(n_279),
.Y(n_2147)
);

OAI221xp5_ASAP7_75t_L g2148 ( 
.A1(n_2105),
.A2(n_1904),
.B1(n_277),
.B2(n_278),
.C(n_280),
.Y(n_2148)
);

NOR2xp33_ASAP7_75t_L g2149 ( 
.A(n_2116),
.B(n_275),
.Y(n_2149)
);

A2O1A1Ixp33_ASAP7_75t_L g2150 ( 
.A1(n_2120),
.A2(n_277),
.B(n_280),
.C(n_281),
.Y(n_2150)
);

NOR3xp33_ASAP7_75t_L g2151 ( 
.A(n_2120),
.B(n_281),
.C(n_282),
.Y(n_2151)
);

OAI221xp5_ASAP7_75t_L g2152 ( 
.A1(n_2105),
.A2(n_282),
.B1(n_284),
.B2(n_285),
.C(n_286),
.Y(n_2152)
);

AOI221xp5_ASAP7_75t_L g2153 ( 
.A1(n_2120),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.C(n_287),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2120),
.B(n_1952),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2120),
.Y(n_2155)
);

NOR2xp67_ASAP7_75t_L g2156 ( 
.A(n_2103),
.B(n_288),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_2105),
.B(n_289),
.Y(n_2157)
);

NAND2x1_ASAP7_75t_L g2158 ( 
.A(n_2126),
.B(n_2154),
.Y(n_2158)
);

NAND4xp75_ASAP7_75t_L g2159 ( 
.A(n_2144),
.B(n_289),
.C(n_290),
.D(n_291),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2149),
.B(n_1952),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2157),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_2131),
.B(n_1952),
.Y(n_2162)
);

AND2x4_ASAP7_75t_L g2163 ( 
.A(n_2156),
.B(n_290),
.Y(n_2163)
);

NOR3xp33_ASAP7_75t_L g2164 ( 
.A(n_2155),
.B(n_2132),
.C(n_2151),
.Y(n_2164)
);

AND2x4_ASAP7_75t_L g2165 ( 
.A(n_2129),
.B(n_291),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2146),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2152),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2150),
.Y(n_2168)
);

NAND4xp25_ASAP7_75t_L g2169 ( 
.A(n_2128),
.B(n_292),
.C(n_293),
.D(n_294),
.Y(n_2169)
);

INVxp33_ASAP7_75t_SL g2170 ( 
.A(n_2133),
.Y(n_2170)
);

CKINVDCx5p33_ASAP7_75t_R g2171 ( 
.A(n_2127),
.Y(n_2171)
);

NAND3xp33_ASAP7_75t_SL g2172 ( 
.A(n_2135),
.B(n_293),
.C(n_294),
.Y(n_2172)
);

INVxp67_ASAP7_75t_L g2173 ( 
.A(n_2139),
.Y(n_2173)
);

NOR3xp33_ASAP7_75t_L g2174 ( 
.A(n_2124),
.B(n_295),
.C(n_296),
.Y(n_2174)
);

NAND3xp33_ASAP7_75t_SL g2175 ( 
.A(n_2136),
.B(n_295),
.C(n_296),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2148),
.Y(n_2176)
);

NAND3xp33_ASAP7_75t_L g2177 ( 
.A(n_2125),
.B(n_297),
.C(n_298),
.Y(n_2177)
);

NOR3xp33_ASAP7_75t_L g2178 ( 
.A(n_2153),
.B(n_297),
.C(n_298),
.Y(n_2178)
);

NOR3xp33_ASAP7_75t_L g2179 ( 
.A(n_2140),
.B(n_299),
.C(n_300),
.Y(n_2179)
);

NOR2xp33_ASAP7_75t_L g2180 ( 
.A(n_2147),
.B(n_299),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_SL g2181 ( 
.A(n_2145),
.B(n_1721),
.Y(n_2181)
);

OAI31xp33_ASAP7_75t_L g2182 ( 
.A1(n_2130),
.A2(n_302),
.A3(n_303),
.B(n_304),
.Y(n_2182)
);

NAND4xp75_ASAP7_75t_L g2183 ( 
.A(n_2141),
.B(n_302),
.C(n_304),
.D(n_305),
.Y(n_2183)
);

NOR3xp33_ASAP7_75t_L g2184 ( 
.A(n_2138),
.B(n_305),
.C(n_306),
.Y(n_2184)
);

NOR2xp67_ASAP7_75t_L g2185 ( 
.A(n_2142),
.B(n_306),
.Y(n_2185)
);

NOR2x1_ASAP7_75t_L g2186 ( 
.A(n_2159),
.B(n_2143),
.Y(n_2186)
);

AOI21xp5_ASAP7_75t_L g2187 ( 
.A1(n_2158),
.A2(n_2180),
.B(n_2173),
.Y(n_2187)
);

INVx3_ASAP7_75t_SL g2188 ( 
.A(n_2171),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2160),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2162),
.Y(n_2190)
);

NAND3xp33_ASAP7_75t_SL g2191 ( 
.A(n_2182),
.B(n_2134),
.C(n_2137),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_2165),
.B(n_2163),
.Y(n_2192)
);

NOR2x1_ASAP7_75t_L g2193 ( 
.A(n_2169),
.B(n_307),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2165),
.Y(n_2194)
);

AOI21xp5_ASAP7_75t_L g2195 ( 
.A1(n_2163),
.A2(n_2175),
.B(n_2172),
.Y(n_2195)
);

NOR3x1_ASAP7_75t_L g2196 ( 
.A(n_2183),
.B(n_308),
.C(n_310),
.Y(n_2196)
);

NOR2xp67_ASAP7_75t_L g2197 ( 
.A(n_2177),
.B(n_308),
.Y(n_2197)
);

NOR2x1_ASAP7_75t_L g2198 ( 
.A(n_2166),
.B(n_310),
.Y(n_2198)
);

NOR4xp75_ASAP7_75t_L g2199 ( 
.A(n_2181),
.B(n_2170),
.C(n_2164),
.D(n_2178),
.Y(n_2199)
);

NOR2x1_ASAP7_75t_L g2200 ( 
.A(n_2168),
.B(n_311),
.Y(n_2200)
);

OR2x2_ASAP7_75t_L g2201 ( 
.A(n_2176),
.B(n_311),
.Y(n_2201)
);

AND2x4_ASAP7_75t_L g2202 ( 
.A(n_2185),
.B(n_312),
.Y(n_2202)
);

NOR2x1_ASAP7_75t_L g2203 ( 
.A(n_2167),
.B(n_2161),
.Y(n_2203)
);

NAND3xp33_ASAP7_75t_SL g2204 ( 
.A(n_2179),
.B(n_312),
.C(n_313),
.Y(n_2204)
);

NAND4xp75_ASAP7_75t_L g2205 ( 
.A(n_2174),
.B(n_314),
.C(n_315),
.D(n_316),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2184),
.B(n_314),
.Y(n_2206)
);

NOR3xp33_ASAP7_75t_L g2207 ( 
.A(n_2158),
.B(n_315),
.C(n_317),
.Y(n_2207)
);

NOR2x1p5_ASAP7_75t_L g2208 ( 
.A(n_2159),
.B(n_317),
.Y(n_2208)
);

NOR2x1_ASAP7_75t_L g2209 ( 
.A(n_2159),
.B(n_318),
.Y(n_2209)
);

NOR2x1_ASAP7_75t_L g2210 ( 
.A(n_2159),
.B(n_318),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2159),
.Y(n_2211)
);

NOR2x1_ASAP7_75t_L g2212 ( 
.A(n_2159),
.B(n_320),
.Y(n_2212)
);

NAND3xp33_ASAP7_75t_SL g2213 ( 
.A(n_2182),
.B(n_321),
.C(n_322),
.Y(n_2213)
);

AND2x4_ASAP7_75t_L g2214 ( 
.A(n_2165),
.B(n_321),
.Y(n_2214)
);

OR2x2_ASAP7_75t_L g2215 ( 
.A(n_2169),
.B(n_322),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_2159),
.Y(n_2216)
);

AND2x2_ASAP7_75t_SL g2217 ( 
.A(n_2179),
.B(n_323),
.Y(n_2217)
);

NOR2x1_ASAP7_75t_L g2218 ( 
.A(n_2159),
.B(n_323),
.Y(n_2218)
);

NOR3x2_ASAP7_75t_L g2219 ( 
.A(n_2159),
.B(n_324),
.C(n_325),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2159),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2159),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2214),
.B(n_2207),
.Y(n_2222)
);

OAI22xp5_ASAP7_75t_L g2223 ( 
.A1(n_2201),
.A2(n_2221),
.B1(n_2220),
.B2(n_2211),
.Y(n_2223)
);

NAND2x1p5_ASAP7_75t_L g2224 ( 
.A(n_2209),
.B(n_1812),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2214),
.Y(n_2225)
);

CKINVDCx5p33_ASAP7_75t_R g2226 ( 
.A(n_2188),
.Y(n_2226)
);

XNOR2x1_ASAP7_75t_L g2227 ( 
.A(n_2186),
.B(n_325),
.Y(n_2227)
);

NOR4xp25_ASAP7_75t_L g2228 ( 
.A(n_2204),
.B(n_2213),
.C(n_2216),
.D(n_2192),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2198),
.B(n_326),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2219),
.Y(n_2230)
);

AOI221xp5_ASAP7_75t_SL g2231 ( 
.A1(n_2187),
.A2(n_327),
.B1(n_328),
.B2(n_329),
.C(n_330),
.Y(n_2231)
);

NAND3x1_ASAP7_75t_L g2232 ( 
.A(n_2200),
.B(n_329),
.C(n_331),
.Y(n_2232)
);

AND2x4_ASAP7_75t_L g2233 ( 
.A(n_2208),
.B(n_2210),
.Y(n_2233)
);

NAND3xp33_ASAP7_75t_SL g2234 ( 
.A(n_2199),
.B(n_331),
.C(n_332),
.Y(n_2234)
);

BUFx2_ASAP7_75t_L g2235 ( 
.A(n_2212),
.Y(n_2235)
);

OAI22xp5_ASAP7_75t_L g2236 ( 
.A1(n_2215),
.A2(n_1986),
.B1(n_1812),
.B2(n_1960),
.Y(n_2236)
);

NOR3xp33_ASAP7_75t_L g2237 ( 
.A(n_2189),
.B(n_333),
.C(n_334),
.Y(n_2237)
);

OAI221xp5_ASAP7_75t_L g2238 ( 
.A1(n_2218),
.A2(n_333),
.B1(n_335),
.B2(n_336),
.C(n_337),
.Y(n_2238)
);

NAND4xp75_ASAP7_75t_L g2239 ( 
.A(n_2203),
.B(n_335),
.C(n_336),
.D(n_337),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2205),
.Y(n_2240)
);

INVxp67_ASAP7_75t_SL g2241 ( 
.A(n_2196),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_2202),
.B(n_338),
.Y(n_2242)
);

BUFx3_ASAP7_75t_L g2243 ( 
.A(n_2194),
.Y(n_2243)
);

NOR3xp33_ASAP7_75t_L g2244 ( 
.A(n_2190),
.B(n_338),
.C(n_339),
.Y(n_2244)
);

CKINVDCx5p33_ASAP7_75t_R g2245 ( 
.A(n_2217),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_2193),
.B(n_2197),
.Y(n_2246)
);

AND4x1_ASAP7_75t_L g2247 ( 
.A(n_2195),
.B(n_339),
.C(n_340),
.D(n_341),
.Y(n_2247)
);

OR2x2_ASAP7_75t_L g2248 ( 
.A(n_2206),
.B(n_340),
.Y(n_2248)
);

NAND4xp75_ASAP7_75t_L g2249 ( 
.A(n_2191),
.B(n_341),
.C(n_342),
.D(n_343),
.Y(n_2249)
);

AND4x2_ASAP7_75t_L g2250 ( 
.A(n_2209),
.B(n_342),
.C(n_344),
.D(n_345),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2247),
.B(n_345),
.Y(n_2251)
);

NOR2xp33_ASAP7_75t_R g2252 ( 
.A(n_2234),
.B(n_346),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2231),
.B(n_347),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_2237),
.B(n_2244),
.Y(n_2254)
);

NOR2xp33_ASAP7_75t_R g2255 ( 
.A(n_2245),
.B(n_348),
.Y(n_2255)
);

NAND2xp33_ASAP7_75t_SL g2256 ( 
.A(n_2227),
.B(n_2229),
.Y(n_2256)
);

NOR2xp33_ASAP7_75t_R g2257 ( 
.A(n_2226),
.B(n_349),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_SL g2258 ( 
.A(n_2233),
.B(n_349),
.Y(n_2258)
);

NOR3xp33_ASAP7_75t_SL g2259 ( 
.A(n_2223),
.B(n_350),
.C(n_351),
.Y(n_2259)
);

NOR2xp33_ASAP7_75t_R g2260 ( 
.A(n_2225),
.B(n_350),
.Y(n_2260)
);

NOR2xp33_ASAP7_75t_R g2261 ( 
.A(n_2235),
.B(n_351),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2249),
.B(n_352),
.Y(n_2262)
);

NAND2xp33_ASAP7_75t_SL g2263 ( 
.A(n_2242),
.B(n_352),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_2233),
.B(n_353),
.Y(n_2264)
);

XNOR2xp5_ASAP7_75t_L g2265 ( 
.A(n_2232),
.B(n_353),
.Y(n_2265)
);

NAND2xp33_ASAP7_75t_SL g2266 ( 
.A(n_2222),
.B(n_354),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_2239),
.B(n_355),
.Y(n_2267)
);

NOR2xp67_ASAP7_75t_L g2268 ( 
.A(n_2238),
.B(n_356),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_SL g2269 ( 
.A(n_2228),
.B(n_2243),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2241),
.B(n_356),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_SL g2271 ( 
.A(n_2230),
.B(n_357),
.Y(n_2271)
);

NOR2xp33_ASAP7_75t_R g2272 ( 
.A(n_2240),
.B(n_357),
.Y(n_2272)
);

NOR2xp33_ASAP7_75t_R g2273 ( 
.A(n_2246),
.B(n_358),
.Y(n_2273)
);

NAND3xp33_ASAP7_75t_L g2274 ( 
.A(n_2248),
.B(n_358),
.C(n_359),
.Y(n_2274)
);

XNOR2xp5_ASAP7_75t_L g2275 ( 
.A(n_2224),
.B(n_359),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2236),
.B(n_360),
.Y(n_2276)
);

NOR2xp33_ASAP7_75t_R g2277 ( 
.A(n_2250),
.B(n_360),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_SL g2278 ( 
.A(n_2231),
.B(n_361),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_SL g2279 ( 
.A(n_2231),
.B(n_361),
.Y(n_2279)
);

NAND3xp33_ASAP7_75t_L g2280 ( 
.A(n_2231),
.B(n_362),
.C(n_363),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2275),
.Y(n_2281)
);

BUFx2_ASAP7_75t_L g2282 ( 
.A(n_2277),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2265),
.Y(n_2283)
);

AO22x2_ASAP7_75t_L g2284 ( 
.A1(n_2269),
.A2(n_362),
.B1(n_363),
.B2(n_364),
.Y(n_2284)
);

HB1xp67_ASAP7_75t_L g2285 ( 
.A(n_2260),
.Y(n_2285)
);

AND2x4_ASAP7_75t_L g2286 ( 
.A(n_2259),
.B(n_365),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2264),
.Y(n_2287)
);

AND2x2_ASAP7_75t_L g2288 ( 
.A(n_2251),
.B(n_366),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2267),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2262),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2270),
.Y(n_2291)
);

HB1xp67_ASAP7_75t_L g2292 ( 
.A(n_2257),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2258),
.Y(n_2293)
);

OAI22xp5_ASAP7_75t_L g2294 ( 
.A1(n_2280),
.A2(n_1960),
.B1(n_1928),
.B2(n_1920),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2253),
.Y(n_2295)
);

AO22x2_ASAP7_75t_L g2296 ( 
.A1(n_2278),
.A2(n_2279),
.B1(n_2271),
.B2(n_2274),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2261),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2276),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2272),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2284),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2284),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2282),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2288),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2286),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2285),
.Y(n_2305)
);

AO22x2_ASAP7_75t_L g2306 ( 
.A1(n_2297),
.A2(n_2254),
.B1(n_2256),
.B2(n_2266),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2296),
.Y(n_2307)
);

OAI22xp5_ASAP7_75t_L g2308 ( 
.A1(n_2293),
.A2(n_2268),
.B1(n_2252),
.B2(n_2273),
.Y(n_2308)
);

OAI22xp5_ASAP7_75t_L g2309 ( 
.A1(n_2283),
.A2(n_2263),
.B1(n_2255),
.B2(n_369),
.Y(n_2309)
);

CKINVDCx20_ASAP7_75t_R g2310 ( 
.A(n_2281),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2292),
.Y(n_2311)
);

NOR2xp33_ASAP7_75t_L g2312 ( 
.A(n_2309),
.B(n_2302),
.Y(n_2312)
);

INVx1_ASAP7_75t_SL g2313 ( 
.A(n_2300),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2301),
.Y(n_2314)
);

OAI21x1_ASAP7_75t_L g2315 ( 
.A1(n_2308),
.A2(n_2299),
.B(n_2295),
.Y(n_2315)
);

CKINVDCx20_ASAP7_75t_R g2316 ( 
.A(n_2310),
.Y(n_2316)
);

HB1xp67_ASAP7_75t_L g2317 ( 
.A(n_2307),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2306),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_2303),
.Y(n_2319)
);

XNOR2xp5_ASAP7_75t_L g2320 ( 
.A(n_2306),
.B(n_2296),
.Y(n_2320)
);

XNOR2xp5_ASAP7_75t_L g2321 ( 
.A(n_2316),
.B(n_2320),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2317),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2318),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_2314),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2322),
.B(n_2313),
.Y(n_2325)
);

NAND2xp33_ASAP7_75t_R g2326 ( 
.A(n_2324),
.B(n_2304),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2321),
.B(n_2287),
.Y(n_2327)
);

AOI22xp33_ASAP7_75t_SL g2328 ( 
.A1(n_2323),
.A2(n_2311),
.B1(n_2305),
.B2(n_2319),
.Y(n_2328)
);

AO21x2_ASAP7_75t_L g2329 ( 
.A1(n_2325),
.A2(n_2312),
.B(n_2315),
.Y(n_2329)
);

NOR3xp33_ASAP7_75t_L g2330 ( 
.A(n_2328),
.B(n_2289),
.C(n_2290),
.Y(n_2330)
);

NOR3xp33_ASAP7_75t_SL g2331 ( 
.A(n_2326),
.B(n_2291),
.C(n_2298),
.Y(n_2331)
);

AOI22xp33_ASAP7_75t_SL g2332 ( 
.A1(n_2329),
.A2(n_2327),
.B1(n_2294),
.B2(n_369),
.Y(n_2332)
);

XNOR2xp5_ASAP7_75t_L g2333 ( 
.A(n_2331),
.B(n_367),
.Y(n_2333)
);

NOR2xp33_ASAP7_75t_L g2334 ( 
.A(n_2333),
.B(n_2330),
.Y(n_2334)
);

AOI21xp33_ASAP7_75t_L g2335 ( 
.A1(n_2332),
.A2(n_367),
.B(n_368),
.Y(n_2335)
);

OR2x6_ASAP7_75t_L g2336 ( 
.A(n_2334),
.B(n_368),
.Y(n_2336)
);

AOI22xp33_ASAP7_75t_L g2337 ( 
.A1(n_2336),
.A2(n_2335),
.B1(n_371),
.B2(n_372),
.Y(n_2337)
);

OR2x6_ASAP7_75t_L g2338 ( 
.A(n_2337),
.B(n_370),
.Y(n_2338)
);

AOI221xp5_ASAP7_75t_L g2339 ( 
.A1(n_2338),
.A2(n_372),
.B1(n_373),
.B2(n_374),
.C(n_375),
.Y(n_2339)
);

AOI211xp5_ASAP7_75t_L g2340 ( 
.A1(n_2339),
.A2(n_376),
.B(n_378),
.C(n_379),
.Y(n_2340)
);


endmodule