module fake_jpeg_27013_n_74 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_74);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_74;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_73;
wire n_71;
wire n_35;
wire n_59;
wire n_68;
wire n_52;
wire n_48;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_28;
wire n_38;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_7),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_0),
.B(n_19),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_1),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_1),
.Y(n_51)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

AO22x2_ASAP7_75t_L g41 ( 
.A1(n_27),
.A2(n_12),
.B1(n_25),
.B2(n_24),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_31),
.B1(n_2),
.B2(n_3),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_41),
.A2(n_32),
.B1(n_27),
.B2(n_13),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_46),
.B1(n_47),
.B2(n_50),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_41),
.B(n_32),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_4),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_10),
.B1(n_22),
.B2(n_21),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_5),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_26),
.B1(n_20),
.B2(n_17),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_51),
.B(n_9),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_3),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_52),
.B(n_4),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_54),
.A2(n_43),
.B1(n_46),
.B2(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_11),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_56),
.C(n_64),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

AOI322xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_61),
.A3(n_64),
.B1(n_63),
.B2(n_66),
.C1(n_51),
.C2(n_62),
.Y(n_71)
);

AOI322xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_59),
.A3(n_65),
.B1(n_42),
.B2(n_60),
.C1(n_48),
.C2(n_8),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_65),
.B(n_60),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_67),
.B1(n_48),
.B2(n_9),
.Y(n_74)
);


endmodule