module real_jpeg_5658_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_288;
wire n_78;
wire n_83;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_0),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_0),
.B(n_183),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_0),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_0),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_0),
.B(n_288),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_0),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_0),
.B(n_377),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_0),
.B(n_106),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_1),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_1),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_1),
.Y(n_262)
);

INVx8_ASAP7_75t_L g313 ( 
.A(n_1),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_1),
.Y(n_333)
);

BUFx5_ASAP7_75t_L g350 ( 
.A(n_1),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_2),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_2),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_2),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_2),
.B(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g178 ( 
.A(n_2),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_2),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_2),
.B(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_3),
.Y(n_163)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_3),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g238 ( 
.A(n_3),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_4),
.B(n_35),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_4),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_4),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_4),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_4),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_4),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_4),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_4),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_5),
.B(n_66),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_5),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_5),
.B(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_5),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_5),
.B(n_221),
.Y(n_220)
);

AND2x2_ASAP7_75t_SL g285 ( 
.A(n_5),
.B(n_201),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_5),
.B(n_374),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_5),
.B(n_194),
.Y(n_414)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_6),
.Y(n_87)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_6),
.Y(n_141)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_6),
.Y(n_233)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_7),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_8),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_8),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_8),
.B(n_308),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_8),
.B(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_8),
.B(n_354),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_8),
.B(n_97),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_8),
.B(n_293),
.Y(n_399)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_9),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_9),
.Y(n_181)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_9),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_9),
.Y(n_317)
);

BUFx5_ASAP7_75t_L g371 ( 
.A(n_9),
.Y(n_371)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_11),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_11),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_11),
.Y(n_273)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_13),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_13),
.B(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_13),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_13),
.B(n_293),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_13),
.B(n_333),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_13),
.B(n_348),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_13),
.B(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_14),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_14),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_14),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_14),
.B(n_311),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_14),
.B(n_330),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_14),
.B(n_181),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_14),
.B(n_386),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_14),
.B(n_357),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_15),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_15),
.B(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_15),
.B(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_15),
.B(n_341),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_15),
.B(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_15),
.B(n_389),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_15),
.B(n_401),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_16),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_17),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_17),
.B(n_59),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_17),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_17),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_17),
.B(n_97),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_17),
.B(n_271),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_17),
.B(n_290),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_17),
.B(n_311),
.Y(n_415)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_19),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_19),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_19),
.B(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_19),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_19),
.B(n_194),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_526),
.B(n_529),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_76),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_75),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_48),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_24),
.B(n_48),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_38),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.C(n_34),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_26),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_26),
.A2(n_30),
.B1(n_39),
.B2(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_28),
.Y(n_222)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_28),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_30),
.A2(n_52),
.B1(n_56),
.B2(n_57),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_30),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_30),
.B(n_52),
.C(n_58),
.Y(n_72)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_32),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_33),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_34),
.B(n_74),
.Y(n_73)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_37),
.Y(n_150)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_71),
.C(n_73),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_49),
.B(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_60),
.C(n_61),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_50),
.B(n_116),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_58),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_52),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_52),
.A2(n_57),
.B1(n_67),
.B2(n_109),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_54),
.Y(n_146)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_54),
.Y(n_276)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_55),
.Y(n_133)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_55),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_62),
.C(n_67),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_60),
.B(n_61),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_62),
.A2(n_63),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_65),
.Y(n_284)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_67),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_67),
.A2(n_104),
.B1(n_105),
.B2(n_109),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_69),
.Y(n_206)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_69),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_69),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_69),
.Y(n_410)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_71),
.A2(n_72),
.B1(n_73),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

AO21x1_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_120),
.B(n_525),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_117),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_78),
.B(n_117),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_114),
.C(n_115),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_79),
.A2(n_80),
.B1(n_521),
.B2(n_522),
.Y(n_520)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_102),
.C(n_110),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_81),
.A2(n_82),
.B1(n_502),
.B2(n_504),
.Y(n_501)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_91),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_88),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_88),
.C(n_91),
.Y(n_114)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_90),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_90),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_90),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_90),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.C(n_98),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_92),
.B(n_492),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_93),
.A2(n_94),
.B1(n_98),
.B2(n_99),
.Y(n_492)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx6_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_102),
.A2(n_110),
.B1(n_111),
.B2(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_102),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.C(n_109),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_103),
.B(n_498),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_104),
.A2(n_105),
.B1(n_193),
.B2(n_196),
.Y(n_192)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_105),
.B(n_189),
.C(n_193),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_108),
.Y(n_291)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_114),
.B(n_115),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_519),
.B(n_524),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_485),
.B(n_516),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_296),
.B(n_484),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_246),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_124),
.B(n_246),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_186),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_125),
.B(n_187),
.C(n_223),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_160),
.C(n_169),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_126),
.B(n_249),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_137),
.C(n_147),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_127),
.B(n_469),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_131),
.C(n_134),
.Y(n_168)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_129),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.Y(n_130)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_137),
.A2(n_138),
.B1(n_147),
.B2(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.C(n_145),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_139),
.B(n_145),
.Y(n_459)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_142),
.B(n_459),
.Y(n_458)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_147),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_148),
.B(n_152),
.C(n_157),
.Y(n_243)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_156),
.B1(n_157),
.B2(n_159),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_152),
.Y(n_159)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_155),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_155),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_156),
.B(n_193),
.C(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_156),
.A2(n_157),
.B1(n_193),
.B2(n_196),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_160),
.B(n_169),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_168),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_161)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_162),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_164),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_164),
.B(n_166),
.C(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_164),
.A2(n_167),
.B1(n_235),
.B2(n_239),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_167),
.B(n_228),
.C(n_239),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_168),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_180),
.C(n_182),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_170),
.B(n_279),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.C(n_178),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_171),
.B(n_258),
.Y(n_257)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_175),
.B(n_178),
.Y(n_258)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_180),
.B(n_182),
.Y(n_279)
);

INVx4_ASAP7_75t_SL g183 ( 
.A(n_184),
.Y(n_183)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_223),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_197),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_188),
.B(n_198),
.C(n_207),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_193),
.Y(n_196)
);

BUFx8_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_207),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.C(n_204),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_199),
.B(n_204),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_200),
.B(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_202),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx8_ASAP7_75t_L g354 ( 
.A(n_206),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_220),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_215),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_209),
.B(n_215),
.C(n_220),
.Y(n_500)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_214),
.Y(n_358)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx5_ASAP7_75t_L g288 ( 
.A(n_219),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_240),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_225),
.B(n_227),
.C(n_240),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_234),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_229),
.B(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_233),
.Y(n_268)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_235),
.Y(n_239)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.C(n_244),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_244),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_250),
.C(n_253),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_248),
.B(n_251),
.Y(n_479)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_253),
.B(n_479),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_277),
.C(n_280),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_255),
.B(n_472),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_259),
.C(n_265),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_256),
.A2(n_257),
.B1(n_450),
.B2(n_451),
.Y(n_449)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_259),
.A2(n_260),
.B(n_263),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_259),
.B(n_265),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_263),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

MAJx2_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_269),
.C(n_274),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_266),
.A2(n_267),
.B1(n_269),
.B2(n_270),
.Y(n_427)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_273),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_273),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_274),
.B(n_427),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_275),
.B(n_370),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g472 ( 
.A1(n_277),
.A2(n_278),
.B1(n_280),
.B2(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_280),
.Y(n_473)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_289),
.C(n_292),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_282),
.B(n_461),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_285),
.C(n_286),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_283),
.B(n_439),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_285),
.Y(n_440)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_289),
.B(n_292),
.Y(n_461)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx6_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

AOI21x1_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_477),
.B(n_483),
.Y(n_296)
);

OAI21x1_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_464),
.B(n_476),
.Y(n_297)
);

AOI21x1_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_446),
.B(n_463),
.Y(n_298)
);

OAI21x1_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_420),
.B(n_445),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_394),
.B(n_419),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_362),
.B(n_393),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_343),
.B(n_361),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_324),
.B(n_342),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_318),
.B(n_323),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_314),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_306),
.B(n_314),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_310),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_319),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_307),
.B(n_310),
.Y(n_325)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx8_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_313),
.Y(n_322)
);

INVx4_ASAP7_75t_L g374 ( 
.A(n_313),
.Y(n_374)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_325),
.B(n_326),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_327),
.A2(n_328),
.B1(n_334),
.B2(n_335),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_327),
.B(n_337),
.C(n_339),
.Y(n_360)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_329),
.B(n_332),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_329),
.B(n_332),
.Y(n_351)
);

INVx8_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_336),
.A2(n_337),
.B1(n_339),
.B2(n_340),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_360),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_344),
.B(n_360),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_352),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_351),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_346),
.B(n_351),
.C(n_364),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_349),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_347),
.B(n_349),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_352),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_355),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_353),
.B(n_382),
.C(n_383),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_359),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_356),
.Y(n_382)
);

INVx6_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_359),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_365),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_363),
.B(n_365),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_380),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_366),
.B(n_381),
.C(n_384),
.Y(n_418)
);

XOR2x2_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_367),
.B(n_369),
.C(n_372),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_372),
.Y(n_368)
);

INVx4_ASAP7_75t_SL g370 ( 
.A(n_371),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_373),
.A2(n_375),
.B1(n_376),
.B2(n_379),
.Y(n_372)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_373),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_375),
.B(n_379),
.Y(n_403)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_384),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_387),
.Y(n_384)
);

MAJx2_ASAP7_75t_L g417 ( 
.A(n_385),
.B(n_390),
.C(n_391),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_388),
.A2(n_390),
.B1(n_391),
.B2(n_392),
.Y(n_387)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_388),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_390),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_395),
.B(n_418),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_395),
.B(n_418),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_396),
.B(n_405),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_404),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_397),
.B(n_404),
.C(n_444),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_403),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_399),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_400),
.Y(n_435)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_403),
.B(n_434),
.C(n_435),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_405),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_411),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_406),
.B(n_413),
.C(n_416),
.Y(n_423)
);

BUFx24_ASAP7_75t_SL g533 ( 
.A(n_406),
.Y(n_533)
);

FAx1_ASAP7_75t_SL g406 ( 
.A(n_407),
.B(n_408),
.CI(n_409),
.CON(n_406),
.SN(n_406)
);

MAJx2_ASAP7_75t_L g431 ( 
.A(n_407),
.B(n_408),
.C(n_409),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_412),
.A2(n_413),
.B1(n_416),
.B2(n_417),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_415),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_414),
.B(n_415),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_417),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_421),
.B(n_443),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_421),
.B(n_443),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_432),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_423),
.B(n_424),
.C(n_432),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_425),
.A2(n_426),
.B1(n_428),
.B2(n_429),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_425),
.B(n_455),
.C(n_456),
.Y(n_454)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.Y(n_429)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_430),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_431),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g432 ( 
.A(n_433),
.B(n_436),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_433),
.B(n_437),
.C(n_442),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_437),
.A2(n_438),
.B1(n_441),
.B2(n_442),
.Y(n_436)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_437),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_438),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_447),
.B(n_462),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_447),
.B(n_462),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_448),
.B(n_453),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_452),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_449),
.B(n_452),
.C(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_450),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_453),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_454),
.B(n_457),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_454),
.B(n_458),
.C(n_460),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_460),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_465),
.B(n_474),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_474),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_467),
.Y(n_465)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_466),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_471),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_468),
.B(n_481),
.C(n_482),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_471),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_478),
.B(n_480),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_478),
.B(n_480),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_513),
.Y(n_485)
);

OAI21xp33_ASAP7_75t_L g516 ( 
.A1(n_486),
.A2(n_517),
.B(n_518),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_487),
.B(n_506),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_487),
.B(n_506),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_488),
.A2(n_489),
.B1(n_495),
.B2(n_505),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_488),
.B(n_496),
.C(n_501),
.Y(n_523)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_491),
.C(n_493),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_490),
.B(n_508),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_491),
.A2(n_493),
.B1(n_494),
.B2(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_491),
.Y(n_509)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_495),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_501),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_499),
.C(n_500),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_497),
.B(n_511),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_499),
.B(n_500),
.Y(n_511)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_502),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_510),
.C(n_512),
.Y(n_506)
);

FAx1_ASAP7_75t_SL g514 ( 
.A(n_507),
.B(n_510),
.CI(n_512),
.CON(n_514),
.SN(n_514)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_514),
.B(n_515),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_514),
.B(n_515),
.Y(n_517)
);

BUFx24_ASAP7_75t_SL g535 ( 
.A(n_514),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_523),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_520),
.B(n_523),
.Y(n_524)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_521),
.Y(n_522)
);

BUFx12f_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx13_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx5_ASAP7_75t_L g531 ( 
.A(n_528),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_530),
.B(n_532),
.Y(n_529)
);

BUFx12f_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);


endmodule