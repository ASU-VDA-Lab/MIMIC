module fake_netlist_6_393_n_1049 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_186, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1049);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_186;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1049;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_209;
wire n_465;
wire n_367;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_1033;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_248;
wire n_517;
wire n_718;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_544;
wire n_468;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_886;
wire n_448;
wire n_953;
wire n_844;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_986;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_870;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_551;
wire n_258;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_594;
wire n_565;
wire n_228;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_981;
wire n_476;
wire n_880;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_928;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_956;
wire n_960;
wire n_841;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_194;
wire n_664;
wire n_949;
wire n_678;
wire n_192;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_139),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g189 ( 
.A(n_55),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_79),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_7),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_138),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_166),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_42),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_4),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_49),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_6),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_71),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_51),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_142),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_144),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_96),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_178),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_124),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_4),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_61),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_90),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_14),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_101),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_119),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_62),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_87),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_6),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_131),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_9),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_3),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_187),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_33),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_153),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_107),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_26),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_92),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_23),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_5),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_30),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_39),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_20),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_135),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_175),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_176),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_32),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_116),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_179),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_100),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_168),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_15),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_118),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_93),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_146),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_60),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_81),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_22),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_91),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_8),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_171),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_37),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_173),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_38),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_97),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_46),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_148),
.Y(n_253)
);

BUFx8_ASAP7_75t_SL g254 ( 
.A(n_121),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_67),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_129),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_113),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_68),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_186),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_226),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_238),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_191),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_207),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_196),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_210),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_238),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_198),
.Y(n_268)
);

INVxp33_ASAP7_75t_L g269 ( 
.A(n_215),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_218),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_223),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_227),
.Y(n_272)
);

INVxp33_ASAP7_75t_L g273 ( 
.A(n_194),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_231),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_188),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_217),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_190),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_231),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_220),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_216),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_225),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_216),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_239),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_189),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_229),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_239),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_250),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_250),
.Y(n_288)
);

INVxp33_ASAP7_75t_SL g289 ( 
.A(n_233),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_189),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_259),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_244),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_259),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_199),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_248),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_212),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_193),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_213),
.Y(n_298)
);

INVxp33_ASAP7_75t_SL g299 ( 
.A(n_197),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_246),
.Y(n_300)
);

INVxp33_ASAP7_75t_L g301 ( 
.A(n_254),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_214),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_221),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_230),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_203),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_235),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_242),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_254),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_237),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_237),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_306),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_273),
.B(n_192),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_195),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_294),
.Y(n_314)
);

NAND2xp33_ASAP7_75t_L g315 ( 
.A(n_280),
.B(n_189),
.Y(n_315)
);

AND2x4_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_202),
.Y(n_316)
);

AND2x4_ASAP7_75t_L g317 ( 
.A(n_282),
.B(n_202),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_284),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_263),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_265),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_264),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_284),
.Y(n_322)
);

INVxp33_ASAP7_75t_SL g323 ( 
.A(n_308),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_308),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_305),
.B(n_248),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_290),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_268),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_283),
.B(n_195),
.Y(n_328)
);

AND2x2_ASAP7_75t_SL g329 ( 
.A(n_285),
.B(n_209),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_290),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_286),
.B(n_209),
.Y(n_331)
);

INVx5_ASAP7_75t_L g332 ( 
.A(n_296),
.Y(n_332)
);

AOI22x1_ASAP7_75t_SL g333 ( 
.A1(n_274),
.A2(n_255),
.B1(n_252),
.B2(n_247),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_298),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_287),
.B(n_240),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_270),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_289),
.B(n_240),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_302),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_303),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_288),
.B(n_291),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_271),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_304),
.Y(n_342)
);

AND2x4_ASAP7_75t_L g343 ( 
.A(n_293),
.B(n_249),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_275),
.B(n_251),
.Y(n_344)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_277),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_307),
.B(n_257),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_297),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_272),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_260),
.Y(n_349)
);

BUFx8_ASAP7_75t_L g350 ( 
.A(n_261),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_264),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_292),
.Y(n_352)
);

OAI21x1_ASAP7_75t_L g353 ( 
.A1(n_269),
.A2(n_189),
.B(n_200),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_300),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_266),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_266),
.B(n_201),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_276),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_276),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_279),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_279),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_281),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_281),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_274),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_318),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_318),
.Y(n_365)
);

AND2x6_ASAP7_75t_L g366 ( 
.A(n_356),
.B(n_189),
.Y(n_366)
);

INVx5_ASAP7_75t_L g367 ( 
.A(n_326),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_326),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_322),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_322),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_311),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_326),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_326),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_312),
.B(n_301),
.Y(n_374)
);

CKINVDCx6p67_ASAP7_75t_R g375 ( 
.A(n_351),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_328),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_326),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_342),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_342),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_344),
.B(n_352),
.Y(n_380)
);

BUFx10_ASAP7_75t_L g381 ( 
.A(n_313),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_329),
.B(n_252),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_329),
.B(n_255),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_330),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_342),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_330),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_330),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_352),
.B(n_278),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_338),
.Y(n_389)
);

INVxp33_ASAP7_75t_SL g390 ( 
.A(n_325),
.Y(n_390)
);

AND3x2_ASAP7_75t_L g391 ( 
.A(n_309),
.B(n_310),
.C(n_337),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_311),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_330),
.Y(n_393)
);

INVxp33_ASAP7_75t_L g394 ( 
.A(n_354),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_331),
.B(n_204),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_338),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_351),
.B(n_205),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_340),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_330),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_334),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_334),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_334),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_334),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_334),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_339),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_339),
.Y(n_406)
);

INVx11_ASAP7_75t_L g407 ( 
.A(n_350),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_339),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_328),
.B(n_206),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_339),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_339),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_355),
.A2(n_236),
.B1(n_208),
.B2(n_211),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_314),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_333),
.B(n_278),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_319),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_319),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_320),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_320),
.Y(n_418)
);

INVx4_ASAP7_75t_L g419 ( 
.A(n_332),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_327),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_327),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_336),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_336),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_341),
.Y(n_424)
);

NAND3xp33_ASAP7_75t_L g425 ( 
.A(n_315),
.B(n_335),
.C(n_331),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_341),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_351),
.B(n_219),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_349),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_348),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_349),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_335),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_340),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_346),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_343),
.B(n_222),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_351),
.B(n_224),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_362),
.B(n_295),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_317),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_425),
.A2(n_353),
.B(n_355),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_394),
.B(n_354),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_371),
.B(n_343),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_392),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_392),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_420),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_414),
.B(n_295),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_431),
.B(n_353),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_414),
.B(n_262),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_364),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_380),
.B(n_363),
.Y(n_448)
);

INVx2_ASAP7_75t_SL g449 ( 
.A(n_395),
.Y(n_449)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_432),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_420),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_376),
.B(n_360),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_391),
.B(n_360),
.Y(n_453)
);

AOI21x1_ASAP7_75t_L g454 ( 
.A1(n_401),
.A2(n_343),
.B(n_346),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_423),
.Y(n_455)
);

AND2x2_ASAP7_75t_SL g456 ( 
.A(n_436),
.B(n_359),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_423),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_415),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_415),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_416),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_376),
.B(n_360),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_416),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_374),
.B(n_347),
.Y(n_463)
);

XNOR2x2_ASAP7_75t_L g464 ( 
.A(n_382),
.B(n_363),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_412),
.B(n_347),
.Y(n_465)
);

INVxp33_ASAP7_75t_L g466 ( 
.A(n_388),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_417),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_417),
.Y(n_468)
);

OR2x2_ASAP7_75t_L g469 ( 
.A(n_383),
.B(n_359),
.Y(n_469)
);

INVx4_ASAP7_75t_SL g470 ( 
.A(n_366),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_412),
.B(n_345),
.Y(n_471)
);

NOR2xp67_ASAP7_75t_L g472 ( 
.A(n_425),
.B(n_345),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_418),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_390),
.B(n_262),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_418),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_398),
.B(n_351),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_421),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_371),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_421),
.Y(n_479)
);

AND2x6_ASAP7_75t_L g480 ( 
.A(n_433),
.B(n_357),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_422),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_381),
.B(n_345),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_422),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_424),
.Y(n_484)
);

NAND2xp33_ASAP7_75t_R g485 ( 
.A(n_395),
.B(n_324),
.Y(n_485)
);

NOR2xp67_ASAP7_75t_L g486 ( 
.A(n_428),
.B(n_332),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_424),
.Y(n_487)
);

BUFx5_ASAP7_75t_L g488 ( 
.A(n_366),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_426),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_371),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_426),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_381),
.B(n_357),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_397),
.B(n_267),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_430),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_430),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_381),
.B(n_357),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_398),
.B(n_357),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_431),
.B(n_346),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_398),
.B(n_357),
.Y(n_499)
);

INVxp33_ASAP7_75t_L g500 ( 
.A(n_432),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_413),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_437),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_437),
.Y(n_503)
);

INVx8_ASAP7_75t_L g504 ( 
.A(n_366),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_429),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_429),
.Y(n_506)
);

NOR2xp67_ASAP7_75t_L g507 ( 
.A(n_389),
.B(n_332),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_427),
.B(n_267),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_378),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_381),
.B(n_358),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_378),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_409),
.B(n_358),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_379),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_435),
.B(n_358),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_370),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_434),
.B(n_321),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_379),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_450),
.B(n_433),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_512),
.A2(n_366),
.B1(n_375),
.B2(n_358),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_450),
.B(n_476),
.Y(n_520)
);

INVxp33_ASAP7_75t_L g521 ( 
.A(n_439),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_471),
.A2(n_366),
.B1(n_375),
.B2(n_358),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_485),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_502),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_445),
.A2(n_366),
.B1(n_315),
.B2(n_385),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_500),
.B(n_452),
.Y(n_526)
);

A2O1A1Ixp33_ASAP7_75t_L g527 ( 
.A1(n_465),
.A2(n_385),
.B(n_396),
.C(n_389),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_503),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_497),
.B(n_366),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_472),
.A2(n_361),
.B1(n_356),
.B2(n_372),
.Y(n_530)
);

NAND2xp33_ASAP7_75t_L g531 ( 
.A(n_488),
.B(n_400),
.Y(n_531)
);

AND2x6_ASAP7_75t_SL g532 ( 
.A(n_463),
.B(n_333),
.Y(n_532)
);

BUFx12f_ASAP7_75t_L g533 ( 
.A(n_448),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_509),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_511),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_516),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_478),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_499),
.B(n_461),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_488),
.B(n_402),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_440),
.B(n_396),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_447),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_443),
.B(n_372),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_451),
.B(n_373),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_L g544 ( 
.A1(n_438),
.A2(n_377),
.B(n_373),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_455),
.B(n_377),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_472),
.A2(n_514),
.B1(n_449),
.B2(n_453),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_457),
.B(n_384),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_490),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_488),
.B(n_402),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_466),
.B(n_323),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_490),
.Y(n_551)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_469),
.B(n_324),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_445),
.A2(n_317),
.B1(n_369),
.B2(n_365),
.Y(n_553)
);

A2O1A1Ixp33_ASAP7_75t_SL g554 ( 
.A1(n_438),
.A2(n_403),
.B(n_408),
.C(n_404),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_490),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_456),
.B(n_510),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_482),
.B(n_316),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_494),
.B(n_386),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_495),
.B(n_386),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_513),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_441),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_501),
.B(n_387),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_498),
.B(n_393),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_517),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_458),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_498),
.B(n_393),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_492),
.B(n_399),
.Y(n_567)
);

INVxp67_ASAP7_75t_SL g568 ( 
.A(n_488),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_496),
.B(n_399),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_459),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_442),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_464),
.B(n_505),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_515),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_488),
.B(n_404),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_506),
.B(n_368),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g576 ( 
.A1(n_504),
.A2(n_400),
.B(n_367),
.Y(n_576)
);

OR2x6_ASAP7_75t_L g577 ( 
.A(n_440),
.B(n_317),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_460),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_462),
.B(n_368),
.Y(n_579)
);

BUFx2_ASAP7_75t_L g580 ( 
.A(n_533),
.Y(n_580)
);

NAND3xp33_ASAP7_75t_L g581 ( 
.A(n_536),
.B(n_474),
.C(n_493),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_571),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_524),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_526),
.B(n_508),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_541),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_SL g586 ( 
.A(n_523),
.B(n_323),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_520),
.B(n_538),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_541),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_528),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_556),
.B(n_470),
.Y(n_590)
);

AO21x2_ASAP7_75t_L g591 ( 
.A1(n_554),
.A2(n_527),
.B(n_544),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_540),
.B(n_467),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_518),
.B(n_480),
.Y(n_593)
);

NAND2xp33_ASAP7_75t_SL g594 ( 
.A(n_525),
.B(n_504),
.Y(n_594)
);

INVx1_ASAP7_75t_SL g595 ( 
.A(n_561),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_534),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_560),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_521),
.B(n_480),
.Y(n_598)
);

NOR3xp33_ASAP7_75t_SL g599 ( 
.A(n_550),
.B(n_444),
.C(n_232),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_564),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_521),
.B(n_480),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_550),
.B(n_468),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_578),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_552),
.B(n_446),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_555),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_555),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_578),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_565),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_537),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_561),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_546),
.B(n_470),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_537),
.B(n_316),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_572),
.A2(n_473),
.B1(n_477),
.B2(n_475),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_530),
.A2(n_480),
.B1(n_481),
.B2(n_479),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_572),
.A2(n_483),
.B1(n_487),
.B2(n_484),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_522),
.A2(n_491),
.B1(n_489),
.B2(n_504),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_570),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_535),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_555),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_555),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_540),
.B(n_470),
.Y(n_621)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_577),
.B(n_316),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_573),
.Y(n_623)
);

BUFx4f_ASAP7_75t_L g624 ( 
.A(n_577),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_577),
.B(n_454),
.Y(n_625)
);

INVx5_ASAP7_75t_L g626 ( 
.A(n_548),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_573),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_548),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_551),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_551),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_557),
.B(n_407),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_562),
.Y(n_632)
);

INVx3_ASAP7_75t_SL g633 ( 
.A(n_539),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_542),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_543),
.Y(n_635)
);

BUFx2_ASAP7_75t_L g636 ( 
.A(n_532),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_545),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_529),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_547),
.Y(n_639)
);

OAI21xp5_ASAP7_75t_L g640 ( 
.A1(n_587),
.A2(n_527),
.B(n_525),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_583),
.Y(n_641)
);

XOR2xp5_ASAP7_75t_L g642 ( 
.A(n_582),
.B(n_519),
.Y(n_642)
);

BUFx2_ASAP7_75t_L g643 ( 
.A(n_609),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_594),
.A2(n_531),
.B(n_568),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_594),
.A2(n_611),
.B(n_569),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_584),
.B(n_553),
.Y(n_646)
);

OAI21x1_ASAP7_75t_L g647 ( 
.A1(n_638),
.A2(n_611),
.B(n_576),
.Y(n_647)
);

AOI21x1_ASAP7_75t_L g648 ( 
.A1(n_593),
.A2(n_567),
.B(n_566),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_589),
.Y(n_649)
);

OR2x6_ASAP7_75t_L g650 ( 
.A(n_609),
.B(n_558),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_602),
.B(n_563),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_612),
.B(n_553),
.Y(n_652)
);

BUFx4f_ASAP7_75t_L g653 ( 
.A(n_580),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g654 ( 
.A1(n_613),
.A2(n_559),
.B1(n_574),
.B2(n_539),
.Y(n_654)
);

OAI21x1_ASAP7_75t_L g655 ( 
.A1(n_638),
.A2(n_579),
.B(n_575),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_602),
.B(n_554),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_L g657 ( 
.A1(n_616),
.A2(n_574),
.B(n_549),
.Y(n_657)
);

OAI21xp5_ASAP7_75t_L g658 ( 
.A1(n_638),
.A2(n_549),
.B(n_405),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_610),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_632),
.A2(n_400),
.B(n_486),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_635),
.A2(n_400),
.B(n_486),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_581),
.B(n_407),
.Y(n_662)
);

OAI21x1_ASAP7_75t_L g663 ( 
.A1(n_585),
.A2(n_368),
.B(n_403),
.Y(n_663)
);

NAND2x1_ASAP7_75t_L g664 ( 
.A(n_605),
.B(n_368),
.Y(n_664)
);

BUFx12f_ASAP7_75t_L g665 ( 
.A(n_610),
.Y(n_665)
);

AND2x2_ASAP7_75t_SL g666 ( 
.A(n_624),
.B(n_350),
.Y(n_666)
);

NOR2xp67_ASAP7_75t_L g667 ( 
.A(n_582),
.B(n_618),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_637),
.A2(n_400),
.B(n_367),
.Y(n_668)
);

O2A1O1Ixp5_ASAP7_75t_L g669 ( 
.A1(n_590),
.A2(n_411),
.B(n_410),
.C(n_403),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_SL g670 ( 
.A(n_586),
.B(n_350),
.Y(n_670)
);

AOI21x1_ASAP7_75t_L g671 ( 
.A1(n_590),
.A2(n_405),
.B(n_401),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_637),
.A2(n_367),
.B(n_507),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_614),
.A2(n_411),
.B(n_410),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_639),
.A2(n_367),
.B(n_507),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_585),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_634),
.B(n_406),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_L g677 ( 
.A1(n_613),
.A2(n_406),
.B(n_234),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_588),
.Y(n_678)
);

AOI221xp5_ASAP7_75t_SL g679 ( 
.A1(n_608),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.C(n_3),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_634),
.B(n_228),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_603),
.B(n_241),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_596),
.B(n_243),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_621),
.Y(n_683)
);

A2O1A1Ixp33_ASAP7_75t_L g684 ( 
.A1(n_631),
.A2(n_245),
.B(n_253),
.C(n_256),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_L g685 ( 
.A1(n_615),
.A2(n_258),
.B(n_332),
.Y(n_685)
);

AOI21x1_ASAP7_75t_L g686 ( 
.A1(n_598),
.A2(n_189),
.B(n_332),
.Y(n_686)
);

NAND2xp33_ASAP7_75t_L g687 ( 
.A(n_601),
.B(n_189),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_592),
.B(n_419),
.Y(n_688)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_595),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_591),
.A2(n_419),
.B(n_34),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_597),
.B(n_0),
.Y(n_691)
);

OAI21xp5_ASAP7_75t_L g692 ( 
.A1(n_615),
.A2(n_419),
.B(n_36),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_SL g693 ( 
.A(n_624),
.B(n_419),
.Y(n_693)
);

NOR2xp67_ASAP7_75t_L g694 ( 
.A(n_631),
.B(n_35),
.Y(n_694)
);

O2A1O1Ixp33_ASAP7_75t_L g695 ( 
.A1(n_692),
.A2(n_604),
.B(n_599),
.C(n_636),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_641),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_646),
.B(n_592),
.Y(n_697)
);

OAI21x1_ASAP7_75t_L g698 ( 
.A1(n_663),
.A2(n_627),
.B(n_623),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_640),
.A2(n_644),
.B(n_692),
.Y(n_699)
);

AOI221xp5_ASAP7_75t_L g700 ( 
.A1(n_679),
.A2(n_600),
.B1(n_617),
.B2(n_592),
.C(n_607),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_662),
.A2(n_625),
.B1(n_622),
.B2(n_630),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_651),
.B(n_627),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_643),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_649),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_SL g705 ( 
.A(n_659),
.B(n_621),
.Y(n_705)
);

OR2x6_ASAP7_75t_L g706 ( 
.A(n_665),
.B(n_621),
.Y(n_706)
);

AO21x2_ASAP7_75t_L g707 ( 
.A1(n_640),
.A2(n_645),
.B(n_690),
.Y(n_707)
);

NAND2x1p5_ASAP7_75t_L g708 ( 
.A(n_653),
.B(n_626),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_652),
.B(n_628),
.Y(n_709)
);

AO31x2_ASAP7_75t_L g710 ( 
.A1(n_656),
.A2(n_591),
.A3(n_633),
.B(n_625),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_689),
.Y(n_711)
);

O2A1O1Ixp33_ASAP7_75t_L g712 ( 
.A1(n_691),
.A2(n_633),
.B(n_625),
.C(n_629),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_642),
.A2(n_629),
.B1(n_620),
.B2(n_619),
.Y(n_713)
);

OAI21xp5_ASAP7_75t_SL g714 ( 
.A1(n_684),
.A2(n_606),
.B(n_605),
.Y(n_714)
);

OAI21x1_ASAP7_75t_L g715 ( 
.A1(n_655),
.A2(n_606),
.B(n_605),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_667),
.B(n_619),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_675),
.Y(n_717)
);

OA21x2_ASAP7_75t_L g718 ( 
.A1(n_648),
.A2(n_626),
.B(n_40),
.Y(n_718)
);

OAI21x1_ASAP7_75t_L g719 ( 
.A1(n_686),
.A2(n_626),
.B(n_41),
.Y(n_719)
);

O2A1O1Ixp33_ASAP7_75t_SL g720 ( 
.A1(n_657),
.A2(n_1),
.B(n_2),
.C(n_5),
.Y(n_720)
);

NOR2xp67_ASAP7_75t_L g721 ( 
.A(n_680),
.B(n_43),
.Y(n_721)
);

AO31x2_ASAP7_75t_L g722 ( 
.A1(n_654),
.A2(n_7),
.A3(n_8),
.B(n_9),
.Y(n_722)
);

OAI21x1_ASAP7_75t_SL g723 ( 
.A1(n_671),
.A2(n_10),
.B(n_11),
.Y(n_723)
);

AOI221x1_ASAP7_75t_L g724 ( 
.A1(n_654),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_670),
.B(n_12),
.Y(n_725)
);

BUFx12f_ASAP7_75t_L g726 ( 
.A(n_666),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_678),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_657),
.A2(n_185),
.B(n_45),
.Y(n_728)
);

OAI21x1_ASAP7_75t_L g729 ( 
.A1(n_673),
.A2(n_47),
.B(n_44),
.Y(n_729)
);

A2O1A1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_694),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_683),
.B(n_16),
.Y(n_731)
);

AOI21x1_ASAP7_75t_L g732 ( 
.A1(n_672),
.A2(n_50),
.B(n_48),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_674),
.A2(n_114),
.B(n_184),
.Y(n_733)
);

NAND3xp33_ASAP7_75t_L g734 ( 
.A(n_687),
.B(n_682),
.C(n_681),
.Y(n_734)
);

CKINVDCx6p67_ASAP7_75t_R g735 ( 
.A(n_650),
.Y(n_735)
);

O2A1O1Ixp33_ASAP7_75t_SL g736 ( 
.A1(n_688),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_660),
.A2(n_661),
.B(n_693),
.Y(n_737)
);

OAI21x1_ASAP7_75t_L g738 ( 
.A1(n_673),
.A2(n_115),
.B(n_183),
.Y(n_738)
);

OAI21x1_ASAP7_75t_L g739 ( 
.A1(n_668),
.A2(n_112),
.B(n_182),
.Y(n_739)
);

OAI21x1_ASAP7_75t_L g740 ( 
.A1(n_669),
.A2(n_111),
.B(n_181),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_SL g741 ( 
.A(n_653),
.B(n_52),
.Y(n_741)
);

AO31x2_ASAP7_75t_L g742 ( 
.A1(n_676),
.A2(n_17),
.A3(n_18),
.B(n_19),
.Y(n_742)
);

OAI22xp33_ASAP7_75t_L g743 ( 
.A1(n_650),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_681),
.B(n_21),
.Y(n_744)
);

BUFx8_ASAP7_75t_L g745 ( 
.A(n_650),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_677),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_746)
);

OAI21x1_ASAP7_75t_L g747 ( 
.A1(n_658),
.A2(n_123),
.B(n_180),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_658),
.A2(n_122),
.B(n_177),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_664),
.B(n_53),
.Y(n_749)
);

O2A1O1Ixp33_ASAP7_75t_L g750 ( 
.A1(n_685),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_685),
.Y(n_751)
);

AO31x2_ASAP7_75t_L g752 ( 
.A1(n_645),
.A2(n_25),
.A3(n_27),
.B(n_28),
.Y(n_752)
);

OAI21x1_ASAP7_75t_L g753 ( 
.A1(n_647),
.A2(n_126),
.B(n_174),
.Y(n_753)
);

OAI22xp33_ASAP7_75t_L g754 ( 
.A1(n_741),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_754)
);

INVx5_ASAP7_75t_L g755 ( 
.A(n_703),
.Y(n_755)
);

INVx8_ASAP7_75t_L g756 ( 
.A(n_706),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_746),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_708),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_699),
.A2(n_128),
.B(n_172),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_717),
.Y(n_760)
);

BUFx12f_ASAP7_75t_L g761 ( 
.A(n_726),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_703),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_725),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_763)
);

OAI22xp33_ASAP7_75t_L g764 ( 
.A1(n_724),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_SL g765 ( 
.A1(n_751),
.A2(n_58),
.B1(n_59),
.B2(n_63),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_734),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_766)
);

OAI22xp33_ASAP7_75t_L g767 ( 
.A1(n_701),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_697),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_696),
.Y(n_769)
);

BUFx4f_ASAP7_75t_SL g770 ( 
.A(n_703),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_704),
.Y(n_771)
);

CKINVDCx11_ASAP7_75t_R g772 ( 
.A(n_706),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_727),
.Y(n_773)
);

BUFx4_ASAP7_75t_R g774 ( 
.A(n_705),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_709),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_721),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_776)
);

INVx1_ASAP7_75t_SL g777 ( 
.A(n_735),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_SL g778 ( 
.A1(n_728),
.A2(n_80),
.B1(n_82),
.B2(n_83),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_SL g779 ( 
.A1(n_744),
.A2(n_745),
.B1(n_748),
.B2(n_707),
.Y(n_779)
);

BUFx4f_ASAP7_75t_SL g780 ( 
.A(n_711),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_722),
.Y(n_781)
);

OAI22x1_ASAP7_75t_L g782 ( 
.A1(n_713),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_SL g783 ( 
.A1(n_750),
.A2(n_745),
.B1(n_720),
.B2(n_723),
.Y(n_783)
);

INVx6_ASAP7_75t_L g784 ( 
.A(n_731),
.Y(n_784)
);

CKINVDCx11_ASAP7_75t_R g785 ( 
.A(n_695),
.Y(n_785)
);

BUFx12f_ASAP7_75t_L g786 ( 
.A(n_716),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_743),
.A2(n_88),
.B1(n_89),
.B2(n_94),
.Y(n_787)
);

INVxp67_ASAP7_75t_SL g788 ( 
.A(n_702),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_749),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_700),
.A2(n_95),
.B1(n_98),
.B2(n_99),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_710),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_733),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_792)
);

OAI22xp33_ASAP7_75t_SL g793 ( 
.A1(n_730),
.A2(n_105),
.B1(n_106),
.B2(n_108),
.Y(n_793)
);

BUFx8_ASAP7_75t_SL g794 ( 
.A(n_732),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_710),
.B(n_109),
.Y(n_795)
);

BUFx4f_ASAP7_75t_L g796 ( 
.A(n_718),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_710),
.Y(n_797)
);

BUFx2_ASAP7_75t_L g798 ( 
.A(n_742),
.Y(n_798)
);

BUFx2_ASAP7_75t_L g799 ( 
.A(n_742),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_722),
.Y(n_800)
);

CKINVDCx14_ASAP7_75t_R g801 ( 
.A(n_712),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_714),
.A2(n_110),
.B1(n_117),
.B2(n_120),
.Y(n_802)
);

OAI22xp33_ASAP7_75t_L g803 ( 
.A1(n_737),
.A2(n_125),
.B1(n_127),
.B2(n_130),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_698),
.Y(n_804)
);

NAND2x1p5_ASAP7_75t_L g805 ( 
.A(n_718),
.B(n_132),
.Y(n_805)
);

BUFx8_ASAP7_75t_L g806 ( 
.A(n_742),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_729),
.A2(n_133),
.B1(n_134),
.B2(n_136),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_722),
.Y(n_808)
);

INVx6_ASAP7_75t_L g809 ( 
.A(n_736),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_SL g810 ( 
.A1(n_764),
.A2(n_752),
.B(n_738),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_775),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_804),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_781),
.Y(n_813)
);

CKINVDCx14_ASAP7_75t_R g814 ( 
.A(n_761),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_800),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_808),
.Y(n_816)
);

OAI21xp33_ASAP7_75t_SL g817 ( 
.A1(n_802),
.A2(n_747),
.B(n_753),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_769),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_771),
.Y(n_819)
);

OA21x2_ASAP7_75t_L g820 ( 
.A1(n_795),
.A2(n_798),
.B(n_799),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_755),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_791),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_791),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_760),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_797),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_773),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_788),
.B(n_752),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_806),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_780),
.B(n_789),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_806),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_796),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_796),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_795),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_805),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_805),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_794),
.Y(n_836)
);

OAI21x1_ASAP7_75t_L g837 ( 
.A1(n_759),
.A2(n_719),
.B(n_740),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_801),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_755),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_784),
.B(n_715),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_755),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_755),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_762),
.Y(n_843)
);

NAND2x1p5_ASAP7_75t_L g844 ( 
.A(n_758),
.B(n_739),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_784),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_777),
.Y(n_846)
);

INVx1_ASAP7_75t_SL g847 ( 
.A(n_770),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_779),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_756),
.Y(n_849)
);

BUFx3_ASAP7_75t_L g850 ( 
.A(n_756),
.Y(n_850)
);

OAI21x1_ASAP7_75t_L g851 ( 
.A1(n_807),
.A2(n_137),
.B(n_140),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_758),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_809),
.Y(n_853)
);

AO21x2_ASAP7_75t_L g854 ( 
.A1(n_810),
.A2(n_754),
.B(n_803),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_818),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_850),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_818),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_818),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_833),
.B(n_785),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_812),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_833),
.B(n_783),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_819),
.Y(n_862)
);

AND2x6_ASAP7_75t_L g863 ( 
.A(n_832),
.B(n_774),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_822),
.B(n_783),
.Y(n_864)
);

AO21x2_ASAP7_75t_L g865 ( 
.A1(n_810),
.A2(n_767),
.B(n_776),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_820),
.B(n_777),
.Y(n_866)
);

BUFx3_ASAP7_75t_L g867 ( 
.A(n_850),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_848),
.B(n_838),
.Y(n_868)
);

AO21x2_ASAP7_75t_L g869 ( 
.A1(n_813),
.A2(n_793),
.B(n_809),
.Y(n_869)
);

OR2x6_ASAP7_75t_L g870 ( 
.A(n_831),
.B(n_756),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_813),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_822),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_822),
.B(n_782),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_823),
.Y(n_874)
);

OAI21xp5_ASAP7_75t_L g875 ( 
.A1(n_817),
.A2(n_793),
.B(n_757),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_819),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_831),
.Y(n_877)
);

AO21x2_ASAP7_75t_L g878 ( 
.A1(n_815),
.A2(n_778),
.B(n_765),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_831),
.Y(n_879)
);

OAI21x1_ASAP7_75t_L g880 ( 
.A1(n_837),
.A2(n_792),
.B(n_766),
.Y(n_880)
);

INVx4_ASAP7_75t_L g881 ( 
.A(n_849),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_820),
.Y(n_882)
);

OR2x2_ASAP7_75t_L g883 ( 
.A(n_866),
.B(n_820),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_860),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_866),
.B(n_820),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_877),
.B(n_838),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_871),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_871),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_877),
.B(n_833),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_879),
.B(n_830),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_866),
.B(n_830),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_855),
.Y(n_892)
);

NOR2x1_ASAP7_75t_SL g893 ( 
.A(n_869),
.B(n_830),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_856),
.B(n_832),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_859),
.B(n_811),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_879),
.B(n_840),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_855),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_864),
.B(n_840),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_864),
.B(n_823),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_856),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_859),
.B(n_824),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_865),
.A2(n_854),
.B1(n_875),
.B2(n_848),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_857),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_864),
.B(n_823),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_887),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_887),
.B(n_862),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_894),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_901),
.B(n_868),
.Y(n_908)
);

INVx1_ASAP7_75t_SL g909 ( 
.A(n_886),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_898),
.B(n_868),
.Y(n_910)
);

INVx5_ASAP7_75t_L g911 ( 
.A(n_891),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_902),
.B(n_861),
.Y(n_912)
);

OR2x2_ASAP7_75t_L g913 ( 
.A(n_895),
.B(n_861),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_888),
.B(n_862),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_888),
.B(n_876),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_898),
.B(n_856),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_890),
.Y(n_917)
);

INVxp67_ASAP7_75t_L g918 ( 
.A(n_886),
.Y(n_918)
);

OAI221xp5_ASAP7_75t_L g919 ( 
.A1(n_883),
.A2(n_875),
.B1(n_836),
.B2(n_828),
.C(n_853),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_892),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_907),
.B(n_891),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_907),
.B(n_891),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_916),
.Y(n_923)
);

OR2x2_ASAP7_75t_L g924 ( 
.A(n_913),
.B(n_883),
.Y(n_924)
);

INVx4_ASAP7_75t_L g925 ( 
.A(n_911),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_920),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_918),
.B(n_885),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_911),
.B(n_909),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_906),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_906),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_911),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_928),
.B(n_911),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_926),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_923),
.B(n_912),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_925),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_925),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_925),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_931),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_928),
.B(n_910),
.Y(n_939)
);

AO221x2_ASAP7_75t_L g940 ( 
.A1(n_934),
.A2(n_836),
.B1(n_931),
.B2(n_929),
.C(n_930),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_933),
.Y(n_941)
);

AO221x2_ASAP7_75t_L g942 ( 
.A1(n_936),
.A2(n_853),
.B1(n_908),
.B2(n_845),
.C(n_905),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_939),
.B(n_936),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_938),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_932),
.A2(n_919),
.B1(n_865),
.B2(n_854),
.Y(n_945)
);

NAND2x1p5_ASAP7_75t_L g946 ( 
.A(n_944),
.B(n_935),
.Y(n_946)
);

AOI33xp33_ASAP7_75t_L g947 ( 
.A1(n_945),
.A2(n_935),
.A3(n_937),
.B1(n_932),
.B2(n_763),
.B3(n_922),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_943),
.B(n_937),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_941),
.Y(n_949)
);

AOI22xp33_ASAP7_75t_SL g950 ( 
.A1(n_940),
.A2(n_865),
.B1(n_854),
.B2(n_893),
.Y(n_950)
);

NAND2x1p5_ASAP7_75t_L g951 ( 
.A(n_942),
.B(n_847),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_944),
.Y(n_952)
);

OR2x2_ASAP7_75t_L g953 ( 
.A(n_943),
.B(n_938),
.Y(n_953)
);

NOR2x1p5_ASAP7_75t_L g954 ( 
.A(n_943),
.B(n_938),
.Y(n_954)
);

INVx2_ASAP7_75t_SL g955 ( 
.A(n_940),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_950),
.A2(n_927),
.B(n_846),
.Y(n_956)
);

OR2x2_ASAP7_75t_L g957 ( 
.A(n_953),
.B(n_924),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_946),
.Y(n_958)
);

OAI221xp5_ASAP7_75t_L g959 ( 
.A1(n_955),
.A2(n_900),
.B1(n_829),
.B2(n_885),
.C(n_921),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_948),
.B(n_921),
.Y(n_960)
);

AOI221x1_ASAP7_75t_L g961 ( 
.A1(n_952),
.A2(n_922),
.B1(n_915),
.B2(n_914),
.C(n_894),
.Y(n_961)
);

AOI21xp33_ASAP7_75t_L g962 ( 
.A1(n_949),
.A2(n_865),
.B(n_854),
.Y(n_962)
);

HB1xp67_ASAP7_75t_L g963 ( 
.A(n_954),
.Y(n_963)
);

OR2x2_ASAP7_75t_L g964 ( 
.A(n_957),
.B(n_952),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_960),
.Y(n_965)
);

NOR3xp33_ASAP7_75t_L g966 ( 
.A(n_958),
.B(n_947),
.C(n_814),
.Y(n_966)
);

AOI221xp5_ASAP7_75t_L g967 ( 
.A1(n_962),
.A2(n_963),
.B1(n_956),
.B2(n_959),
.C(n_951),
.Y(n_967)
);

OAI31xp33_ASAP7_75t_SL g968 ( 
.A1(n_961),
.A2(n_890),
.A3(n_894),
.B(n_845),
.Y(n_968)
);

OA21x2_ASAP7_75t_L g969 ( 
.A1(n_961),
.A2(n_915),
.B(n_914),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_959),
.A2(n_900),
.B1(n_882),
.B2(n_917),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_963),
.B(n_899),
.Y(n_971)
);

NAND4xp25_ASAP7_75t_L g972 ( 
.A(n_966),
.B(n_850),
.C(n_772),
.D(n_867),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_964),
.B(n_899),
.Y(n_973)
);

AOI221xp5_ASAP7_75t_L g974 ( 
.A1(n_967),
.A2(n_882),
.B1(n_843),
.B2(n_787),
.C(n_817),
.Y(n_974)
);

AOI21xp33_ASAP7_75t_L g975 ( 
.A1(n_965),
.A2(n_786),
.B(n_835),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_971),
.B(n_896),
.Y(n_976)
);

OAI322xp33_ASAP7_75t_L g977 ( 
.A1(n_970),
.A2(n_827),
.A3(n_903),
.B1(n_897),
.B2(n_892),
.C1(n_841),
.C2(n_904),
.Y(n_977)
);

BUFx3_ASAP7_75t_L g978 ( 
.A(n_973),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_976),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_972),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_977),
.Y(n_981)
);

INVx1_ASAP7_75t_SL g982 ( 
.A(n_975),
.Y(n_982)
);

INVxp67_ASAP7_75t_L g983 ( 
.A(n_974),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_976),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_973),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_973),
.Y(n_986)
);

NAND3xp33_ASAP7_75t_L g987 ( 
.A(n_980),
.B(n_968),
.C(n_969),
.Y(n_987)
);

NOR2x1_ASAP7_75t_L g988 ( 
.A(n_978),
.B(n_969),
.Y(n_988)
);

NOR2x1p5_ASAP7_75t_L g989 ( 
.A(n_984),
.B(n_867),
.Y(n_989)
);

INVxp67_ASAP7_75t_L g990 ( 
.A(n_980),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_L g991 ( 
.A1(n_982),
.A2(n_867),
.B1(n_881),
.B2(n_863),
.Y(n_991)
);

NAND4xp25_ASAP7_75t_L g992 ( 
.A(n_979),
.B(n_768),
.C(n_881),
.D(n_790),
.Y(n_992)
);

OAI211xp5_ASAP7_75t_L g993 ( 
.A1(n_983),
.A2(n_881),
.B(n_849),
.C(n_841),
.Y(n_993)
);

NOR3x1_ASAP7_75t_L g994 ( 
.A(n_981),
.B(n_851),
.C(n_821),
.Y(n_994)
);

AO22x2_ASAP7_75t_L g995 ( 
.A1(n_986),
.A2(n_881),
.B1(n_903),
.B2(n_897),
.Y(n_995)
);

NAND2xp33_ASAP7_75t_L g996 ( 
.A(n_988),
.B(n_985),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_989),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_SL g998 ( 
.A(n_990),
.B(n_983),
.Y(n_998)
);

NOR4xp75_ASAP7_75t_L g999 ( 
.A(n_987),
.B(n_994),
.C(n_993),
.D(n_991),
.Y(n_999)
);

OAI221xp5_ASAP7_75t_L g1000 ( 
.A1(n_992),
.A2(n_849),
.B1(n_881),
.B2(n_834),
.C(n_835),
.Y(n_1000)
);

NAND4xp25_ASAP7_75t_L g1001 ( 
.A(n_995),
.B(n_834),
.C(n_873),
.D(n_832),
.Y(n_1001)
);

OAI221xp5_ASAP7_75t_L g1002 ( 
.A1(n_988),
.A2(n_849),
.B1(n_870),
.B2(n_821),
.C(n_832),
.Y(n_1002)
);

AND4x2_ASAP7_75t_L g1003 ( 
.A(n_999),
.B(n_893),
.C(n_849),
.D(n_863),
.Y(n_1003)
);

NAND4xp25_ASAP7_75t_L g1004 ( 
.A(n_998),
.B(n_1002),
.C(n_1000),
.D(n_1001),
.Y(n_1004)
);

NAND2x1p5_ASAP7_75t_L g1005 ( 
.A(n_997),
.B(n_849),
.Y(n_1005)
);

NOR2x1_ASAP7_75t_L g1006 ( 
.A(n_996),
.B(n_869),
.Y(n_1006)
);

NOR2x1_ASAP7_75t_L g1007 ( 
.A(n_996),
.B(n_869),
.Y(n_1007)
);

INVxp33_ASAP7_75t_SL g1008 ( 
.A(n_998),
.Y(n_1008)
);

NAND5xp2_ASAP7_75t_L g1009 ( 
.A(n_998),
.B(n_873),
.C(n_844),
.D(n_904),
.E(n_896),
.Y(n_1009)
);

OAI21xp33_ASAP7_75t_L g1010 ( 
.A1(n_998),
.A2(n_873),
.B(n_870),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_998),
.B(n_842),
.Y(n_1011)
);

OAI221xp5_ASAP7_75t_SL g1012 ( 
.A1(n_1002),
.A2(n_870),
.B1(n_842),
.B2(n_839),
.C(n_889),
.Y(n_1012)
);

AOI321xp33_ASAP7_75t_L g1013 ( 
.A1(n_1011),
.A2(n_842),
.A3(n_852),
.B1(n_839),
.B2(n_826),
.C(n_824),
.Y(n_1013)
);

NOR2xp67_ASAP7_75t_L g1014 ( 
.A(n_1004),
.B(n_141),
.Y(n_1014)
);

AOI32xp33_ASAP7_75t_L g1015 ( 
.A1(n_1006),
.A2(n_1007),
.A3(n_1010),
.B1(n_1003),
.B2(n_1008),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_1005),
.B(n_852),
.Y(n_1016)
);

NOR3xp33_ASAP7_75t_L g1017 ( 
.A(n_1012),
.B(n_851),
.C(n_880),
.Y(n_1017)
);

NAND3xp33_ASAP7_75t_SL g1018 ( 
.A(n_1009),
.B(n_844),
.C(n_889),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_SL g1019 ( 
.A1(n_1008),
.A2(n_870),
.B1(n_839),
.B2(n_852),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_1008),
.B(n_884),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_1005),
.Y(n_1021)
);

NOR2x1_ASAP7_75t_L g1022 ( 
.A(n_1014),
.B(n_839),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_1015),
.B(n_884),
.Y(n_1023)
);

OR3x2_ASAP7_75t_L g1024 ( 
.A(n_1020),
.B(n_143),
.C(n_145),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1016),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1018),
.Y(n_1026)
);

NOR3xp33_ASAP7_75t_SL g1027 ( 
.A(n_1019),
.B(n_1017),
.C(n_1013),
.Y(n_1027)
);

INVx4_ASAP7_75t_L g1028 ( 
.A(n_1021),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_1028),
.B(n_878),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1022),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_1023),
.A2(n_878),
.B(n_837),
.Y(n_1031)
);

AOI22x1_ASAP7_75t_L g1032 ( 
.A1(n_1026),
.A2(n_147),
.B1(n_149),
.B2(n_150),
.Y(n_1032)
);

AOI221xp5_ASAP7_75t_L g1033 ( 
.A1(n_1027),
.A2(n_858),
.B1(n_857),
.B2(n_816),
.C(n_815),
.Y(n_1033)
);

AND2x2_ASAP7_75t_SL g1034 ( 
.A(n_1025),
.B(n_151),
.Y(n_1034)
);

NOR3xp33_ASAP7_75t_L g1035 ( 
.A(n_1024),
.B(n_152),
.C(n_154),
.Y(n_1035)
);

AOI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_1035),
.A2(n_1029),
.B1(n_1033),
.B2(n_1031),
.Y(n_1036)
);

INVxp67_ASAP7_75t_L g1037 ( 
.A(n_1034),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1032),
.Y(n_1038)
);

AO22x2_ASAP7_75t_L g1039 ( 
.A1(n_1030),
.A2(n_872),
.B1(n_874),
.B2(n_858),
.Y(n_1039)
);

OAI22x1_ASAP7_75t_L g1040 ( 
.A1(n_1038),
.A2(n_874),
.B1(n_816),
.B2(n_825),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_1037),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1041),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1042),
.B(n_1036),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1043),
.Y(n_1044)
);

AO22x2_ASAP7_75t_L g1045 ( 
.A1(n_1044),
.A2(n_1040),
.B1(n_1039),
.B2(n_156),
.Y(n_1045)
);

XNOR2xp5_ASAP7_75t_L g1046 ( 
.A(n_1045),
.B(n_157),
.Y(n_1046)
);

OAI31xp33_ASAP7_75t_SL g1047 ( 
.A1(n_1046),
.A2(n_158),
.A3(n_159),
.B(n_160),
.Y(n_1047)
);

AOI221xp5_ASAP7_75t_L g1048 ( 
.A1(n_1047),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.C(n_164),
.Y(n_1048)
);

AOI211xp5_ASAP7_75t_L g1049 ( 
.A1(n_1048),
.A2(n_165),
.B(n_167),
.C(n_170),
.Y(n_1049)
);


endmodule