module fake_netlist_6_3134_n_1013 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1013);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1013;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_760;
wire n_741;
wire n_1008;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1009;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_222;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_795;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_886;
wire n_448;
wire n_953;
wire n_844;
wire n_1004;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_998;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_928;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_722;
wire n_688;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_25),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_62),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_149),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_94),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_70),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_3),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_55),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_106),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_98),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_124),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_161),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_66),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_155),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_31),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_119),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_173),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_30),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_150),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_2),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_24),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_177),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_63),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_60),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_10),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_78),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_158),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_146),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_185),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_88),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_180),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_189),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_118),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_44),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_90),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_190),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_145),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_100),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_157),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_76),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_203),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_11),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_89),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_52),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_164),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_84),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_201),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_12),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_49),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_82),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_132),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_64),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_14),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_196),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_11),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_39),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_97),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_24),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_40),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_95),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_125),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_176),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_35),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_102),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_103),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_85),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_23),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_16),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_122),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_198),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_53),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_199),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_156),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_80),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_48),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_16),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_151),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_73),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_17),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_105),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_152),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_61),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_282),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_244),
.B(n_0),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_282),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_206),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_208),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_270),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_210),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_209),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_270),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_270),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_215),
.B(n_0),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_270),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_213),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_261),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_214),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_239),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_223),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_218),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_271),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_204),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_224),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_228),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_219),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_251),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_256),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_220),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_222),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_211),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_211),
.Y(n_314)
);

INVxp33_ASAP7_75t_SL g315 ( 
.A(n_258),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_235),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_235),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_274),
.Y(n_318)
);

INVxp33_ASAP7_75t_SL g319 ( 
.A(n_279),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_226),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_273),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_205),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_207),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_272),
.B(n_1),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_245),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_229),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_227),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_216),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_221),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_225),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_272),
.B(n_1),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_231),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_237),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_278),
.B(n_2),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_273),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_230),
.Y(n_336)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_243),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_238),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_249),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_295),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_327),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_327),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_306),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_295),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_291),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_294),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_297),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_313),
.B(n_212),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_302),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_307),
.Y(n_350)
);

NAND2xp33_ASAP7_75t_SL g351 ( 
.A(n_324),
.B(n_250),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_289),
.B(n_217),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_290),
.B(n_217),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_310),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_314),
.Y(n_355)
);

AND2x4_ASAP7_75t_L g356 ( 
.A(n_331),
.B(n_248),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_321),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_293),
.B(n_248),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_322),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_328),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_330),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_336),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_338),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_301),
.B(n_233),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_316),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_317),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_286),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_288),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_298),
.B(n_253),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_300),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_296),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_318),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_334),
.Y(n_373)
);

AND2x4_ASAP7_75t_L g374 ( 
.A(n_287),
.B(n_253),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_325),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_321),
.B(n_281),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_305),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_323),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_303),
.B(n_281),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_306),
.A2(n_252),
.B1(n_236),
.B2(n_283),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_308),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_311),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_315),
.B(n_242),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_312),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_320),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_326),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_315),
.A2(n_319),
.B1(n_309),
.B2(n_335),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_319),
.B(n_227),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_332),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_337),
.B(n_234),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_309),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_323),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_329),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_329),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_333),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_333),
.B(n_246),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_360),
.Y(n_397)
);

OR2x2_ASAP7_75t_L g398 ( 
.A(n_375),
.B(n_255),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_360),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_361),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_344),
.Y(n_401)
);

NOR2x1p5_ASAP7_75t_L g402 ( 
.A(n_370),
.B(n_240),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_344),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_L g404 ( 
.A1(n_374),
.A2(n_285),
.B1(n_275),
.B2(n_268),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_361),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_356),
.B(n_264),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_355),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_349),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_363),
.Y(n_409)
);

INVx6_ASAP7_75t_L g410 ( 
.A(n_356),
.Y(n_410)
);

NAND2xp33_ASAP7_75t_L g411 ( 
.A(n_373),
.B(n_227),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_357),
.Y(n_412)
);

AND2x6_ASAP7_75t_L g413 ( 
.A(n_374),
.B(n_227),
.Y(n_413)
);

AND2x2_ASAP7_75t_SL g414 ( 
.A(n_374),
.B(n_232),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_356),
.B(n_276),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_355),
.B(n_241),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_363),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_344),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_378),
.Y(n_419)
);

INVx5_ASAP7_75t_L g420 ( 
.A(n_344),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_344),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_352),
.B(n_247),
.Y(n_422)
);

BUFx6f_ASAP7_75t_SL g423 ( 
.A(n_392),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_367),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_343),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_367),
.Y(n_426)
);

OAI22x1_ASAP7_75t_L g427 ( 
.A1(n_387),
.A2(n_304),
.B1(n_299),
.B2(n_292),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_341),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_341),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_L g430 ( 
.A1(n_374),
.A2(n_232),
.B1(n_263),
.B2(n_266),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_343),
.Y(n_431)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_370),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_392),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_349),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_L g435 ( 
.A1(n_373),
.A2(n_232),
.B1(n_263),
.B2(n_267),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_341),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_350),
.Y(n_437)
);

INVx4_ASAP7_75t_L g438 ( 
.A(n_356),
.Y(n_438)
);

AOI22xp33_ASAP7_75t_L g439 ( 
.A1(n_371),
.A2(n_232),
.B1(n_263),
.B2(n_265),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_371),
.B(n_340),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_340),
.B(n_263),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_372),
.B(n_254),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_382),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_392),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_372),
.B(n_257),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_342),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_350),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_342),
.Y(n_448)
);

INVx2_ASAP7_75t_SL g449 ( 
.A(n_377),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_375),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_354),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_348),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_348),
.B(n_259),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_354),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_365),
.Y(n_455)
);

BUFx10_ASAP7_75t_L g456 ( 
.A(n_396),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_342),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_365),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_353),
.B(n_260),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_366),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_366),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_359),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_347),
.B(n_262),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_383),
.A2(n_284),
.B1(n_277),
.B2(n_280),
.Y(n_464)
);

BUFx10_ASAP7_75t_L g465 ( 
.A(n_396),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_347),
.B(n_345),
.Y(n_466)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_376),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_345),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_346),
.B(n_269),
.Y(n_469)
);

NAND2xp33_ASAP7_75t_SL g470 ( 
.A(n_380),
.B(n_339),
.Y(n_470)
);

A2O1A1Ixp33_ASAP7_75t_L g471 ( 
.A1(n_430),
.A2(n_351),
.B(n_379),
.C(n_358),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_410),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_450),
.Y(n_473)
);

AO22x2_ASAP7_75t_L g474 ( 
.A1(n_433),
.A2(n_396),
.B1(n_395),
.B2(n_394),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_452),
.Y(n_475)
);

AO22x2_ASAP7_75t_L g476 ( 
.A1(n_425),
.A2(n_396),
.B1(n_395),
.B2(n_394),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_408),
.B(n_390),
.Y(n_477)
);

OAI221xp5_ASAP7_75t_L g478 ( 
.A1(n_404),
.A2(n_369),
.B1(n_388),
.B2(n_368),
.C(n_362),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_436),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_414),
.B(n_381),
.Y(n_480)
);

AO22x2_ASAP7_75t_L g481 ( 
.A1(n_431),
.A2(n_391),
.B1(n_393),
.B2(n_364),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_407),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_410),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_436),
.Y(n_484)
);

NAND2x1p5_ASAP7_75t_L g485 ( 
.A(n_432),
.B(n_381),
.Y(n_485)
);

AO22x2_ASAP7_75t_L g486 ( 
.A1(n_449),
.A2(n_391),
.B1(n_393),
.B2(n_385),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_410),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_414),
.B(n_384),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_422),
.B(n_438),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_424),
.Y(n_490)
);

BUFx8_ASAP7_75t_L g491 ( 
.A(n_419),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_430),
.A2(n_384),
.B1(n_386),
.B2(n_389),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_426),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_446),
.Y(n_494)
);

NAND2x1p5_ASAP7_75t_L g495 ( 
.A(n_432),
.B(n_467),
.Y(n_495)
);

BUFx8_ASAP7_75t_L g496 ( 
.A(n_423),
.Y(n_496)
);

AO22x2_ASAP7_75t_L g497 ( 
.A1(n_398),
.A2(n_385),
.B1(n_376),
.B2(n_386),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_397),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_399),
.B(n_389),
.Y(n_499)
);

AO22x2_ASAP7_75t_L g500 ( 
.A1(n_412),
.A2(n_376),
.B1(n_390),
.B2(n_304),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_438),
.B(n_376),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_446),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_422),
.B(n_359),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_462),
.Y(n_504)
);

AO22x2_ASAP7_75t_L g505 ( 
.A1(n_470),
.A2(n_292),
.B1(n_299),
.B2(n_368),
.Y(n_505)
);

AO22x2_ASAP7_75t_L g506 ( 
.A1(n_408),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_400),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_405),
.B(n_362),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_442),
.B(n_392),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_409),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_417),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_434),
.B(n_392),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_467),
.B(n_346),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_444),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_423),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_437),
.Y(n_516)
);

NAND2xp33_ASAP7_75t_L g517 ( 
.A(n_413),
.B(n_435),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_462),
.Y(n_518)
);

NAND2xp33_ASAP7_75t_L g519 ( 
.A(n_413),
.B(n_339),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_447),
.Y(n_520)
);

NOR2xp67_ASAP7_75t_L g521 ( 
.A(n_443),
.B(n_202),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_451),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_404),
.B(n_29),
.Y(n_523)
);

INVx5_ASAP7_75t_L g524 ( 
.A(n_413),
.Y(n_524)
);

NOR2x2_ASAP7_75t_L g525 ( 
.A(n_427),
.B(n_4),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_454),
.Y(n_526)
);

AO22x2_ASAP7_75t_L g527 ( 
.A1(n_453),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_428),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_466),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_440),
.B(n_32),
.Y(n_530)
);

BUFx8_ASAP7_75t_L g531 ( 
.A(n_416),
.Y(n_531)
);

AO22x2_ASAP7_75t_L g532 ( 
.A1(n_459),
.A2(n_406),
.B1(n_415),
.B2(n_445),
.Y(n_532)
);

NAND2x1p5_ASAP7_75t_L g533 ( 
.A(n_458),
.B(n_33),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_440),
.B(n_34),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_466),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_455),
.Y(n_536)
);

NAND3xp33_ASAP7_75t_L g537 ( 
.A(n_464),
.B(n_6),
.C(n_7),
.Y(n_537)
);

AO22x2_ASAP7_75t_L g538 ( 
.A1(n_459),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_538)
);

AO22x2_ASAP7_75t_L g539 ( 
.A1(n_406),
.A2(n_8),
.B1(n_9),
.B2(n_12),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_429),
.Y(n_540)
);

AND2x6_ASAP7_75t_L g541 ( 
.A(n_415),
.B(n_401),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_442),
.B(n_13),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_460),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_445),
.A2(n_114),
.B1(n_197),
.B2(n_195),
.Y(n_544)
);

NAND2x1p5_ASAP7_75t_L g545 ( 
.A(n_458),
.B(n_36),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_461),
.Y(n_546)
);

AO22x2_ASAP7_75t_L g547 ( 
.A1(n_435),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_547)
);

AO22x2_ASAP7_75t_L g548 ( 
.A1(n_416),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_458),
.B(n_37),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_439),
.B(n_38),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_439),
.B(n_41),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_464),
.A2(n_117),
.B1(n_194),
.B2(n_193),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_468),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_448),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_477),
.B(n_456),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_509),
.B(n_456),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_492),
.B(n_465),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_SL g558 ( 
.A(n_515),
.B(n_402),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_499),
.B(n_465),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_529),
.B(n_469),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_499),
.B(n_469),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_535),
.B(n_463),
.Y(n_562)
);

NAND2xp33_ASAP7_75t_SL g563 ( 
.A(n_514),
.B(n_463),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_480),
.B(n_418),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_488),
.B(n_521),
.Y(n_565)
);

XNOR2x2_ASAP7_75t_L g566 ( 
.A(n_548),
.B(n_18),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_512),
.B(n_418),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_485),
.B(n_418),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_503),
.B(n_421),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_475),
.B(n_421),
.Y(n_570)
);

NAND2xp33_ASAP7_75t_SL g571 ( 
.A(n_523),
.B(n_403),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_542),
.B(n_421),
.Y(n_572)
);

NAND2xp33_ASAP7_75t_SL g573 ( 
.A(n_550),
.B(n_441),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_473),
.B(n_457),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_471),
.B(n_420),
.Y(n_575)
);

NAND2xp33_ASAP7_75t_SL g576 ( 
.A(n_551),
.B(n_441),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_489),
.B(n_420),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_490),
.B(n_413),
.Y(n_578)
);

NAND2xp33_ASAP7_75t_SL g579 ( 
.A(n_493),
.B(n_411),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_498),
.B(n_413),
.Y(n_580)
);

NAND2xp33_ASAP7_75t_SL g581 ( 
.A(n_507),
.B(n_19),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_553),
.B(n_420),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_508),
.B(n_420),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_482),
.B(n_42),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_508),
.B(n_43),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_524),
.B(n_45),
.Y(n_586)
);

NAND2xp33_ASAP7_75t_SL g587 ( 
.A(n_510),
.B(n_19),
.Y(n_587)
);

NAND2xp33_ASAP7_75t_SL g588 ( 
.A(n_511),
.B(n_20),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_524),
.B(n_46),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_524),
.B(n_47),
.Y(n_590)
);

NAND2xp33_ASAP7_75t_SL g591 ( 
.A(n_516),
.B(n_20),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_495),
.B(n_50),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_520),
.B(n_51),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_522),
.B(n_54),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_526),
.B(n_56),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_536),
.B(n_21),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_472),
.B(n_57),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_543),
.B(n_21),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_546),
.B(n_22),
.Y(n_599)
);

NAND2xp33_ASAP7_75t_SL g600 ( 
.A(n_530),
.B(n_22),
.Y(n_600)
);

AND2x2_ASAP7_75t_SL g601 ( 
.A(n_517),
.B(n_58),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_483),
.B(n_59),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_487),
.B(n_65),
.Y(n_603)
);

AND2x4_ASAP7_75t_SL g604 ( 
.A(n_479),
.B(n_484),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_500),
.B(n_23),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_SL g606 ( 
.A(n_534),
.B(n_25),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_504),
.B(n_67),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_518),
.B(n_68),
.Y(n_608)
);

NAND2xp33_ASAP7_75t_SL g609 ( 
.A(n_501),
.B(n_26),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_532),
.B(n_26),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_532),
.B(n_27),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_513),
.B(n_69),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_494),
.B(n_71),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_497),
.B(n_27),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_502),
.B(n_72),
.Y(n_615)
);

NAND2xp33_ASAP7_75t_SL g616 ( 
.A(n_549),
.B(n_28),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_537),
.B(n_74),
.Y(n_617)
);

NAND2xp33_ASAP7_75t_SL g618 ( 
.A(n_496),
.B(n_28),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_554),
.B(n_75),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_552),
.B(n_77),
.Y(n_620)
);

AO31x2_ASAP7_75t_L g621 ( 
.A1(n_610),
.A2(n_528),
.A3(n_540),
.B(n_497),
.Y(n_621)
);

OAI21xp33_ASAP7_75t_L g622 ( 
.A1(n_560),
.A2(n_547),
.B(n_527),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_584),
.Y(n_623)
);

AO31x2_ASAP7_75t_L g624 ( 
.A1(n_611),
.A2(n_541),
.A3(n_474),
.B(n_476),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_565),
.A2(n_519),
.B(n_478),
.Y(n_625)
);

OAI21x1_ASAP7_75t_L g626 ( 
.A1(n_575),
.A2(n_564),
.B(n_569),
.Y(n_626)
);

BUFx10_ASAP7_75t_L g627 ( 
.A(n_584),
.Y(n_627)
);

CKINVDCx16_ASAP7_75t_R g628 ( 
.A(n_558),
.Y(n_628)
);

OA21x2_ASAP7_75t_L g629 ( 
.A1(n_577),
.A2(n_544),
.B(n_541),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_562),
.A2(n_533),
.B(n_545),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_561),
.B(n_531),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_595),
.B(n_474),
.Y(n_632)
);

BUFx2_ASAP7_75t_L g633 ( 
.A(n_595),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_573),
.A2(n_576),
.B(n_620),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_601),
.Y(n_635)
);

INVxp67_ASAP7_75t_SL g636 ( 
.A(n_567),
.Y(n_636)
);

OAI21x1_ASAP7_75t_L g637 ( 
.A1(n_578),
.A2(n_541),
.B(n_476),
.Y(n_637)
);

OAI21x1_ASAP7_75t_L g638 ( 
.A1(n_580),
.A2(n_486),
.B(n_500),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_563),
.B(n_491),
.Y(n_639)
);

AO21x1_ASAP7_75t_L g640 ( 
.A1(n_557),
.A2(n_538),
.B(n_547),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_601),
.Y(n_641)
);

NAND3xp33_ASAP7_75t_L g642 ( 
.A(n_581),
.B(n_525),
.C(n_481),
.Y(n_642)
);

AOI21xp33_ASAP7_75t_L g643 ( 
.A1(n_555),
.A2(n_481),
.B(n_486),
.Y(n_643)
);

OAI21x1_ASAP7_75t_L g644 ( 
.A1(n_583),
.A2(n_79),
.B(n_81),
.Y(n_644)
);

OAI21x1_ASAP7_75t_L g645 ( 
.A1(n_612),
.A2(n_83),
.B(n_86),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_574),
.B(n_505),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_571),
.A2(n_548),
.B(n_538),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_596),
.B(n_527),
.Y(n_648)
);

OAI21x1_ASAP7_75t_L g649 ( 
.A1(n_592),
.A2(n_87),
.B(n_91),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_559),
.B(n_505),
.Y(n_650)
);

NAND3xp33_ASAP7_75t_L g651 ( 
.A(n_587),
.B(n_506),
.C(n_539),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_568),
.A2(n_539),
.B(n_506),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_613),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_613),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_598),
.B(n_200),
.Y(n_655)
);

AO31x2_ASAP7_75t_L g656 ( 
.A1(n_614),
.A2(n_92),
.A3(n_93),
.B(n_96),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_616),
.Y(n_657)
);

OAI21xp5_ASAP7_75t_L g658 ( 
.A1(n_617),
.A2(n_99),
.B(n_101),
.Y(n_658)
);

NAND2x1_ASAP7_75t_L g659 ( 
.A(n_599),
.B(n_104),
.Y(n_659)
);

BUFx12f_ASAP7_75t_L g660 ( 
.A(n_605),
.Y(n_660)
);

OAI21x1_ASAP7_75t_L g661 ( 
.A1(n_572),
.A2(n_107),
.B(n_108),
.Y(n_661)
);

AO21x1_ASAP7_75t_L g662 ( 
.A1(n_609),
.A2(n_109),
.B(n_110),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_556),
.B(n_111),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_L g664 ( 
.A1(n_585),
.A2(n_112),
.B1(n_113),
.B2(n_115),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_570),
.B(n_116),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_604),
.B(n_120),
.Y(n_666)
);

OAI21x1_ASAP7_75t_SL g667 ( 
.A1(n_566),
.A2(n_121),
.B(n_123),
.Y(n_667)
);

INVx4_ASAP7_75t_SL g668 ( 
.A(n_618),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_582),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_579),
.B(n_126),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_615),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_593),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_594),
.B(n_192),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_607),
.Y(n_674)
);

INVx4_ASAP7_75t_L g675 ( 
.A(n_588),
.Y(n_675)
);

OAI21x1_ASAP7_75t_L g676 ( 
.A1(n_626),
.A2(n_619),
.B(n_608),
.Y(n_676)
);

INVxp67_ASAP7_75t_SL g677 ( 
.A(n_654),
.Y(n_677)
);

OAI21x1_ASAP7_75t_L g678 ( 
.A1(n_634),
.A2(n_597),
.B(n_603),
.Y(n_678)
);

OAI21x1_ASAP7_75t_L g679 ( 
.A1(n_637),
.A2(n_602),
.B(n_590),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_644),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_636),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_675),
.B(n_635),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_653),
.Y(n_683)
);

AOI21xp33_ASAP7_75t_L g684 ( 
.A1(n_648),
.A2(n_589),
.B(n_586),
.Y(n_684)
);

OAI21x1_ASAP7_75t_L g685 ( 
.A1(n_661),
.A2(n_606),
.B(n_600),
.Y(n_685)
);

OAI21x1_ASAP7_75t_L g686 ( 
.A1(n_625),
.A2(n_591),
.B(n_128),
.Y(n_686)
);

OAI221xp5_ASAP7_75t_L g687 ( 
.A1(n_642),
.A2(n_127),
.B1(n_129),
.B2(n_130),
.C(n_131),
.Y(n_687)
);

OA21x2_ASAP7_75t_L g688 ( 
.A1(n_635),
.A2(n_133),
.B(n_134),
.Y(n_688)
);

OAI21x1_ASAP7_75t_L g689 ( 
.A1(n_645),
.A2(n_135),
.B(n_136),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_653),
.Y(n_690)
);

BUFx12f_ASAP7_75t_L g691 ( 
.A(n_660),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_628),
.Y(n_692)
);

OAI21xp5_ASAP7_75t_L g693 ( 
.A1(n_630),
.A2(n_137),
.B(n_138),
.Y(n_693)
);

OAI21x1_ASAP7_75t_SL g694 ( 
.A1(n_640),
.A2(n_139),
.B(n_140),
.Y(n_694)
);

A2O1A1Ixp33_ASAP7_75t_L g695 ( 
.A1(n_622),
.A2(n_647),
.B(n_670),
.C(n_651),
.Y(n_695)
);

OAI21xp5_ASAP7_75t_L g696 ( 
.A1(n_655),
.A2(n_638),
.B(n_672),
.Y(n_696)
);

OAI21x1_ASAP7_75t_L g697 ( 
.A1(n_649),
.A2(n_141),
.B(n_142),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_SL g698 ( 
.A1(n_675),
.A2(n_143),
.B1(n_144),
.B2(n_147),
.Y(n_698)
);

NAND2x1p5_ASAP7_75t_L g699 ( 
.A(n_654),
.B(n_148),
.Y(n_699)
);

OAI21x1_ASAP7_75t_L g700 ( 
.A1(n_659),
.A2(n_153),
.B(n_154),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_633),
.B(n_160),
.Y(n_701)
);

OAI21xp5_ASAP7_75t_L g702 ( 
.A1(n_641),
.A2(n_162),
.B(n_163),
.Y(n_702)
);

OAI21x1_ASAP7_75t_L g703 ( 
.A1(n_629),
.A2(n_165),
.B(n_166),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_623),
.B(n_666),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_657),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_641),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_SL g707 ( 
.A1(n_628),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_707)
);

OAI21xp5_ASAP7_75t_L g708 ( 
.A1(n_663),
.A2(n_174),
.B(n_175),
.Y(n_708)
);

OAI21xp5_ASAP7_75t_L g709 ( 
.A1(n_658),
.A2(n_178),
.B(n_179),
.Y(n_709)
);

OAI21x1_ASAP7_75t_L g710 ( 
.A1(n_629),
.A2(n_181),
.B(n_182),
.Y(n_710)
);

OAI21xp5_ASAP7_75t_L g711 ( 
.A1(n_652),
.A2(n_183),
.B(n_184),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_646),
.Y(n_712)
);

BUFx8_ASAP7_75t_SL g713 ( 
.A(n_666),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_627),
.B(n_186),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_L g715 ( 
.A1(n_632),
.A2(n_187),
.B1(n_188),
.B2(n_191),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_621),
.Y(n_716)
);

BUFx2_ASAP7_75t_L g717 ( 
.A(n_668),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_669),
.B(n_639),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_621),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_SL g720 ( 
.A1(n_667),
.A2(n_631),
.B1(n_650),
.B2(n_627),
.Y(n_720)
);

HB1xp67_ASAP7_75t_L g721 ( 
.A(n_624),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_621),
.Y(n_722)
);

OAI21x1_ASAP7_75t_L g723 ( 
.A1(n_673),
.A2(n_674),
.B(n_671),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_665),
.Y(n_724)
);

OA21x2_ASAP7_75t_L g725 ( 
.A1(n_622),
.A2(n_662),
.B(n_643),
.Y(n_725)
);

OAI22xp5_ASAP7_75t_L g726 ( 
.A1(n_664),
.A2(n_624),
.B1(n_668),
.B2(n_656),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_624),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_716),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_704),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_716),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_717),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_719),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_719),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_713),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_722),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_722),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_727),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_727),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_695),
.B(n_656),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_721),
.Y(n_740)
);

INVxp67_ASAP7_75t_SL g741 ( 
.A(n_681),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_683),
.Y(n_742)
);

BUFx4f_ASAP7_75t_SL g743 ( 
.A(n_691),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_712),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_690),
.Y(n_745)
);

BUFx4f_ASAP7_75t_SL g746 ( 
.A(n_691),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_692),
.Y(n_747)
);

OAI21x1_ASAP7_75t_L g748 ( 
.A1(n_703),
.A2(n_656),
.B(n_710),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_723),
.Y(n_749)
);

INVx4_ASAP7_75t_L g750 ( 
.A(n_718),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_725),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_725),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_713),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_725),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_723),
.Y(n_755)
);

OAI21x1_ASAP7_75t_L g756 ( 
.A1(n_703),
.A2(n_710),
.B(n_676),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_686),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_686),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_688),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_724),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_689),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_695),
.B(n_726),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_724),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_696),
.B(n_682),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_688),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_680),
.Y(n_766)
);

INVx4_ASAP7_75t_SL g767 ( 
.A(n_724),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_688),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_685),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_685),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_689),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_680),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_697),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_682),
.B(n_718),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_704),
.B(n_718),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_700),
.Y(n_776)
);

INVx4_ASAP7_75t_L g777 ( 
.A(n_724),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_697),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_720),
.A2(n_692),
.B1(n_704),
.B2(n_711),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_700),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_679),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_679),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_676),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_678),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_701),
.B(n_677),
.Y(n_785)
);

INVxp67_ASAP7_75t_SL g786 ( 
.A(n_699),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_705),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_699),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_767),
.B(n_714),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_745),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_774),
.B(n_707),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_764),
.B(n_684),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_774),
.B(n_702),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_744),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_747),
.Y(n_795)
);

CKINVDCx20_ASAP7_75t_R g796 ( 
.A(n_743),
.Y(n_796)
);

HB1xp67_ASAP7_75t_L g797 ( 
.A(n_744),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_742),
.Y(n_798)
);

AND2x4_ASAP7_75t_L g799 ( 
.A(n_767),
.B(n_693),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_R g800 ( 
.A(n_747),
.B(n_698),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_775),
.B(n_708),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_R g802 ( 
.A(n_746),
.B(n_731),
.Y(n_802)
);

NAND2xp33_ASAP7_75t_R g803 ( 
.A(n_785),
.B(n_709),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_764),
.B(n_694),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_R g805 ( 
.A(n_731),
.B(n_729),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_R g806 ( 
.A(n_729),
.B(n_687),
.Y(n_806)
);

NAND2xp33_ASAP7_75t_R g807 ( 
.A(n_788),
.B(n_739),
.Y(n_807)
);

NAND2xp33_ASAP7_75t_R g808 ( 
.A(n_788),
.B(n_678),
.Y(n_808)
);

BUFx10_ASAP7_75t_L g809 ( 
.A(n_760),
.Y(n_809)
);

INVxp33_ASAP7_75t_L g810 ( 
.A(n_787),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_734),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_742),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_787),
.B(n_715),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_767),
.B(n_706),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_760),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_750),
.B(n_745),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_732),
.Y(n_817)
);

NAND2xp33_ASAP7_75t_R g818 ( 
.A(n_739),
.B(n_762),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_R g819 ( 
.A(n_734),
.B(n_753),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_750),
.B(n_763),
.Y(n_820)
);

XNOR2xp5_ASAP7_75t_L g821 ( 
.A(n_753),
.B(n_779),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_750),
.B(n_760),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_R g823 ( 
.A(n_760),
.B(n_763),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_732),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_R g825 ( 
.A(n_760),
.B(n_763),
.Y(n_825)
);

OR2x6_ASAP7_75t_L g826 ( 
.A(n_762),
.B(n_750),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_763),
.Y(n_827)
);

OR2x4_ASAP7_75t_L g828 ( 
.A(n_763),
.B(n_740),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_777),
.B(n_741),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_777),
.B(n_767),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_740),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_777),
.B(n_786),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_728),
.B(n_730),
.Y(n_833)
);

NAND2xp33_ASAP7_75t_SL g834 ( 
.A(n_777),
.B(n_751),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_R g835 ( 
.A(n_766),
.B(n_772),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_736),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_737),
.B(n_738),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_728),
.B(n_730),
.Y(n_838)
);

INVxp67_ASAP7_75t_L g839 ( 
.A(n_733),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_733),
.Y(n_840)
);

NAND2xp33_ASAP7_75t_R g841 ( 
.A(n_776),
.B(n_780),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_798),
.B(n_752),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_812),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_833),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_792),
.B(n_735),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_828),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_833),
.Y(n_847)
);

INVxp67_ASAP7_75t_SL g848 ( 
.A(n_797),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_838),
.Y(n_849)
);

INVxp67_ASAP7_75t_SL g850 ( 
.A(n_794),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_817),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_824),
.Y(n_852)
);

NOR2xp67_ASAP7_75t_L g853 ( 
.A(n_792),
.B(n_784),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_793),
.B(n_752),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_826),
.Y(n_855)
);

BUFx8_ASAP7_75t_SL g856 ( 
.A(n_796),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_836),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_838),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_816),
.B(n_754),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_794),
.B(n_801),
.Y(n_860)
);

INVxp67_ASAP7_75t_SL g861 ( 
.A(n_808),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_829),
.B(n_735),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_831),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_839),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_790),
.B(n_737),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_826),
.B(n_839),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_840),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_840),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_821),
.B(n_780),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_826),
.B(n_751),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_828),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_837),
.B(n_754),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_820),
.B(n_822),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_804),
.B(n_769),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_834),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_803),
.A2(n_776),
.B1(n_758),
.B2(n_757),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_832),
.B(n_769),
.Y(n_877)
);

INVxp33_ASAP7_75t_L g878 ( 
.A(n_802),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_804),
.Y(n_879)
);

INVxp67_ASAP7_75t_L g880 ( 
.A(n_848),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_854),
.B(n_770),
.Y(n_881)
);

HB1xp67_ASAP7_75t_L g882 ( 
.A(n_879),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_854),
.B(n_879),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_870),
.B(n_770),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_863),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_863),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_843),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_870),
.B(n_783),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_843),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_843),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_860),
.B(n_810),
.Y(n_891)
);

INVx5_ASAP7_75t_L g892 ( 
.A(n_855),
.Y(n_892)
);

OR2x2_ASAP7_75t_L g893 ( 
.A(n_874),
.B(n_755),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_874),
.B(n_783),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_869),
.A2(n_813),
.B1(n_799),
.B2(n_818),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_850),
.B(n_755),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_864),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_859),
.B(n_749),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_864),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_846),
.Y(n_900)
);

OAI211xp5_ASAP7_75t_L g901 ( 
.A1(n_876),
.A2(n_800),
.B(n_806),
.C(n_805),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_845),
.B(n_847),
.Y(n_902)
);

OAI221xp5_ASAP7_75t_L g903 ( 
.A1(n_876),
.A2(n_807),
.B1(n_841),
.B2(n_811),
.C(n_791),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_887),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_880),
.B(n_853),
.Y(n_905)
);

BUFx3_ASAP7_75t_L g906 ( 
.A(n_900),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_893),
.B(n_859),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_883),
.B(n_861),
.Y(n_908)
);

INVx4_ASAP7_75t_L g909 ( 
.A(n_900),
.Y(n_909)
);

OR2x2_ASAP7_75t_L g910 ( 
.A(n_893),
.B(n_867),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_885),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_882),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_892),
.B(n_846),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_883),
.B(n_888),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_898),
.B(n_894),
.Y(n_915)
);

INVx1_ASAP7_75t_SL g916 ( 
.A(n_891),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_887),
.Y(n_917)
);

NOR2x1p5_ASAP7_75t_L g918 ( 
.A(n_902),
.B(n_846),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_897),
.B(n_853),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_892),
.Y(n_920)
);

NAND2xp33_ASAP7_75t_SL g921 ( 
.A(n_918),
.B(n_819),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_916),
.A2(n_901),
.B1(n_903),
.B2(n_895),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_919),
.B(n_888),
.Y(n_923)
);

NAND2xp33_ASAP7_75t_SL g924 ( 
.A(n_909),
.B(n_878),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_905),
.B(n_884),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_913),
.A2(n_855),
.B1(n_799),
.B2(n_866),
.Y(n_926)
);

AO221x2_ASAP7_75t_L g927 ( 
.A1(n_911),
.A2(n_899),
.B1(n_886),
.B2(n_875),
.C(n_889),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_908),
.B(n_884),
.Y(n_928)
);

OAI221xp5_ASAP7_75t_L g929 ( 
.A1(n_920),
.A2(n_871),
.B1(n_855),
.B2(n_892),
.C(n_875),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_906),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_926),
.B(n_913),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_930),
.B(n_856),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_927),
.B(n_908),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_928),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_923),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_922),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_925),
.Y(n_937)
);

INVx4_ASAP7_75t_L g938 ( 
.A(n_924),
.Y(n_938)
);

NOR2x1_ASAP7_75t_L g939 ( 
.A(n_929),
.B(n_909),
.Y(n_939)
);

NAND2x1p5_ASAP7_75t_L g940 ( 
.A(n_938),
.B(n_909),
.Y(n_940)
);

OAI311xp33_ASAP7_75t_L g941 ( 
.A1(n_933),
.A2(n_896),
.A3(n_910),
.B1(n_862),
.C1(n_855),
.Y(n_941)
);

INVxp33_ASAP7_75t_L g942 ( 
.A(n_932),
.Y(n_942)
);

OAI21xp33_ASAP7_75t_L g943 ( 
.A1(n_936),
.A2(n_939),
.B(n_935),
.Y(n_943)
);

INVx2_ASAP7_75t_SL g944 ( 
.A(n_940),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_943),
.B(n_935),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_942),
.B(n_937),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_946),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_944),
.Y(n_948)
);

INVx1_ASAP7_75t_SL g949 ( 
.A(n_945),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_946),
.B(n_934),
.Y(n_950)
);

OA211x2_ASAP7_75t_L g951 ( 
.A1(n_950),
.A2(n_949),
.B(n_948),
.C(n_938),
.Y(n_951)
);

NOR4xp25_ASAP7_75t_L g952 ( 
.A(n_947),
.B(n_941),
.C(n_948),
.D(n_917),
.Y(n_952)
);

AOI211xp5_ASAP7_75t_SL g953 ( 
.A1(n_947),
.A2(n_931),
.B(n_913),
.C(n_912),
.Y(n_953)
);

AOI211xp5_ASAP7_75t_L g954 ( 
.A1(n_949),
.A2(n_921),
.B(n_931),
.C(n_795),
.Y(n_954)
);

NAND4xp25_ASAP7_75t_L g955 ( 
.A(n_947),
.B(n_920),
.C(n_906),
.D(n_789),
.Y(n_955)
);

NAND4xp25_ASAP7_75t_L g956 ( 
.A(n_947),
.B(n_789),
.C(n_827),
.D(n_814),
.Y(n_956)
);

NOR3xp33_ASAP7_75t_L g957 ( 
.A(n_947),
.B(n_871),
.C(n_830),
.Y(n_957)
);

NOR2x1_ASAP7_75t_L g958 ( 
.A(n_948),
.B(n_917),
.Y(n_958)
);

OAI21xp33_ASAP7_75t_L g959 ( 
.A1(n_955),
.A2(n_866),
.B(n_868),
.Y(n_959)
);

OAI211xp5_ASAP7_75t_SL g960 ( 
.A1(n_953),
.A2(n_910),
.B(n_915),
.C(n_907),
.Y(n_960)
);

OAI21xp5_ASAP7_75t_SL g961 ( 
.A1(n_957),
.A2(n_814),
.B(n_832),
.Y(n_961)
);

XNOR2xp5_ASAP7_75t_L g962 ( 
.A(n_954),
.B(n_951),
.Y(n_962)
);

AOI21xp33_ASAP7_75t_L g963 ( 
.A1(n_958),
.A2(n_896),
.B(n_892),
.Y(n_963)
);

AO22x2_ASAP7_75t_L g964 ( 
.A1(n_952),
.A2(n_904),
.B1(n_914),
.B2(n_915),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_SL g965 ( 
.A1(n_956),
.A2(n_914),
.B(n_868),
.Y(n_965)
);

XNOR2xp5_ASAP7_75t_L g966 ( 
.A(n_962),
.B(n_873),
.Y(n_966)
);

INVx1_ASAP7_75t_SL g967 ( 
.A(n_964),
.Y(n_967)
);

INVxp67_ASAP7_75t_L g968 ( 
.A(n_963),
.Y(n_968)
);

OR2x2_ASAP7_75t_L g969 ( 
.A(n_965),
.B(n_907),
.Y(n_969)
);

NAND4xp75_ASAP7_75t_L g970 ( 
.A(n_960),
.B(n_894),
.C(n_867),
.D(n_873),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_961),
.B(n_959),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_962),
.B(n_892),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_962),
.A2(n_877),
.B1(n_904),
.B2(n_881),
.Y(n_973)
);

NAND3xp33_ASAP7_75t_L g974 ( 
.A(n_968),
.B(n_815),
.C(n_849),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_966),
.B(n_815),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_967),
.B(n_890),
.Y(n_976)
);

NAND3xp33_ASAP7_75t_L g977 ( 
.A(n_972),
.B(n_815),
.C(n_849),
.Y(n_977)
);

XNOR2x1_ASAP7_75t_L g978 ( 
.A(n_971),
.B(n_877),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_R g979 ( 
.A(n_969),
.B(n_809),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_R g980 ( 
.A(n_970),
.B(n_809),
.Y(n_980)
);

NAND3xp33_ASAP7_75t_L g981 ( 
.A(n_973),
.B(n_844),
.C(n_847),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_R g982 ( 
.A(n_966),
.B(n_844),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_972),
.B(n_825),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_972),
.B(n_823),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_981),
.A2(n_890),
.B1(n_898),
.B2(n_858),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_975),
.A2(n_858),
.B1(n_877),
.B2(n_857),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_978),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_982),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_976),
.B(n_881),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_979),
.Y(n_990)
);

OAI211xp5_ASAP7_75t_SL g991 ( 
.A1(n_983),
.A2(n_865),
.B(n_758),
.C(n_757),
.Y(n_991)
);

AOI221xp5_ASAP7_75t_SL g992 ( 
.A1(n_984),
.A2(n_857),
.B1(n_852),
.B2(n_851),
.C(n_842),
.Y(n_992)
);

INVx1_ASAP7_75t_SL g993 ( 
.A(n_980),
.Y(n_993)
);

XNOR2x1_ASAP7_75t_L g994 ( 
.A(n_974),
.B(n_877),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_988),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_990),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_993),
.A2(n_987),
.B1(n_977),
.B2(n_989),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_L g998 ( 
.A1(n_994),
.A2(n_857),
.B1(n_852),
.B2(n_851),
.Y(n_998)
);

OR2x2_ASAP7_75t_SL g999 ( 
.A(n_992),
.B(n_851),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_986),
.A2(n_852),
.B1(n_765),
.B2(n_768),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_996),
.A2(n_991),
.B(n_985),
.Y(n_1001)
);

AOI22xp33_ASAP7_75t_SL g1002 ( 
.A1(n_995),
.A2(n_835),
.B1(n_842),
.B2(n_784),
.Y(n_1002)
);

INVxp67_ASAP7_75t_L g1003 ( 
.A(n_997),
.Y(n_1003)
);

AOI31xp33_ASAP7_75t_L g1004 ( 
.A1(n_1003),
.A2(n_998),
.A3(n_1000),
.B(n_999),
.Y(n_1004)
);

AOI22xp33_ASAP7_75t_L g1005 ( 
.A1(n_1002),
.A2(n_872),
.B1(n_784),
.B2(n_771),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_1005),
.A2(n_1001),
.B1(n_771),
.B2(n_778),
.Y(n_1006)
);

XOR2xp5_ASAP7_75t_L g1007 ( 
.A(n_1004),
.B(n_778),
.Y(n_1007)
);

AOI222xp33_ASAP7_75t_SL g1008 ( 
.A1(n_1006),
.A2(n_768),
.B1(n_765),
.B2(n_759),
.C1(n_784),
.C2(n_781),
.Y(n_1008)
);

AOI222xp33_ASAP7_75t_SL g1009 ( 
.A1(n_1007),
.A2(n_759),
.B1(n_782),
.B2(n_781),
.C1(n_761),
.C2(n_773),
.Y(n_1009)
);

AOI22xp33_ASAP7_75t_L g1010 ( 
.A1(n_1007),
.A2(n_872),
.B1(n_773),
.B2(n_761),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_1009),
.Y(n_1011)
);

OAI221xp5_ASAP7_75t_R g1012 ( 
.A1(n_1011),
.A2(n_1010),
.B1(n_1008),
.B2(n_748),
.C(n_756),
.Y(n_1012)
);

AOI211xp5_ASAP7_75t_L g1013 ( 
.A1(n_1012),
.A2(n_782),
.B(n_748),
.C(n_749),
.Y(n_1013)
);


endmodule