module fake_jpeg_31451_n_168 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_168);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_36),
.Y(n_59)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_15),
.B(n_7),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_37),
.B(n_41),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

INVxp67_ASAP7_75t_SL g55 ( 
.A(n_39),
.Y(n_55)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2x1_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_26),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_51),
.B(n_68),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_27),
.B1(n_24),
.B2(n_29),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_61),
.B1(n_64),
.B2(n_66),
.Y(n_76)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_27),
.B1(n_29),
.B2(n_26),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_34),
.A2(n_31),
.B1(n_28),
.B2(n_23),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_41),
.B1(n_46),
.B2(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_35),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_36),
.B(n_21),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_39),
.B(n_25),
.C(n_16),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_71),
.B(n_72),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_23),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_38),
.C(n_32),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_70),
.C(n_69),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_86),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_56),
.A2(n_25),
.B1(n_31),
.B2(n_28),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_91),
.B1(n_69),
.B2(n_33),
.Y(n_104)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_17),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_55),
.Y(n_95)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_21),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_54),
.A2(n_32),
.B1(n_38),
.B2(n_22),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_35),
.B1(n_33),
.B2(n_76),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_48),
.B(n_15),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_90),
.Y(n_112)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_61),
.A2(n_18),
.B1(n_17),
.B2(n_19),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_66),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_93),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_95),
.B(n_71),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_78),
.A2(n_49),
.B1(n_54),
.B2(n_50),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_104),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_83),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_18),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_108),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_77),
.A2(n_48),
.B1(n_52),
.B2(n_22),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_105),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_19),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_19),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_110),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_19),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_7),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_13),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_106),
.Y(n_131)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_91),
.C(n_75),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_123),
.C(n_96),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_94),
.A2(n_84),
.B(n_90),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_125),
.Y(n_135)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_84),
.B(n_93),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_124),
.A2(n_104),
.B(n_101),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_11),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_81),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_116),
.Y(n_139)
);

AOI221xp5_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_133),
.B1(n_127),
.B2(n_117),
.C(n_113),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_131),
.C(n_136),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_112),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_132),
.Y(n_146)
);

NAND3xp33_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_106),
.C(n_112),
.Y(n_132)
);

OAI321xp33_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_104),
.A3(n_9),
.B1(n_6),
.B2(n_13),
.C(n_99),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_104),
.C(n_85),
.Y(n_136)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_137),
.A2(n_124),
.B(n_121),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_141),
.A2(n_145),
.B(n_148),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_138),
.Y(n_143)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_144),
.A2(n_129),
.B1(n_102),
.B2(n_6),
.Y(n_151)
);

A2O1A1O1Ixp25_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_126),
.B(n_114),
.C(n_113),
.D(n_122),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_137),
.A2(n_115),
.B1(n_107),
.B2(n_74),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_147),
.A2(n_107),
.B1(n_134),
.B2(n_98),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_102),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_151),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_135),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_142),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_140),
.A2(n_107),
.B1(n_3),
.B2(n_5),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_147),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_157),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_146),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_148),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_158),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_159),
.A2(n_149),
.B1(n_154),
.B2(n_145),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_2),
.Y(n_164)
);

OAI21x1_ASAP7_75t_L g163 ( 
.A1(n_160),
.A2(n_156),
.B(n_159),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_163),
.A2(n_164),
.B(n_162),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_161),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_3),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_167),
.B(n_5),
.Y(n_168)
);


endmodule