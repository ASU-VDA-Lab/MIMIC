module fake_netlist_6_1683_n_110 (n_16, n_1, n_9, n_8, n_18, n_10, n_6, n_15, n_3, n_14, n_0, n_4, n_13, n_11, n_17, n_12, n_7, n_2, n_5, n_19, n_110);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_13;
input n_11;
input n_17;
input n_12;
input n_7;
input n_2;
input n_5;
input n_19;

output n_110;

wire n_52;
wire n_91;
wire n_46;
wire n_21;
wire n_88;
wire n_98;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_23;
wire n_20;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_109;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_97;
wire n_94;
wire n_108;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVxp67_ASAP7_75t_SL g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVxp67_ASAP7_75t_SL g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_9),
.B(n_13),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_1),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_24),
.Y(n_38)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_R g44 ( 
.A(n_21),
.B(n_1),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_25),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_22),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_22),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

AND2x4_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_20),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

AO22x2_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_35),
.B1(n_30),
.B2(n_28),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

AO22x2_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_30),
.B1(n_28),
.B2(n_27),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_45),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_47),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_20),
.B(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_46),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_61),
.A2(n_40),
.B1(n_37),
.B2(n_42),
.Y(n_64)
);

OAI21x1_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_52),
.B(n_50),
.Y(n_65)
);

NOR2x1_ASAP7_75t_SL g66 ( 
.A(n_61),
.B(n_26),
.Y(n_66)
);

OAI21x1_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_50),
.B(n_52),
.Y(n_67)
);

AOI221xp5_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_37),
.B1(n_34),
.B2(n_23),
.C(n_42),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

OR2x6_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_58),
.Y(n_70)
);

BUFx8_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_64),
.Y(n_72)
);

AOI211xp5_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_60),
.B(n_40),
.C(n_53),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_69),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

OAI211xp5_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_68),
.B(n_44),
.C(n_31),
.Y(n_78)
);

AND2x4_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_65),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_56),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_56),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_67),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_78),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_80),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_79),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_81),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_56),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

OAI221xp5_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_75),
.B1(n_27),
.B2(n_26),
.C(n_82),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_82),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_86),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_86),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_84),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_88),
.Y(n_97)
);

NOR4xp25_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_88),
.C(n_44),
.D(n_4),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_93),
.A2(n_72),
.B(n_71),
.Y(n_99)
);

AOI211xp5_ASAP7_75t_L g100 ( 
.A1(n_95),
.A2(n_57),
.B(n_3),
.C(n_5),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_96),
.A2(n_57),
.B(n_71),
.C(n_55),
.Y(n_101)
);

NOR3xp33_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_94),
.C(n_65),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

OAI22x1_ASAP7_75t_SL g104 ( 
.A1(n_103),
.A2(n_99),
.B1(n_101),
.B2(n_6),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_105),
.Y(n_106)
);

AO22x2_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_104),
.B1(n_105),
.B2(n_7),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_56),
.B1(n_54),
.B2(n_7),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_54),
.B1(n_5),
.B2(n_8),
.Y(n_109)
);

AOI221xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_2),
.B1(n_8),
.B2(n_10),
.C(n_107),
.Y(n_110)
);


endmodule