module fake_jpeg_6805_n_109 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_109);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_109;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_4),
.B(n_8),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_12),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_24),
.B(n_25),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_0),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_37),
.Y(n_44)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2x1_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_25),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_45),
.A2(n_22),
.B(n_19),
.C(n_18),
.Y(n_58)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_42),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_16),
.B1(n_13),
.B2(n_12),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_54),
.B1(n_38),
.B2(n_40),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_25),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_11),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_22),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_18),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_16),
.B1(n_21),
.B2(n_13),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_35),
.B(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_55),
.B(n_19),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_56),
.B(n_60),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_52),
.B(n_45),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_45),
.B(n_16),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_62),
.B(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_27),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_55),
.B(n_42),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_66),
.A2(n_49),
.B1(n_50),
.B2(n_48),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_68),
.B(n_11),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_54),
.B(n_50),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_71),
.A2(n_58),
.B(n_67),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_47),
.B1(n_38),
.B2(n_43),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_51),
.C(n_48),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_77),
.C(n_27),
.Y(n_81)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_27),
.C(n_46),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_57),
.B1(n_66),
.B2(n_53),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_83),
.B1(n_84),
.B2(n_38),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_77),
.C(n_68),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_11),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_43),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_73),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_89),
.C(n_91),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_20),
.B(n_3),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_85),
.A2(n_76),
.B1(n_69),
.B2(n_70),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_88),
.A2(n_20),
.B1(n_3),
.B2(n_4),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_72),
.C(n_34),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_40),
.C(n_34),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_80),
.B1(n_78),
.B2(n_84),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_34),
.C(n_20),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_96),
.B(n_98),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_97),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_9),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g102 ( 
.A1(n_99),
.A2(n_87),
.B1(n_94),
.B2(n_95),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_5),
.Y(n_105)
);

O2A1O1Ixp5_ASAP7_75t_L g104 ( 
.A1(n_102),
.A2(n_101),
.B(n_6),
.C(n_7),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_104),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

BUFx24_ASAP7_75t_SL g108 ( 
.A(n_107),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_106),
.Y(n_109)
);


endmodule