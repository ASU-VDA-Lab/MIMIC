module real_aes_17554_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g117 ( .A(n_0), .B(n_118), .Y(n_117) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_1), .A2(n_4), .B1(n_215), .B2(n_600), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g152 ( .A1(n_2), .A2(n_44), .B1(n_153), .B2(n_155), .Y(n_152) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_3), .A2(n_25), .B1(n_155), .B2(n_179), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_5), .A2(n_16), .B1(n_196), .B2(n_233), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_6), .A2(n_61), .B1(n_181), .B2(n_253), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_7), .A2(n_17), .B1(n_153), .B2(n_200), .Y(n_523) );
INVx1_ASAP7_75t_L g118 ( .A(n_8), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g585 ( .A(n_9), .Y(n_585) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_10), .Y(n_269) );
AOI22xp5_ASAP7_75t_L g251 ( .A1(n_11), .A2(n_18), .B1(n_198), .B2(n_252), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g823 ( .A1(n_12), .A2(n_65), .B1(n_824), .B2(n_825), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_12), .Y(n_824) );
BUFx2_ASAP7_75t_L g110 ( .A(n_13), .Y(n_110) );
OR2x2_ASAP7_75t_L g134 ( .A(n_13), .B(n_39), .Y(n_134) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_14), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_15), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g214 ( .A1(n_19), .A2(n_101), .B1(n_196), .B2(n_215), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g828 ( .A1(n_20), .A2(n_489), .B(n_829), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_21), .A2(n_40), .B1(n_229), .B2(n_230), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_22), .B(n_197), .Y(n_270) );
OAI22x1_ASAP7_75t_SL g821 ( .A1(n_23), .A2(n_822), .B1(n_823), .B2(n_826), .Y(n_821) );
CKINVDCx5p33_ASAP7_75t_R g826 ( .A(n_23), .Y(n_826) );
OAI21x1_ASAP7_75t_L g169 ( .A1(n_24), .A2(n_59), .B(n_170), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_26), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g593 ( .A(n_27), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_28), .B(n_159), .Y(n_547) );
INVx4_ASAP7_75t_R g536 ( .A(n_29), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g160 ( .A1(n_30), .A2(n_48), .B1(n_161), .B2(n_163), .Y(n_160) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_31), .A2(n_55), .B1(n_163), .B2(n_196), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_32), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_33), .B(n_229), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_34), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_35), .B(n_155), .Y(n_554) );
INVx1_ASAP7_75t_L g602 ( .A(n_36), .Y(n_602) );
A2O1A1Ixp33_ASAP7_75t_SL g583 ( .A1(n_37), .A2(n_153), .B(n_165), .C(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_38), .A2(n_56), .B1(n_153), .B2(n_163), .Y(n_591) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_39), .Y(n_109) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_41), .A2(n_88), .B1(n_153), .B2(n_178), .Y(n_177) );
OAI22xp5_ASAP7_75t_SL g137 ( .A1(n_42), .A2(n_54), .B1(n_138), .B2(n_139), .Y(n_137) );
INVx1_ASAP7_75t_L g139 ( .A(n_42), .Y(n_139) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_43), .A2(n_47), .B1(n_153), .B2(n_200), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_45), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_46), .A2(n_60), .B1(n_196), .B2(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g551 ( .A(n_49), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_50), .B(n_153), .Y(n_553) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_51), .Y(n_564) );
INVx2_ASAP7_75t_L g123 ( .A(n_52), .Y(n_123) );
INVx1_ASAP7_75t_L g113 ( .A(n_53), .Y(n_113) );
BUFx3_ASAP7_75t_L g499 ( .A(n_53), .Y(n_499) );
INVx1_ASAP7_75t_L g138 ( .A(n_54), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_57), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_58), .A2(n_89), .B1(n_153), .B2(n_163), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_62), .A2(n_77), .B1(n_161), .B2(n_218), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g526 ( .A(n_63), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_64), .A2(n_79), .B1(n_153), .B2(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g825 ( .A(n_65), .Y(n_825) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_66), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_67), .A2(n_100), .B1(n_196), .B2(n_198), .Y(n_195) );
AND2x4_ASAP7_75t_L g149 ( .A(n_68), .B(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g170 ( .A(n_69), .Y(n_170) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_70), .A2(n_91), .B1(n_161), .B2(n_163), .Y(n_598) );
AO22x1_ASAP7_75t_L g512 ( .A1(n_71), .A2(n_78), .B1(n_230), .B2(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g150 ( .A(n_72), .Y(n_150) );
AND2x2_ASAP7_75t_L g586 ( .A(n_73), .B(n_167), .Y(n_586) );
CKINVDCx14_ASAP7_75t_R g127 ( .A(n_74), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_74), .B(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_75), .B(n_181), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g579 ( .A(n_76), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_80), .B(n_155), .Y(n_565) );
INVx2_ASAP7_75t_L g159 ( .A(n_81), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_82), .B(n_167), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_83), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g180 ( .A1(n_84), .A2(n_99), .B1(n_163), .B2(n_181), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_85), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_86), .B(n_188), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_87), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_90), .B(n_167), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_92), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_93), .B(n_167), .Y(n_561) );
INVx1_ASAP7_75t_L g116 ( .A(n_94), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_94), .B(n_132), .Y(n_131) );
NAND2xp33_ASAP7_75t_L g273 ( .A(n_95), .B(n_197), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g837 ( .A(n_96), .Y(n_837) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_97), .A2(n_181), .B(n_183), .C(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g538 ( .A(n_98), .B(n_539), .Y(n_538) );
NAND2xp33_ASAP7_75t_L g569 ( .A(n_102), .B(n_162), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_119), .B(n_836), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx3_ASAP7_75t_L g839 ( .A(n_106), .Y(n_839) );
AND2x4_ASAP7_75t_L g106 ( .A(n_107), .B(n_111), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
NOR2x1p5_ASAP7_75t_L g111 ( .A(n_112), .B(n_114), .Y(n_111) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g132 ( .A(n_113), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_117), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g819 ( .A(n_116), .Y(n_819) );
OR2x6_ASAP7_75t_L g119 ( .A(n_120), .B(n_492), .Y(n_119) );
NOR2x1_ASAP7_75t_L g120 ( .A(n_121), .B(n_124), .Y(n_120) );
BUFx8_ASAP7_75t_SL g121 ( .A(n_122), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g496 ( .A(n_123), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_123), .B(n_833), .Y(n_832) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_484), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_135), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
INVx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
CKINVDCx8_ASAP7_75t_R g129 ( .A(n_130), .Y(n_129) );
INVx4_ASAP7_75t_L g488 ( .A(n_130), .Y(n_488) );
INVx5_ASAP7_75t_L g491 ( .A(n_130), .Y(n_491) );
AND2x6_ASAP7_75t_SL g130 ( .A(n_131), .B(n_133), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_133), .B(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NOR2x1_ASAP7_75t_L g835 ( .A(n_134), .B(n_499), .Y(n_835) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AOI21xp33_ASAP7_75t_SL g484 ( .A1(n_136), .A2(n_485), .B(n_489), .Y(n_484) );
XNOR2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_140), .Y(n_136) );
OAI22x1_ASAP7_75t_L g502 ( .A1(n_140), .A2(n_503), .B1(n_817), .B2(n_820), .Y(n_502) );
NOR2x1p5_ASAP7_75t_L g140 ( .A(n_141), .B(n_394), .Y(n_140) );
NAND4xp75_ASAP7_75t_L g141 ( .A(n_142), .B(n_339), .C(n_359), .D(n_375), .Y(n_141) );
NOR2x1p5_ASAP7_75t_SL g142 ( .A(n_143), .B(n_309), .Y(n_142) );
NAND4xp75_ASAP7_75t_L g143 ( .A(n_144), .B(n_245), .C(n_286), .D(n_295), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_145), .B(n_206), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_173), .Y(n_145) );
AND2x4_ASAP7_75t_L g419 ( .A(n_146), .B(n_346), .Y(n_419) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_147), .Y(n_262) );
INVx2_ASAP7_75t_L g280 ( .A(n_147), .Y(n_280) );
AND2x2_ASAP7_75t_L g303 ( .A(n_147), .B(n_265), .Y(n_303) );
OR2x2_ASAP7_75t_L g358 ( .A(n_147), .B(n_174), .Y(n_358) );
AO31x2_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_151), .A3(n_166), .B(n_171), .Y(n_147) );
INVx2_ASAP7_75t_L g203 ( .A(n_148), .Y(n_203) );
AO31x2_ASAP7_75t_L g226 ( .A1(n_148), .A2(n_175), .A3(n_227), .B(n_235), .Y(n_226) );
AO31x2_ASAP7_75t_L g249 ( .A1(n_148), .A2(n_192), .A3(n_250), .B(n_256), .Y(n_249) );
AO31x2_ASAP7_75t_L g521 ( .A1(n_148), .A2(n_223), .A3(n_522), .B(n_525), .Y(n_521) );
BUFx10_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g185 ( .A(n_149), .Y(n_185) );
INVx1_ASAP7_75t_L g519 ( .A(n_149), .Y(n_519) );
BUFx10_ASAP7_75t_L g556 ( .A(n_149), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_156), .B1(n_160), .B2(n_164), .Y(n_151) );
INVx1_ASAP7_75t_L g198 ( .A(n_153), .Y(n_198) );
INVx4_ASAP7_75t_L g200 ( .A(n_153), .Y(n_200) );
INVx1_ASAP7_75t_L g218 ( .A(n_153), .Y(n_218) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_154), .Y(n_155) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_154), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_154), .Y(n_163) );
INVx2_ASAP7_75t_L g179 ( .A(n_154), .Y(n_179) );
INVx1_ASAP7_75t_L g181 ( .A(n_154), .Y(n_181) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_154), .Y(n_197) );
INVx1_ASAP7_75t_L g216 ( .A(n_154), .Y(n_216) );
INVx1_ASAP7_75t_L g231 ( .A(n_154), .Y(n_231) );
INVx1_ASAP7_75t_L g234 ( .A(n_154), .Y(n_234) );
INVx1_ASAP7_75t_L g254 ( .A(n_154), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_155), .B(n_579), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g213 ( .A1(n_156), .A2(n_164), .B1(n_214), .B2(n_217), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g227 ( .A1(n_156), .A2(n_164), .B1(n_228), .B2(n_232), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_156), .A2(n_164), .B1(n_241), .B2(n_242), .Y(n_240) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g515 ( .A(n_157), .Y(n_515) );
BUFx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g567 ( .A(n_158), .Y(n_567) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
BUFx8_ASAP7_75t_L g165 ( .A(n_159), .Y(n_165) );
INVx1_ASAP7_75t_L g183 ( .A(n_159), .Y(n_183) );
INVx1_ASAP7_75t_L g550 ( .A(n_159), .Y(n_550) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g229 ( .A(n_162), .Y(n_229) );
OAI22xp33_ASAP7_75t_L g535 ( .A1(n_162), .A2(n_234), .B1(n_536), .B2(n_537), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_163), .B(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g600 ( .A(n_163), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g176 ( .A1(n_164), .A2(n_177), .B1(n_180), .B2(n_182), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g194 ( .A1(n_164), .A2(n_195), .B1(n_199), .B2(n_201), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_164), .A2(n_201), .B1(n_251), .B2(n_255), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_164), .A2(n_272), .B(n_273), .Y(n_271) );
OAI22x1_ASAP7_75t_L g522 ( .A1(n_164), .A2(n_182), .B1(n_523), .B2(n_524), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_164), .A2(n_515), .B1(n_590), .B2(n_591), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_164), .A2(n_182), .B1(n_598), .B2(n_599), .Y(n_597) );
INVx6_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
O2A1O1Ixp5_ASAP7_75t_L g268 ( .A1(n_165), .A2(n_200), .B(n_269), .C(n_270), .Y(n_268) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_165), .A2(n_512), .B(n_514), .C(n_518), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_165), .A2(n_569), .B(n_570), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_165), .B(n_512), .Y(n_614) );
AO31x2_ASAP7_75t_L g588 ( .A1(n_166), .A2(n_556), .A3(n_589), .B(n_592), .Y(n_588) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2x1_ASAP7_75t_L g571 ( .A(n_167), .B(n_572), .Y(n_571) );
INVx4_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_168), .B(n_172), .Y(n_171) );
BUFx3_ASAP7_75t_L g175 ( .A(n_168), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_168), .B(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_168), .B(n_236), .Y(n_235) );
INVx2_ASAP7_75t_SL g266 ( .A(n_168), .Y(n_266) );
AND2x2_ASAP7_75t_L g555 ( .A(n_168), .B(n_556), .Y(n_555) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g188 ( .A(n_169), .Y(n_188) );
AND2x2_ASAP7_75t_L g276 ( .A(n_173), .B(n_277), .Y(n_276) );
AND2x4_ASAP7_75t_L g426 ( .A(n_173), .B(n_303), .Y(n_426) );
AND2x4_ASAP7_75t_L g173 ( .A(n_174), .B(n_190), .Y(n_173) );
OR2x2_ASAP7_75t_L g263 ( .A(n_174), .B(n_264), .Y(n_263) );
BUFx2_ASAP7_75t_L g294 ( .A(n_174), .Y(n_294) );
AND2x2_ASAP7_75t_L g300 ( .A(n_174), .B(n_191), .Y(n_300) );
INVx1_ASAP7_75t_L g318 ( .A(n_174), .Y(n_318) );
INVx2_ASAP7_75t_L g347 ( .A(n_174), .Y(n_347) );
AO31x2_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .A3(n_184), .B(n_186), .Y(n_174) );
INVx2_ASAP7_75t_SL g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_179), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_182), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_SL g201 ( .A(n_183), .Y(n_201) );
AO31x2_ASAP7_75t_L g239 ( .A1(n_184), .A2(n_219), .A3(n_240), .B(n_243), .Y(n_239) );
AO31x2_ASAP7_75t_L g596 ( .A1(n_184), .A2(n_192), .A3(n_597), .B(n_601), .Y(n_596) );
INVx2_ASAP7_75t_SL g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_SL g274 ( .A(n_185), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_187), .B(n_189), .Y(n_186) );
INVx2_ASAP7_75t_L g220 ( .A(n_187), .Y(n_220) );
NOR2xp33_ASAP7_75t_SL g256 ( .A(n_187), .B(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g193 ( .A(n_188), .Y(n_193) );
INVx2_ASAP7_75t_L g223 ( .A(n_188), .Y(n_223) );
OAI21xp33_ASAP7_75t_L g518 ( .A1(n_188), .A2(n_517), .B(n_519), .Y(n_518) );
INVx3_ASAP7_75t_L g323 ( .A(n_190), .Y(n_323) );
INVx2_ASAP7_75t_L g328 ( .A(n_190), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_190), .B(n_279), .Y(n_333) );
AND2x2_ASAP7_75t_L g356 ( .A(n_190), .B(n_335), .Y(n_356) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_190), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_190), .B(n_411), .Y(n_410) );
INVx3_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
BUFx2_ASAP7_75t_L g345 ( .A(n_191), .Y(n_345) );
AND2x2_ASAP7_75t_L g393 ( .A(n_191), .B(n_347), .Y(n_393) );
AO31x2_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_194), .A3(n_202), .B(n_204), .Y(n_191) );
AOI21x1_ASAP7_75t_L g575 ( .A1(n_192), .A2(n_576), .B(n_586), .Y(n_575) );
BUFx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_193), .B(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g539 ( .A(n_193), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_193), .B(n_593), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_193), .B(n_602), .Y(n_601) );
INVx3_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVxp67_ASAP7_75t_SL g513 ( .A(n_197), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g563 ( .A1(n_200), .A2(n_564), .B(n_565), .C(n_566), .Y(n_563) );
AO31x2_ASAP7_75t_L g212 ( .A1(n_202), .A2(n_213), .A3(n_219), .B(n_221), .Y(n_212) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_203), .A2(n_531), .B(n_534), .Y(n_530) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_208), .B(n_224), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_208), .B(n_337), .Y(n_384) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2x1p5_ASAP7_75t_L g381 ( .A(n_209), .B(n_337), .Y(n_381) );
INVx1_ASAP7_75t_L g482 ( .A(n_209), .Y(n_482) );
INVx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g432 ( .A(n_210), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g285 ( .A(n_211), .Y(n_285) );
OR2x2_ASAP7_75t_L g366 ( .A(n_211), .B(n_238), .Y(n_366) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g308 ( .A(n_212), .Y(n_308) );
AND2x4_ASAP7_75t_L g314 ( .A(n_212), .B(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_216), .B(n_581), .Y(n_580) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_219), .A2(n_530), .B(n_538), .Y(n_529) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_222), .B(n_223), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_223), .B(n_244), .Y(n_243) );
AOI32xp33_ASAP7_75t_L g452 ( .A1(n_224), .A2(n_355), .A3(n_453), .B1(n_455), .B2(n_456), .Y(n_452) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
OR2x2_ASAP7_75t_L g401 ( .A(n_225), .B(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_226), .B(n_237), .Y(n_225) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_226), .Y(n_247) );
OR2x2_ASAP7_75t_L g283 ( .A(n_226), .B(n_239), .Y(n_283) );
INVx1_ASAP7_75t_L g298 ( .A(n_226), .Y(n_298) );
AND2x2_ASAP7_75t_L g307 ( .A(n_226), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g313 ( .A(n_226), .Y(n_313) );
INVx2_ASAP7_75t_L g338 ( .A(n_226), .Y(n_338) );
AND2x2_ASAP7_75t_L g457 ( .A(n_226), .B(n_249), .Y(n_457) );
OAI21xp33_ASAP7_75t_SL g546 ( .A1(n_230), .A2(n_547), .B(n_548), .Y(n_546) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_237), .B(n_290), .Y(n_377) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g248 ( .A(n_239), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g306 ( .A(n_239), .Y(n_306) );
INVx2_ASAP7_75t_L g315 ( .A(n_239), .Y(n_315) );
AND2x4_ASAP7_75t_L g337 ( .A(n_239), .B(n_338), .Y(n_337) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_239), .Y(n_429) );
AOI22x1_ASAP7_75t_SL g245 ( .A1(n_246), .A2(n_258), .B1(n_276), .B2(n_281), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
NAND4xp25_ASAP7_75t_L g406 ( .A(n_248), .B(n_407), .C(n_408), .D(n_409), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_248), .B(n_307), .Y(n_437) );
INVx4_ASAP7_75t_SL g290 ( .A(n_249), .Y(n_290) );
BUFx2_ASAP7_75t_L g353 ( .A(n_249), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_249), .B(n_298), .Y(n_416) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_254), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g378 ( .A(n_260), .B(n_327), .Y(n_378) );
NOR2x1_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x4_ASAP7_75t_L g301 ( .A(n_264), .B(n_279), .Y(n_301) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_265), .B(n_280), .Y(n_325) );
OAI21x1_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_267), .B(n_275), .Y(n_265) );
OAI21x1_ASAP7_75t_L g320 ( .A1(n_266), .A2(n_267), .B(n_275), .Y(n_320) );
OAI21x1_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_271), .B(n_274), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_277), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g343 ( .A(n_277), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g382 ( .A(n_278), .B(n_300), .Y(n_382) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g425 ( .A(n_280), .B(n_335), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_281), .A2(n_398), .B1(n_400), .B2(n_403), .C(n_405), .Y(n_397) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx2_ASAP7_75t_L g291 ( .A(n_283), .Y(n_291) );
OR2x2_ASAP7_75t_L g391 ( .A(n_283), .B(n_330), .Y(n_391) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_292), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_287), .A2(n_413), .B1(n_417), .B2(n_420), .Y(n_412) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_291), .Y(n_287) );
AND2x4_ASAP7_75t_L g336 ( .A(n_288), .B(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g448 ( .A(n_288), .B(n_366), .Y(n_448) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x4_ASAP7_75t_L g296 ( .A(n_290), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g312 ( .A(n_290), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g371 ( .A(n_290), .B(n_308), .Y(n_371) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_290), .Y(n_388) );
INVx1_ASAP7_75t_L g402 ( .A(n_290), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_290), .B(n_315), .Y(n_445) );
AND2x4_ASAP7_75t_L g352 ( .A(n_291), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g350 ( .A(n_293), .Y(n_350) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_294), .B(n_335), .Y(n_334) );
NAND2x1_ASAP7_75t_L g454 ( .A(n_294), .B(n_356), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_299), .B1(n_302), .B2(n_304), .Y(n_295) );
AND2x2_ASAP7_75t_L g321 ( .A(n_296), .B(n_314), .Y(n_321) );
INVx1_ASAP7_75t_L g362 ( .A(n_296), .Y(n_362) );
AND2x2_ASAP7_75t_L g469 ( .A(n_296), .B(n_330), .Y(n_469) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x4_ASAP7_75t_SL g299 ( .A(n_300), .B(n_301), .Y(n_299) );
AND2x2_ASAP7_75t_L g302 ( .A(n_300), .B(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g442 ( .A(n_300), .Y(n_442) );
AND2x2_ASAP7_75t_L g459 ( .A(n_300), .B(n_319), .Y(n_459) );
AND2x2_ASAP7_75t_L g475 ( .A(n_300), .B(n_425), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_301), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g398 ( .A(n_301), .B(n_399), .Y(n_398) );
OAI22xp33_ASAP7_75t_L g405 ( .A1(n_301), .A2(n_391), .B1(n_406), .B2(n_410), .Y(n_405) );
INVx1_ASAP7_75t_L g361 ( .A(n_303), .Y(n_361) );
AND2x2_ASAP7_75t_L g392 ( .A(n_303), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_303), .B(n_399), .Y(n_421) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g427 ( .A(n_307), .B(n_428), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_307), .A2(n_331), .B1(n_436), .B2(n_438), .Y(n_435) );
INVx3_ASAP7_75t_L g330 ( .A(n_308), .Y(n_330) );
AND2x2_ASAP7_75t_L g462 ( .A(n_308), .B(n_315), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_326), .Y(n_309) );
AOI32xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_316), .A3(n_319), .B1(n_321), .B2(n_322), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_313), .Y(n_408) );
INVx1_ASAP7_75t_L g433 ( .A(n_313), .Y(n_433) );
INVx3_ASAP7_75t_L g389 ( .A(n_314), .Y(n_389) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OAI221xp5_ASAP7_75t_L g464 ( .A1(n_317), .A2(n_465), .B1(n_466), .B2(n_467), .C(n_468), .Y(n_464) );
BUFx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g441 ( .A(n_319), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g477 ( .A(n_319), .B(n_438), .Y(n_477) );
BUFx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g335 ( .A(n_320), .Y(n_335) );
NAND2x1p5_ASAP7_75t_L g349 ( .A(n_322), .B(n_350), .Y(n_349) );
AO22x1_ASAP7_75t_L g379 ( .A1(n_322), .A2(n_380), .B1(n_382), .B2(n_383), .Y(n_379) );
NAND2x1p5_ASAP7_75t_L g483 ( .A(n_322), .B(n_350), .Y(n_483) );
AND2x4_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx2_ASAP7_75t_L g399 ( .A(n_323), .Y(n_399) );
INVx1_ASAP7_75t_L g409 ( .A(n_323), .Y(n_409) );
AND2x2_ASAP7_75t_L g329 ( .A(n_324), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVxp67_ASAP7_75t_SL g411 ( .A(n_325), .Y(n_411) );
INVx1_ASAP7_75t_L g451 ( .A(n_325), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_329), .B(n_331), .C(n_336), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NOR2x1p5_ASAP7_75t_L g438 ( .A(n_328), .B(n_358), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_329), .B(n_388), .Y(n_465) );
AOI31xp33_ASAP7_75t_L g348 ( .A1(n_330), .A2(n_349), .A3(n_351), .B(n_354), .Y(n_348) );
INVx4_ASAP7_75t_L g407 ( .A(n_330), .Y(n_407) );
OR2x2_ASAP7_75t_L g444 ( .A(n_330), .B(n_445), .Y(n_444) );
INVx2_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
AND2x4_ASAP7_75t_L g346 ( .A(n_335), .B(n_347), .Y(n_346) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_337), .Y(n_342) );
AND2x2_ASAP7_75t_L g373 ( .A(n_337), .B(n_371), .Y(n_373) );
NOR2xp67_ASAP7_75t_L g339 ( .A(n_340), .B(n_348), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVx1_ASAP7_75t_L g466 ( .A(n_343), .Y(n_466) );
INVx1_ASAP7_75t_L g374 ( .A(n_344), .Y(n_374) );
AND2x4_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
INVx1_ASAP7_75t_L g404 ( .A(n_345), .Y(n_404) );
AND2x2_ASAP7_75t_L g403 ( .A(n_346), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OAI322xp33_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_362), .A3(n_363), .B1(n_367), .B2(n_370), .C1(n_372), .C2(n_374), .Y(n_360) );
INVxp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AOI211x1_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_378), .B(n_379), .C(n_385), .Y(n_375) );
INVx1_ASAP7_75t_L g480 ( .A(n_376), .Y(n_480) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g434 ( .A(n_378), .Y(n_434) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OA21x2_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_390), .B(n_392), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx2_ASAP7_75t_L g455 ( .A(n_389), .Y(n_455) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND2xp33_ASAP7_75t_L g450 ( .A(n_393), .B(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_463), .Y(n_394) );
NOR3xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_430), .C(n_446), .Y(n_395) );
NAND3xp33_ASAP7_75t_L g396 ( .A(n_397), .B(n_412), .C(n_422), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_399), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OAI21xp33_ASAP7_75t_L g458 ( .A1(n_403), .A2(n_459), .B(n_460), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_407), .B(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_407), .B(n_457), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_408), .B(n_482), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_409), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OAI21xp5_ASAP7_75t_L g468 ( .A1(n_419), .A2(n_469), .B(n_470), .Y(n_468) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OAI21xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_426), .B(n_427), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OAI211xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_434), .B(n_435), .C(n_439), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_440), .B(n_443), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_SL g449 ( .A(n_441), .B(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_445), .Y(n_467) );
OAI211xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_449), .B(n_452), .C(n_458), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_457), .B(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g478 ( .A(n_457), .Y(n_478) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g474 ( .A(n_462), .Y(n_474) );
NOR3xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_472), .C(n_479), .Y(n_463) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AOI21xp33_ASAP7_75t_SL g472 ( .A1(n_473), .A2(n_476), .B(n_478), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AOI21xp33_ASAP7_75t_R g479 ( .A1(n_480), .A2(n_481), .B(n_483), .Y(n_479) );
INVx4_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx12f_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
OAI21xp33_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_500), .B(n_828), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_494), .Y(n_493) );
BUFx12f_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x6_ASAP7_75t_SL g495 ( .A(n_496), .B(n_497), .Y(n_495) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_502), .B1(n_821), .B2(n_827), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x4_ASAP7_75t_L g503 ( .A(n_504), .B(n_727), .Y(n_503) );
NOR3xp33_ASAP7_75t_L g504 ( .A(n_505), .B(n_656), .C(n_698), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_630), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_540), .B1(n_605), .B2(n_616), .Y(n_506) );
INVx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_527), .Y(n_508) );
AOI21xp33_ASAP7_75t_L g649 ( .A1(n_509), .A2(n_650), .B(n_652), .Y(n_649) );
AOI21xp33_ASAP7_75t_L g722 ( .A1(n_509), .A2(n_723), .B(n_724), .Y(n_722) );
OR2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_520), .Y(n_509) );
INVx2_ASAP7_75t_L g642 ( .A(n_510), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_510), .B(n_521), .Y(n_672) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g613 ( .A(n_514), .Y(n_613) );
OAI21x1_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_517), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_515), .A2(n_553), .B(n_554), .Y(n_552) );
INVx1_ASAP7_75t_L g615 ( .A(n_518), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_519), .A2(n_577), .B(n_583), .Y(n_576) );
AND2x2_ASAP7_75t_L g712 ( .A(n_520), .B(n_559), .Y(n_712) );
INVx1_ASAP7_75t_L g745 ( .A(n_520), .Y(n_745) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g607 ( .A(n_521), .B(n_560), .Y(n_607) );
AND2x2_ASAP7_75t_L g638 ( .A(n_521), .B(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g647 ( .A(n_521), .Y(n_647) );
OR2x2_ASAP7_75t_L g666 ( .A(n_521), .B(n_529), .Y(n_666) );
AND2x2_ASAP7_75t_L g681 ( .A(n_521), .B(n_529), .Y(n_681) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_528), .B(n_680), .Y(n_723) );
OR2x2_ASAP7_75t_L g811 ( .A(n_528), .B(n_672), .Y(n_811) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g639 ( .A(n_529), .Y(n_639) );
AND2x2_ASAP7_75t_L g648 ( .A(n_529), .B(n_611), .Y(n_648) );
AND2x2_ASAP7_75t_L g651 ( .A(n_529), .B(n_560), .Y(n_651) );
AND2x2_ASAP7_75t_L g670 ( .A(n_529), .B(n_559), .Y(n_670) );
AND2x4_ASAP7_75t_L g689 ( .A(n_529), .B(n_612), .Y(n_689) );
OAI21xp33_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_557), .B(n_594), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_541), .B(n_684), .Y(n_787) );
CKINVDCx14_ASAP7_75t_R g541 ( .A(n_542), .Y(n_541) );
BUFx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_543), .B(n_604), .Y(n_603) );
INVx3_ASAP7_75t_L g620 ( .A(n_543), .Y(n_620) );
OR2x2_ASAP7_75t_L g628 ( .A(n_543), .B(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_543), .B(n_621), .Y(n_653) );
AND2x2_ASAP7_75t_L g678 ( .A(n_543), .B(n_596), .Y(n_678) );
AND2x2_ASAP7_75t_L g696 ( .A(n_543), .B(n_626), .Y(n_696) );
INVx1_ASAP7_75t_L g735 ( .A(n_543), .Y(n_735) );
AND2x2_ASAP7_75t_L g737 ( .A(n_543), .B(n_738), .Y(n_737) );
NAND2x1p5_ASAP7_75t_SL g756 ( .A(n_543), .B(n_677), .Y(n_756) );
AND2x4_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
OAI21xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_552), .B(n_555), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
BUFx4f_ASAP7_75t_L g582 ( .A(n_550), .Y(n_582) );
INVx1_ASAP7_75t_L g572 ( .A(n_556), .Y(n_572) );
OAI32xp33_ASAP7_75t_L g640 ( .A1(n_557), .A2(n_632), .A3(n_641), .B1(n_643), .B2(n_645), .Y(n_640) );
OR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_573), .Y(n_557) );
INVx1_ASAP7_75t_L g680 ( .A(n_558), .Y(n_680) );
AND2x2_ASAP7_75t_L g688 ( .A(n_558), .B(n_689), .Y(n_688) );
BUFx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g687 ( .A(n_559), .B(n_611), .Y(n_687) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
BUFx3_ASAP7_75t_L g637 ( .A(n_560), .Y(n_637) );
AND2x2_ASAP7_75t_L g646 ( .A(n_560), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g752 ( .A(n_560), .Y(n_752) );
NAND2x1p5_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
OAI21x1_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_568), .B(n_571), .Y(n_562) );
INVx2_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g622 ( .A(n_573), .Y(n_622) );
OR2x2_ASAP7_75t_L g632 ( .A(n_573), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g754 ( .A(n_573), .Y(n_754) );
OR2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_587), .Y(n_573) );
AND2x2_ASAP7_75t_L g655 ( .A(n_574), .B(n_588), .Y(n_655) );
INVx2_ASAP7_75t_L g677 ( .A(n_574), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_574), .B(n_596), .Y(n_697) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g604 ( .A(n_575), .Y(n_604) );
OAI21xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_580), .B(n_582), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_587), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g686 ( .A(n_587), .Y(n_686) );
INVx2_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
BUFx2_ASAP7_75t_L g626 ( .A(n_588), .Y(n_626) );
OR2x2_ASAP7_75t_L g692 ( .A(n_588), .B(n_596), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_588), .B(n_596), .Y(n_725) );
INVx2_ASAP7_75t_L g673 ( .A(n_594), .Y(n_673) );
OR2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_603), .Y(n_594) );
OR2x2_ASAP7_75t_L g660 ( .A(n_595), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g738 ( .A(n_595), .Y(n_738) );
INVx1_ASAP7_75t_L g621 ( .A(n_596), .Y(n_621) );
INVx1_ASAP7_75t_L g629 ( .A(n_596), .Y(n_629) );
INVx1_ASAP7_75t_L g644 ( .A(n_596), .Y(n_644) );
OR2x2_ASAP7_75t_L g748 ( .A(n_603), .B(n_725), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_604), .B(n_620), .Y(n_661) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_604), .Y(n_663) );
OR2x2_ASAP7_75t_L g762 ( .A(n_604), .B(n_686), .Y(n_762) );
INVxp67_ASAP7_75t_L g786 ( .A(n_604), .Y(n_786) );
INVx2_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
NAND2x1_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_607), .B(n_648), .Y(n_715) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g664 ( .A(n_609), .B(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g777 ( .A(n_610), .Y(n_777) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g806 ( .A(n_611), .B(n_639), .Y(n_806) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g732 ( .A(n_612), .B(n_639), .Y(n_732) );
AOI21x1_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_614), .B(n_615), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_623), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_622), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_619), .B(n_655), .Y(n_769) );
AND2x4_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
INVx2_ASAP7_75t_L g633 ( .A(n_620), .Y(n_633) );
AND2x2_ASAP7_75t_L g683 ( .A(n_620), .B(n_684), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_620), .B(n_677), .Y(n_726) );
OR2x2_ASAP7_75t_L g798 ( .A(n_620), .B(n_685), .Y(n_798) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g718 ( .A(n_624), .B(n_719), .Y(n_718) );
AND2x4_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx2_ASAP7_75t_L g709 ( .A(n_625), .Y(n_709) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g699 ( .A(n_628), .B(n_700), .Y(n_699) );
INVxp67_ASAP7_75t_SL g710 ( .A(n_628), .Y(n_710) );
OR2x2_ASAP7_75t_L g761 ( .A(n_628), .B(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g816 ( .A(n_628), .Y(n_816) );
AOI211xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_634), .B(n_640), .C(n_649), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g705 ( .A(n_633), .B(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_633), .B(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_L g778 ( .A(n_633), .B(n_655), .Y(n_778) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_638), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_636), .B(n_681), .Y(n_703) );
NAND2x1p5_ASAP7_75t_L g720 ( .A(n_636), .B(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g788 ( .A(n_636), .B(n_789), .Y(n_788) );
INVx3_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
BUFx2_ASAP7_75t_L g731 ( .A(n_637), .Y(n_731) );
AND2x2_ASAP7_75t_L g759 ( .A(n_638), .B(n_687), .Y(n_759) );
INVx2_ASAP7_75t_L g782 ( .A(n_638), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_638), .B(n_680), .Y(n_814) );
AND2x4_ASAP7_75t_SL g768 ( .A(n_641), .B(n_646), .Y(n_768) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g721 ( .A(n_642), .B(n_647), .Y(n_721) );
OR2x2_ASAP7_75t_L g773 ( .A(n_642), .B(n_666), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_643), .B(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_643), .B(n_655), .Y(n_809) );
BUFx3_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g757 ( .A(n_644), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_648), .Y(n_645) );
INVx1_ASAP7_75t_L g740 ( .A(n_646), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_646), .B(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g790 ( .A(n_647), .Y(n_790) );
BUFx2_ASAP7_75t_L g658 ( .A(n_648), .Y(n_658) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g776 ( .A(n_651), .B(n_777), .Y(n_776) );
OR2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g700 ( .A(n_655), .Y(n_700) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_655), .Y(n_717) );
NAND3xp33_ASAP7_75t_SL g656 ( .A(n_657), .B(n_667), .C(n_682), .Y(n_656) );
AOI22xp33_ASAP7_75t_SL g657 ( .A1(n_658), .A2(n_659), .B1(n_662), .B2(n_664), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AOI222xp33_ASAP7_75t_L g770 ( .A1(n_664), .A2(n_690), .B1(n_771), .B2(n_774), .C1(n_776), .C2(n_778), .Y(n_770) );
AND2x2_ASAP7_75t_L g802 ( .A(n_665), .B(n_751), .Y(n_802) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OR2x2_ASAP7_75t_L g750 ( .A(n_666), .B(n_751), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_673), .B1(n_674), .B2(n_679), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
INVx2_ASAP7_75t_SL g746 ( .A(n_670), .Y(n_746) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_678), .Y(n_674) );
AND2x2_ASAP7_75t_L g733 ( .A(n_675), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g691 ( .A(n_676), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OR2x2_ASAP7_75t_L g685 ( .A(n_677), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g800 ( .A(n_678), .Y(n_800) );
AND2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_681), .B(n_777), .Y(n_796) );
INVx1_ASAP7_75t_L g813 ( .A(n_681), .Y(n_813) );
AOI222xp33_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_687), .B1(n_688), .B2(n_690), .C1(n_693), .C2(n_694), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_689), .Y(n_693) );
AND2x2_ASAP7_75t_L g711 ( .A(n_689), .B(n_712), .Y(n_711) );
INVx3_ASAP7_75t_L g742 ( .A(n_689), .Y(n_742) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx2_ASAP7_75t_L g706 ( .A(n_692), .Y(n_706) );
OR2x2_ASAP7_75t_L g775 ( .A(n_692), .B(n_756), .Y(n_775) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
OAI211xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_701), .B(n_704), .C(n_713), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
OAI21xp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_707), .B(n_711), .Y(n_704) );
AOI221xp5_ASAP7_75t_L g791 ( .A1(n_705), .A2(n_743), .B1(n_792), .B2(n_795), .C(n_797), .Y(n_791) );
AND2x4_ASAP7_75t_L g734 ( .A(n_706), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
INVx1_ASAP7_75t_L g765 ( .A(n_712), .Y(n_765) );
AOI211x1_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_716), .B(n_718), .C(n_722), .Y(n_713) );
INVxp67_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g783 ( .A(n_721), .Y(n_783) );
NAND3xp33_ASAP7_75t_L g771 ( .A(n_724), .B(n_772), .C(n_773), .Y(n_771) );
OR2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
INVx1_ASAP7_75t_L g807 ( .A(n_725), .Y(n_807) );
NOR2x1_ASAP7_75t_L g727 ( .A(n_728), .B(n_779), .Y(n_727) );
NAND4xp25_ASAP7_75t_L g728 ( .A(n_729), .B(n_736), .C(n_758), .D(n_770), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_733), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
AND2x2_ASAP7_75t_L g789 ( .A(n_732), .B(n_790), .Y(n_789) );
AOI221x1_ASAP7_75t_L g758 ( .A1(n_734), .A2(n_759), .B1(n_760), .B2(n_763), .C(n_766), .Y(n_758) );
AND2x2_ASAP7_75t_L g784 ( .A(n_734), .B(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g794 ( .A(n_735), .Y(n_794) );
AOI221xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_739), .B1(n_743), .B2(n_747), .C(n_749), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_741), .B(n_765), .Y(n_764) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
OR2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_746), .A2(n_750), .B1(n_753), .B2(n_755), .Y(n_749) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g766 ( .A1(n_750), .A2(n_767), .B(n_769), .Y(n_766) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g772 ( .A(n_752), .Y(n_772) );
OR2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVxp67_ASAP7_75t_L g793 ( .A(n_762), .Y(n_793) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
OAI22xp33_ASAP7_75t_L g812 ( .A1(n_775), .A2(n_813), .B1(n_814), .B2(n_815), .Y(n_812) );
NAND3xp33_ASAP7_75t_L g779 ( .A(n_780), .B(n_791), .C(n_803), .Y(n_779) );
AOI22xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_784), .B1(n_787), .B2(n_788), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_782), .B(n_783), .Y(n_781) );
INVxp67_ASAP7_75t_SL g785 ( .A(n_786), .Y(n_785) );
OR2x2_ASAP7_75t_L g799 ( .A(n_786), .B(n_800), .Y(n_799) );
NAND2x1_ASAP7_75t_L g815 ( .A(n_786), .B(n_816), .Y(n_815) );
AND2x2_ASAP7_75t_L g792 ( .A(n_793), .B(n_794), .Y(n_792) );
INVx2_ASAP7_75t_SL g795 ( .A(n_796), .Y(n_795) );
AOI21xp5_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_799), .B(n_801), .Y(n_797) );
INVx1_ASAP7_75t_SL g801 ( .A(n_802), .Y(n_801) );
AOI221xp5_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_807), .B1(n_808), .B2(n_810), .C(n_812), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx3_ASAP7_75t_R g810 ( .A(n_811), .Y(n_810) );
INVx4_ASAP7_75t_L g820 ( .A(n_817), .Y(n_820) );
BUFx12f_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
CKINVDCx5p33_ASAP7_75t_R g818 ( .A(n_819), .Y(n_818) );
AND2x2_ASAP7_75t_L g834 ( .A(n_819), .B(n_835), .Y(n_834) );
CKINVDCx5p33_ASAP7_75t_R g827 ( .A(n_821), .Y(n_827) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
BUFx10_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
NOR2xp33_ASAP7_75t_L g836 ( .A(n_837), .B(n_838), .Y(n_836) );
BUFx6f_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
endmodule