module fake_jpeg_27572_n_287 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_287);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_287;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_21;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx13_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_29),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_31),
.Y(n_44)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_33),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_25),
.B(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_46),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_39),
.A2(n_42),
.B(n_45),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_13),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_25),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_46),
.B(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_49),
.B(n_61),
.Y(n_82)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_55),
.Y(n_68)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_33),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_58),
.Y(n_70)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_23),
.Y(n_61)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_44),
.B(n_23),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_64),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_15),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_45),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_67),
.B1(n_43),
.B2(n_36),
.Y(n_77)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_31),
.B1(n_29),
.B2(n_26),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_69),
.A2(n_84),
.B1(n_55),
.B2(n_85),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_62),
.B(n_39),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_71),
.B(n_73),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_37),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_37),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_74),
.B(n_79),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_77),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_59),
.B(n_26),
.Y(n_78)
);

AO21x1_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_86),
.B(n_45),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_42),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_51),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_31),
.B1(n_29),
.B2(n_35),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_45),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_67),
.A2(n_20),
.B1(n_13),
.B2(n_18),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_87),
.A2(n_14),
.B1(n_36),
.B2(n_16),
.Y(n_95)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_88),
.B(n_94),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_42),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_90),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_93),
.Y(n_118)
);

NOR2x1_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_34),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_57),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_101),
.B1(n_78),
.B2(n_85),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_96),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_71),
.A2(n_32),
.B(n_12),
.C(n_17),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_99),
.A2(n_100),
.B(n_78),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_71),
.A2(n_32),
.B(n_12),
.C(n_17),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_52),
.Y(n_102)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

AO22x1_ASAP7_75t_SL g103 ( 
.A1(n_69),
.A2(n_16),
.B1(n_34),
.B2(n_41),
.Y(n_103)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_52),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_104),
.B(n_106),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_72),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_107),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_73),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_22),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_98),
.A2(n_74),
.B1(n_80),
.B2(n_86),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_119),
.B1(n_120),
.B2(n_97),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_86),
.B1(n_78),
.B2(n_84),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_92),
.B1(n_89),
.B2(n_107),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_91),
.A2(n_80),
.B1(n_15),
.B2(n_25),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_112),
.A2(n_114),
.B(n_115),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_117),
.B(n_124),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_98),
.A2(n_91),
.B1(n_106),
.B2(n_88),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_96),
.A2(n_68),
.B1(n_75),
.B2(n_83),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_127),
.Y(n_134)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_96),
.B(n_72),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_83),
.B(n_75),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_81),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_128),
.Y(n_138)
);

INVx4_ASAP7_75t_SL g127 ( 
.A(n_103),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_97),
.C(n_92),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_118),
.C(n_129),
.Y(n_156)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_136),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_133),
.B(n_140),
.Y(n_159)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_137),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_171)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_109),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_144),
.Y(n_165)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_90),
.Y(n_145)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_100),
.B(n_99),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_146),
.A2(n_129),
.B(n_25),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_100),
.Y(n_147)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_151),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_99),
.Y(n_149)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_150),
.A2(n_25),
.B(n_34),
.Y(n_163)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_127),
.A2(n_81),
.B1(n_14),
.B2(n_15),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_112),
.B1(n_128),
.B2(n_126),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_155),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_164),
.C(n_173),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_SL g193 ( 
.A(n_158),
.B(n_162),
.C(n_168),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_163),
.A2(n_175),
.B(n_139),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_41),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_138),
.A2(n_16),
.B1(n_15),
.B2(n_72),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_166),
.A2(n_38),
.B1(n_17),
.B2(n_19),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_23),
.B1(n_20),
.B2(n_13),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_135),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_171),
.A2(n_146),
.B1(n_150),
.B2(n_12),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_41),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_145),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_174),
.B(n_178),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_144),
.A2(n_12),
.B(n_13),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_SL g176 ( 
.A1(n_154),
.A2(n_155),
.B(n_138),
.C(n_153),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_176),
.A2(n_139),
.B(n_66),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_141),
.B(n_143),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_149),
.Y(n_181)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_184),
.Y(n_203)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_187),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_161),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_186),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_169),
.B(n_135),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_160),
.B(n_147),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_188),
.B(n_199),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_151),
.Y(n_189)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_180),
.B(n_159),
.C(n_172),
.Y(n_190)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_198),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_192),
.A2(n_179),
.B1(n_193),
.B2(n_183),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_194),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_195),
.A2(n_200),
.B(n_201),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_54),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_157),
.B(n_177),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_173),
.B(n_11),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_163),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_175),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_192),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_204),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_196),
.B(n_156),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_205),
.B(n_41),
.Y(n_235)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_195),
.A2(n_179),
.B1(n_176),
.B2(n_164),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_210),
.A2(n_181),
.B1(n_189),
.B2(n_193),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_176),
.C(n_162),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_216),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_176),
.C(n_54),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_51),
.C(n_41),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_220),
.B(n_194),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_222),
.A2(n_225),
.B1(n_234),
.B2(n_212),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_224),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_206),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_210),
.A2(n_190),
.B1(n_198),
.B2(n_185),
.Y(n_225)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_201),
.Y(n_229)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_218),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_232),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_219),
.A2(n_213),
.B(n_217),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_207),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_51),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_235),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_221),
.A2(n_18),
.B1(n_21),
.B2(n_20),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_227),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_241),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_225),
.A2(n_203),
.B1(n_208),
.B2(n_217),
.Y(n_239)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_239),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_216),
.C(n_220),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_214),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_247),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_245),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_212),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_19),
.C(n_21),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_21),
.C(n_18),
.Y(n_256)
);

OAI21xp33_ASAP7_75t_L g252 ( 
.A1(n_238),
.A2(n_228),
.B(n_223),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_255),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_248),
.A2(n_8),
.B(n_10),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_253),
.A2(n_4),
.B(n_9),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_19),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_257),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_21),
.C(n_18),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_237),
.C(n_242),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_260),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_239),
.C(n_24),
.Y(n_260)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_261),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_254),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_265),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_250),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_260),
.B(n_4),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_267),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_5),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_5),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_269),
.B(n_0),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_268),
.B(n_5),
.C(n_9),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_274),
.C(n_272),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_263),
.A2(n_6),
.B1(n_10),
.B2(n_2),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_0),
.C(n_1),
.Y(n_278)
);

OAI21x1_ASAP7_75t_L g276 ( 
.A1(n_275),
.A2(n_262),
.B(n_261),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_277),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_272),
.C(n_273),
.Y(n_279)
);

FAx1_ASAP7_75t_SL g281 ( 
.A(n_279),
.B(n_0),
.CI(n_1),
.CON(n_281),
.SN(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_280),
.C(n_1),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_281),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_283),
.A2(n_0),
.B(n_1),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_284),
.A2(n_2),
.B(n_3),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_2),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_286),
.A2(n_3),
.B(n_263),
.Y(n_287)
);


endmodule