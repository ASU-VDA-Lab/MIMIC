module fake_jpeg_6856_n_228 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_228);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_7),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_33),
.B(n_36),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_7),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_7),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_42),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_45),
.B(n_50),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_29),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_28),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_55),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_18),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_64),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_19),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_27),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_22),
.B1(n_26),
.B2(n_25),
.Y(n_59)
);

NAND2xp33_ASAP7_75t_SL g85 ( 
.A(n_59),
.B(n_60),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_26),
.B1(n_22),
.B2(n_20),
.Y(n_60)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_22),
.B1(n_26),
.B2(n_15),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_20),
.B1(n_23),
.B2(n_28),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_19),
.Y(n_64)
);

AOI21xp33_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_37),
.B(n_24),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_66),
.A2(n_82),
.B(n_21),
.Y(n_100)
);

NAND3xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_32),
.C(n_23),
.Y(n_68)
);

OR2x4_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_63),
.Y(n_93)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_79),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_49),
.B1(n_60),
.B2(n_48),
.Y(n_90)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_31),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_72),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_31),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_74),
.Y(n_99)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_76),
.B(n_83),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_31),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_77),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_54),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_32),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_75),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_27),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_17),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_84),
.B(n_44),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_90),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_75),
.B(n_44),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_75),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_81),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_78),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_59),
.B(n_52),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_94),
.A2(n_100),
.B(n_84),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_85),
.A2(n_53),
.B1(n_58),
.B2(n_52),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_103),
.Y(n_114)
);

AO22x1_ASAP7_75t_SL g97 ( 
.A1(n_66),
.A2(n_38),
.B1(n_61),
.B2(n_47),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_97),
.A2(n_98),
.B1(n_101),
.B2(n_105),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_70),
.A2(n_61),
.B1(n_58),
.B2(n_62),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_70),
.A2(n_61),
.B1(n_58),
.B2(n_43),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_43),
.C(n_53),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_77),
.C(n_74),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_80),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_69),
.A2(n_53),
.B1(n_38),
.B2(n_47),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_78),
.A2(n_47),
.B1(n_27),
.B2(n_24),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_106),
.A2(n_76),
.B1(n_71),
.B2(n_83),
.Y(n_122)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_47),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_122),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_117),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_89),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_115),
.B(n_73),
.Y(n_134)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_121),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_102),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_82),
.Y(n_118)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

OAI22x1_ASAP7_75t_SL g120 ( 
.A1(n_97),
.A2(n_68),
.B1(n_82),
.B2(n_78),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_120),
.A2(n_129),
.B1(n_94),
.B2(n_91),
.Y(n_132)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_97),
.A2(n_76),
.B1(n_80),
.B2(n_72),
.Y(n_123)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_128),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_73),
.Y(n_125)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_126),
.B(n_106),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_107),
.C(n_87),
.Y(n_142)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_129),
.A2(n_100),
.B(n_108),
.Y(n_133)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_107),
.Y(n_139)
);

NOR3xp33_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_133),
.C(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_144),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_114),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_140),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_143),
.C(n_127),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_87),
.C(n_99),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_148),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_121),
.B(n_104),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_150),
.Y(n_167)
);

OAI32xp33_ASAP7_75t_L g150 ( 
.A1(n_111),
.A2(n_110),
.A3(n_128),
.B1(n_130),
.B2(n_123),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_99),
.B(n_98),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_151),
.A2(n_119),
.B1(n_124),
.B2(n_109),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_158),
.C(n_162),
.Y(n_176)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_165),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_139),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_143),
.C(n_112),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_159),
.A2(n_168),
.B1(n_147),
.B2(n_149),
.Y(n_173)
);

AO221x1_ASAP7_75t_L g161 ( 
.A1(n_134),
.A2(n_67),
.B1(n_24),
.B2(n_27),
.C(n_21),
.Y(n_161)
);

AO221x1_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_148),
.B1(n_135),
.B2(n_17),
.C(n_3),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_109),
.C(n_122),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_126),
.C(n_90),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_164),
.C(n_78),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_142),
.C(n_137),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_137),
.A2(n_126),
.B1(n_65),
.B2(n_103),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_131),
.A2(n_79),
.B1(n_65),
.B2(n_24),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_140),
.B1(n_131),
.B2(n_141),
.Y(n_175)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_174),
.Y(n_185)
);

O2A1O1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_171),
.A2(n_175),
.B(n_178),
.C(n_183),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_154),
.B(n_150),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_172),
.A2(n_173),
.B(n_6),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_180),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_167),
.A2(n_144),
.B1(n_146),
.B2(n_141),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_0),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_165),
.B(n_135),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_182),
.C(n_155),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_13),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_167),
.A2(n_163),
.B1(n_162),
.B2(n_164),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_152),
.Y(n_187)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_187),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_192),
.C(n_1),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_189),
.B(n_170),
.Y(n_198)
);

NAND3xp33_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_168),
.C(n_160),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_190),
.A2(n_196),
.B(n_179),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_153),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_191),
.A2(n_194),
.B(n_195),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_166),
.C(n_153),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_0),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_198),
.B(n_200),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_193),
.A2(n_183),
.B1(n_173),
.B2(n_181),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_201),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_195),
.A2(n_180),
.B1(n_176),
.B2(n_182),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_202),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_193),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_204),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_190),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_8),
.C(n_12),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_204),
.B(n_185),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_207),
.A2(n_197),
.B(n_203),
.Y(n_214)
);

AOI31xp67_ASAP7_75t_L g210 ( 
.A1(n_200),
.A2(n_8),
.A3(n_12),
.B(n_11),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_5),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_211),
.B(n_5),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_212),
.A2(n_205),
.B(n_10),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_206),
.B(n_199),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_213),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_214),
.A2(n_215),
.B(n_212),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_208),
.A2(n_201),
.B1(n_4),
.B2(n_3),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_216),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_217),
.A2(n_218),
.B(n_209),
.Y(n_219)
);

AOI322xp5_ASAP7_75t_L g223 ( 
.A1(n_219),
.A2(n_222),
.A3(n_207),
.B1(n_216),
.B2(n_9),
.C1(n_10),
.C2(n_12),
.Y(n_223)
);

OAI21x1_ASAP7_75t_L g226 ( 
.A1(n_223),
.A2(n_224),
.B(n_13),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_6),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_220),
.Y(n_225)
);

O2A1O1Ixp33_ASAP7_75t_SL g227 ( 
.A1(n_225),
.A2(n_4),
.B(n_13),
.C(n_211),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_227),
.Y(n_228)
);


endmodule