module fake_jpeg_7745_n_204 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_5),
.B(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_32),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_35),
.Y(n_59)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_27),
.Y(n_34)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_22),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_18),
.B(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_39),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_46),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_31),
.A2(n_20),
.B1(n_27),
.B2(n_23),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_53),
.B1(n_57),
.B2(n_38),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_51),
.Y(n_73)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_31),
.A2(n_27),
.B1(n_23),
.B2(n_22),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_32),
.A2(n_26),
.B1(n_30),
.B2(n_28),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_41),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_41),
.B1(n_40),
.B2(n_29),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_60),
.A2(n_33),
.B1(n_15),
.B2(n_28),
.Y(n_69)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_74),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_57),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_66),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_64),
.B(n_67),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_33),
.B1(n_54),
.B2(n_47),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_65),
.A2(n_69),
.B1(n_72),
.B2(n_15),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_35),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_59),
.B(n_50),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_70),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_56),
.A2(n_21),
.B1(n_16),
.B2(n_19),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_63),
.A2(n_43),
.B(n_55),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_82),
.B(n_73),
.Y(n_111)
);

BUFx10_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_55),
.B(n_60),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_89),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_65),
.A2(n_60),
.B1(n_54),
.B2(n_47),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_86),
.B1(n_70),
.B2(n_45),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_60),
.B1(n_54),
.B2(n_52),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_87),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_90),
.A2(n_91),
.B1(n_58),
.B2(n_75),
.Y(n_108)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

AO21x1_ASAP7_75t_L g102 ( 
.A1(n_94),
.A2(n_95),
.B(n_96),
.Y(n_102)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

NAND3xp33_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_51),
.C(n_14),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_62),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_107),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_74),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_21),
.C(n_30),
.Y(n_130)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_99),
.B(n_104),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_91),
.Y(n_127)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_64),
.Y(n_107)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_109),
.A2(n_110),
.B1(n_112),
.B2(n_93),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_78),
.A2(n_75),
.B1(n_16),
.B2(n_19),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_111),
.A2(n_104),
.B(n_107),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_82),
.A2(n_73),
.B1(n_71),
.B2(n_49),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_113),
.B(n_114),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_88),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_92),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_129),
.C(n_130),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_118),
.B(n_103),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_119),
.A2(n_121),
.B(n_99),
.Y(n_137)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_120),
.B(n_125),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_111),
.A2(n_112),
.B(n_105),
.Y(n_121)
);

NAND3xp33_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_95),
.C(n_92),
.Y(n_122)
);

OAI322xp33_ASAP7_75t_L g144 ( 
.A1(n_122),
.A2(n_124),
.A3(n_42),
.B1(n_29),
.B2(n_25),
.C1(n_6),
.C2(n_7),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_83),
.C(n_93),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_106),
.Y(n_125)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_131),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_49),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_113),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_133),
.B(n_137),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_103),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_147),
.C(n_2),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_135),
.A2(n_140),
.B(n_123),
.Y(n_156)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_143),
.Y(n_161)
);

A2O1A1O1Ixp25_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_102),
.B(n_42),
.C(n_29),
.D(n_25),
.Y(n_140)
);

OAI32xp33_ASAP7_75t_L g141 ( 
.A1(n_132),
.A2(n_102),
.A3(n_29),
.B1(n_25),
.B2(n_5),
.Y(n_141)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_117),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_144),
.B(n_148),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_25),
.Y(n_146)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_146),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_42),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_129),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_150),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_119),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_123),
.B1(n_100),
.B2(n_90),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_151),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_135),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_156),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_130),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_142),
.C(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_158),
.A2(n_162),
.B1(n_136),
.B2(n_146),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_145),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_165),
.Y(n_177)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_164),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_172),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_161),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_171),
.Y(n_182)
);

XNOR2x1_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_142),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_169),
.A2(n_173),
.B(n_149),
.Y(n_180)
);

NAND3xp33_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_2),
.C(n_3),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_101),
.C(n_100),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_174),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_163),
.A2(n_160),
.B1(n_150),
.B2(n_100),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_170),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_8),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_181),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_80),
.B(n_6),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_167),
.C(n_7),
.Y(n_184)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

AOI322xp5_ASAP7_75t_L g186 ( 
.A1(n_175),
.A2(n_170),
.A3(n_166),
.B1(n_172),
.B2(n_80),
.C1(n_11),
.C2(n_4),
.Y(n_186)
);

AOI21xp33_ASAP7_75t_L g192 ( 
.A1(n_186),
.A2(n_182),
.B(n_183),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_187),
.A2(n_189),
.B(n_177),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_4),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_190),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_8),
.C(n_9),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_192),
.A2(n_188),
.B(n_10),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_9),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_179),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_194),
.C(n_186),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_196),
.A2(n_197),
.B(n_199),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_198),
.B(n_12),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_10),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_13),
.Y(n_203)
);

AO21x1_ASAP7_75t_L g202 ( 
.A1(n_201),
.A2(n_195),
.B(n_13),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_203),
.Y(n_204)
);


endmodule