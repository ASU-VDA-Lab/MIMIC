module fake_jpeg_15983_n_24 (n_3, n_2, n_1, n_0, n_4, n_24);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_24;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g5 ( 
.A(n_4),
.Y(n_5)
);

INVx4_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_0),
.Y(n_7)
);

INVx6_ASAP7_75t_SL g8 ( 
.A(n_3),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_6),
.B(n_1),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_10),
.B(n_11),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_6),
.B(n_2),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_12),
.B(n_13),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g13 ( 
.A1(n_5),
.A2(n_2),
.B1(n_3),
.B2(n_9),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_16),
.A2(n_5),
.B1(n_11),
.B2(n_10),
.Y(n_18)
);

BUFx24_ASAP7_75t_SL g20 ( 
.A(n_18),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_20),
.B(n_15),
.Y(n_21)
);

BUFx24_ASAP7_75t_SL g23 ( 
.A(n_21),
.Y(n_23)
);

AOI322xp5_ASAP7_75t_L g22 ( 
.A1(n_19),
.A2(n_7),
.A3(n_8),
.B1(n_14),
.B2(n_17),
.C1(n_20),
.C2(n_18),
.Y(n_22)
);

NOR2x1_ASAP7_75t_L g24 ( 
.A(n_23),
.B(n_22),
.Y(n_24)
);


endmodule