module fake_jpeg_19763_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_24),
.B(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_31),
.Y(n_48)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_24),
.B1(n_17),
.B2(n_18),
.Y(n_46)
);

OAI21xp33_ASAP7_75t_L g92 ( 
.A1(n_46),
.A2(n_23),
.B(n_20),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_48),
.Y(n_66)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_18),
.B1(n_17),
.B2(n_27),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_51),
.A2(n_33),
.B1(n_34),
.B2(n_21),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_55),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_25),
.C(n_21),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_65),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_22),
.B1(n_27),
.B2(n_21),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_59),
.A2(n_53),
.B1(n_64),
.B2(n_60),
.Y(n_85)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_38),
.B(n_33),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_34),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_22),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_44),
.B1(n_39),
.B2(n_35),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_70),
.A2(n_76),
.B1(n_79),
.B2(n_83),
.Y(n_118)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_65),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_80),
.Y(n_105)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_53),
.A2(n_44),
.B1(n_36),
.B2(n_40),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_77),
.B(n_81),
.Y(n_95)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_55),
.A2(n_40),
.B1(n_42),
.B2(n_41),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_65),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_48),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_92),
.B1(n_62),
.B2(n_52),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_52),
.A2(n_42),
.B1(n_41),
.B2(n_43),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_84),
.B(n_87),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_46),
.B1(n_52),
.B2(n_62),
.Y(n_102)
);

INVxp33_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_58),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_99),
.B(n_106),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

INVxp67_ASAP7_75t_SL g131 ( 
.A(n_101),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_83),
.B1(n_78),
.B2(n_89),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_60),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_0),
.B(n_1),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_0),
.B(n_1),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_113),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_62),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_110),
.B(n_112),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_80),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_67),
.Y(n_113)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_66),
.B(n_81),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_23),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_47),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_91),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_69),
.A2(n_20),
.B1(n_16),
.B2(n_61),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_120),
.A2(n_87),
.B1(n_84),
.B2(n_89),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_123),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_110),
.B(n_66),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_128),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_126),
.A2(n_137),
.B1(n_144),
.B2(n_148),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_127),
.A2(n_134),
.B1(n_116),
.B2(n_96),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_93),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_97),
.A2(n_75),
.B1(n_74),
.B2(n_71),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_129),
.A2(n_133),
.B(n_100),
.Y(n_161)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_135),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_102),
.A2(n_83),
.B1(n_90),
.B2(n_68),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_98),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_136),
.B(n_142),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_83),
.B1(n_47),
.B2(n_45),
.Y(n_137)
);

NOR2x1_ASAP7_75t_SL g138 ( 
.A(n_112),
.B(n_23),
.Y(n_138)
);

XOR2x2_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_120),
.Y(n_157)
);

OA21x2_ASAP7_75t_L g139 ( 
.A1(n_105),
.A2(n_45),
.B(n_47),
.Y(n_139)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_118),
.A2(n_43),
.B1(n_41),
.B2(n_45),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_23),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_107),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_121),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_118),
.A2(n_43),
.B1(n_56),
.B2(n_32),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_61),
.B1(n_32),
.B2(n_30),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_94),
.B1(n_114),
.B2(n_3),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_140),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_151),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_105),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_152),
.A2(n_157),
.B(n_139),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_106),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_153),
.B(n_162),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_95),
.C(n_108),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_167),
.C(n_172),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_134),
.A2(n_95),
.B1(n_119),
.B2(n_111),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_160),
.A2(n_170),
.B1(n_173),
.B2(n_141),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_182),
.B(n_147),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_111),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_143),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_166),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_113),
.C(n_115),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_125),
.Y(n_168)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_171),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_115),
.C(n_103),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_127),
.A2(n_114),
.B1(n_103),
.B2(n_96),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_115),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_4),
.C(n_5),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_94),
.C(n_114),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_181),
.C(n_141),
.Y(n_192)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_123),
.Y(n_176)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_176),
.Y(n_202)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_179),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_211)
);

AOI22x1_ASAP7_75t_L g180 ( 
.A1(n_138),
.A2(n_23),
.B1(n_30),
.B2(n_32),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_180),
.A2(n_28),
.B1(n_3),
.B2(n_4),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_129),
.B(n_142),
.C(n_139),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_130),
.A2(n_133),
.B(n_131),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_144),
.Y(n_190)
);

NAND3xp33_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_15),
.C(n_14),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_184),
.B(n_190),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_161),
.A2(n_126),
.B(n_136),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_185),
.A2(n_188),
.B(n_193),
.Y(n_225)
);

OAI32xp33_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_137),
.A3(n_150),
.B1(n_139),
.B2(n_148),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_208),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_189),
.A2(n_152),
.B(n_178),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_212),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_157),
.A2(n_135),
.B(n_132),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_169),
.A2(n_159),
.B1(n_181),
.B2(n_167),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_194),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_153),
.C(n_162),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_154),
.C(n_175),
.Y(n_219)
);

BUFx24_ASAP7_75t_SL g198 ( 
.A(n_174),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_168),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_199),
.A2(n_201),
.B1(n_203),
.B2(n_179),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_170),
.A2(n_14),
.B1(n_2),
.B2(n_3),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_173),
.A2(n_14),
.B1(n_2),
.B2(n_3),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_169),
.A2(n_30),
.B1(n_25),
.B2(n_26),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_172),
.A2(n_28),
.B1(n_26),
.B2(n_16),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_163),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_152),
.B(n_1),
.Y(n_210)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_210),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_211),
.Y(n_229)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_209),
.B(n_155),
.Y(n_216)
);

XNOR2x1_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_224),
.Y(n_241)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_217),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_234),
.Y(n_240)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_197),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_221),
.Y(n_244)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

OAI21xp33_ASAP7_75t_SL g224 ( 
.A1(n_210),
.A2(n_182),
.B(n_180),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_186),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_230),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_227),
.A2(n_194),
.B1(n_205),
.B2(n_187),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_186),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_232),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_202),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_202),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_235),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_183),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_200),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_238),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_191),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_199),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_200),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_158),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_239),
.B(n_238),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_230),
.Y(n_243)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_246),
.A2(n_247),
.B1(n_214),
.B2(n_201),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_218),
.A2(n_227),
.B1(n_229),
.B2(n_222),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_191),
.C(n_192),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_254),
.C(n_256),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_225),
.A2(n_185),
.B(n_193),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_258),
.Y(n_264)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_252),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_188),
.C(n_189),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_180),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_206),
.C(n_212),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_219),
.B(n_195),
.C(n_190),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_260),
.C(n_216),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_214),
.B(n_195),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_164),
.C(n_208),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_225),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_263),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_248),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_255),
.A2(n_218),
.B1(n_231),
.B2(n_226),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_266),
.A2(n_246),
.B1(n_244),
.B2(n_241),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_203),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_215),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_271),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_241),
.B(n_222),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_274),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_253),
.B(n_223),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_276),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_232),
.Y(n_273)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_217),
.C(n_220),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_260),
.C(n_267),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_221),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_156),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_4),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_245),
.Y(n_278)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_282),
.C(n_265),
.Y(n_294)
);

INVx3_ASAP7_75t_SL g281 ( 
.A(n_264),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_285),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_244),
.C(n_251),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_247),
.Y(n_283)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_283),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_268),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_262),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_270),
.A2(n_249),
.B(n_242),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_287),
.A2(n_274),
.B(n_7),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_279),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_6),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_295),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_265),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_298),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_263),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_302),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_6),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_301),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_288),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_303),
.A2(n_305),
.B1(n_7),
.B2(n_8),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_282),
.C(n_284),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_290),
.C(n_287),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_284),
.Y(n_306)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_306),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_295),
.Y(n_308)
);

A2O1A1Ixp33_ASAP7_75t_L g318 ( 
.A1(n_308),
.A2(n_300),
.B(n_293),
.C(n_296),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_310),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_304),
.A2(n_289),
.B(n_279),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_10),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_7),
.C(n_9),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_9),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_321),
.B(n_306),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_9),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_319),
.B(n_320),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_312),
.Y(n_321)
);

OAI21xp33_ASAP7_75t_L g324 ( 
.A1(n_322),
.A2(n_307),
.B(n_11),
.Y(n_324)
);

O2A1O1Ixp33_ASAP7_75t_SL g326 ( 
.A1(n_324),
.A2(n_325),
.B(n_314),
.C(n_320),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_316),
.C(n_309),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_327),
.A2(n_317),
.B(n_323),
.Y(n_328)
);

NOR3xp33_ASAP7_75t_SL g329 ( 
.A(n_328),
.B(n_311),
.C(n_11),
.Y(n_329)
);

AOI33xp33_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_311),
.B3(n_286),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_11),
.B(n_12),
.Y(n_331)
);


endmodule