module fake_jpeg_16110_n_290 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_290);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_102;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_7),
.B(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_7),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_18),
.B1(n_19),
.B2(n_22),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_53),
.B1(n_31),
.B2(n_34),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_38),
.Y(n_64)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_17),
.C(n_18),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_30),
.Y(n_73)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_34),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_31),
.A2(n_18),
.B1(n_19),
.B2(n_22),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_38),
.B(n_24),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_55),
.B(n_24),
.Y(n_77)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_58),
.A2(n_37),
.B1(n_40),
.B2(n_50),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_60),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_61),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_48),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_67),
.B1(n_73),
.B2(n_79),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_28),
.B1(n_20),
.B2(n_22),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_55),
.A2(n_31),
.B1(n_34),
.B2(n_38),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_51),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_69),
.B(n_71),
.Y(n_88)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_56),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_24),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_20),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_74),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_77),
.B(n_30),
.Y(n_95)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_47),
.A2(n_31),
.B1(n_34),
.B2(n_37),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_85),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_39),
.C(n_35),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_39),
.C(n_35),
.Y(n_89)
);

FAx1_ASAP7_75t_SL g128 ( 
.A(n_89),
.B(n_101),
.CI(n_32),
.CON(n_128),
.SN(n_128)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_73),
.A2(n_28),
.B1(n_20),
.B2(n_16),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_0),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_91),
.A2(n_100),
.B(n_30),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_92),
.A2(n_57),
.B1(n_78),
.B2(n_54),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_104),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_77),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_40),
.B1(n_49),
.B2(n_37),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_96),
.A2(n_37),
.B1(n_54),
.B2(n_32),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_0),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_39),
.C(n_35),
.Y(n_101)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_65),
.B1(n_64),
.B2(n_40),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_110),
.B1(n_112),
.B2(n_122),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_59),
.B1(n_62),
.B2(n_80),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_111),
.B(n_113),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_62),
.B1(n_80),
.B2(n_37),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_84),
.B(n_66),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_114),
.B(n_118),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_83),
.B(n_23),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_115),
.B(n_121),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_81),
.A2(n_39),
.B(n_0),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_119),
.B(n_120),
.Y(n_147)
);

OAI32xp33_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_62),
.A3(n_26),
.B1(n_23),
.B2(n_29),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_88),
.A2(n_16),
.B(n_29),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_39),
.B(n_1),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_87),
.Y(n_121)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_103),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_126),
.Y(n_136)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_127),
.A2(n_94),
.B1(n_98),
.B2(n_86),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_101),
.Y(n_138)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_89),
.A2(n_54),
.B1(n_33),
.B2(n_32),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_132),
.A2(n_33),
.B1(n_52),
.B2(n_43),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_85),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_138),
.C(n_140),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_128),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_143),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_139),
.A2(n_148),
.B1(n_159),
.B2(n_160),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_90),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_118),
.Y(n_143)
);

XNOR2x2_ASAP7_75t_SL g144 ( 
.A(n_116),
.B(n_91),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_119),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_112),
.A2(n_110),
.B1(n_107),
.B2(n_132),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_145),
.A2(n_149),
.B1(n_155),
.B2(n_61),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_131),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_146),
.B(n_156),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_126),
.A2(n_104),
.B1(n_97),
.B2(n_82),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_107),
.A2(n_82),
.B1(n_33),
.B2(n_106),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_108),
.B(n_76),
.C(n_39),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_61),
.C(n_21),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_91),
.Y(n_152)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_127),
.A2(n_33),
.B1(n_97),
.B2(n_52),
.Y(n_155)
);

INVx13_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_161),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_100),
.B1(n_16),
.B2(n_15),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_120),
.A2(n_27),
.B1(n_26),
.B2(n_23),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_109),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_136),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_168),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_188),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_165),
.B(n_160),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_158),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_39),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_182),
.C(n_186),
.Y(n_197)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_172),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_189),
.Y(n_201)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_134),
.A2(n_27),
.B1(n_26),
.B2(n_15),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_176),
.A2(n_187),
.B(n_147),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_139),
.A2(n_29),
.B1(n_27),
.B2(n_15),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_177),
.A2(n_183),
.B1(n_21),
.B2(n_3),
.Y(n_209)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_179),
.Y(n_212)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_39),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_143),
.A2(n_21),
.B1(n_52),
.B2(n_68),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_184),
.Y(n_191)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_185),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_137),
.A2(n_1),
.B(n_61),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_141),
.B(n_152),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_21),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_133),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_200),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_198),
.A2(n_166),
.B(n_163),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_147),
.C(n_144),
.Y(n_200)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_188),
.A2(n_159),
.B1(n_1),
.B2(n_3),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_203),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_21),
.Y(n_205)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_205),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_208),
.A2(n_187),
.B(n_164),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_210),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_2),
.C(n_3),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_2),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

NOR2x1_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_176),
.Y(n_215)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_171),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_219),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_218),
.B(n_198),
.Y(n_235)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_192),
.A2(n_190),
.B(n_173),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_220),
.A2(n_228),
.B(n_212),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_204),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_222),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_206),
.B(n_165),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_203),
.A2(n_186),
.B1(n_182),
.B2(n_168),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_225),
.A2(n_229),
.B1(n_230),
.B2(n_215),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_174),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_205),
.Y(n_238)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_207),
.A2(n_5),
.B(n_9),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_195),
.C(n_197),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_232),
.C(n_239),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_197),
.C(n_200),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_210),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_235),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_216),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_242),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_238),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_202),
.Y(n_239)
);

FAx1_ASAP7_75t_SL g240 ( 
.A(n_227),
.B(n_211),
.CI(n_191),
.CON(n_240),
.SN(n_240)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_240),
.B(n_214),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_196),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_238),
.C(n_241),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_243),
.A2(n_230),
.B1(n_228),
.B2(n_194),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_251),
.C(n_256),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_253),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_248),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

AO21x1_ASAP7_75t_L g250 ( 
.A1(n_237),
.A2(n_207),
.B(n_226),
.Y(n_250)
);

AOI21x1_ASAP7_75t_SL g258 ( 
.A1(n_250),
.A2(n_240),
.B(n_10),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_213),
.C(n_214),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_232),
.C(n_239),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_219),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_9),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_244),
.A2(n_224),
.B1(n_213),
.B2(n_229),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_257),
.B(n_260),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_258),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_9),
.C(n_10),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_263),
.B(n_265),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_255),
.A2(n_10),
.B(n_11),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_12),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_12),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_250),
.Y(n_269)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_269),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_270),
.B(n_274),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_266),
.B(n_251),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_273),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_245),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_258),
.B(n_252),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_261),
.Y(n_276)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_276),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_267),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_278),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_268),
.B(n_260),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_279),
.A2(n_257),
.B(n_13),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_282),
.B(n_277),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_284),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_283),
.B(n_280),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_285),
.C(n_275),
.Y(n_287)
);

OAI21x1_ASAP7_75t_SL g288 ( 
.A1(n_287),
.A2(n_281),
.B(n_13),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_12),
.C(n_13),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_14),
.Y(n_290)
);


endmodule