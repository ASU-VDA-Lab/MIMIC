module real_jpeg_10983_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_15;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_4),
.A2(n_27),
.B1(n_41),
.B2(n_42),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_4),
.A2(n_27),
.B1(n_68),
.B2(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_4),
.B(n_64),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_4),
.A2(n_64),
.B(n_92),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g148 ( 
.A1(n_4),
.A2(n_5),
.B(n_25),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_4),
.B(n_97),
.Y(n_171)
);

O2A1O1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_4),
.A2(n_9),
.B(n_68),
.C(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_4),
.B(n_105),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

O2A1O1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_5),
.A2(n_38),
.B(n_41),
.C(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_5),
.B(n_41),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_6),
.A2(n_33),
.B1(n_41),
.B2(n_42),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_6),
.A2(n_11),
.B1(n_33),
.B2(n_64),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_6),
.A2(n_33),
.B1(n_68),
.B2(n_69),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_8),
.A2(n_41),
.B1(n_42),
.B2(n_45),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_45),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_9),
.A2(n_68),
.B(n_78),
.C(n_79),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_9),
.B(n_68),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_9),
.A2(n_41),
.B1(n_42),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_9),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_10),
.A2(n_11),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_10),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_10),
.A2(n_65),
.B1(n_68),
.B2(n_69),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_65),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_10),
.A2(n_41),
.B1(n_42),
.B2(n_65),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_11),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_132),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_131),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_111),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_16),
.B(n_111),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_83),
.B2(n_110),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_50),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_29),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_21),
.B(n_157),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_28),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_22),
.B(n_158),
.Y(n_161)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_23),
.A2(n_34),
.B(n_35),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_24),
.B(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_35),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_27),
.A2(n_39),
.B(n_42),
.C(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_27),
.B(n_37),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_27),
.B(n_35),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g184 ( 
.A1(n_27),
.A2(n_41),
.B(n_80),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_28),
.B(n_32),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_28),
.B(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_29),
.A2(n_35),
.B(n_53),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_30),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

INVxp33_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_53),
.B(n_54),
.Y(n_52)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_34),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_40),
.B(n_46),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_37),
.A2(n_122),
.B(n_123),
.Y(n_121)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_47),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_38),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_38),
.B(n_58),
.Y(n_210)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_46),
.B(n_151),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_48),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_48),
.B(n_152),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_59),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_52),
.B(n_55),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_54),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_54),
.B(n_161),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_56),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_57),
.B(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_58),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_75),
.B2(n_76),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_71),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_62),
.B(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_63),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_64),
.A2(n_66),
.B(n_67),
.C(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_67),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_66),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_66)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_70),
.Y(n_90)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_90),
.B1(n_91),
.B2(n_93),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_72),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_73),
.B(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_74),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_79),
.B(n_81),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_77),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_79),
.B(n_130),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_82),
.B(n_128),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_83),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_94),
.C(n_102),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_84),
.A2(n_85),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_94),
.A2(n_95),
.B1(n_102),
.B2(n_103),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_101),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_99),
.B(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.C(n_116),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_112),
.B(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_115),
.B(n_116),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.C(n_124),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_117),
.B(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_120),
.A2(n_121),
.B1(n_124),
.B2(n_125),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_126),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_232),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_228),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_215),
.B(n_227),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_195),
.B(n_214),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_177),
.B(n_194),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_166),
.B(n_176),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_153),
.B(n_165),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_145),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_145),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_149),
.B2(n_150),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_147),
.B(n_149),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_159),
.B(n_164),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_156),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_168),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_175),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_173),
.C(n_175),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_179),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_186),
.B1(n_187),
.B2(n_193),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_180),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_183),
.B2(n_185),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_183),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_183),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_192),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_188),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_192),
.C(n_193),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_196),
.B(n_197),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_207),
.B2(n_208),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_209),
.C(n_213),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_204),
.C(n_205),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_209),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_211),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_216),
.B(n_217),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_226),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_222),
.C(n_225),
.Y(n_229)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_221),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_224),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_230),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);


endmodule