module fake_jpeg_23800_n_112 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_112);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_112;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_10),
.B(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_27),
.A2(n_22),
.B1(n_23),
.B2(n_14),
.Y(n_42)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_29),
.Y(n_36)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_23),
.B1(n_22),
.B2(n_13),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_12),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_21),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_14),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_30),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_19),
.B1(n_24),
.B2(n_25),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_27),
.A2(n_19),
.B1(n_15),
.B2(n_13),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_45),
.A2(n_30),
.B1(n_33),
.B2(n_9),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_47),
.A2(n_40),
.B1(n_35),
.B2(n_44),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_SL g48 ( 
.A(n_43),
.B(n_20),
.C(n_25),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_54),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_26),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_3),
.Y(n_51)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_4),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_58),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_35),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_62),
.B(n_65),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_50),
.B(n_58),
.C(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_53),
.B(n_55),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_68),
.Y(n_74)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_73),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_50),
.B(n_36),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_82),
.B(n_71),
.Y(n_90)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_80),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_46),
.B1(n_44),
.B2(n_35),
.Y(n_79)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_66),
.B(n_53),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_70),
.A2(n_39),
.B(n_55),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_70),
.C(n_72),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_88),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_63),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_86),
.B(n_87),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_63),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_70),
.C(n_72),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_90),
.B(n_88),
.Y(n_96)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_92),
.A2(n_95),
.B1(n_96),
.B2(n_94),
.Y(n_100)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

NOR2x1p5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_91),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_98),
.Y(n_102)
);

NOR3xp33_ASAP7_75t_SL g98 ( 
.A(n_94),
.B(n_89),
.C(n_64),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_64),
.C(n_62),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_95),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_75),
.C(n_61),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_103),
.A2(n_81),
.B(n_73),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_101),
.C(n_81),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_102),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_7),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_107),
.C(n_33),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_109),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_110),
.A2(n_39),
.B(n_8),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_10),
.Y(n_112)
);


endmodule