module fake_jpeg_25357_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_1),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

INVx11_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_16),
.B(n_20),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_9),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_18),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_8),
.Y(n_19)
);

AND2x2_ASAP7_75t_SL g22 ( 
.A(n_19),
.B(n_18),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_18),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_16),
.A2(n_14),
.B1(n_15),
.B2(n_13),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_24),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_11),
.B1(n_14),
.B2(n_13),
.Y(n_24)
);

NOR2x1_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_19),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_30),
.Y(n_33)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_19),
.Y(n_30)
);

AND2x6_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_35),
.Y(n_39)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_10),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_37),
.B(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_42),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_31),
.B1(n_29),
.B2(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_32),
.C(n_8),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_12),
.Y(n_47)
);

AOI21xp33_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_32),
.B(n_8),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_47),
.C(n_43),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_49),
.A2(n_50),
.B1(n_46),
.B2(n_2),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_48),
.A2(n_41),
.B1(n_44),
.B2(n_10),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_52),
.A2(n_3),
.B(n_5),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_55),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_51),
.C(n_5),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_58),
.A2(n_1),
.B1(n_6),
.B2(n_52),
.Y(n_59)
);


endmodule