module fake_jpeg_24031_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_48;
wire n_35;
wire n_71;
wire n_52;
wire n_68;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx1_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx5_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_7),
.B(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_20),
.Y(n_36)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_29),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_26)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_17),
.B1(n_11),
.B2(n_14),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_12),
.A2(n_0),
.B1(n_5),
.B2(n_8),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_9),
.C(n_18),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_8),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_25),
.B1(n_32),
.B2(n_37),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_29),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_37),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_16),
.B1(n_18),
.B2(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_9),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_21),
.B(n_11),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_48),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_31),
.A2(n_23),
.B1(n_22),
.B2(n_27),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_33),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_25),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_33),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_30),
.A2(n_34),
.B(n_38),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_34),
.C(n_39),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_50),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_34),
.B(n_39),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_54),
.C(n_56),
.Y(n_58)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

BUFx24_ASAP7_75t_SL g59 ( 
.A(n_55),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_61),
.Y(n_65)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_57),
.A2(n_45),
.B1(n_44),
.B2(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

AOI322xp5_ASAP7_75t_SL g63 ( 
.A1(n_59),
.A2(n_35),
.A3(n_43),
.B1(n_49),
.B2(n_51),
.C1(n_57),
.C2(n_60),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_58),
.Y(n_66)
);

OAI21x1_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_65),
.B(n_64),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_64),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_68),
.Y(n_72)
);


endmodule