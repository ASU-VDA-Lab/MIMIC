module fake_jpeg_3913_n_44 (n_3, n_2, n_1, n_0, n_4, n_5, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_4),
.Y(n_6)
);

BUFx16f_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

INVx8_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_2),
.B(n_5),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_18),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_7),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_20),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_7),
.A2(n_0),
.B(n_1),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_8),
.C(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_19),
.B(n_9),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_6),
.B(n_5),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_6),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_26),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_10),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_28),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_17),
.B1(n_20),
.B2(n_16),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_SL g35 ( 
.A(n_30),
.B(n_32),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_14),
.C(n_18),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_22),
.B(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_34),
.B(n_19),
.Y(n_39)
);

OAI21xp33_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_22),
.B(n_23),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_15),
.B(n_13),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_37),
.A2(n_33),
.B(n_32),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_40),
.C(n_35),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_19),
.Y(n_42)
);

AOI322xp5_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_42),
.A3(n_9),
.B1(n_11),
.B2(n_13),
.C1(n_36),
.C2(n_30),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_43),
.A2(n_9),
.B(n_13),
.Y(n_44)
);


endmodule