module fake_netlist_6_2638_n_1117 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1117);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1117;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_1008;
wire n_465;
wire n_367;
wire n_680;
wire n_741;
wire n_760;
wire n_1027;
wire n_875;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_462;
wire n_1033;
wire n_607;
wire n_671;
wire n_726;
wire n_1052;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_988;
wire n_969;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1099;
wire n_1026;
wire n_443;
wire n_1101;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_222;
wire n_718;
wire n_248;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_901;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_1078;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_1116;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_772;
wire n_656;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_886;
wire n_448;
wire n_844;
wire n_1017;
wire n_1004;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_1084;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_870;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_982;
wire n_964;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_959;
wire n_879;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_518;
wire n_299;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_1001;
wire n_827;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_143),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_61),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_112),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_125),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_194),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_117),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_128),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_25),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_126),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_83),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_101),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_54),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_65),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_169),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_132),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_150),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_91),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_16),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_26),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_168),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_146),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_78),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_47),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_139),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_192),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_1),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_185),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_207),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_92),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_129),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_12),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_32),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_50),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_134),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_190),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_100),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_20),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_17),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_59),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_4),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_195),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_189),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_200),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_160),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_204),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_151),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_177),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_212),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_1),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_153),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_66),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_88),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_34),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_99),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_84),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_199),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_103),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_165),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_90),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_69),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_73),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_55),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_107),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_119),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_26),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_196),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_148),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_9),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_170),
.Y(n_281)
);

INVxp33_ASAP7_75t_R g282 ( 
.A(n_41),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_16),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_238),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_238),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_277),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_244),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

INVx4_ASAP7_75t_R g289 ( 
.A(n_222),
.Y(n_289)
);

INVxp33_ASAP7_75t_SL g290 ( 
.A(n_230),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_244),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_231),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_261),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_261),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_277),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_277),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_277),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_223),
.Y(n_298)
);

BUFx2_ASAP7_75t_SL g299 ( 
.A(n_219),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_283),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_214),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_218),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_249),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_213),
.Y(n_304)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_224),
.Y(n_305)
);

INVxp33_ASAP7_75t_SL g306 ( 
.A(n_243),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_216),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_226),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_250),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_233),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_249),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_266),
.Y(n_312)
);

BUFx5_ASAP7_75t_L g313 ( 
.A(n_271),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_219),
.Y(n_314)
);

INVxp33_ASAP7_75t_L g315 ( 
.A(n_220),
.Y(n_315)
);

INVxp33_ASAP7_75t_SL g316 ( 
.A(n_252),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_272),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_221),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_215),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_215),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_245),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_245),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_247),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_225),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_227),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_228),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_280),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_217),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_247),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_217),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_253),
.Y(n_331)
);

INVxp33_ASAP7_75t_L g332 ( 
.A(n_220),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_274),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_284),
.B(n_263),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_304),
.B(n_253),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_290),
.A2(n_274),
.B1(n_279),
.B2(n_251),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_286),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_286),
.Y(n_338)
);

INVx5_ASAP7_75t_L g339 ( 
.A(n_313),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_285),
.B(n_257),
.Y(n_340)
);

AND2x2_ASAP7_75t_SL g341 ( 
.A(n_298),
.B(n_246),
.Y(n_341)
);

INVx5_ASAP7_75t_L g342 ( 
.A(n_313),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_292),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_295),
.Y(n_344)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_313),
.Y(n_345)
);

BUFx12f_ASAP7_75t_L g346 ( 
.A(n_307),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_296),
.Y(n_347)
);

AND2x2_ASAP7_75t_SL g348 ( 
.A(n_301),
.B(n_246),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_297),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_319),
.Y(n_350)
);

OA21x2_ASAP7_75t_L g351 ( 
.A1(n_320),
.A2(n_251),
.B(n_232),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_323),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_313),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_290),
.A2(n_279),
.B1(n_234),
.B2(n_235),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_292),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_329),
.Y(n_356)
);

AND2x2_ASAP7_75t_SL g357 ( 
.A(n_302),
.B(n_246),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_299),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_313),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_314),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_287),
.B(n_257),
.Y(n_361)
);

AND2x4_ASAP7_75t_L g362 ( 
.A(n_321),
.B(n_246),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_331),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_308),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_313),
.Y(n_365)
);

AND2x4_ASAP7_75t_L g366 ( 
.A(n_322),
.B(n_229),
.Y(n_366)
);

NAND2x1p5_ASAP7_75t_L g367 ( 
.A(n_312),
.B(n_257),
.Y(n_367)
);

AND2x2_ASAP7_75t_SL g368 ( 
.A(n_317),
.B(n_282),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_300),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_313),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_291),
.Y(n_371)
);

AOI22x1_ASAP7_75t_SL g372 ( 
.A1(n_314),
.A2(n_281),
.B1(n_278),
.B2(n_276),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_293),
.Y(n_373)
);

OAI22x1_ASAP7_75t_SL g374 ( 
.A1(n_303),
.A2(n_275),
.B1(n_273),
.B2(n_270),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_306),
.A2(n_255),
.B1(n_268),
.B2(n_267),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_318),
.Y(n_376)
);

NOR2x1_ASAP7_75t_L g377 ( 
.A(n_294),
.B(n_236),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_305),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_310),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_288),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_328),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_324),
.B(n_269),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_315),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_332),
.B(n_237),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_328),
.B(n_330),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_306),
.A2(n_254),
.B1(n_262),
.B2(n_260),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_325),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_326),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_341),
.B(n_330),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_344),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_341),
.A2(n_316),
.B1(n_309),
.B2(n_327),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_341),
.B(n_316),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_373),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_383),
.B(n_309),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_360),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_350),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_383),
.B(n_327),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_373),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_344),
.Y(n_399)
);

AND2x6_ASAP7_75t_L g400 ( 
.A(n_377),
.B(n_289),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_373),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_344),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_350),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_384),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_350),
.Y(n_405)
);

NAND2xp33_ASAP7_75t_L g406 ( 
.A(n_335),
.B(n_239),
.Y(n_406)
);

NAND2xp33_ASAP7_75t_SL g407 ( 
.A(n_334),
.B(n_333),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_347),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_347),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_347),
.Y(n_410)
);

NAND2xp33_ASAP7_75t_SL g411 ( 
.A(n_334),
.B(n_333),
.Y(n_411)
);

AND2x6_ASAP7_75t_L g412 ( 
.A(n_377),
.B(n_45),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_349),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_371),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_378),
.B(n_240),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_371),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_350),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_388),
.B(n_241),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_355),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_349),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_336),
.B(n_303),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_336),
.A2(n_311),
.B1(n_264),
.B2(n_259),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_369),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_384),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_350),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_349),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_337),
.Y(n_427)
);

BUFx6f_ASAP7_75t_SL g428 ( 
.A(n_368),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_364),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_337),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_369),
.Y(n_431)
);

AND3x1_ASAP7_75t_L g432 ( 
.A(n_385),
.B(n_311),
.C(n_0),
.Y(n_432)
);

OAI21x1_ASAP7_75t_L g433 ( 
.A1(n_351),
.A2(n_248),
.B(n_242),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_338),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_380),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_364),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_367),
.B(n_256),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_350),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_364),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_352),
.Y(n_440)
);

INVx8_ASAP7_75t_L g441 ( 
.A(n_366),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_338),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_352),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_378),
.B(n_258),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_385),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_338),
.Y(n_446)
);

OA21x2_ASAP7_75t_L g447 ( 
.A1(n_362),
.A2(n_48),
.B(n_46),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_352),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_352),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_388),
.B(n_2),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_352),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_352),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_338),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_356),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_355),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_356),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_348),
.B(n_49),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_356),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_378),
.B(n_51),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_356),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_380),
.B(n_52),
.Y(n_461)
);

BUFx6f_ASAP7_75t_SL g462 ( 
.A(n_368),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_404),
.B(n_381),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_395),
.B(n_381),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_391),
.B(n_381),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_429),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_459),
.B(n_348),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_441),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_418),
.B(n_381),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_459),
.B(n_348),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_429),
.B(n_357),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_441),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_415),
.B(n_387),
.Y(n_473)
);

AO221x1_ASAP7_75t_L g474 ( 
.A1(n_422),
.A2(n_387),
.B1(n_379),
.B2(n_380),
.C(n_374),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_389),
.B(n_387),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_415),
.B(n_357),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_415),
.B(n_357),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_444),
.B(n_366),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_434),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_444),
.B(n_366),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_444),
.B(n_366),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_392),
.B(n_376),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_461),
.B(n_424),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_461),
.B(n_379),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_394),
.B(n_382),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_397),
.B(n_358),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_434),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_435),
.B(n_375),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_436),
.B(n_362),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_439),
.B(n_354),
.Y(n_490)
);

NAND3xp33_ASAP7_75t_L g491 ( 
.A(n_450),
.B(n_386),
.C(n_375),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_423),
.B(n_362),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_437),
.B(n_386),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_431),
.B(n_367),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_414),
.B(n_343),
.Y(n_495)
);

NAND2x1_ASAP7_75t_L g496 ( 
.A(n_396),
.B(n_362),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_416),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_419),
.B(n_367),
.Y(n_498)
);

A2O1A1Ixp33_ASAP7_75t_L g499 ( 
.A1(n_457),
.A2(n_361),
.B(n_340),
.C(n_368),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_427),
.Y(n_500)
);

AO221x1_ASAP7_75t_L g501 ( 
.A1(n_432),
.A2(n_374),
.B1(n_372),
.B2(n_351),
.C(n_356),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_441),
.B(n_400),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_427),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_430),
.Y(n_504)
);

INVxp33_ASAP7_75t_L g505 ( 
.A(n_421),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_407),
.B(n_346),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_406),
.B(n_346),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_428),
.B(n_346),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_430),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_406),
.B(n_351),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_400),
.B(n_351),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_442),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_441),
.B(n_353),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_400),
.B(n_353),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_393),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_403),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_393),
.Y(n_517)
);

NAND2xp33_ASAP7_75t_SL g518 ( 
.A(n_428),
.B(n_340),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_398),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_407),
.B(n_361),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_411),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_411),
.B(n_356),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_400),
.B(n_353),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_445),
.B(n_363),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_455),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_400),
.B(n_359),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_421),
.B(n_372),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_398),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_401),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_400),
.B(n_363),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_401),
.B(n_359),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_440),
.B(n_363),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_396),
.B(n_359),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_442),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_440),
.B(n_363),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_446),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_402),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_396),
.B(n_370),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_417),
.B(n_425),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_SL g540 ( 
.A(n_428),
.B(n_363),
.Y(n_540)
);

NOR3xp33_ASAP7_75t_L g541 ( 
.A(n_402),
.B(n_345),
.C(n_365),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_417),
.B(n_370),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_417),
.B(n_370),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_446),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_425),
.B(n_365),
.Y(n_545)
);

NOR2xp67_ASAP7_75t_L g546 ( 
.A(n_456),
.B(n_53),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_443),
.B(n_363),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_484),
.B(n_425),
.Y(n_548)
);

CKINVDCx16_ASAP7_75t_R g549 ( 
.A(n_508),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_500),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_525),
.Y(n_551)
);

BUFx8_ASAP7_75t_L g552 ( 
.A(n_464),
.Y(n_552)
);

NAND2x1p5_ASAP7_75t_L g553 ( 
.A(n_468),
.B(n_447),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_483),
.B(n_438),
.Y(n_554)
);

AO22x2_ASAP7_75t_L g555 ( 
.A1(n_491),
.A2(n_462),
.B1(n_455),
.B2(n_5),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_463),
.B(n_438),
.Y(n_556)
);

AO22x2_ASAP7_75t_L g557 ( 
.A1(n_493),
.A2(n_462),
.B1(n_4),
.B2(n_5),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_475),
.A2(n_462),
.B1(n_412),
.B2(n_448),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_463),
.B(n_467),
.Y(n_559)
);

INVxp67_ASAP7_75t_SL g560 ( 
.A(n_516),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_518),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_503),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_504),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_509),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_466),
.Y(n_565)
);

BUFx8_ASAP7_75t_L g566 ( 
.A(n_497),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_515),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_473),
.B(n_456),
.Y(n_568)
);

AO22x2_ASAP7_75t_L g569 ( 
.A1(n_465),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_517),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_519),
.Y(n_571)
);

OR2x6_ASAP7_75t_SL g572 ( 
.A(n_527),
.B(n_412),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_470),
.A2(n_447),
.B1(n_443),
.B2(n_460),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_528),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_482),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_529),
.Y(n_576)
);

NAND2x1p5_ASAP7_75t_L g577 ( 
.A(n_468),
.B(n_472),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_485),
.B(n_438),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_537),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_516),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_476),
.A2(n_447),
.B1(n_448),
.B2(n_460),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_479),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_487),
.Y(n_583)
);

AO22x2_ASAP7_75t_L g584 ( 
.A1(n_520),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_584)
);

AO22x2_ASAP7_75t_L g585 ( 
.A1(n_488),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_585)
);

BUFx8_ASAP7_75t_L g586 ( 
.A(n_474),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_469),
.B(n_449),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_478),
.B(n_449),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_477),
.A2(n_412),
.B1(n_420),
.B2(n_451),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_494),
.B(n_458),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_512),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_480),
.B(n_451),
.Y(n_592)
);

NAND2x1p5_ASAP7_75t_L g593 ( 
.A(n_468),
.B(n_447),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_481),
.B(n_420),
.Y(n_594)
);

BUFx8_ASAP7_75t_L g595 ( 
.A(n_468),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_534),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_536),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_544),
.Y(n_598)
);

AO22x2_ASAP7_75t_L g599 ( 
.A1(n_521),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_599)
);

AO22x2_ASAP7_75t_L g600 ( 
.A1(n_506),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_489),
.Y(n_601)
);

AO22x2_ASAP7_75t_L g602 ( 
.A1(n_498),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_492),
.B(n_458),
.Y(n_603)
);

AO22x2_ASAP7_75t_L g604 ( 
.A1(n_501),
.A2(n_524),
.B1(n_522),
.B2(n_499),
.Y(n_604)
);

AO22x2_ASAP7_75t_L g605 ( 
.A1(n_505),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_539),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_490),
.B(n_390),
.Y(n_607)
);

NOR2xp67_ASAP7_75t_L g608 ( 
.A(n_486),
.B(n_507),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_495),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_495),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_533),
.Y(n_611)
);

AND2x6_ASAP7_75t_L g612 ( 
.A(n_511),
.B(n_452),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_471),
.B(n_390),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_496),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_538),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_542),
.Y(n_616)
);

INVx4_ASAP7_75t_L g617 ( 
.A(n_551),
.Y(n_617)
);

O2A1O1Ixp33_ASAP7_75t_L g618 ( 
.A1(n_609),
.A2(n_507),
.B(n_510),
.C(n_511),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_594),
.A2(n_513),
.B(n_472),
.Y(n_619)
);

AND2x6_ASAP7_75t_L g620 ( 
.A(n_558),
.B(n_502),
.Y(n_620)
);

O2A1O1Ixp5_ASAP7_75t_L g621 ( 
.A1(n_573),
.A2(n_510),
.B(n_530),
.C(n_526),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_565),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_610),
.B(n_530),
.Y(n_623)
);

NAND2x1p5_ASAP7_75t_L g624 ( 
.A(n_580),
.B(n_472),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_L g625 ( 
.A1(n_559),
.A2(n_541),
.B(n_523),
.Y(n_625)
);

INVxp67_ASAP7_75t_L g626 ( 
.A(n_552),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_588),
.A2(n_472),
.B(n_516),
.Y(n_627)
);

AOI21x1_ASAP7_75t_L g628 ( 
.A1(n_556),
.A2(n_514),
.B(n_531),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_592),
.A2(n_516),
.B(n_543),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_548),
.A2(n_545),
.B(n_540),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_575),
.B(n_532),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_567),
.Y(n_632)
);

O2A1O1Ixp33_ASAP7_75t_L g633 ( 
.A1(n_607),
.A2(n_541),
.B(n_532),
.C(n_547),
.Y(n_633)
);

NAND2x1p5_ASAP7_75t_L g634 ( 
.A(n_570),
.B(n_546),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_578),
.A2(n_345),
.B(n_535),
.Y(n_635)
);

O2A1O1Ixp33_ASAP7_75t_L g636 ( 
.A1(n_601),
.A2(n_547),
.B(n_535),
.C(n_413),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_571),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_577),
.Y(n_638)
);

INVxp33_ASAP7_75t_SL g639 ( 
.A(n_608),
.Y(n_639)
);

A2O1A1Ixp33_ASAP7_75t_L g640 ( 
.A1(n_589),
.A2(n_433),
.B(n_399),
.C(n_409),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_604),
.A2(n_412),
.B1(n_433),
.B2(n_403),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_574),
.B(n_412),
.Y(n_642)
);

AO21x1_ASAP7_75t_L g643 ( 
.A1(n_581),
.A2(n_408),
.B(n_399),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_L g644 ( 
.A1(n_613),
.A2(n_409),
.B(n_408),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_L g645 ( 
.A1(n_615),
.A2(n_413),
.B(n_410),
.Y(n_645)
);

AOI21x1_ASAP7_75t_L g646 ( 
.A1(n_603),
.A2(n_426),
.B(n_410),
.Y(n_646)
);

OR2x6_ASAP7_75t_SL g647 ( 
.A(n_550),
.B(n_412),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_553),
.A2(n_345),
.B(n_403),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_549),
.B(n_18),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_576),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_604),
.A2(n_426),
.B1(n_453),
.B2(n_454),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_579),
.B(n_453),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_562),
.Y(n_653)
);

NOR2x1p5_ASAP7_75t_L g654 ( 
.A(n_551),
.B(n_403),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_593),
.A2(n_345),
.B(n_403),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g656 ( 
.A(n_552),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_561),
.B(n_606),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_616),
.B(n_611),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_595),
.B(n_405),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_568),
.B(n_405),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_554),
.A2(n_454),
.B(n_405),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_563),
.B(n_405),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_564),
.B(n_405),
.Y(n_663)
);

NOR3xp33_ASAP7_75t_L g664 ( 
.A(n_614),
.B(n_365),
.C(n_19),
.Y(n_664)
);

NAND2xp33_ASAP7_75t_L g665 ( 
.A(n_612),
.B(n_583),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_555),
.B(n_19),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_560),
.A2(n_454),
.B(n_342),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_595),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_582),
.Y(n_669)
);

A2O1A1Ixp33_ASAP7_75t_L g670 ( 
.A1(n_590),
.A2(n_454),
.B(n_342),
.C(n_339),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_587),
.A2(n_454),
.B(n_342),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_568),
.B(n_20),
.Y(n_672)
);

AOI33xp33_ASAP7_75t_L g673 ( 
.A1(n_591),
.A2(n_21),
.A3(n_22),
.B1(n_23),
.B2(n_24),
.B3(n_25),
.Y(n_673)
);

BUFx8_ASAP7_75t_L g674 ( 
.A(n_566),
.Y(n_674)
);

CKINVDCx8_ASAP7_75t_R g675 ( 
.A(n_590),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_596),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_612),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_597),
.A2(n_342),
.B(n_339),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_623),
.B(n_585),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_631),
.B(n_586),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_674),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_658),
.B(n_585),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_674),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_639),
.B(n_586),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_666),
.B(n_557),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_622),
.B(n_632),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_657),
.B(n_637),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_664),
.A2(n_555),
.B1(n_557),
.B2(n_569),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_677),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_650),
.B(n_660),
.Y(n_690)
);

OAI21xp5_ASAP7_75t_L g691 ( 
.A1(n_618),
.A2(n_598),
.B(n_612),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_660),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_653),
.B(n_569),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_654),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_676),
.B(n_572),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_SL g696 ( 
.A1(n_649),
.A2(n_566),
.B1(n_605),
.B2(n_600),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_669),
.B(n_584),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_646),
.Y(n_698)
);

INVxp67_ASAP7_75t_L g699 ( 
.A(n_668),
.Y(n_699)
);

NAND2x1_ASAP7_75t_L g700 ( 
.A(n_677),
.B(n_638),
.Y(n_700)
);

OR2x2_ASAP7_75t_L g701 ( 
.A(n_672),
.B(n_21),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_675),
.B(n_602),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_625),
.B(n_602),
.Y(n_703)
);

NAND2x1p5_ASAP7_75t_L g704 ( 
.A(n_638),
.B(n_584),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_652),
.Y(n_705)
);

AND3x1_ASAP7_75t_SL g706 ( 
.A(n_673),
.B(n_605),
.C(n_599),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_617),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_617),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_665),
.A2(n_600),
.B1(n_599),
.B2(n_342),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_625),
.B(n_342),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_662),
.Y(n_711)
);

CKINVDCx16_ASAP7_75t_R g712 ( 
.A(n_656),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_626),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_620),
.A2(n_339),
.B1(n_23),
.B2(n_24),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_628),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_663),
.Y(n_716)
);

NAND3xp33_ASAP7_75t_L g717 ( 
.A(n_641),
.B(n_339),
.C(n_22),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_651),
.B(n_56),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_624),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_645),
.B(n_57),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_659),
.B(n_58),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_SL g722 ( 
.A1(n_620),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_627),
.B(n_60),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_624),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_645),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_642),
.Y(n_726)
);

NAND2xp33_ASAP7_75t_L g727 ( 
.A(n_620),
.B(n_339),
.Y(n_727)
);

NAND2x1p5_ASAP7_75t_L g728 ( 
.A(n_619),
.B(n_339),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_647),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_729)
);

CKINVDCx16_ASAP7_75t_R g730 ( 
.A(n_620),
.Y(n_730)
);

AND2x6_ASAP7_75t_L g731 ( 
.A(n_670),
.B(n_62),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_621),
.Y(n_732)
);

AOI22x1_ASAP7_75t_L g733 ( 
.A1(n_634),
.A2(n_135),
.B1(n_210),
.B2(n_209),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_634),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_633),
.B(n_30),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_629),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_643),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_682),
.B(n_636),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_690),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_707),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_685),
.B(n_644),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_686),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_707),
.Y(n_743)
);

OR2x6_ASAP7_75t_L g744 ( 
.A(n_721),
.B(n_630),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_692),
.B(n_661),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_686),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_727),
.A2(n_635),
.B(n_640),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_708),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_708),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_685),
.B(n_644),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_692),
.B(n_667),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_713),
.Y(n_752)
);

BUFx10_ASAP7_75t_L g753 ( 
.A(n_681),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_694),
.B(n_648),
.Y(n_754)
);

OA21x2_ASAP7_75t_L g755 ( 
.A1(n_732),
.A2(n_671),
.B(n_655),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_727),
.A2(n_736),
.B(n_710),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_687),
.B(n_680),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_682),
.B(n_678),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_694),
.B(n_690),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_697),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_734),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_705),
.B(n_31),
.Y(n_762)
);

NAND2x1p5_ASAP7_75t_L g763 ( 
.A(n_689),
.B(n_723),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_695),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_705),
.B(n_679),
.Y(n_765)
);

AO21x1_ASAP7_75t_L g766 ( 
.A1(n_735),
.A2(n_33),
.B(n_34),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_689),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_689),
.Y(n_768)
);

AND2x6_ASAP7_75t_L g769 ( 
.A(n_718),
.B(n_63),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_697),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_736),
.A2(n_691),
.B(n_725),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_679),
.B(n_33),
.Y(n_772)
);

CKINVDCx16_ASAP7_75t_R g773 ( 
.A(n_712),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_693),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_736),
.A2(n_137),
.B(n_208),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_693),
.B(n_701),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_684),
.B(n_64),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_716),
.Y(n_778)
);

BUFx2_ASAP7_75t_L g779 ( 
.A(n_699),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_732),
.A2(n_138),
.B(n_206),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_713),
.Y(n_781)
);

HB1xp67_ASAP7_75t_L g782 ( 
.A(n_702),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_711),
.B(n_35),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_709),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_784)
);

A2O1A1Ixp33_ASAP7_75t_SL g785 ( 
.A1(n_737),
.A2(n_36),
.B(n_37),
.C(n_38),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_721),
.B(n_38),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_700),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_716),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_703),
.B(n_39),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_701),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_726),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_721),
.B(n_67),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_688),
.B(n_39),
.Y(n_793)
);

INVx4_ASAP7_75t_L g794 ( 
.A(n_681),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_719),
.B(n_68),
.Y(n_795)
);

AO21x2_ASAP7_75t_L g796 ( 
.A1(n_715),
.A2(n_142),
.B(n_205),
.Y(n_796)
);

A2O1A1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_717),
.A2(n_40),
.B(n_41),
.C(n_42),
.Y(n_797)
);

AOI21xp33_ASAP7_75t_SL g798 ( 
.A1(n_696),
.A2(n_683),
.B(n_730),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_726),
.B(n_40),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_724),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_722),
.B(n_42),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_723),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_715),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_718),
.B(n_43),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_704),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_803),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_791),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_778),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_779),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_774),
.B(n_704),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_774),
.B(n_720),
.Y(n_811)
);

O2A1O1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_785),
.A2(n_729),
.B(n_720),
.C(n_723),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_741),
.B(n_714),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_750),
.B(n_698),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_757),
.A2(n_706),
.B1(n_683),
.B2(n_731),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_739),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_SL g817 ( 
.A1(n_792),
.A2(n_731),
.B(n_728),
.Y(n_817)
);

A2O1A1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_797),
.A2(n_698),
.B(n_733),
.C(n_731),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_747),
.A2(n_728),
.B(n_731),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_790),
.B(n_731),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_776),
.B(n_731),
.Y(n_821)
);

O2A1O1Ixp5_ASAP7_75t_L g822 ( 
.A1(n_784),
.A2(n_43),
.B(n_44),
.C(n_70),
.Y(n_822)
);

NOR2xp67_ASAP7_75t_L g823 ( 
.A(n_743),
.B(n_71),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_747),
.A2(n_147),
.B(n_72),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_760),
.B(n_44),
.Y(n_825)
);

BUFx2_ASAP7_75t_L g826 ( 
.A(n_744),
.Y(n_826)
);

NAND2x1p5_ASAP7_75t_L g827 ( 
.A(n_802),
.B(n_74),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_765),
.B(n_75),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_770),
.B(n_76),
.Y(n_829)
);

INVx1_ASAP7_75t_SL g830 ( 
.A(n_740),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_765),
.B(n_77),
.Y(n_831)
);

O2A1O1Ixp5_ASAP7_75t_L g832 ( 
.A1(n_784),
.A2(n_79),
.B(n_80),
.C(n_81),
.Y(n_832)
);

HB1xp67_ASAP7_75t_L g833 ( 
.A(n_742),
.Y(n_833)
);

OR2x2_ASAP7_75t_L g834 ( 
.A(n_738),
.B(n_211),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_804),
.A2(n_82),
.B(n_85),
.C(n_86),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_746),
.B(n_738),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_788),
.Y(n_837)
);

OR2x2_ASAP7_75t_L g838 ( 
.A(n_789),
.B(n_203),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_800),
.Y(n_839)
);

O2A1O1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_786),
.A2(n_87),
.B(n_89),
.C(n_93),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_782),
.B(n_202),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_772),
.B(n_94),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_762),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_804),
.B(n_95),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_748),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_767),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_756),
.A2(n_96),
.B(n_97),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_789),
.B(n_98),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_758),
.B(n_201),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_762),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_758),
.B(n_102),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_748),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_793),
.B(n_198),
.Y(n_853)
);

INVx3_ASAP7_75t_SL g854 ( 
.A(n_773),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_SL g855 ( 
.A(n_794),
.B(n_104),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_802),
.B(n_105),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_799),
.Y(n_857)
);

BUFx12f_ASAP7_75t_L g858 ( 
.A(n_753),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_799),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_764),
.B(n_106),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_802),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_764),
.B(n_197),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_764),
.B(n_108),
.Y(n_863)
);

CKINVDCx20_ASAP7_75t_R g864 ( 
.A(n_753),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_SL g865 ( 
.A1(n_777),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_763),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_865),
.A2(n_769),
.B1(n_801),
.B2(n_766),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_815),
.A2(n_798),
.B1(n_792),
.B2(n_805),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_SL g869 ( 
.A1(n_855),
.A2(n_769),
.B1(n_744),
.B2(n_780),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_808),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_866),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_813),
.A2(n_769),
.B1(n_744),
.B2(n_751),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_813),
.A2(n_769),
.B1(n_826),
.B2(n_820),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_826),
.A2(n_751),
.B1(n_754),
.B2(n_745),
.Y(n_874)
);

OAI22xp5_ASAP7_75t_SL g875 ( 
.A1(n_854),
.A2(n_794),
.B1(n_752),
.B2(n_781),
.Y(n_875)
);

OAI21xp33_ASAP7_75t_L g876 ( 
.A1(n_838),
.A2(n_783),
.B(n_780),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_849),
.A2(n_754),
.B1(n_759),
.B2(n_795),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_830),
.B(n_761),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_849),
.A2(n_759),
.B1(n_795),
.B2(n_775),
.Y(n_879)
);

OAI21xp5_ASAP7_75t_SL g880 ( 
.A1(n_812),
.A2(n_771),
.B(n_761),
.Y(n_880)
);

INVx6_ASAP7_75t_L g881 ( 
.A(n_861),
.Y(n_881)
);

OAI222xp33_ASAP7_75t_L g882 ( 
.A1(n_834),
.A2(n_749),
.B1(n_756),
.B2(n_767),
.C1(n_768),
.C2(n_796),
.Y(n_882)
);

BUFx3_ASAP7_75t_L g883 ( 
.A(n_852),
.Y(n_883)
);

BUFx12f_ASAP7_75t_L g884 ( 
.A(n_858),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_808),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_839),
.Y(n_886)
);

OAI22xp33_ASAP7_75t_L g887 ( 
.A1(n_823),
.A2(n_761),
.B1(n_748),
.B2(n_787),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_851),
.A2(n_796),
.B1(n_768),
.B2(n_787),
.Y(n_888)
);

AOI22xp33_ASAP7_75t_L g889 ( 
.A1(n_851),
.A2(n_787),
.B1(n_755),
.B2(n_115),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_821),
.A2(n_755),
.B1(n_114),
.B2(n_116),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_866),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_843),
.B(n_113),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_837),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_853),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_806),
.Y(n_895)
);

BUFx4f_ASAP7_75t_SL g896 ( 
.A(n_858),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_836),
.B(n_122),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_853),
.A2(n_123),
.B1(n_124),
.B2(n_127),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_806),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_809),
.A2(n_130),
.B1(n_131),
.B2(n_133),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_850),
.B(n_136),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_L g902 ( 
.A1(n_864),
.A2(n_140),
.B1(n_141),
.B2(n_144),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_L g903 ( 
.A1(n_854),
.A2(n_857),
.B1(n_859),
.B2(n_848),
.Y(n_903)
);

OAI21xp5_ASAP7_75t_SL g904 ( 
.A1(n_840),
.A2(n_835),
.B(n_824),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_860),
.B(n_838),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_807),
.Y(n_906)
);

CKINVDCx20_ASAP7_75t_R g907 ( 
.A(n_864),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_866),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_848),
.A2(n_145),
.B1(n_149),
.B2(n_152),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_818),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_886),
.B(n_836),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_908),
.B(n_871),
.Y(n_912)
);

OR2x2_ASAP7_75t_L g913 ( 
.A(n_886),
.B(n_816),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_903),
.B(n_814),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_871),
.B(n_852),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_908),
.B(n_811),
.Y(n_916)
);

AO21x2_ASAP7_75t_L g917 ( 
.A1(n_882),
.A2(n_819),
.B(n_847),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_893),
.B(n_811),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_904),
.A2(n_822),
.B(n_832),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_893),
.B(n_905),
.Y(n_920)
);

O2A1O1Ixp33_ASAP7_75t_SL g921 ( 
.A1(n_907),
.A2(n_887),
.B(n_868),
.C(n_902),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_871),
.B(n_845),
.Y(n_922)
);

INVx5_ASAP7_75t_L g923 ( 
.A(n_881),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_870),
.Y(n_924)
);

OAI211xp5_ASAP7_75t_L g925 ( 
.A1(n_876),
.A2(n_844),
.B(n_825),
.C(n_841),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_891),
.B(n_810),
.Y(n_926)
);

OR2x6_ASAP7_75t_L g927 ( 
.A(n_880),
.B(n_817),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_899),
.B(n_833),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_870),
.B(n_810),
.Y(n_929)
);

INVx2_ASAP7_75t_SL g930 ( 
.A(n_883),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_885),
.Y(n_931)
);

OR2x2_ASAP7_75t_L g932 ( 
.A(n_885),
.B(n_846),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_904),
.A2(n_831),
.B(n_828),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_876),
.A2(n_863),
.B(n_862),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_869),
.A2(n_863),
.B(n_862),
.Y(n_935)
);

OA21x2_ASAP7_75t_L g936 ( 
.A1(n_888),
.A2(n_841),
.B(n_825),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_895),
.B(n_861),
.Y(n_937)
);

NOR2xp67_ASAP7_75t_L g938 ( 
.A(n_891),
.B(n_861),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_916),
.B(n_891),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_916),
.B(n_895),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_920),
.B(n_911),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_924),
.Y(n_942)
);

OR2x6_ASAP7_75t_L g943 ( 
.A(n_927),
.B(n_817),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_911),
.B(n_906),
.Y(n_944)
);

AND2x4_ASAP7_75t_SL g945 ( 
.A(n_927),
.B(n_915),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_924),
.Y(n_946)
);

OR2x2_ASAP7_75t_L g947 ( 
.A(n_913),
.B(n_906),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_918),
.B(n_883),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_931),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_918),
.B(n_897),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_932),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_926),
.B(n_878),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_929),
.B(n_897),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_932),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_923),
.B(n_874),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_923),
.B(n_872),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_923),
.B(n_938),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_926),
.B(n_873),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_926),
.B(n_881),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_937),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_926),
.B(n_881),
.Y(n_961)
);

OAI21xp33_ASAP7_75t_L g962 ( 
.A1(n_958),
.A2(n_925),
.B(n_919),
.Y(n_962)
);

NOR3xp33_ASAP7_75t_L g963 ( 
.A(n_958),
.B(n_933),
.C(n_921),
.Y(n_963)
);

INVx4_ASAP7_75t_SL g964 ( 
.A(n_943),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_943),
.A2(n_927),
.B(n_917),
.Y(n_965)
);

INVx1_ASAP7_75t_SL g966 ( 
.A(n_952),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_945),
.B(n_957),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_942),
.Y(n_968)
);

INVx1_ASAP7_75t_SL g969 ( 
.A(n_952),
.Y(n_969)
);

O2A1O1Ixp5_ASAP7_75t_L g970 ( 
.A1(n_956),
.A2(n_934),
.B(n_935),
.C(n_914),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_959),
.B(n_923),
.Y(n_971)
);

OA21x2_ASAP7_75t_L g972 ( 
.A1(n_942),
.A2(n_938),
.B(n_912),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_957),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_949),
.Y(n_974)
);

CKINVDCx16_ASAP7_75t_R g975 ( 
.A(n_957),
.Y(n_975)
);

OR2x6_ASAP7_75t_L g976 ( 
.A(n_943),
.B(n_927),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_946),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_962),
.B(n_941),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_972),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_975),
.B(n_959),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_975),
.B(n_961),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_972),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_977),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_963),
.B(n_957),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_977),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_966),
.B(n_954),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_968),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_967),
.B(n_961),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_967),
.B(n_945),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_983),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_983),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_979),
.Y(n_992)
);

INVx4_ASAP7_75t_L g993 ( 
.A(n_979),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_979),
.Y(n_994)
);

BUFx2_ASAP7_75t_L g995 ( 
.A(n_989),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_989),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_985),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_990),
.Y(n_998)
);

OR2x2_ASAP7_75t_L g999 ( 
.A(n_995),
.B(n_978),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_995),
.B(n_984),
.Y(n_1000)
);

INVx1_ASAP7_75t_SL g1001 ( 
.A(n_996),
.Y(n_1001)
);

NAND3xp33_ASAP7_75t_L g1002 ( 
.A(n_997),
.B(n_996),
.C(n_970),
.Y(n_1002)
);

OAI21xp33_ASAP7_75t_L g1003 ( 
.A1(n_990),
.A2(n_965),
.B(n_976),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_999),
.B(n_980),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_1001),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_998),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_1000),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_1002),
.Y(n_1008)
);

BUFx2_ASAP7_75t_L g1009 ( 
.A(n_1003),
.Y(n_1009)
);

AOI22xp33_ASAP7_75t_L g1010 ( 
.A1(n_1002),
.A2(n_867),
.B1(n_917),
.B2(n_991),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_1001),
.B(n_988),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_1002),
.A2(n_917),
.B1(n_991),
.B2(n_976),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_999),
.B(n_884),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_1007),
.B(n_884),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_1005),
.Y(n_1015)
);

AOI32xp33_ASAP7_75t_L g1016 ( 
.A1(n_1008),
.A2(n_982),
.A3(n_993),
.B1(n_980),
.B2(n_981),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1011),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_1007),
.B(n_907),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_1006),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_1004),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_1010),
.A2(n_976),
.B1(n_964),
.B2(n_981),
.Y(n_1021)
);

NAND2x1_ASAP7_75t_SL g1022 ( 
.A(n_1018),
.B(n_1013),
.Y(n_1022)
);

XNOR2xp5_ASAP7_75t_L g1023 ( 
.A(n_1021),
.B(n_1009),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_1020),
.B(n_1010),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_1015),
.B(n_1012),
.Y(n_1025)
);

NOR2x1_ASAP7_75t_L g1026 ( 
.A(n_1014),
.B(n_993),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_1017),
.B(n_988),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_1019),
.B(n_896),
.Y(n_1028)
);

NOR2x1_ASAP7_75t_L g1029 ( 
.A(n_1016),
.B(n_993),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_1027),
.B(n_1012),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_1028),
.B(n_973),
.Y(n_1031)
);

NOR3x1_ASAP7_75t_L g1032 ( 
.A(n_1024),
.B(n_1025),
.C(n_1023),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_1026),
.B(n_973),
.Y(n_1033)
);

NOR2x1_ASAP7_75t_L g1034 ( 
.A(n_1029),
.B(n_993),
.Y(n_1034)
);

AOI222xp33_ASAP7_75t_L g1035 ( 
.A1(n_1022),
.A2(n_982),
.B1(n_994),
.B2(n_992),
.C1(n_875),
.C2(n_964),
.Y(n_1035)
);

OAI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_1030),
.A2(n_994),
.B1(n_992),
.B2(n_973),
.Y(n_1036)
);

NAND2xp33_ASAP7_75t_L g1037 ( 
.A(n_1034),
.B(n_875),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1035),
.B(n_969),
.Y(n_1038)
);

CKINVDCx16_ASAP7_75t_R g1039 ( 
.A(n_1031),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1033),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_1032),
.B(n_992),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_1031),
.B(n_967),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1035),
.B(n_987),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_1041),
.A2(n_994),
.B(n_992),
.C(n_987),
.Y(n_1044)
);

AOI22xp33_ASAP7_75t_L g1045 ( 
.A1(n_1042),
.A2(n_1040),
.B1(n_1037),
.B2(n_1038),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_1043),
.A2(n_994),
.B(n_986),
.Y(n_1046)
);

AOI211xp5_ASAP7_75t_L g1047 ( 
.A1(n_1036),
.A2(n_910),
.B(n_900),
.C(n_842),
.Y(n_1047)
);

AOI211xp5_ASAP7_75t_L g1048 ( 
.A1(n_1039),
.A2(n_842),
.B(n_971),
.C(n_892),
.Y(n_1048)
);

NAND3xp33_ASAP7_75t_L g1049 ( 
.A(n_1041),
.B(n_901),
.C(n_909),
.Y(n_1049)
);

AOI221xp5_ASAP7_75t_L g1050 ( 
.A1(n_1041),
.A2(n_974),
.B1(n_894),
.B2(n_898),
.C(n_971),
.Y(n_1050)
);

AOI211xp5_ASAP7_75t_SL g1051 ( 
.A1(n_1041),
.A2(n_856),
.B(n_956),
.C(n_964),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_1049),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1046),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1045),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_1051),
.B(n_968),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1044),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1054),
.Y(n_1057)
);

AOI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_1052),
.A2(n_1050),
.B1(n_1048),
.B2(n_1047),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_1056),
.A2(n_976),
.B1(n_972),
.B2(n_943),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_1053),
.A2(n_972),
.B1(n_943),
.B2(n_930),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1055),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_1054),
.B(n_964),
.Y(n_1062)
);

NAND2x1_ASAP7_75t_L g1063 ( 
.A(n_1053),
.B(n_856),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_1054),
.B(n_930),
.Y(n_1064)
);

INVxp67_ASAP7_75t_L g1065 ( 
.A(n_1054),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_1062),
.B(n_948),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1064),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_1065),
.Y(n_1068)
);

OAI21xp33_ASAP7_75t_L g1069 ( 
.A1(n_1057),
.A2(n_956),
.B(n_949),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_1061),
.A2(n_856),
.B(n_827),
.Y(n_1070)
);

AOI322xp5_ASAP7_75t_L g1071 ( 
.A1(n_1058),
.A2(n_956),
.A3(n_948),
.B1(n_955),
.B2(n_939),
.C1(n_890),
.C2(n_889),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_1063),
.A2(n_923),
.B1(n_954),
.B2(n_960),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_1059),
.B(n_960),
.Y(n_1073)
);

NOR3xp33_ASAP7_75t_L g1074 ( 
.A(n_1060),
.B(n_829),
.C(n_950),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1067),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1068),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1066),
.Y(n_1077)
);

INVx2_ASAP7_75t_SL g1078 ( 
.A(n_1073),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_1072),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_1069),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1070),
.Y(n_1081)
);

OR2x2_ASAP7_75t_L g1082 ( 
.A(n_1074),
.B(n_951),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1071),
.Y(n_1083)
);

INVx3_ASAP7_75t_L g1084 ( 
.A(n_1067),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1067),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1066),
.Y(n_1086)
);

OAI211xp5_ASAP7_75t_L g1087 ( 
.A1(n_1067),
.A2(n_923),
.B(n_829),
.C(n_946),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1084),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1084),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1075),
.A2(n_827),
.B(n_953),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_1085),
.A2(n_827),
.B1(n_951),
.B2(n_881),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1086),
.B(n_939),
.Y(n_1092)
);

NAND4xp75_ASAP7_75t_L g1093 ( 
.A(n_1076),
.B(n_936),
.C(n_158),
.D(n_159),
.Y(n_1093)
);

OR5x1_ASAP7_75t_L g1094 ( 
.A(n_1087),
.B(n_157),
.C(n_161),
.D(n_162),
.E(n_163),
.Y(n_1094)
);

AND3x4_ASAP7_75t_L g1095 ( 
.A(n_1080),
.B(n_955),
.C(n_915),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_1077),
.Y(n_1096)
);

AOI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_1096),
.A2(n_1076),
.B1(n_1078),
.B2(n_1083),
.Y(n_1097)
);

NOR4xp25_ASAP7_75t_L g1098 ( 
.A(n_1088),
.B(n_1079),
.C(n_1081),
.D(n_1082),
.Y(n_1098)
);

XOR2xp5_ASAP7_75t_L g1099 ( 
.A(n_1089),
.B(n_164),
.Y(n_1099)
);

OAI322xp33_ASAP7_75t_L g1100 ( 
.A1(n_1092),
.A2(n_1090),
.A3(n_1091),
.B1(n_1094),
.B2(n_1095),
.C1(n_1093),
.C2(n_913),
.Y(n_1100)
);

OAI221xp5_ASAP7_75t_L g1101 ( 
.A1(n_1088),
.A2(n_936),
.B1(n_879),
.B2(n_947),
.C(n_877),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1096),
.A2(n_955),
.B1(n_915),
.B2(n_940),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_1096),
.A2(n_955),
.B1(n_915),
.B2(n_940),
.Y(n_1103)
);

OAI221xp5_ASAP7_75t_L g1104 ( 
.A1(n_1097),
.A2(n_936),
.B1(n_947),
.B2(n_944),
.C(n_928),
.Y(n_1104)
);

AOI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1098),
.A2(n_1099),
.B1(n_1102),
.B2(n_1103),
.Y(n_1105)
);

AOI211xp5_ASAP7_75t_L g1106 ( 
.A1(n_1100),
.A2(n_166),
.B(n_167),
.C(n_171),
.Y(n_1106)
);

OA21x2_ASAP7_75t_L g1107 ( 
.A1(n_1105),
.A2(n_1101),
.B(n_922),
.Y(n_1107)
);

NOR3xp33_ASAP7_75t_L g1108 ( 
.A(n_1107),
.B(n_1106),
.C(n_1104),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1108),
.B(n_172),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1108),
.B(n_173),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_1109),
.Y(n_1111)
);

AOI331xp33_ASAP7_75t_L g1112 ( 
.A1(n_1110),
.A2(n_174),
.A3(n_175),
.B1(n_176),
.B2(n_178),
.B3(n_179),
.C1(n_180),
.Y(n_1112)
);

NAND2xp33_ASAP7_75t_L g1113 ( 
.A(n_1109),
.B(n_861),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1111),
.A2(n_181),
.B(n_182),
.Y(n_1114)
);

AO21x2_ASAP7_75t_L g1115 ( 
.A1(n_1113),
.A2(n_183),
.B(n_184),
.Y(n_1115)
);

AOI221xp5_ASAP7_75t_L g1116 ( 
.A1(n_1115),
.A2(n_1112),
.B1(n_186),
.B2(n_187),
.C(n_188),
.Y(n_1116)
);

AOI211xp5_ASAP7_75t_L g1117 ( 
.A1(n_1116),
.A2(n_1114),
.B(n_191),
.C(n_193),
.Y(n_1117)
);


endmodule