module fake_netlist_1_10384_n_48 (n_11, n_1, n_2, n_13, n_16, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_48);
input n_11;
input n_1;
input n_2;
input n_13;
input n_16;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_48;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_47;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_46;
wire n_25;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
OAI21x1_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_5), .B(n_15), .Y(n_17) );
BUFx6f_ASAP7_75t_L g18 ( .A(n_8), .Y(n_18) );
OAI22xp5_ASAP7_75t_L g19 ( .A1(n_3), .A2(n_6), .B1(n_11), .B2(n_8), .Y(n_19) );
CKINVDCx20_ASAP7_75t_R g20 ( .A(n_2), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_9), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_7), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_6), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_7), .B(n_0), .Y(n_24) );
AND3x1_ASAP7_75t_L g25 ( .A(n_21), .B(n_0), .C(n_1), .Y(n_25) );
HB1xp67_ASAP7_75t_L g26 ( .A(n_21), .Y(n_26) );
HB1xp67_ASAP7_75t_L g27 ( .A(n_23), .Y(n_27) );
OAI21x1_ASAP7_75t_SL g28 ( .A1(n_25), .A2(n_19), .B(n_22), .Y(n_28) );
AOI22xp33_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_23), .B1(n_22), .B2(n_24), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
AOI22xp33_ASAP7_75t_SL g31 ( .A1(n_28), .A2(n_20), .B1(n_19), .B2(n_27), .Y(n_31) );
AND2x2_ASAP7_75t_L g32 ( .A(n_31), .B(n_29), .Y(n_32) );
AOI221xp5_ASAP7_75t_L g33 ( .A1(n_30), .A2(n_20), .B1(n_24), .B2(n_22), .C(n_18), .Y(n_33) );
OAI22xp5_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_30), .B1(n_24), .B2(n_18), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_32), .Y(n_36) );
OAI22xp5_ASAP7_75t_L g37 ( .A1(n_35), .A2(n_18), .B1(n_2), .B2(n_3), .Y(n_37) );
OAI211xp5_ASAP7_75t_L g38 ( .A1(n_35), .A2(n_18), .B(n_17), .C(n_5), .Y(n_38) );
AOI21xp5_ASAP7_75t_L g39 ( .A1(n_34), .A2(n_17), .B(n_18), .Y(n_39) );
OAI22xp5_ASAP7_75t_SL g40 ( .A1(n_37), .A2(n_36), .B1(n_18), .B2(n_9), .Y(n_40) );
NOR2x1_ASAP7_75t_L g41 ( .A(n_38), .B(n_18), .Y(n_41) );
OAI22xp5_ASAP7_75t_SL g42 ( .A1(n_39), .A2(n_1), .B1(n_4), .B2(n_10), .Y(n_42) );
NOR2x1_ASAP7_75t_L g43 ( .A(n_37), .B(n_17), .Y(n_43) );
AND2x4_ASAP7_75t_L g44 ( .A(n_41), .B(n_13), .Y(n_44) );
CKINVDCx20_ASAP7_75t_R g45 ( .A(n_42), .Y(n_45) );
INVx1_ASAP7_75t_L g46 ( .A(n_40), .Y(n_46) );
OAI22xp33_ASAP7_75t_L g47 ( .A1(n_45), .A2(n_43), .B1(n_10), .B2(n_11), .Y(n_47) );
AOI322xp5_ASAP7_75t_L g48 ( .A1(n_47), .A2(n_4), .A3(n_12), .B1(n_14), .B2(n_44), .C1(n_45), .C2(n_46), .Y(n_48) );
endmodule