module fake_jpeg_15077_n_393 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_393);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_393;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

CKINVDCx6p67_ASAP7_75t_R g105 ( 
.A(n_38),
.Y(n_105)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_18),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_56),
.Y(n_71)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_51),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_17),
.B(n_7),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_52),
.B(n_57),
.Y(n_74)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_14),
.B(n_6),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_54),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_23),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_27),
.B(n_6),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_23),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_33),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_16),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_75),
.B(n_84),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_41),
.A2(n_37),
.B1(n_34),
.B2(n_29),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_78),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_17),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_81),
.B(n_88),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_46),
.A2(n_16),
.B1(n_35),
.B2(n_19),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_19),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_45),
.A2(n_34),
.B1(n_29),
.B2(n_36),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_53),
.A2(n_19),
.B1(n_35),
.B2(n_30),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_30),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_89),
.B(n_15),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_40),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_90),
.B(n_9),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_20),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_93),
.B(n_99),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_60),
.Y(n_94)
);

INVx3_ASAP7_75t_SL g150 ( 
.A(n_94),
.Y(n_150)
);

NAND2xp33_ASAP7_75t_SL g96 ( 
.A(n_49),
.B(n_20),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_31),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_32),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_42),
.B(n_32),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_100),
.B(n_106),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_48),
.A2(n_21),
.B1(n_35),
.B2(n_24),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_102),
.A2(n_115),
.B1(n_117),
.B2(n_15),
.Y(n_127)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_51),
.B(n_32),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_107),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_39),
.A2(n_21),
.B1(n_24),
.B2(n_26),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_108),
.A2(n_15),
.B1(n_6),
.B2(n_3),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_55),
.B(n_32),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_111),
.B(n_116),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_43),
.A2(n_21),
.B1(n_24),
.B2(n_26),
.Y(n_113)
);

AO22x1_ASAP7_75t_SL g120 ( 
.A1(n_113),
.A2(n_59),
.B1(n_44),
.B2(n_50),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_38),
.A2(n_26),
.B1(n_28),
.B2(n_36),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_61),
.B(n_31),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_38),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_71),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_118),
.B(n_121),
.Y(n_174)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_119),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_120),
.A2(n_73),
.B1(n_98),
.B2(n_109),
.Y(n_172)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_75),
.B(n_49),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_122),
.B(n_135),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_123),
.A2(n_136),
.B1(n_165),
.B2(n_95),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_97),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_124),
.B(n_126),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_127),
.A2(n_12),
.B(n_101),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_81),
.B(n_64),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_129),
.B(n_139),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_97),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_131),
.B(n_138),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_88),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_132),
.B(n_143),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_134),
.A2(n_114),
.B(n_105),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_84),
.B(n_15),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_104),
.A2(n_8),
.B1(n_13),
.B2(n_3),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_137),
.A2(n_109),
.B1(n_79),
.B2(n_73),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_74),
.B(n_5),
.Y(n_139)
);

XOR2x2_ASAP7_75t_L g140 ( 
.A(n_96),
.B(n_5),
.Y(n_140)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_9),
.C(n_10),
.Y(n_170)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_142),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_85),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_68),
.B(n_8),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_144),
.B(n_146),
.Y(n_192)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_69),
.Y(n_145)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_68),
.B(n_8),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_91),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_148),
.B(n_149),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_77),
.Y(n_149)
);

AO22x1_ASAP7_75t_L g151 ( 
.A1(n_79),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_151)
);

O2A1O1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_98),
.B(n_112),
.C(n_1),
.Y(n_176)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_67),
.Y(n_152)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_91),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_L g195 ( 
.A1(n_153),
.A2(n_105),
.B(n_12),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_70),
.B(n_8),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_167),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_107),
.Y(n_157)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_77),
.Y(n_159)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_159),
.Y(n_203)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_70),
.Y(n_160)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_160),
.Y(n_198)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_80),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_161),
.Y(n_191)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_80),
.Y(n_163)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_72),
.B(n_3),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_164),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_101),
.A2(n_4),
.B1(n_9),
.B2(n_10),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_114),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_72),
.B(n_4),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_113),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_170),
.A2(n_176),
.B(n_178),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_171),
.A2(n_175),
.B1(n_199),
.B2(n_121),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_172),
.A2(n_189),
.B1(n_200),
.B2(n_150),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_122),
.B(n_105),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_181),
.B(n_197),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_141),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_184),
.B(n_204),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_168),
.A2(n_110),
.B1(n_95),
.B2(n_94),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_140),
.A2(n_105),
.B(n_110),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_194),
.A2(n_151),
.B(n_148),
.Y(n_232)
);

OA21x2_ASAP7_75t_L g257 ( 
.A1(n_195),
.A2(n_176),
.B(n_194),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_135),
.B(n_92),
.C(n_82),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_132),
.B(n_82),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_212),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_141),
.Y(n_204)
);

BUFx24_ASAP7_75t_SL g205 ( 
.A(n_125),
.Y(n_205)
);

BUFx24_ASAP7_75t_SL g235 ( 
.A(n_205),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_158),
.A2(n_12),
.B1(n_1),
.B2(n_0),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_206),
.A2(n_209),
.B1(n_210),
.B2(n_169),
.Y(n_220)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_145),
.Y(n_207)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_207),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_125),
.A2(n_12),
.B1(n_1),
.B2(n_0),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_162),
.A2(n_0),
.B1(n_92),
.B2(n_133),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_144),
.B(n_146),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_154),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_214),
.B(n_153),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_155),
.B(n_167),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_215),
.A2(n_142),
.B1(n_157),
.B2(n_147),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_134),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_217),
.A2(n_232),
.B(n_241),
.Y(n_260)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_198),
.Y(n_218)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_218),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_220),
.A2(n_227),
.B1(n_230),
.B2(n_231),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_130),
.Y(n_221)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_221),
.Y(n_279)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_222),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_223),
.A2(n_252),
.B1(n_185),
.B2(n_191),
.Y(n_268)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_225),
.B(n_244),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_173),
.B(n_169),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_226),
.B(n_228),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_174),
.B(n_156),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_169),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_254),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_200),
.A2(n_120),
.B1(n_152),
.B2(n_160),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_215),
.A2(n_120),
.B1(n_126),
.B2(n_137),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_233),
.B(n_234),
.Y(n_272)
);

NOR2x1_ASAP7_75t_L g234 ( 
.A(n_170),
.B(n_151),
.Y(n_234)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_180),
.Y(n_236)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_236),
.Y(n_265)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_180),
.Y(n_237)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_237),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_198),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_238),
.B(n_243),
.Y(n_274)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_182),
.Y(n_239)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_239),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_202),
.B(n_154),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_182),
.Y(n_243)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_185),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_208),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_246),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_215),
.A2(n_119),
.B1(n_161),
.B2(n_166),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_247),
.A2(n_191),
.B1(n_183),
.B2(n_203),
.Y(n_286)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_196),
.Y(n_248)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_248),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_249),
.B(n_201),
.Y(n_290)
);

AND2x4_ASAP7_75t_L g250 ( 
.A(n_178),
.B(n_150),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_250),
.A2(n_257),
.B(n_216),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_196),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_251),
.B(n_253),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_172),
.A2(n_163),
.B1(n_131),
.B2(n_124),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_190),
.B(n_149),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_192),
.B(n_150),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_187),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_255),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_179),
.B(n_128),
.Y(n_256)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_256),
.Y(n_284)
);

AO22x2_ASAP7_75t_L g258 ( 
.A1(n_250),
.A2(n_171),
.B1(n_175),
.B2(n_189),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_258),
.A2(n_286),
.B1(n_241),
.B2(n_232),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_SL g307 ( 
.A(n_262),
.B(n_268),
.C(n_270),
.Y(n_307)
);

OAI32xp33_ASAP7_75t_L g266 ( 
.A1(n_250),
.A2(n_177),
.A3(n_212),
.B1(n_193),
.B2(n_213),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_266),
.B(n_278),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_177),
.C(n_197),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_269),
.B(n_291),
.C(n_245),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_250),
.A2(n_204),
.B(n_188),
.Y(n_270)
);

XNOR2x1_ASAP7_75t_L g278 ( 
.A(n_234),
.B(n_193),
.Y(n_278)
);

OAI32xp33_ASAP7_75t_L g280 ( 
.A1(n_224),
.A2(n_211),
.A3(n_188),
.B1(n_191),
.B2(n_201),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_280),
.B(n_247),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_248),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_283),
.B(n_219),
.Y(n_308)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_218),
.Y(n_285)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_285),
.Y(n_297)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_236),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_287),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_245),
.A2(n_211),
.B(n_183),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_288),
.A2(n_231),
.B(n_230),
.Y(n_309)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_237),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_289),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_290),
.A2(n_235),
.B1(n_291),
.B2(n_288),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_242),
.B(n_159),
.C(n_203),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_292),
.A2(n_294),
.B1(n_296),
.B2(n_304),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_273),
.A2(n_241),
.B1(n_217),
.B2(n_257),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_259),
.B(n_225),
.Y(n_295)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_295),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_258),
.A2(n_217),
.B1(n_257),
.B2(n_224),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_298),
.B(n_314),
.C(n_260),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_261),
.B(n_254),
.Y(n_299)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_299),
.Y(n_327)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_279),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_300),
.B(n_308),
.Y(n_333)
);

AOI21x1_ASAP7_75t_SL g301 ( 
.A1(n_258),
.A2(n_270),
.B(n_262),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_301),
.Y(n_321)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_264),
.Y(n_302)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_302),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_282),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_303),
.B(n_312),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_258),
.A2(n_244),
.B1(n_222),
.B2(n_239),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_264),
.B(n_246),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_306),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_309),
.B(n_310),
.Y(n_334)
);

NOR2x1_ASAP7_75t_L g311 ( 
.A(n_258),
.B(n_249),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_311),
.B(n_316),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_261),
.B(n_229),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_260),
.A2(n_220),
.B1(n_227),
.B2(n_252),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_313),
.A2(n_315),
.B1(n_317),
.B2(n_284),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_269),
.B(n_240),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_277),
.B(n_267),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_268),
.A2(n_272),
.B1(n_278),
.B2(n_290),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_266),
.B(n_280),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_263),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_302),
.Y(n_320)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_320),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_323),
.B(n_336),
.C(n_337),
.Y(n_343)
);

MAJx2_ASAP7_75t_L g324 ( 
.A(n_305),
.B(n_275),
.C(n_274),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_324),
.B(n_332),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_292),
.Y(n_326)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_326),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_303),
.Y(n_328)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_328),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_329),
.A2(n_330),
.B1(n_309),
.B2(n_294),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_313),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_299),
.B(n_281),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_331),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_314),
.B(n_289),
.C(n_265),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_298),
.B(n_287),
.C(n_265),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_305),
.B(n_271),
.C(n_276),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_341),
.B(n_336),
.C(n_334),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_330),
.A2(n_311),
.B1(n_301),
.B2(n_318),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_342),
.A2(n_346),
.B1(n_350),
.B2(n_359),
.Y(n_362)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_338),
.Y(n_344)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_344),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_333),
.B(n_284),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_345),
.B(n_351),
.C(n_352),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_326),
.A2(n_307),
.B1(n_310),
.B2(n_317),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_340),
.B(n_322),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_337),
.B(n_296),
.C(n_312),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_353),
.B(n_354),
.C(n_325),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_323),
.B(n_319),
.C(n_293),
.Y(n_354)
);

INVx5_ASAP7_75t_L g355 ( 
.A(n_328),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_355),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_341),
.B(n_307),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_356),
.B(n_332),
.C(n_325),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_329),
.A2(n_319),
.B1(n_293),
.B2(n_297),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_356),
.B(n_334),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_363),
.B(n_360),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_357),
.A2(n_321),
.B1(n_335),
.B2(n_339),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_364),
.A2(n_350),
.B1(n_355),
.B2(n_358),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_347),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_365),
.B(n_344),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_366),
.B(n_368),
.C(n_371),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_354),
.A2(n_321),
.B1(n_320),
.B2(n_327),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_367),
.B(n_369),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_343),
.B(n_297),
.C(n_324),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_343),
.B(n_352),
.C(n_353),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_372),
.B(n_373),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_374),
.B(n_378),
.C(n_362),
.Y(n_379)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_370),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_375),
.A2(n_281),
.B1(n_263),
.B2(n_285),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_366),
.B(n_349),
.C(n_331),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_379),
.B(n_378),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_381),
.B(n_348),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_377),
.A2(n_342),
.B(n_365),
.Y(n_382)
);

AOI32xp33_ASAP7_75t_L g385 ( 
.A1(n_382),
.A2(n_349),
.A3(n_376),
.B1(n_361),
.B2(n_327),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_383),
.B(n_384),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_385),
.B(n_379),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_387),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_388),
.B(n_384),
.C(n_386),
.Y(n_389)
);

AOI31xp33_ASAP7_75t_L g390 ( 
.A1(n_389),
.A2(n_376),
.A3(n_380),
.B(n_361),
.Y(n_390)
);

BUFx24_ASAP7_75t_SL g391 ( 
.A(n_390),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_391),
.B(n_271),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_392),
.B(n_276),
.Y(n_393)
);


endmodule