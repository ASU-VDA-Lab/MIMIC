module fake_jpeg_29657_n_308 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_308);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_61),
.Y(n_76)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

BUFx8_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_1),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_51),
.B(n_67),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_19),
.B(n_1),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_52),
.B(n_70),
.Y(n_100)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_18),
.B(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_21),
.B(n_2),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_64),
.Y(n_90)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g82 ( 
.A(n_66),
.B(n_27),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_21),
.B(n_3),
.Y(n_67)
);

BUFx4f_ASAP7_75t_SL g68 ( 
.A(n_35),
.Y(n_68)
);

CKINVDCx12_ASAP7_75t_R g103 ( 
.A(n_68),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_30),
.B(n_16),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_69),
.B(n_71),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_35),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_35),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_84),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_27),
.C(n_42),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_79),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_78),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_50),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_66),
.C(n_45),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_113),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_30),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_44),
.A2(n_22),
.B1(n_34),
.B2(n_28),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_85),
.A2(n_86),
.B1(n_104),
.B2(n_105),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_58),
.A2(n_42),
.B1(n_38),
.B2(n_20),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_36),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_95),
.Y(n_131)
);

NAND2xp33_ASAP7_75t_SL g94 ( 
.A(n_53),
.B(n_55),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_94),
.A2(n_24),
.B(n_6),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_36),
.Y(n_95)
);

NAND2x2_ASAP7_75t_SL g99 ( 
.A(n_68),
.B(n_34),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_99),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_65),
.A2(n_38),
.B1(n_42),
.B2(n_40),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_70),
.A2(n_38),
.B1(n_41),
.B2(n_20),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_46),
.A2(n_41),
.B1(n_32),
.B2(n_29),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_106),
.A2(n_112),
.B1(n_12),
.B2(n_13),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_64),
.A2(n_22),
.B1(n_39),
.B2(n_34),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_108),
.A2(n_114),
.B1(n_8),
.B2(n_9),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_40),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_8),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_47),
.A2(n_32),
.B1(n_29),
.B2(n_24),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_68),
.A2(n_56),
.B(n_39),
.C(n_34),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_44),
.A2(n_39),
.B1(n_28),
.B2(n_24),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_100),
.A2(n_39),
.B(n_28),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_117),
.A2(n_98),
.B(n_113),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_99),
.A2(n_24),
.B1(n_28),
.B2(n_7),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_120),
.A2(n_105),
.B1(n_86),
.B2(n_94),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_130),
.Y(n_156)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_123),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_139),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_5),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_128),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_5),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_83),
.B(n_5),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_135),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_100),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_130)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

BUFx4f_ASAP7_75t_SL g133 ( 
.A(n_103),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_134),
.B(n_142),
.Y(n_181)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_80),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_138),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_93),
.B(n_10),
.Y(n_138)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_99),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_143),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_10),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_147),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_96),
.B(n_13),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_149),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_141),
.B(n_148),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_84),
.B(n_14),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_88),
.B(n_16),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_95),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_75),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_99),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_151),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_92),
.B(n_109),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_172),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_126),
.B(n_72),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_155),
.B(n_184),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_73),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_179),
.C(n_182),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_163),
.A2(n_165),
.B1(n_166),
.B2(n_180),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_150),
.A2(n_82),
.B1(n_111),
.B2(n_79),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_131),
.A2(n_97),
.B1(n_89),
.B2(n_102),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_167),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_131),
.B(n_147),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_118),
.B(n_81),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_137),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_119),
.A2(n_121),
.B1(n_142),
.B2(n_144),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_175),
.A2(n_183),
.B1(n_139),
.B2(n_145),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_119),
.B(n_87),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_121),
.A2(n_89),
.B1(n_97),
.B2(n_102),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_119),
.B(n_91),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_134),
.A2(n_77),
.B1(n_107),
.B2(n_130),
.Y(n_183)
);

NOR3xp33_ASAP7_75t_SL g184 ( 
.A(n_146),
.B(n_77),
.C(n_122),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_156),
.A2(n_149),
.B(n_133),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_185),
.A2(n_207),
.B(n_156),
.Y(n_218)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_188),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

AND2x6_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_117),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_190),
.A2(n_213),
.B(n_187),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_152),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_133),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_192),
.Y(n_235)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_193),
.Y(n_215)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_194),
.B(n_195),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_132),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_196),
.A2(n_205),
.B1(n_162),
.B2(n_160),
.Y(n_231)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_201),
.Y(n_220)
);

AOI22x1_ASAP7_75t_L g198 ( 
.A1(n_175),
.A2(n_125),
.B1(n_116),
.B2(n_123),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_177),
.B1(n_180),
.B2(n_160),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_135),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_200),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_168),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_115),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_208),
.Y(n_226)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_203),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_181),
.A2(n_124),
.B1(n_179),
.B2(n_154),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_176),
.A2(n_165),
.B(n_170),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_157),
.B(n_155),
.Y(n_208)
);

INVx13_ASAP7_75t_L g209 ( 
.A(n_169),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_210),
.Y(n_230)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_166),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_153),
.B(n_181),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_186),
.Y(n_233)
);

AND2x6_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_181),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_171),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_227),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_218),
.A2(n_229),
.B(n_206),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_204),
.A2(n_163),
.B1(n_174),
.B2(n_153),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_221),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_204),
.A2(n_174),
.B1(n_161),
.B2(n_156),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_222),
.A2(n_196),
.B1(n_198),
.B2(n_210),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_183),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_177),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_228),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_206),
.A2(n_207),
.B(n_185),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_236),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_232),
.B(n_233),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_212),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_248),
.Y(n_263)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_214),
.Y(n_240)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_240),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_202),
.Y(n_241)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_241),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_220),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_242),
.B(n_247),
.Y(n_264)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_234),
.Y(n_244)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_244),
.Y(n_267)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_230),
.Y(n_246)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_203),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

AOI221xp5_ASAP7_75t_L g261 ( 
.A1(n_249),
.A2(n_235),
.B1(n_217),
.B2(n_221),
.C(n_219),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_253),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_229),
.A2(n_190),
.B(n_201),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_224),
.Y(n_255)
);

NOR3xp33_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_211),
.C(n_223),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_216),
.C(n_236),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_254),
.C(n_243),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_228),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_262),
.Y(n_279)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_261),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_227),
.Y(n_262)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_265),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_249),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_274),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_275),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_258),
.A2(n_251),
.B(n_253),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_218),
.B(n_258),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_225),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_254),
.C(n_232),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_252),
.C(n_256),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_240),
.C(n_187),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_277),
.B(n_278),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_269),
.B(n_186),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_267),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_215),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_262),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_284),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_283),
.A2(n_287),
.B(n_289),
.Y(n_291)
);

OAI21x1_ASAP7_75t_L g284 ( 
.A1(n_273),
.A2(n_252),
.B(n_226),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_285),
.A2(n_271),
.B(n_226),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_259),
.C(n_238),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_244),
.Y(n_294)
);

O2A1O1Ixp33_ASAP7_75t_SL g290 ( 
.A1(n_281),
.A2(n_263),
.B(n_276),
.C(n_259),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_290),
.A2(n_296),
.B(n_231),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_293),
.Y(n_298)
);

AOI322xp5_ASAP7_75t_L g293 ( 
.A1(n_286),
.A2(n_272),
.A3(n_213),
.B1(n_248),
.B2(n_246),
.C1(n_268),
.C2(n_245),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_287),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_188),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_194),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_289),
.C(n_282),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_294),
.C(n_198),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_300),
.A2(n_301),
.B1(n_215),
.B2(n_222),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_295),
.A2(n_233),
.B(n_201),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_303),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_298),
.C(n_193),
.Y(n_305)
);

AOI221xp5_ASAP7_75t_L g307 ( 
.A1(n_305),
.A2(n_304),
.B1(n_302),
.B2(n_197),
.C(n_209),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_306),
.Y(n_308)
);


endmodule