module fake_jpeg_14351_n_647 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_647);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_647;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_538;
wire n_47;
wire n_312;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_63),
.Y(n_145)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_65),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_66),
.Y(n_163)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_68),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_69),
.Y(n_190)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_71),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_73),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_74),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_75),
.Y(n_205)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_77),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_19),
.B(n_8),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_78),
.B(n_91),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_80),
.Y(n_161)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_82),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_83),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_84),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_85),
.Y(n_208)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

BUFx2_ASAP7_75t_SL g184 ( 
.A(n_86),
.Y(n_184)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

INVx3_ASAP7_75t_SL g165 ( 
.A(n_89),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_19),
.B(n_8),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_92),
.Y(n_164)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

BUFx12_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_95),
.Y(n_158)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_96),
.Y(n_194)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_98),
.Y(n_167)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_26),
.Y(n_99)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_99),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_100),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_101),
.Y(n_212)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_103),
.Y(n_177)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_104),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_105),
.Y(n_206)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_26),
.Y(n_106)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_106),
.Y(n_182)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_107),
.Y(n_185)
);

BUFx24_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

NAND2xp33_ASAP7_75t_SL g178 ( 
.A(n_108),
.B(n_109),
.Y(n_178)
);

HAxp5_ASAP7_75t_SL g109 ( 
.A(n_24),
.B(n_0),
.CON(n_109),
.SN(n_109)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_110),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_27),
.B(n_17),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_60),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_116),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_113),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_114),
.Y(n_195)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_46),
.Y(n_115)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_115),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_27),
.B(n_17),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_31),
.Y(n_153)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_46),
.Y(n_118)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_24),
.Y(n_119)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_46),
.Y(n_121)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_46),
.Y(n_122)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_36),
.Y(n_124)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_124),
.Y(n_172)
);

BUFx12_ASAP7_75t_L g125 ( 
.A(n_24),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_125),
.Y(n_152)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_36),
.Y(n_126)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

BUFx4f_ASAP7_75t_L g127 ( 
.A(n_36),
.Y(n_127)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_127),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_36),
.Y(n_128)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_128),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_36),
.Y(n_129)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_129),
.Y(n_199)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_42),
.Y(n_130)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_130),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_133),
.B(n_153),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_81),
.B(n_39),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_134),
.B(n_148),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_39),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_109),
.A2(n_36),
.B1(n_20),
.B2(n_57),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_150),
.A2(n_191),
.B(n_200),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_92),
.A2(n_31),
.B1(n_43),
.B2(n_35),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_160),
.A2(n_173),
.B1(n_183),
.B2(n_30),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_98),
.A2(n_43),
.B1(n_35),
.B2(n_29),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_115),
.B(n_29),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_179),
.B(n_188),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_112),
.B(n_44),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_180),
.B(n_186),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_100),
.A2(n_101),
.B1(n_65),
.B2(n_66),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_112),
.B(n_44),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_82),
.B(n_21),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_108),
.A2(n_123),
.B1(n_95),
.B2(n_116),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_108),
.A2(n_62),
.B1(n_57),
.B2(n_52),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_125),
.B(n_21),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_201),
.B(n_204),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_63),
.B(n_38),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_68),
.A2(n_38),
.B1(n_48),
.B2(n_52),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_209),
.A2(n_213),
.B1(n_214),
.B2(n_56),
.Y(n_265)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_127),
.Y(n_210)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_82),
.B(n_48),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_211),
.B(n_215),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_75),
.A2(n_20),
.B1(n_57),
.B2(n_52),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_114),
.A2(n_62),
.B1(n_37),
.B2(n_40),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_69),
.B(n_45),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_216),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_145),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_218),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_219),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_L g220 ( 
.A1(n_209),
.A2(n_89),
.B1(n_77),
.B2(n_79),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_220),
.A2(n_227),
.B1(n_265),
.B2(n_276),
.Y(n_335)
);

AND2x2_ASAP7_75t_SL g221 ( 
.A(n_178),
.B(n_121),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_221),
.B(n_236),
.Y(n_299)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_222),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_149),
.Y(n_223)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_223),
.Y(n_296)
);

BUFx6f_ASAP7_75t_SL g224 ( 
.A(n_131),
.Y(n_224)
);

INVx13_ASAP7_75t_L g314 ( 
.A(n_224),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_202),
.A2(n_74),
.B1(n_126),
.B2(n_20),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_225),
.A2(n_226),
.B1(n_238),
.B2(n_259),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_194),
.A2(n_37),
.B1(n_40),
.B2(n_50),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_L g227 ( 
.A1(n_150),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_169),
.Y(n_228)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_228),
.Y(n_301)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_151),
.Y(n_229)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_229),
.Y(n_305)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_137),
.Y(n_230)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_230),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_145),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_232),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_144),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_233),
.B(n_255),
.Y(n_342)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_151),
.Y(n_237)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_237),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_158),
.A2(n_37),
.B1(n_40),
.B2(n_50),
.Y(n_238)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_239),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_132),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_240),
.B(n_250),
.Y(n_297)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_177),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_241),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_159),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_242),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_161),
.A2(n_90),
.B1(n_129),
.B2(n_128),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_243),
.A2(n_251),
.B1(n_252),
.B2(n_280),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_159),
.Y(n_245)
);

INVx5_ASAP7_75t_L g306 ( 
.A(n_245),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_191),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_246),
.Y(n_332)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_138),
.Y(n_247)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_247),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_152),
.B(n_122),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_248),
.Y(n_351)
);

INVx11_ASAP7_75t_L g249 ( 
.A(n_184),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_249),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_146),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_208),
.A2(n_30),
.B1(n_113),
.B2(n_103),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_208),
.A2(n_105),
.B1(n_156),
.B2(n_62),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_139),
.Y(n_253)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_253),
.Y(n_311)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_155),
.Y(n_254)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_254),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_147),
.B(n_50),
.Y(n_255)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_171),
.Y(n_257)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_257),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_131),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_258),
.B(n_267),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_158),
.A2(n_45),
.B1(n_59),
.B2(n_56),
.Y(n_259)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_163),
.Y(n_260)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_260),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_203),
.Y(n_261)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_261),
.Y(n_345)
);

AOI22x1_ASAP7_75t_L g262 ( 
.A1(n_135),
.A2(n_94),
.B1(n_59),
.B2(n_56),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_262),
.A2(n_287),
.B(n_141),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_136),
.B(n_59),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_263),
.B(n_278),
.Y(n_344)
);

INVx8_ASAP7_75t_L g264 ( 
.A(n_163),
.Y(n_264)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_264),
.Y(n_348)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_182),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_266),
.B(n_271),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_195),
.A2(n_51),
.B1(n_32),
.B2(n_47),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_172),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_268),
.B(n_269),
.Y(n_315)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_193),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_197),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_270),
.B(n_272),
.Y(n_320)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_199),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_198),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_177),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_273),
.B(n_274),
.Y(n_350)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_206),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_214),
.A2(n_51),
.B1(n_32),
.B2(n_47),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_206),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_277),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_170),
.B(n_51),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_156),
.A2(n_32),
.B1(n_47),
.B2(n_9),
.Y(n_280)
);

NAND2x1_ASAP7_75t_L g281 ( 
.A(n_136),
.B(n_47),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_281),
.B(n_176),
.C(n_187),
.Y(n_322)
);

OAI22xp33_ASAP7_75t_L g282 ( 
.A1(n_200),
.A2(n_47),
.B1(n_16),
.B2(n_14),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_282),
.A2(n_165),
.B1(n_140),
.B2(n_190),
.Y(n_298)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_175),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_283),
.B(n_285),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_142),
.B(n_16),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_284),
.B(n_290),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_165),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_143),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_286),
.B(n_288),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_190),
.A2(n_16),
.B1(n_12),
.B2(n_11),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_154),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_157),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_289),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_140),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_174),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_291),
.B(n_162),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_298),
.A2(n_304),
.B1(n_319),
.B2(n_321),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_246),
.A2(n_212),
.B1(n_181),
.B2(n_167),
.Y(n_302)
);

AO21x2_ASAP7_75t_L g357 ( 
.A1(n_302),
.A2(n_325),
.B(n_258),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_256),
.A2(n_162),
.B1(n_196),
.B2(n_135),
.Y(n_304)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_316),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_256),
.A2(n_192),
.B1(n_196),
.B2(n_205),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_236),
.A2(n_235),
.B1(n_217),
.B2(n_220),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_322),
.A2(n_328),
.B(n_222),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_243),
.A2(n_174),
.B1(n_207),
.B2(n_205),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_324),
.A2(n_330),
.B1(n_333),
.B2(n_340),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_276),
.A2(n_212),
.B1(n_164),
.B2(n_181),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_227),
.A2(n_231),
.B1(n_221),
.B2(n_255),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_279),
.B(n_167),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_341),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_244),
.A2(n_207),
.B1(n_164),
.B2(n_168),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_262),
.A2(n_185),
.B1(n_141),
.B2(n_2),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_223),
.B(n_0),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_262),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_343),
.A2(n_346),
.B1(n_264),
.B2(n_291),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_221),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_281),
.B(n_16),
.C(n_12),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_347),
.B(n_230),
.C(n_228),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_275),
.B(n_12),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_349),
.B(n_12),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_329),
.B(n_234),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_355),
.B(n_363),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_335),
.A2(n_282),
.B1(n_229),
.B2(n_237),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_356),
.A2(n_298),
.B1(n_310),
.B2(n_350),
.Y(n_410)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_357),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_341),
.B(n_248),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_358),
.B(n_359),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_344),
.B(n_248),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_331),
.B(n_247),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_360),
.B(n_362),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_308),
.Y(n_361)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_361),
.Y(n_420)
);

A2O1A1Ixp33_ASAP7_75t_L g362 ( 
.A1(n_299),
.A2(n_224),
.B(n_249),
.C(n_253),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_299),
.B(n_266),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_299),
.B(n_322),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_364),
.B(n_358),
.Y(n_419)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_296),
.Y(n_365)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_365),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_329),
.B(n_257),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_366),
.B(n_375),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_308),
.A2(n_239),
.B(n_261),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_367),
.A2(n_372),
.B(n_392),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_297),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_368),
.B(n_379),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_332),
.A2(n_273),
.B1(n_241),
.B2(n_274),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_369),
.A2(n_378),
.B(n_388),
.Y(n_432)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_296),
.Y(n_370)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_370),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_308),
.A2(n_289),
.B(n_283),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_301),
.Y(n_373)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_373),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_342),
.B(n_216),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_376),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_377),
.A2(n_387),
.B1(n_390),
.B2(n_393),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_349),
.B(n_271),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_380),
.B(n_381),
.Y(n_408)
);

O2A1O1Ixp33_ASAP7_75t_SL g381 ( 
.A1(n_330),
.A2(n_277),
.B(n_270),
.C(n_219),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_313),
.B(n_260),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_382),
.B(n_385),
.Y(n_427)
);

INVx6_ASAP7_75t_L g383 ( 
.A(n_292),
.Y(n_383)
);

INVx5_ASAP7_75t_L g400 ( 
.A(n_383),
.Y(n_400)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_306),
.Y(n_384)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_384),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_351),
.B(n_10),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_320),
.Y(n_386)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_386),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_321),
.A2(n_245),
.B1(n_242),
.B2(n_232),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_313),
.B(n_218),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_315),
.Y(n_389)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_389),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_319),
.A2(n_11),
.B1(n_10),
.B2(n_4),
.Y(n_390)
);

CKINVDCx14_ASAP7_75t_R g391 ( 
.A(n_350),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_391),
.B(n_398),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_328),
.A2(n_10),
.B(n_3),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_304),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_295),
.A2(n_340),
.B1(n_335),
.B2(n_324),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_394),
.A2(n_352),
.B1(n_311),
.B2(n_309),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_351),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_395),
.A2(n_300),
.B1(n_348),
.B2(n_317),
.Y(n_412)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_301),
.Y(n_396)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_396),
.Y(n_437)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_337),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_397),
.Y(n_424)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_300),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_334),
.A2(n_6),
.B(n_7),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_399),
.A2(n_392),
.B(n_367),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_394),
.A2(n_295),
.B1(n_316),
.B2(n_343),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_402),
.A2(n_421),
.B1(n_433),
.B2(n_436),
.Y(n_449)
);

AOI32xp33_ASAP7_75t_L g409 ( 
.A1(n_378),
.A2(n_346),
.A3(n_317),
.B1(n_310),
.B2(n_333),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_409),
.A2(n_418),
.B(n_385),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_410),
.A2(n_412),
.B1(n_430),
.B2(n_434),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_361),
.A2(n_347),
.B(n_350),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_414),
.A2(n_435),
.B(n_362),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_356),
.A2(n_326),
.B1(n_348),
.B2(n_323),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_415),
.A2(n_416),
.B1(n_417),
.B2(n_438),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_354),
.A2(n_326),
.B1(n_323),
.B2(n_305),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_354),
.A2(n_305),
.B1(n_339),
.B2(n_352),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_419),
.B(n_376),
.C(n_398),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_374),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_361),
.A2(n_339),
.B1(n_306),
.B2(n_293),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_364),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_372),
.A2(n_303),
.B(n_345),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_374),
.A2(n_294),
.B1(n_307),
.B2(n_318),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_364),
.A2(n_371),
.B1(n_360),
.B2(n_397),
.Y(n_438)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_407),
.Y(n_440)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_440),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_419),
.B(n_359),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_441),
.B(n_452),
.C(n_454),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_404),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_442),
.B(n_467),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_424),
.B(n_353),
.Y(n_443)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_443),
.Y(n_494)
);

A2O1A1O1Ixp25_ASAP7_75t_L g444 ( 
.A1(n_423),
.A2(n_363),
.B(n_353),
.C(n_366),
.D(n_375),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_444),
.A2(n_451),
.B(n_453),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_432),
.Y(n_445)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_445),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_418),
.A2(n_399),
.B(n_391),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_446),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_424),
.B(n_368),
.Y(n_447)
);

CKINVDCx14_ASAP7_75t_R g498 ( 
.A(n_447),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_448),
.A2(n_455),
.B(n_464),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_418),
.A2(n_369),
.B(n_370),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_426),
.B(n_365),
.C(n_355),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_431),
.A2(n_420),
.B(n_423),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_432),
.Y(n_456)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_456),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_402),
.A2(n_371),
.B1(n_381),
.B2(n_377),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_457),
.A2(n_466),
.B1(n_475),
.B2(n_412),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_404),
.B(n_382),
.Y(n_458)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_458),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_417),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_459),
.B(n_474),
.Y(n_482)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_407),
.Y(n_460)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_460),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_438),
.A2(n_387),
.B1(n_393),
.B2(n_357),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_461),
.A2(n_465),
.B1(n_470),
.B2(n_429),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_419),
.B(n_379),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_462),
.B(n_463),
.C(n_472),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_401),
.B(n_338),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_431),
.A2(n_362),
.B(n_381),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_408),
.A2(n_357),
.B1(n_390),
.B2(n_388),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_429),
.A2(n_433),
.B1(n_405),
.B2(n_436),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_434),
.B(n_396),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_408),
.A2(n_357),
.B(n_373),
.Y(n_469)
);

NAND2x1_ASAP7_75t_L g505 ( 
.A(n_469),
.B(n_437),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_410),
.A2(n_357),
.B1(n_384),
.B2(n_383),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_434),
.B(n_395),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_471),
.B(n_473),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_401),
.B(n_414),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_411),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_411),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_413),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_413),
.B(n_384),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_476),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_480),
.A2(n_500),
.B1(n_430),
.B2(n_357),
.Y(n_541)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_447),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_481),
.B(n_484),
.Y(n_529)
);

CKINVDCx16_ASAP7_75t_R g484 ( 
.A(n_458),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_452),
.B(n_414),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_485),
.B(n_488),
.Y(n_518)
);

XNOR2x2_ASAP7_75t_SL g487 ( 
.A(n_472),
.B(n_403),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_487),
.B(n_465),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_462),
.B(n_403),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_466),
.A2(n_405),
.B1(n_420),
.B2(n_409),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_490),
.A2(n_496),
.B1(n_461),
.B2(n_470),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_SL g491 ( 
.A(n_441),
.B(n_425),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_SL g527 ( 
.A(n_491),
.B(n_502),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_454),
.B(n_425),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_492),
.B(n_495),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_463),
.B(n_427),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_451),
.B(n_403),
.C(n_435),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_499),
.B(n_503),
.C(n_504),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_468),
.A2(n_421),
.B1(n_435),
.B2(n_439),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_SL g502 ( 
.A(n_443),
.B(n_427),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_442),
.B(n_428),
.C(n_437),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_455),
.B(n_448),
.C(n_446),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_505),
.A2(n_464),
.B(n_453),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_444),
.B(n_469),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_507),
.B(n_488),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_510),
.B(n_406),
.Y(n_511)
);

CKINVDCx14_ASAP7_75t_R g547 ( 
.A(n_511),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_478),
.A2(n_505),
.B(n_501),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_512),
.A2(n_517),
.B(n_514),
.Y(n_553)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_483),
.Y(n_513)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_513),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_L g564 ( 
.A1(n_514),
.A2(n_474),
.B(n_473),
.Y(n_564)
);

CKINVDCx16_ASAP7_75t_R g515 ( 
.A(n_483),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_515),
.B(n_516),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_480),
.A2(n_449),
.B1(n_457),
.B2(n_459),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_478),
.A2(n_505),
.B(n_501),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_498),
.B(n_406),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_519),
.B(n_533),
.Y(n_565)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_506),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_520),
.A2(n_525),
.B1(n_530),
.B2(n_532),
.Y(n_550)
);

XNOR2x1_ASAP7_75t_L g543 ( 
.A(n_521),
.B(n_528),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_494),
.B(n_467),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_524),
.B(n_537),
.Y(n_542)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_506),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_486),
.B(n_468),
.C(n_450),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_526),
.B(n_531),
.C(n_534),
.Y(n_544)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_477),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_486),
.B(n_450),
.C(n_471),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_508),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_494),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_485),
.B(n_449),
.C(n_476),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_482),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_535),
.A2(n_536),
.B(n_540),
.Y(n_554)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_510),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_509),
.B(n_475),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_538),
.B(n_490),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_500),
.A2(n_415),
.B1(n_412),
.B2(n_444),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_539),
.A2(n_541),
.B1(n_499),
.B2(n_439),
.Y(n_557)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_503),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_523),
.B(n_489),
.C(n_492),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_545),
.B(n_548),
.C(n_555),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_546),
.A2(n_541),
.B1(n_535),
.B2(n_513),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_523),
.B(n_489),
.C(n_479),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_522),
.B(n_504),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_549),
.B(n_345),
.Y(n_585)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_518),
.B(n_507),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_551),
.B(n_552),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_518),
.B(n_491),
.Y(n_552)
);

OAI21xp5_ASAP7_75t_L g580 ( 
.A1(n_553),
.A2(n_559),
.B(n_564),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_540),
.B(n_493),
.C(n_497),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_531),
.B(n_497),
.C(n_487),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_556),
.B(n_560),
.C(n_527),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_557),
.A2(n_566),
.B1(n_561),
.B2(n_564),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_522),
.B(n_495),
.Y(n_558)
);

XOR2xp5_ASAP7_75t_L g577 ( 
.A(n_558),
.B(n_562),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_512),
.A2(n_517),
.B(n_521),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_526),
.B(n_502),
.C(n_460),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_528),
.B(n_534),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_539),
.A2(n_440),
.B1(n_428),
.B2(n_422),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_567),
.B(n_580),
.Y(n_588)
);

CKINVDCx14_ASAP7_75t_R g568 ( 
.A(n_565),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_568),
.A2(n_575),
.B1(n_581),
.B2(n_551),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_570),
.B(n_585),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_547),
.B(n_511),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_571),
.B(n_572),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_560),
.B(n_525),
.C(n_520),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_544),
.B(n_533),
.C(n_536),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_574),
.B(n_578),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_566),
.A2(n_538),
.B1(n_529),
.B2(n_537),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_546),
.A2(n_524),
.B1(n_530),
.B2(n_532),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_576),
.A2(n_583),
.B1(n_559),
.B2(n_556),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_544),
.B(n_527),
.C(n_422),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_545),
.B(n_430),
.C(n_416),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_579),
.B(n_584),
.Y(n_598)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_550),
.Y(n_582)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_582),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_563),
.A2(n_400),
.B1(n_383),
.B2(n_303),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_542),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_555),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_586),
.B(n_587),
.Y(n_599)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_554),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_588),
.B(n_600),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_SL g589 ( 
.A1(n_569),
.A2(n_548),
.B(n_553),
.Y(n_589)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_589),
.A2(n_400),
.B(n_300),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_569),
.B(n_574),
.C(n_577),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_591),
.B(n_592),
.Y(n_606)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_585),
.B(n_557),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_572),
.B(n_562),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_594),
.B(n_595),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_577),
.B(n_549),
.C(n_558),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g600 ( 
.A(n_573),
.B(n_543),
.Y(n_600)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_601),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_602),
.A2(n_581),
.B1(n_584),
.B2(n_570),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_579),
.B(n_380),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_603),
.B(n_605),
.Y(n_618)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_573),
.B(n_543),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_L g617 ( 
.A(n_604),
.B(n_311),
.Y(n_617)
);

XNOR2xp5_ASAP7_75t_L g605 ( 
.A(n_580),
.B(n_552),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_591),
.B(n_567),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_608),
.B(n_609),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_596),
.A2(n_576),
.B1(n_578),
.B2(n_542),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_610),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_597),
.B(n_583),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_611),
.B(n_612),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_588),
.B(n_400),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_613),
.A2(n_592),
.B(n_600),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_594),
.B(n_307),
.C(n_309),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_615),
.B(n_590),
.Y(n_625)
);

O2A1O1Ixp33_ASAP7_75t_SL g616 ( 
.A1(n_599),
.A2(n_327),
.B(n_312),
.C(n_314),
.Y(n_616)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_616),
.Y(n_627)
);

XOR2xp5_ASAP7_75t_L g624 ( 
.A(n_617),
.B(n_605),
.Y(n_624)
);

INVxp67_ASAP7_75t_L g622 ( 
.A(n_614),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_622),
.B(n_628),
.Y(n_631)
);

XOR2xp5_ASAP7_75t_L g634 ( 
.A(n_624),
.B(n_625),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_L g626 ( 
.A1(n_618),
.A2(n_593),
.B(n_598),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_626),
.B(n_607),
.Y(n_636)
);

OAI21xp5_ASAP7_75t_SL g628 ( 
.A1(n_606),
.A2(n_595),
.B(n_590),
.Y(n_628)
);

INVxp67_ASAP7_75t_L g633 ( 
.A(n_629),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_619),
.B(n_604),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_630),
.B(n_615),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_SL g639 ( 
.A(n_632),
.B(n_623),
.Y(n_639)
);

OAI321xp33_ASAP7_75t_L g635 ( 
.A1(n_621),
.A2(n_616),
.A3(n_610),
.B1(n_609),
.B2(n_607),
.C(n_617),
.Y(n_635)
);

NOR3xp33_ASAP7_75t_L g638 ( 
.A(n_635),
.B(n_636),
.C(n_623),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_620),
.B(n_318),
.C(n_327),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_637),
.B(n_627),
.C(n_312),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_SL g643 ( 
.A1(n_638),
.A2(n_631),
.B(n_633),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_639),
.B(n_640),
.C(n_641),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_634),
.B(n_627),
.C(n_336),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_SL g644 ( 
.A1(n_643),
.A2(n_631),
.B(n_336),
.Y(n_644)
);

A2O1A1Ixp33_ASAP7_75t_L g645 ( 
.A1(n_644),
.A2(n_642),
.B(n_314),
.C(n_6),
.Y(n_645)
);

XOR2xp5_ASAP7_75t_L g646 ( 
.A(n_645),
.B(n_314),
.Y(n_646)
);

XOR2xp5_ASAP7_75t_L g647 ( 
.A(n_646),
.B(n_6),
.Y(n_647)
);


endmodule