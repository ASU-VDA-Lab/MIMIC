module fake_jpeg_3612_n_675 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_675);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_675;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_11),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_59),
.B(n_71),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_60),
.Y(n_154)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_61),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_62),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_63),
.Y(n_178)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_65),
.Y(n_211)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_68),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_69),
.Y(n_162)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_70),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_44),
.Y(n_71)
);

BUFx2_ASAP7_75t_R g72 ( 
.A(n_50),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_72),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_73),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_31),
.B(n_18),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_74),
.B(n_94),
.Y(n_136)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_75),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_76),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_44),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_77),
.B(n_78),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_41),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_79),
.B(n_98),
.Y(n_160)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_23),
.B(n_0),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_80),
.B(n_4),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_81),
.Y(n_200)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_82),
.Y(n_201)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_83),
.Y(n_212)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_85),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_88),
.Y(n_209)
);

BUFx10_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

CKINVDCx6p67_ASAP7_75t_R g191 ( 
.A(n_89),
.Y(n_191)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_90),
.Y(n_180)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_92),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_93),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_41),
.B(n_0),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_23),
.Y(n_95)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_96),
.Y(n_179)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_97),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_51),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_34),
.Y(n_99)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_99),
.Y(n_202)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_100),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_51),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_101),
.B(n_103),
.Y(n_171)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_27),
.Y(n_102)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_24),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_20),
.Y(n_104)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_104),
.Y(n_158)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_27),
.Y(n_105)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_22),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_106),
.B(n_116),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_28),
.B(n_0),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_107),
.B(n_108),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_30),
.B(n_17),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_34),
.Y(n_109)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_27),
.Y(n_110)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_28),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_42),
.Y(n_112)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_27),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_113),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_114),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_28),
.B(n_2),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_117),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_25),
.B(n_2),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_33),
.B(n_3),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_27),
.Y(n_118)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_118),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_24),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_119),
.B(n_124),
.Y(n_198)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_35),
.Y(n_120)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_120),
.Y(n_214)
);

BUFx12_ASAP7_75t_L g121 ( 
.A(n_42),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_121),
.Y(n_205)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_45),
.Y(n_122)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_122),
.Y(n_188)
);

INVx6_ASAP7_75t_SL g123 ( 
.A(n_42),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_123),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_34),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_35),
.B(n_4),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_53),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_56),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_126),
.B(n_130),
.Y(n_199)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_37),
.Y(n_127)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_127),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_25),
.Y(n_128)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_45),
.Y(n_129)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_129),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_37),
.Y(n_130)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_45),
.Y(n_131)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_42),
.Y(n_132)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_132),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_130),
.B(n_58),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_142),
.B(n_164),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_80),
.A2(n_45),
.B1(n_30),
.B2(n_40),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_144),
.A2(n_93),
.B1(n_111),
.B2(n_121),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_87),
.A2(n_25),
.B1(n_53),
.B2(n_47),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g247 ( 
.A(n_145),
.B(n_166),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_26),
.B1(n_45),
.B2(n_58),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_146),
.A2(n_176),
.B1(n_185),
.B2(n_193),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_66),
.B(n_57),
.C(n_38),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_148),
.B(n_229),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_65),
.A2(n_43),
.B1(n_32),
.B2(n_40),
.Y(n_166)
);

NAND3xp33_ASAP7_75t_SL g168 ( 
.A(n_96),
.B(n_57),
.C(n_48),
.Y(n_168)
);

OA21x2_ASAP7_75t_L g255 ( 
.A1(n_168),
.A2(n_121),
.B(n_89),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_116),
.B(n_48),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_170),
.B(n_173),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_80),
.B(n_38),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_175),
.B(n_221),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_60),
.A2(n_26),
.B1(n_47),
.B2(n_46),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_60),
.A2(n_26),
.B1(n_46),
.B2(n_43),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_104),
.A2(n_32),
.B1(n_22),
.B2(n_52),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_187),
.A2(n_193),
.B1(n_146),
.B2(n_185),
.Y(n_279)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_97),
.Y(n_190)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_190),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_62),
.A2(n_52),
.B1(n_20),
.B2(n_56),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_128),
.B(n_4),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_194),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_102),
.B(n_5),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_195),
.B(n_204),
.Y(n_253)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_105),
.Y(n_197)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_197),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_129),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_203),
.B(n_206),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_118),
.B(n_5),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_100),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_67),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_207),
.A2(n_224),
.B1(n_230),
.B2(n_16),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_92),
.B(n_5),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_208),
.B(n_219),
.Y(n_258)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_64),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_210),
.Y(n_239)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_122),
.Y(n_213)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_213),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_95),
.B(n_7),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_215),
.B(n_226),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_92),
.B(n_114),
.Y(n_219)
);

AND2x2_ASAP7_75t_SL g221 ( 
.A(n_62),
.B(n_7),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_72),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_222)
);

AOI21xp33_ASAP7_75t_L g260 ( 
.A1(n_222),
.A2(n_15),
.B(n_16),
.Y(n_260)
);

INVx11_ASAP7_75t_L g223 ( 
.A(n_112),
.Y(n_223)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_68),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_110),
.B(n_8),
.Y(n_226)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_131),
.Y(n_228)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_228),
.Y(n_286)
);

AO21x1_ASAP7_75t_L g229 ( 
.A1(n_99),
.A2(n_8),
.B(n_12),
.Y(n_229)
);

AO22x1_ASAP7_75t_L g232 ( 
.A1(n_229),
.A2(n_73),
.B1(n_114),
.B2(n_132),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_109),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_63),
.B(n_12),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_231),
.B(n_184),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_232),
.B(n_279),
.Y(n_328)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_135),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_233),
.Y(n_339)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_155),
.Y(n_234)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_234),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_181),
.A2(n_84),
.B1(n_76),
.B2(n_69),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_236),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_135),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_237),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_171),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_238),
.B(n_273),
.Y(n_364)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_159),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g366 ( 
.A(n_240),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_172),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_242),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_175),
.B(n_90),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_243),
.B(n_249),
.Y(n_321)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_163),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_246),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_149),
.B(n_88),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_139),
.A2(n_86),
.B1(n_81),
.B2(n_85),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_251),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_199),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_254),
.B(n_272),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_255),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_257),
.A2(n_270),
.B1(n_280),
.B2(n_313),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_221),
.B(n_15),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_259),
.B(n_264),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_260),
.A2(n_259),
.B(n_261),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_153),
.Y(n_262)
);

INVx6_ASAP7_75t_L g362 ( 
.A(n_262),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_153),
.Y(n_263)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_263),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_150),
.B(n_15),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_265),
.A2(n_282),
.B1(n_141),
.B2(n_281),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_266),
.B(n_267),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_160),
.B(n_16),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_201),
.Y(n_268)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_268),
.Y(n_320)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_212),
.Y(n_269)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_269),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_133),
.A2(n_89),
.B1(n_134),
.B2(n_214),
.Y(n_270)
);

AND2x2_ASAP7_75t_SL g271 ( 
.A(n_140),
.B(n_147),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_271),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_191),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_136),
.B(n_216),
.Y(n_273)
);

BUFx12f_ASAP7_75t_L g274 ( 
.A(n_154),
.Y(n_274)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_274),
.Y(n_358)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_137),
.Y(n_275)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_275),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_198),
.B(n_220),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_276),
.B(n_281),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_211),
.B(n_152),
.Y(n_277)
);

AND2x2_ASAP7_75t_SL g318 ( 
.A(n_277),
.B(n_289),
.Y(n_318)
);

BUFx12_ASAP7_75t_L g278 ( 
.A(n_191),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_278),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_168),
.A2(n_222),
.B1(n_194),
.B2(n_180),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_191),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_139),
.A2(n_158),
.B1(n_179),
.B2(n_211),
.Y(n_282)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_162),
.Y(n_283)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_283),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_217),
.B(n_220),
.Y(n_285)
);

AOI21xp33_ASAP7_75t_L g373 ( 
.A1(n_285),
.A2(n_295),
.B(n_299),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_287),
.B(n_312),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_156),
.B(n_177),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_288),
.B(n_296),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_158),
.B(n_183),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_180),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_290),
.B(n_291),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_225),
.Y(n_291)
);

AND2x2_ASAP7_75t_SL g292 ( 
.A(n_169),
.B(n_188),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_292),
.B(n_243),
.C(n_288),
.Y(n_375)
);

INVx5_ASAP7_75t_L g293 ( 
.A(n_154),
.Y(n_293)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_293),
.Y(n_330)
);

O2A1O1Ixp33_ASAP7_75t_L g294 ( 
.A1(n_176),
.A2(n_205),
.B(n_178),
.C(n_223),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_294),
.A2(n_272),
.B(n_232),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_138),
.B(n_172),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_189),
.B(n_167),
.Y(n_296)
);

INVx5_ASAP7_75t_L g297 ( 
.A(n_196),
.Y(n_297)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_297),
.Y(n_338)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_151),
.Y(n_298)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_298),
.Y(n_342)
);

NOR2x1_ASAP7_75t_R g299 ( 
.A(n_178),
.B(n_230),
.Y(n_299)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_196),
.Y(n_300)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_300),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_162),
.Y(n_301)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_301),
.Y(n_355)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_182),
.Y(n_302)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_302),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_224),
.B(n_161),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_303),
.B(n_316),
.Y(n_340)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_137),
.Y(n_304)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_304),
.Y(n_363)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_182),
.Y(n_305)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_305),
.Y(n_368)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_228),
.Y(n_306)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_306),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_157),
.B(n_143),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_307),
.B(n_308),
.Y(n_369)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_210),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_225),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_309),
.B(n_310),
.Y(n_377)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_143),
.Y(n_310)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_151),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_200),
.A2(n_227),
.B1(n_202),
.B2(n_157),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_174),
.B(n_202),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_314),
.B(n_297),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_L g315 ( 
.A1(n_200),
.A2(n_227),
.B1(n_161),
.B2(n_192),
.Y(n_315)
);

OA22x2_ASAP7_75t_L g354 ( 
.A1(n_315),
.A2(n_233),
.B1(n_283),
.B2(n_301),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_209),
.B(n_174),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_209),
.B(n_186),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_317),
.B(n_292),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_303),
.A2(n_192),
.B1(n_165),
.B2(n_218),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_322),
.A2(n_371),
.B1(n_244),
.B2(n_293),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g325 ( 
.A(n_261),
.B(n_165),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_325),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_247),
.A2(n_141),
.B1(n_186),
.B2(n_218),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_327),
.A2(n_336),
.B1(n_255),
.B2(n_317),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_329),
.Y(n_387)
);

AOI22x1_ASAP7_75t_SL g335 ( 
.A1(n_248),
.A2(n_141),
.B1(n_235),
.B2(n_249),
.Y(n_335)
);

NOR2x1_ASAP7_75t_L g391 ( 
.A(n_335),
.B(n_361),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_247),
.A2(n_280),
.B1(n_257),
.B2(n_287),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_271),
.B(n_277),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_344),
.B(n_346),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_345),
.A2(n_372),
.B(n_244),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_271),
.B(n_277),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_353),
.B(n_356),
.Y(n_401)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_354),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_256),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_289),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_357),
.B(n_379),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_292),
.B(n_289),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_299),
.A2(n_258),
.B1(n_254),
.B2(n_239),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_261),
.A2(n_255),
.B(n_294),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_375),
.B(n_252),
.C(n_239),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_376),
.B(n_284),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_328),
.A2(n_245),
.B1(n_253),
.B2(n_296),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_380),
.A2(n_388),
.B1(n_399),
.B2(n_410),
.Y(n_467)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_342),
.Y(n_381)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_381),
.Y(n_430)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_366),
.Y(n_382)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_382),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_383),
.A2(n_400),
.B(n_414),
.Y(n_431)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_342),
.Y(n_384)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_384),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_364),
.B(n_311),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_385),
.B(n_386),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_331),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_328),
.A2(n_316),
.B1(n_264),
.B2(n_298),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_366),
.Y(n_389)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_389),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_390),
.B(n_318),
.Y(n_439)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_366),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_392),
.B(n_397),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_321),
.B(n_250),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_393),
.B(n_398),
.Y(n_435)
);

FAx1_ASAP7_75t_SL g395 ( 
.A(n_375),
.B(n_241),
.CI(n_284),
.CON(n_395),
.SN(n_395)
);

NOR4xp25_ASAP7_75t_L g449 ( 
.A(n_395),
.B(n_320),
.C(n_323),
.D(n_368),
.Y(n_449)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_352),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_396),
.Y(n_451)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_360),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_321),
.B(n_241),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_328),
.A2(n_312),
.B1(n_237),
.B2(n_262),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_402),
.B(n_421),
.C(n_422),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_377),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_404),
.B(n_407),
.Y(n_437)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_352),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_405),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_347),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_406),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_350),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_367),
.B(n_252),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_410),
.B(n_413),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_336),
.A2(n_304),
.B1(n_275),
.B2(n_263),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_411),
.A2(n_412),
.B1(n_423),
.B2(n_422),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_340),
.A2(n_286),
.B1(n_306),
.B2(n_300),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_367),
.B(n_286),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_372),
.A2(n_278),
.B(n_274),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_415),
.A2(n_426),
.B(n_353),
.Y(n_440)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_360),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_416),
.B(n_418),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_348),
.B(n_278),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_417),
.Y(n_464)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_368),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_340),
.B(n_274),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_419),
.B(n_420),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_332),
.B(n_376),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_332),
.B(n_325),
.C(n_374),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_332),
.B(n_325),
.C(n_318),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_326),
.A2(n_351),
.B1(n_335),
.B2(n_345),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_349),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_424),
.B(n_425),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_349),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_373),
.A2(n_337),
.B(n_341),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_359),
.B(n_333),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_427),
.B(n_393),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_319),
.B(n_365),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_428),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_423),
.A2(n_337),
.B1(n_341),
.B2(n_346),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_429),
.A2(n_433),
.B1(n_434),
.B2(n_438),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_383),
.A2(n_346),
.B1(n_344),
.B2(n_361),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_414),
.A2(n_408),
.B1(n_411),
.B2(n_413),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_408),
.A2(n_344),
.B1(n_361),
.B2(n_318),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_439),
.B(n_380),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_440),
.A2(n_446),
.B(n_449),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_391),
.A2(n_327),
.B(n_324),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_441),
.A2(n_443),
.B(n_440),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_391),
.A2(n_415),
.B(n_426),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_420),
.B(n_325),
.C(n_359),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_445),
.B(n_447),
.C(n_394),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_409),
.A2(n_322),
.B(n_369),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_402),
.B(n_320),
.C(n_323),
.Y(n_447)
);

AO21x1_ASAP7_75t_SL g454 ( 
.A1(n_395),
.A2(n_409),
.B(n_390),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_462),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_394),
.A2(n_387),
.B(n_403),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_457),
.A2(n_458),
.B(n_330),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_401),
.A2(n_343),
.B(n_363),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_388),
.A2(n_354),
.B1(n_355),
.B2(n_338),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_459),
.A2(n_412),
.B1(n_382),
.B2(n_389),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_460),
.B(n_418),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_398),
.B(n_363),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_466),
.B(n_467),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_427),
.B(n_419),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_468),
.B(n_469),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_387),
.A2(n_354),
.B1(n_355),
.B2(n_334),
.Y(n_469)
);

AO22x1_ASAP7_75t_L g470 ( 
.A1(n_394),
.A2(n_354),
.B1(n_343),
.B2(n_338),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_470),
.B(n_358),
.Y(n_509)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_465),
.Y(n_473)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_473),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_437),
.B(n_407),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_474),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_404),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_475),
.B(n_476),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_464),
.B(n_386),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_456),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_477),
.B(n_478),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_456),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_479),
.B(n_492),
.C(n_504),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_480),
.A2(n_508),
.B1(n_470),
.B2(n_434),
.Y(n_523)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_465),
.Y(n_481)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_481),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_467),
.A2(n_421),
.B1(n_395),
.B2(n_399),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_482),
.A2(n_487),
.B1(n_493),
.B2(n_446),
.Y(n_531)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_448),
.Y(n_483)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_483),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_485),
.B(n_442),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_486),
.A2(n_499),
.B(n_502),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_437),
.B(n_425),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_488),
.B(n_491),
.Y(n_511)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_448),
.Y(n_489)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_489),
.Y(n_514)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_430),
.Y(n_490)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_490),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_R g491 ( 
.A1(n_454),
.A2(n_416),
.B1(n_397),
.B2(n_392),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_442),
.B(n_330),
.C(n_378),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_462),
.A2(n_424),
.B1(n_384),
.B2(n_381),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_451),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_494),
.B(n_497),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_461),
.B(n_458),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_495),
.Y(n_533)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_436),
.Y(n_496)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_496),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_461),
.B(n_396),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_436),
.Y(n_498)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_498),
.Y(n_546)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_455),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_500),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_443),
.A2(n_378),
.B(n_370),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_432),
.B(n_405),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_503),
.B(n_506),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_442),
.B(n_370),
.C(n_358),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_455),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_505),
.B(n_509),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_432),
.B(n_334),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_444),
.A2(n_339),
.B1(n_362),
.B2(n_406),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_521),
.B(n_537),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_523),
.A2(n_531),
.B1(n_539),
.B2(n_541),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_486),
.A2(n_441),
.B(n_431),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_524),
.A2(n_484),
.B(n_502),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_492),
.B(n_447),
.C(n_439),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_527),
.B(n_532),
.C(n_542),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_472),
.A2(n_460),
.B1(n_444),
.B2(n_459),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_528),
.A2(n_536),
.B1(n_489),
.B2(n_501),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_491),
.A2(n_429),
.B1(n_433),
.B2(n_438),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_529),
.B(n_544),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_504),
.B(n_479),
.C(n_447),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_488),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_535),
.B(n_538),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_472),
.A2(n_459),
.B1(n_435),
.B2(n_454),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_485),
.B(n_468),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_476),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_475),
.A2(n_457),
.B1(n_435),
.B2(n_466),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_482),
.B(n_445),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_540),
.B(n_543),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_495),
.A2(n_457),
.B1(n_446),
.B2(n_449),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_483),
.B(n_439),
.C(n_445),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_471),
.B(n_453),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_501),
.A2(n_470),
.B1(n_431),
.B2(n_469),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_544),
.A2(n_545),
.B1(n_478),
.B2(n_477),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_474),
.A2(n_463),
.B1(n_450),
.B2(n_430),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_516),
.Y(n_547)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_547),
.Y(n_582)
);

CKINVDCx16_ASAP7_75t_R g548 ( 
.A(n_516),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_548),
.B(n_560),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_525),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_549),
.B(n_552),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_534),
.B(n_487),
.Y(n_550)
);

NAND3xp33_ASAP7_75t_L g594 ( 
.A(n_550),
.B(n_566),
.C(n_496),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_527),
.B(n_471),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_551),
.B(n_563),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_525),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_511),
.Y(n_556)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_556),
.Y(n_597)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_513),
.Y(n_557)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_557),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_519),
.B(n_453),
.C(n_481),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_558),
.B(n_565),
.C(n_572),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_559),
.A2(n_570),
.B1(n_529),
.B2(n_516),
.Y(n_580)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_510),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_510),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_561),
.B(n_564),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_L g562 ( 
.A1(n_530),
.A2(n_484),
.B(n_509),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_SL g578 ( 
.A1(n_562),
.A2(n_567),
.B(n_524),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_521),
.B(n_471),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_518),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_519),
.B(n_473),
.C(n_507),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_533),
.B(n_537),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_532),
.B(n_507),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_569),
.B(n_517),
.Y(n_593)
);

BUFx24_ASAP7_75t_SL g571 ( 
.A(n_512),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_SL g581 ( 
.A(n_571),
.B(n_497),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_540),
.B(n_493),
.C(n_499),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_542),
.B(n_543),
.C(n_514),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_573),
.B(n_494),
.C(n_514),
.Y(n_588)
);

INVxp33_ASAP7_75t_SL g574 ( 
.A(n_515),
.Y(n_574)
);

INVxp33_ASAP7_75t_L g590 ( 
.A(n_574),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_575),
.A2(n_528),
.B1(n_536),
.B2(n_520),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_523),
.A2(n_506),
.B1(n_480),
.B2(n_503),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_577),
.Y(n_598)
);

XOR2xp5_ASAP7_75t_L g606 ( 
.A(n_578),
.B(n_593),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_580),
.A2(n_594),
.B1(n_596),
.B2(n_602),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_581),
.B(n_595),
.Y(n_617)
);

XNOR2xp5_ASAP7_75t_SL g586 ( 
.A(n_568),
.B(n_530),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g605 ( 
.A(n_586),
.B(n_601),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_588),
.B(n_589),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_554),
.B(n_512),
.C(n_522),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_549),
.B(n_517),
.Y(n_591)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_591),
.Y(n_603)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_592),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_576),
.B(n_498),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_559),
.A2(n_546),
.B1(n_526),
.B2(n_522),
.Y(n_596)
);

XNOR2x1_ASAP7_75t_L g599 ( 
.A(n_572),
.B(n_470),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g611 ( 
.A(n_599),
.B(n_562),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_558),
.B(n_452),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_555),
.A2(n_508),
.B1(n_546),
.B2(n_526),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_583),
.B(n_554),
.C(n_565),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_604),
.B(n_609),
.C(n_613),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_583),
.B(n_569),
.C(n_568),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_SL g626 ( 
.A(n_607),
.B(n_610),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_590),
.A2(n_570),
.B(n_567),
.Y(n_608)
);

CKINVDCx14_ASAP7_75t_R g632 ( 
.A(n_608),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_589),
.B(n_553),
.C(n_573),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g610 ( 
.A(n_584),
.B(n_553),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_SL g636 ( 
.A(n_611),
.B(n_579),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_593),
.B(n_551),
.C(n_563),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_588),
.B(n_570),
.C(n_547),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_614),
.B(n_616),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_SL g615 ( 
.A1(n_585),
.A2(n_552),
.B1(n_490),
.B2(n_500),
.Y(n_615)
);

INVxp67_ASAP7_75t_SL g635 ( 
.A(n_615),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_584),
.B(n_505),
.C(n_450),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_590),
.B(n_463),
.C(n_339),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_620),
.B(n_621),
.Y(n_634)
);

A2O1A1Ixp33_ASAP7_75t_SL g621 ( 
.A1(n_585),
.A2(n_347),
.B(n_362),
.C(n_591),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g622 ( 
.A(n_598),
.Y(n_622)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_622),
.Y(n_630)
);

XOR2xp5_ASAP7_75t_L g623 ( 
.A(n_613),
.B(n_586),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g650 ( 
.A(n_623),
.Y(n_650)
);

XOR2xp5_ASAP7_75t_L g624 ( 
.A(n_606),
.B(n_599),
.Y(n_624)
);

INVxp67_ASAP7_75t_L g652 ( 
.A(n_624),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_603),
.A2(n_578),
.B(n_582),
.Y(n_625)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_625),
.Y(n_651)
);

XOR2xp5_ASAP7_75t_L g627 ( 
.A(n_606),
.B(n_580),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_627),
.B(n_628),
.Y(n_649)
);

INVx6_ASAP7_75t_L g628 ( 
.A(n_617),
.Y(n_628)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_615),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_631),
.B(n_633),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_622),
.A2(n_596),
.B1(n_592),
.B2(n_602),
.Y(n_633)
);

NOR2xp67_ASAP7_75t_L g641 ( 
.A(n_636),
.B(n_605),
.Y(n_641)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_618),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_638),
.B(n_639),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_621),
.B(n_600),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_641),
.A2(n_624),
.B(n_627),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_637),
.B(n_612),
.C(n_604),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_642),
.B(n_643),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_637),
.B(n_609),
.C(n_619),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_SL g645 ( 
.A(n_629),
.B(n_597),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_645),
.B(n_646),
.Y(n_657)
);

MAJIxp5_ASAP7_75t_L g646 ( 
.A(n_635),
.B(n_611),
.C(n_621),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_626),
.B(n_628),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_SL g661 ( 
.A(n_647),
.B(n_587),
.Y(n_661)
);

CKINVDCx16_ASAP7_75t_R g648 ( 
.A(n_625),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_648),
.A2(n_632),
.B1(n_630),
.B2(n_639),
.Y(n_653)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_653),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_643),
.B(n_650),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_654),
.B(n_658),
.Y(n_662)
);

OAI21xp5_ASAP7_75t_L g655 ( 
.A1(n_651),
.A2(n_623),
.B(n_634),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_655),
.A2(n_659),
.B(n_661),
.Y(n_667)
);

MAJIxp5_ASAP7_75t_L g658 ( 
.A(n_642),
.B(n_636),
.C(n_633),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g660 ( 
.A(n_649),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_660),
.A2(n_650),
.B1(n_652),
.B2(n_640),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_663),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_656),
.B(n_644),
.Y(n_665)
);

MAJIxp5_ASAP7_75t_L g669 ( 
.A(n_665),
.B(n_662),
.C(n_667),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_SL g666 ( 
.A1(n_657),
.A2(n_652),
.B(n_634),
.Y(n_666)
);

AOI21x1_ASAP7_75t_SL g668 ( 
.A1(n_666),
.A2(n_654),
.B(n_621),
.Y(n_668)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_668),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g672 ( 
.A(n_669),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_672),
.A2(n_670),
.B(n_664),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_L g674 ( 
.A1(n_673),
.A2(n_671),
.B(n_663),
.Y(n_674)
);

XOR2xp5_ASAP7_75t_L g675 ( 
.A(n_674),
.B(n_646),
.Y(n_675)
);


endmodule