module fake_jpeg_2208_n_147 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_147);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_147;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_12),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_34),
.Y(n_58)
);

NAND2xp33_ASAP7_75t_SL g34 ( 
.A(n_23),
.B(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_14),
.Y(n_40)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_43),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_15),
.B(n_0),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_23),
.B1(n_43),
.B2(n_28),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_51),
.B1(n_56),
.B2(n_19),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_17),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_49),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_43),
.B(n_17),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_30),
.B1(n_29),
.B2(n_28),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_35),
.B(n_25),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_30),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_23),
.B1(n_16),
.B2(n_21),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_16),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_24),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_0),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_24),
.B(n_18),
.C(n_29),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_49),
.B(n_42),
.C(n_26),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_61),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_64),
.B(n_75),
.Y(n_97)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_66),
.A2(n_79),
.B(n_80),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_21),
.B1(n_19),
.B2(n_26),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_50),
.B1(n_47),
.B2(n_46),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_68),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_95)
);

NOR2x1_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_15),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_70),
.B(n_74),
.Y(n_85)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_15),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_54),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_52),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_62),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_15),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_81),
.A2(n_1),
.B(n_2),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_48),
.C(n_59),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

OAI32xp33_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_69),
.A3(n_81),
.B1(n_70),
.B2(n_80),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_89),
.Y(n_107)
);

OAI22x1_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_52),
.B1(n_53),
.B2(n_46),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_95),
.B1(n_90),
.B2(n_77),
.Y(n_105)
);

NOR4xp25_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_91),
.C(n_93),
.D(n_2),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_79),
.A2(n_53),
.B1(n_52),
.B2(n_47),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_73),
.B1(n_91),
.B2(n_72),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_63),
.A2(n_60),
.B(n_20),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_65),
.A2(n_76),
.B1(n_71),
.B2(n_78),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_82),
.B1(n_83),
.B2(n_97),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_101),
.Y(n_111)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_100),
.Y(n_116)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_84),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_103),
.Y(n_112)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_84),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_105),
.Y(n_119)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_108),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_109),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_88),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_118),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_107),
.A2(n_87),
.B(n_85),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_86),
.C(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

AOI31xp67_ASAP7_75t_L g122 ( 
.A1(n_118),
.A2(n_85),
.A3(n_107),
.B(n_103),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_122),
.A2(n_111),
.B1(n_120),
.B2(n_116),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_99),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_126),
.C(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_124),
.A2(n_127),
.B1(n_116),
.B2(n_101),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_100),
.B(n_106),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_113),
.C(n_115),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_132),
.Y(n_137)
);

AOI31xp67_ASAP7_75t_L g138 ( 
.A1(n_133),
.A2(n_134),
.A3(n_125),
.B(n_20),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_128),
.B(n_116),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_130),
.A2(n_125),
.B1(n_9),
.B2(n_12),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_131),
.C(n_9),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_134),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_140),
.Y(n_142)
);

AO22x1_ASAP7_75t_L g141 ( 
.A1(n_136),
.A2(n_60),
.B1(n_4),
.B2(n_5),
.Y(n_141)
);

OAI221xp5_ASAP7_75t_L g143 ( 
.A1(n_141),
.A2(n_138),
.B1(n_137),
.B2(n_6),
.C(n_4),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_143),
.B(n_141),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_142),
.B(n_139),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_3),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_60),
.Y(n_147)
);


endmodule