module fake_jpeg_5964_n_18 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_18);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_18;

wire n_13;
wire n_14;
wire n_11;
wire n_17;
wire n_16;
wire n_12;
wire n_15;

INVx2_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

AND2x2_ASAP7_75t_L g12 ( 
.A(n_2),
.B(n_6),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_0),
.A2(n_4),
.B1(n_1),
.B2(n_7),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_8),
.B(n_3),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_14),
.A2(n_9),
.B1(n_10),
.B2(n_0),
.Y(n_15)
);

MAJx2_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_16),
.C(n_12),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_14),
.A2(n_1),
.B1(n_11),
.B2(n_13),
.Y(n_16)
);

HB1xp67_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);


endmodule