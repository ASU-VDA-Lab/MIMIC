module fake_jpeg_29533_n_200 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_200);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_200;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_35),
.B(n_37),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_1),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_18),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_22),
.Y(n_55)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_29),
.B1(n_19),
.B2(n_16),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_49),
.A2(n_63),
.B1(n_38),
.B2(n_44),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_31),
.C(n_23),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_51),
.B(n_65),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_27),
.B1(n_31),
.B2(n_23),
.Y(n_51)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_43),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_54),
.B(n_55),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_29),
.B1(n_19),
.B2(n_16),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_58),
.A2(n_34),
.B1(n_40),
.B2(n_45),
.Y(n_75)
);

CKINVDCx9p33_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_27),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_17),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_29),
.B1(n_21),
.B2(n_26),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_34),
.A2(n_21),
.B1(n_28),
.B2(n_26),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_66),
.B(n_30),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_70),
.B(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_39),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_37),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_30),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_87),
.Y(n_97)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_75),
.A2(n_63),
.B1(n_38),
.B2(n_44),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_17),
.B(n_33),
.C(n_28),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_78),
.B(n_24),
.Y(n_100)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_90),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_59),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_89),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_55),
.Y(n_87)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_92),
.Y(n_104)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_38),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_92),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_65),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_95),
.A2(n_46),
.B1(n_54),
.B2(n_56),
.Y(n_123)
);

OAI32xp33_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_38),
.A3(n_33),
.B1(n_24),
.B2(n_52),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_110),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_100),
.B(n_103),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_83),
.B(n_90),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_46),
.C(n_47),
.Y(n_103)
);

BUFx4f_ASAP7_75t_SL g106 ( 
.A(n_69),
.Y(n_106)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_14),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_107),
.B(n_108),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_79),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_14),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_76),
.B(n_86),
.Y(n_114)
);

AOI21xp33_ASAP7_75t_L g117 ( 
.A1(n_114),
.A2(n_68),
.B(n_67),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_109),
.A2(n_75),
.B1(n_89),
.B2(n_81),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_115),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_117),
.B(n_119),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_99),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_109),
.A2(n_47),
.B1(n_56),
.B2(n_80),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_127),
.Y(n_136)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_123),
.A2(n_131),
.B1(n_133),
.B2(n_94),
.Y(n_135)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_126),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_101),
.A2(n_57),
.B1(n_40),
.B2(n_74),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_96),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_95),
.A2(n_57),
.B1(n_88),
.B2(n_69),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_114),
.A2(n_85),
.B1(n_84),
.B2(n_77),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_143),
.B1(n_127),
.B2(n_132),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_129),
.A2(n_103),
.B(n_108),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_138),
.A2(n_116),
.B(n_100),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_120),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_123),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_130),
.A2(n_93),
.B1(n_98),
.B2(n_97),
.Y(n_143)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_151),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_121),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_124),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_153),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_128),
.C(n_134),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_164),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_142),
.B(n_143),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_159),
.Y(n_166)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_139),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_141),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_112),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_161),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_112),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_137),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_163),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_147),
.Y(n_163)
);

OAI322xp33_ASAP7_75t_L g164 ( 
.A1(n_136),
.A2(n_131),
.A3(n_125),
.B1(n_118),
.B2(n_126),
.C1(n_106),
.C2(n_94),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_157),
.A2(n_139),
.B1(n_135),
.B2(n_136),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_167),
.A2(n_169),
.B1(n_170),
.B2(n_152),
.Y(n_176)
);

AOI221xp5_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_148),
.B1(n_146),
.B2(n_145),
.C(n_105),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_154),
.A2(n_118),
.B(n_113),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_172),
.A2(n_1),
.B(n_2),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_158),
.B(n_153),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_168),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_176),
.B(n_177),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_105),
.C(n_106),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_178),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_184)
);

NOR3xp33_ASAP7_75t_SL g179 ( 
.A(n_166),
.B(n_7),
.C(n_15),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_13),
.Y(n_180)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_180),
.Y(n_185)
);

OAI21x1_ASAP7_75t_L g181 ( 
.A1(n_171),
.A2(n_168),
.B(n_172),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_183),
.A2(n_177),
.B(n_10),
.Y(n_189)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_179),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_188),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_165),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_191),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_10),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_184),
.A2(n_187),
.B(n_183),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_192),
.A2(n_188),
.B1(n_185),
.B2(n_8),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_193),
.A2(n_194),
.B1(n_4),
.B2(n_6),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_1),
.C(n_2),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_195),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_196),
.A2(n_197),
.B1(n_6),
.B2(n_3),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_198),
.A2(n_3),
.B(n_6),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_43),
.Y(n_200)
);


endmodule