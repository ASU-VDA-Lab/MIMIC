module fake_jpeg_14958_n_121 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_121);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_27),
.Y(n_38)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_12),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_24),
.Y(n_37)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_18),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_21),
.B1(n_12),
.B2(n_19),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_41),
.B1(n_33),
.B2(n_15),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_37),
.B(n_11),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_26),
.A2(n_17),
.B1(n_23),
.B2(n_15),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_22),
.B1(n_20),
.B2(n_13),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_17),
.B1(n_23),
.B2(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_44),
.Y(n_65)
);

NOR2x1_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_45),
.B(n_56),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_42),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_57),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_16),
.B1(n_22),
.B2(n_20),
.Y(n_47)
);

NOR3xp33_ASAP7_75t_SL g74 ( 
.A(n_47),
.B(n_45),
.C(n_41),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_24),
.B(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_53),
.Y(n_67)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_43),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_55),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_28),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_13),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_59),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_27),
.C(n_31),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_62),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_63),
.B(n_35),
.Y(n_76)
);

NOR4xp25_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_48),
.C(n_46),
.D(n_57),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_77),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_80),
.B(n_84),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_72),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_86),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_64),
.Y(n_93)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_55),
.B(n_50),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_72),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_60),
.B1(n_50),
.B2(n_51),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_87),
.A2(n_89),
.B1(n_68),
.B2(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_52),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_75),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_58),
.B1(n_61),
.B2(n_0),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_71),
.C(n_69),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_71),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_97),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_91),
.B1(n_85),
.B2(n_79),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_64),
.Y(n_97)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

AO21x1_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_74),
.B(n_66),
.Y(n_100)
);

NOR3xp33_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_75),
.C(n_13),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_87),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_103),
.A2(n_96),
.B1(n_94),
.B2(n_79),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_100),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_102),
.A2(n_89),
.B1(n_66),
.B2(n_92),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_107),
.A2(n_99),
.B1(n_83),
.B2(n_73),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_108),
.B(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_111),
.C(n_104),
.Y(n_113)
);

XOR2x2_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_3),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_112),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_113),
.B(n_114),
.Y(n_116)
);

A2O1A1O1Ixp25_ASAP7_75t_L g117 ( 
.A1(n_115),
.A2(n_112),
.B(n_109),
.C(n_108),
.D(n_8),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_117),
.A2(n_5),
.B(n_6),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_119),
.A2(n_116),
.B(n_3),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_120),
.B(n_3),
.Y(n_121)
);


endmodule