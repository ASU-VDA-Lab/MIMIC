module fake_ariane_1165_n_119 (n_8, n_7, n_22, n_1, n_6, n_13, n_20, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_10, n_119);

input n_8;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_10;

output n_119;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_106;
wire n_53;
wire n_111;
wire n_115;
wire n_66;
wire n_71;
wire n_24;
wire n_109;
wire n_96;
wire n_49;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_107;
wire n_72;
wire n_105;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_117;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_112;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_118;
wire n_93;
wire n_23;
wire n_61;
wire n_108;
wire n_102;
wire n_43;
wire n_87;
wire n_81;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_116;
wire n_104;
wire n_78;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_35;
wire n_54;
wire n_25;

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_15),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_21),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVxp33_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_0),
.Y(n_43)
);

AND2x4_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_1),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_1),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_6),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_7),
.Y(n_47)
);

NAND2x1p5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_27),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_8),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_36),
.B(n_17),
.Y(n_52)
);

OR2x6_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_8),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_50),
.B(n_34),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_50),
.B(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_54),
.B(n_29),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_54),
.B(n_40),
.Y(n_59)
);

NAND2xp33_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_54),
.B(n_28),
.Y(n_61)
);

NAND2xp33_ASAP7_75t_SL g62 ( 
.A(n_44),
.B(n_23),
.Y(n_62)
);

NAND2xp33_ASAP7_75t_SL g63 ( 
.A(n_44),
.B(n_30),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_52),
.B(n_32),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_38),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_42),
.B(n_39),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_42),
.B(n_39),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

AO21x2_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_51),
.B(n_45),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_48),
.B(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_48),
.Y(n_72)
);

AO31x2_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_47),
.A3(n_43),
.B(n_55),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_62),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

OAI211xp5_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_49),
.B(n_53),
.C(n_48),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_53),
.B1(n_10),
.B2(n_9),
.Y(n_77)
);

OAI21x1_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_53),
.B(n_18),
.Y(n_78)
);

OAI21x1_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_53),
.B(n_19),
.Y(n_79)
);

CKINVDCx11_ASAP7_75t_R g80 ( 
.A(n_74),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_9),
.Y(n_82)
);

AND2x4_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_74),
.Y(n_83)
);

OR2x6_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_76),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_R g85 ( 
.A(n_75),
.B(n_72),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_72),
.Y(n_87)
);

AND2x4_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_68),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_69),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_78),
.Y(n_90)
);

NAND2xp33_ASAP7_75t_SL g91 ( 
.A(n_69),
.B(n_71),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_73),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

AOI211xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_78),
.B(n_79),
.C(n_73),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_91),
.C(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

NOR2x1_ASAP7_75t_SL g99 ( 
.A(n_84),
.B(n_69),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_73),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

AOI322xp5_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_70),
.A3(n_73),
.B1(n_78),
.B2(n_79),
.C1(n_87),
.C2(n_80),
.Y(n_102)
);

NOR4xp25_ASAP7_75t_SL g103 ( 
.A(n_98),
.B(n_84),
.C(n_85),
.D(n_79),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_97),
.A2(n_84),
.B1(n_70),
.B2(n_81),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_70),
.B1(n_81),
.B2(n_85),
.Y(n_105)
);

AO221x2_ASAP7_75t_L g106 ( 
.A1(n_102),
.A2(n_73),
.B1(n_98),
.B2(n_96),
.C(n_99),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_SL g107 ( 
.A1(n_104),
.A2(n_95),
.B(n_92),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_106),
.A2(n_92),
.B1(n_100),
.B2(n_95),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_100),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

NAND3xp33_ASAP7_75t_SL g111 ( 
.A(n_110),
.B(n_102),
.C(n_103),
.Y(n_111)
);

OAI211xp5_ASAP7_75t_L g112 ( 
.A1(n_109),
.A2(n_96),
.B(n_93),
.C(n_94),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_R g113 ( 
.A(n_111),
.B(n_93),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_R g114 ( 
.A(n_112),
.B(n_93),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g116 ( 
.A1(n_114),
.A2(n_100),
.B(n_92),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_106),
.B1(n_101),
.B2(n_105),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_117),
.A2(n_115),
.B(n_99),
.Y(n_118)
);

OAI221xp5_ASAP7_75t_R g119 ( 
.A1(n_118),
.A2(n_73),
.B1(n_94),
.B2(n_101),
.C(n_117),
.Y(n_119)
);


endmodule