module fake_jpeg_22283_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_33),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_15),
.B1(n_16),
.B2(n_30),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_42),
.A2(n_27),
.B1(n_19),
.B2(n_20),
.Y(n_74)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_48),
.Y(n_69)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_51),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_34),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_16),
.B1(n_15),
.B2(n_30),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_20),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_18),
.Y(n_75)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_27),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_58),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_65),
.B1(n_73),
.B2(n_74),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_54),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_20),
.B1(n_30),
.B2(n_27),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_75),
.B(n_81),
.Y(n_98)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_82),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_28),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_28),
.Y(n_110)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_0),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_85),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_44),
.B(n_25),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_47),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_90),
.Y(n_118)
);

NOR3xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_19),
.C(n_18),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_92),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_62),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_71),
.A2(n_45),
.B1(n_60),
.B2(n_56),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_94),
.B1(n_103),
.B2(n_65),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_71),
.A2(n_60),
.B1(n_56),
.B2(n_48),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_69),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_96),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_99),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_75),
.B(n_18),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_67),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_102),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_67),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_49),
.B1(n_57),
.B2(n_53),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_84),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_109),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_46),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_66),
.C(n_24),
.Y(n_124)
);

AO21x2_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_86),
.B(n_55),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_111),
.A2(n_117),
.B1(n_128),
.B2(n_130),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_61),
.B1(n_80),
.B2(n_78),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_112),
.A2(n_114),
.B1(n_120),
.B2(n_127),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_113),
.B(n_115),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_80),
.B1(n_78),
.B2(n_77),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_64),
.B1(n_70),
.B2(n_72),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_87),
.A2(n_70),
.B1(n_76),
.B2(n_41),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_134),
.C(n_129),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_107),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_126),
.A2(n_108),
.B1(n_105),
.B2(n_101),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_66),
.B1(n_55),
.B2(n_86),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_91),
.A2(n_94),
.B1(n_93),
.B2(n_87),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_24),
.B(n_25),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_89),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_110),
.A2(n_29),
.B1(n_26),
.B2(n_25),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_135),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_110),
.A2(n_29),
.B1(n_26),
.B2(n_25),
.Y(n_132)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

AND2x2_ASAP7_75t_SL g134 ( 
.A(n_95),
.B(n_43),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_137),
.Y(n_169)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_125),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_138),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_98),
.Y(n_141)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_98),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_143),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_125),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_145),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_99),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_146),
.B(n_152),
.Y(n_162)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_150),
.Y(n_176)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_114),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_108),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_108),
.Y(n_153)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_157),
.Y(n_171)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_156),
.B(n_159),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_132),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_158),
.B(n_130),
.Y(n_164)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_116),
.Y(n_179)
);

NAND3xp33_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_115),
.C(n_134),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_175),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_142),
.C(n_146),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_154),
.B(n_150),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_165),
.A2(n_119),
.B(n_104),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_152),
.B(n_128),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_23),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_111),
.Y(n_174)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_151),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_181),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_144),
.A2(n_155),
.B1(n_148),
.B2(n_135),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_178),
.A2(n_182),
.B1(n_184),
.B2(n_134),
.Y(n_193)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_151),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_144),
.A2(n_111),
.B1(n_122),
.B2(n_126),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_149),
.Y(n_183)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_148),
.A2(n_111),
.B1(n_157),
.B2(n_149),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_136),
.A2(n_113),
.B1(n_117),
.B2(n_111),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_185),
.A2(n_86),
.B1(n_100),
.B2(n_29),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_173),
.B(n_158),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_188),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_169),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_187),
.B(n_201),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_164),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_168),
.B(n_143),
.Y(n_189)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_207),
.C(n_179),
.Y(n_220)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_206),
.Y(n_213)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_183),
.A2(n_111),
.B1(n_134),
.B2(n_102),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_191),
.A2(n_205),
.B1(n_172),
.B2(n_178),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_193),
.A2(n_202),
.B1(n_185),
.B2(n_180),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_196),
.Y(n_221)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_199),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_176),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_171),
.B(n_105),
.C(n_119),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_171),
.C(n_175),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_182),
.A2(n_28),
.B1(n_23),
.B2(n_29),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_100),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_100),
.Y(n_226)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_168),
.B(n_23),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_218),
.C(n_222),
.Y(n_232)
);

BUFx24_ASAP7_75t_SL g210 ( 
.A(n_203),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_223),
.Y(n_233)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_205),
.A2(n_180),
.B1(n_184),
.B2(n_163),
.Y(n_214)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_214),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_215),
.A2(n_217),
.B1(n_192),
.B2(n_195),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_195),
.A2(n_166),
.B1(n_170),
.B2(n_172),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_167),
.C(n_165),
.Y(n_218)
);

XOR2x2_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_167),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_219),
.B(n_220),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_100),
.C(n_26),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_201),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_224),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_227),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_188),
.B(n_28),
.Y(n_227)
);

XNOR2x2_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_26),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_228),
.B(n_191),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_204),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_235),
.Y(n_256)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_234),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_207),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_225),
.B(n_197),
.Y(n_237)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_237),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_194),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_244),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_228),
.Y(n_239)
);

OAI21xp33_ASAP7_75t_SL g250 ( 
.A1(n_239),
.A2(n_241),
.B(n_243),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_212),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_191),
.C(n_1),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_0),
.C(n_2),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_236),
.A2(n_213),
.B1(n_218),
.B2(n_220),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_247),
.A2(n_251),
.B1(n_253),
.B2(n_254),
.Y(n_262)
);

INVxp33_ASAP7_75t_L g248 ( 
.A(n_242),
.Y(n_248)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_230),
.A2(n_222),
.B1(n_216),
.B2(n_14),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_216),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_257),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_253),
.B(n_2),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_14),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_258),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_229),
.C(n_240),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_12),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_242),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_259),
.A2(n_244),
.B1(n_243),
.B2(n_232),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_264),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_249),
.A2(n_255),
.B1(n_246),
.B2(n_250),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_262),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_248),
.A2(n_233),
.B1(n_3),
.B2(n_4),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_13),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_267),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_257),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_271),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_5),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_10),
.Y(n_271)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_272),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_263),
.A2(n_256),
.B(n_11),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_277),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_270),
.A2(n_11),
.B(n_10),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_268),
.A2(n_5),
.B(n_6),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_279),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_262),
.A2(n_5),
.B(n_6),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_5),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_6),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_272),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_281),
.Y(n_285)
);

XNOR2x1_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_287),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_265),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_286),
.A2(n_7),
.B(n_8),
.Y(n_293)
);

NAND2x1p5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_265),
.Y(n_287)
);

AO21x1_ASAP7_75t_L g294 ( 
.A1(n_289),
.A2(n_282),
.B(n_8),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_288),
.A2(n_275),
.B(n_8),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_290),
.A2(n_292),
.B(n_293),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_283),
.B(n_9),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_291),
.C(n_8),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_295),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_297),
.A2(n_7),
.B(n_9),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_298),
.B(n_7),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_9),
.Y(n_300)
);


endmodule