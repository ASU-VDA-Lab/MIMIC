module fake_jpeg_10505_n_109 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_109);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_109;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx6_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx4f_ASAP7_75t_SL g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_21),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_22),
.B(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_28),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g27 ( 
.A(n_12),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_15),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_10),
.B(n_19),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_11),
.B1(n_20),
.B2(n_14),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_31),
.A2(n_38),
.B1(n_29),
.B2(n_14),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g48 ( 
.A1(n_32),
.A2(n_27),
.B(n_3),
.Y(n_48)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_19),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_27),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_25),
.A2(n_11),
.B1(n_10),
.B2(n_16),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_36),
.B(n_22),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_23),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_48),
.B(n_31),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_42),
.B(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_28),
.Y(n_43)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_16),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_46),
.Y(n_61)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_28),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_30),
.B(n_38),
.Y(n_50)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_29),
.Y(n_52)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_20),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_55),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_13),
.B1(n_4),
.B2(n_5),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_2),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_58),
.B(n_65),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_37),
.B(n_31),
.Y(n_58)
);

OAI32xp33_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_17),
.A3(n_26),
.B1(n_13),
.B2(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_26),
.B(n_4),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_26),
.B(n_4),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_2),
.C(n_6),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_8),
.B1(n_7),
.B2(n_2),
.Y(n_81)
);

AOI22x1_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_41),
.B1(n_54),
.B2(n_51),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_79),
.B1(n_81),
.B2(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_74),
.Y(n_83)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_41),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_76),
.Y(n_82)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_53),
.B(n_5),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_80),
.B(n_57),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_46),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_65),
.C(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_84),
.A2(n_85),
.B(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_88),
.Y(n_90)
);

NAND3xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_64),
.C(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_87),
.B(n_89),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_80),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_SL g91 ( 
.A1(n_86),
.A2(n_71),
.B(n_73),
.C(n_66),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_94),
.B1(n_69),
.B2(n_82),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_82),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_88),
.A2(n_75),
.B1(n_56),
.B2(n_66),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_96),
.A2(n_94),
.B(n_91),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_99),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_95),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_78),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_101),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_91),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_102),
.A2(n_69),
.B(n_103),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_99),
.B(n_91),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_105),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_106),
.Y(n_109)
);


endmodule