module fake_netlist_1_9261_n_38 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_38);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
AND2x4_ASAP7_75t_L g12 ( .A(n_10), .B(n_4), .Y(n_12) );
CKINVDCx16_ASAP7_75t_R g13 ( .A(n_8), .Y(n_13) );
BUFx6f_ASAP7_75t_L g14 ( .A(n_3), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_7), .Y(n_15) );
XNOR2x1_ASAP7_75t_L g16 ( .A(n_1), .B(n_3), .Y(n_16) );
NAND2x1p5_ASAP7_75t_L g17 ( .A(n_8), .B(n_9), .Y(n_17) );
BUFx3_ASAP7_75t_L g18 ( .A(n_12), .Y(n_18) );
AOI22xp33_ASAP7_75t_L g19 ( .A1(n_12), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_19) );
INVx3_ASAP7_75t_L g20 ( .A(n_12), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
CKINVDCx11_ASAP7_75t_R g22 ( .A(n_18), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_22), .B(n_13), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_21), .B(n_18), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_23), .B(n_13), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_24), .B(n_21), .Y(n_26) );
AOI221xp5_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_23), .B1(n_19), .B2(n_20), .C(n_18), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_26), .Y(n_28) );
OAI211xp5_ASAP7_75t_L g29 ( .A1(n_27), .A2(n_15), .B(n_20), .C(n_14), .Y(n_29) );
AOI21xp33_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_20), .B(n_16), .Y(n_30) );
OAI22xp5_ASAP7_75t_L g31 ( .A1(n_28), .A2(n_16), .B1(n_17), .B2(n_15), .Y(n_31) );
AOI21xp5_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_17), .B(n_14), .Y(n_32) );
AOI22xp5_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_17), .B1(n_14), .B2(n_4), .Y(n_33) );
OAI22xp5_ASAP7_75t_L g34 ( .A1(n_30), .A2(n_14), .B1(n_2), .B2(n_5), .Y(n_34) );
OAI21x1_ASAP7_75t_SL g35 ( .A1(n_33), .A2(n_0), .B(n_5), .Y(n_35) );
HB1xp67_ASAP7_75t_L g36 ( .A(n_34), .Y(n_36) );
AOI22xp5_ASAP7_75t_L g37 ( .A1(n_36), .A2(n_32), .B1(n_14), .B2(n_7), .Y(n_37) );
AOI22xp5_ASAP7_75t_SL g38 ( .A1(n_37), .A2(n_35), .B1(n_6), .B2(n_11), .Y(n_38) );
endmodule