module fake_jpeg_30726_n_502 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_502);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_502;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_7),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_49),
.B(n_35),
.Y(n_103)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_51),
.B(n_53),
.Y(n_135)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_58),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_59),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_7),
.B1(n_13),
.B2(n_10),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_60),
.A2(n_22),
.B1(n_39),
.B2(n_33),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_30),
.B(n_42),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g143 ( 
.A(n_63),
.B(n_20),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_70),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g119 ( 
.A(n_71),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g147 ( 
.A(n_72),
.Y(n_147)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_30),
.B(n_8),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_76),
.B(n_81),
.Y(n_138)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_35),
.B(n_8),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_15),
.Y(n_87)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_15),
.Y(n_89)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

INVx5_ASAP7_75t_SL g90 ( 
.A(n_47),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_90),
.B(n_43),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_92),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

NAND2xp33_ASAP7_75t_SL g96 ( 
.A(n_18),
.B(n_8),
.Y(n_96)
);

NAND2xp33_ASAP7_75t_SL g132 ( 
.A(n_96),
.B(n_43),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_103),
.B(n_109),
.Y(n_160)
);

HAxp5_ASAP7_75t_SL g108 ( 
.A(n_51),
.B(n_22),
.CON(n_108),
.SN(n_108)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_108),
.B(n_21),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_49),
.B(n_42),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_56),
.A2(n_34),
.B1(n_31),
.B2(n_18),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_111),
.A2(n_117),
.B1(n_140),
.B2(n_152),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_81),
.A2(n_18),
.B1(n_34),
.B2(n_31),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_123),
.A2(n_24),
.B1(n_39),
.B2(n_21),
.Y(n_183)
);

OA22x2_ASAP7_75t_L g125 ( 
.A1(n_53),
.A2(n_29),
.B1(n_38),
.B2(n_20),
.Y(n_125)
);

OA22x2_ASAP7_75t_SL g188 ( 
.A1(n_125),
.A2(n_24),
.B1(n_32),
.B2(n_92),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_149),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_78),
.B(n_33),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_145),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_48),
.A2(n_34),
.B1(n_29),
.B2(n_28),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_26),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_92),
.B(n_26),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_90),
.A2(n_43),
.B1(n_28),
.B2(n_34),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_153),
.B(n_180),
.Y(n_215)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_148),
.Y(n_154)
);

INVx3_ASAP7_75t_SL g204 ( 
.A(n_154),
.Y(n_204)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_156),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_108),
.A2(n_16),
.B1(n_25),
.B2(n_38),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_157),
.Y(n_233)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_158),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_159),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_25),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_162),
.B(n_167),
.Y(n_220)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_113),
.Y(n_163)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_163),
.Y(n_232)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_114),
.Y(n_164)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_164),
.Y(n_237)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_165),
.Y(n_234)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

INVx3_ASAP7_75t_SL g208 ( 
.A(n_166),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_122),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_16),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_168),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_118),
.Y(n_169)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_169),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_135),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_170),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_125),
.A2(n_61),
.B1(n_70),
.B2(n_66),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_171),
.A2(n_173),
.B1(n_194),
.B2(n_119),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_125),
.A2(n_58),
.B1(n_64),
.B2(n_95),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_106),
.A2(n_93),
.B1(n_59),
.B2(n_77),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_174),
.A2(n_183),
.B1(n_147),
.B2(n_119),
.Y(n_206)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_102),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_175),
.Y(n_223)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_120),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_128),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_177),
.Y(n_231)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_100),
.Y(n_178)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_178),
.Y(n_227)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_107),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_179),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_118),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g182 ( 
.A1(n_152),
.A2(n_67),
.B1(n_69),
.B2(n_29),
.Y(n_182)
);

AO22x1_ASAP7_75t_L g222 ( 
.A1(n_182),
.A2(n_188),
.B1(n_189),
.B2(n_140),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_100),
.Y(n_184)
);

INVx3_ASAP7_75t_SL g209 ( 
.A(n_184),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_104),
.Y(n_185)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_101),
.Y(n_186)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_186),
.Y(n_229)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_110),
.B(n_27),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_193),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_141),
.Y(n_191)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_191),
.Y(n_235)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_104),
.Y(n_192)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_192),
.Y(n_238)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_115),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_L g194 ( 
.A1(n_97),
.A2(n_94),
.B1(n_91),
.B2(n_88),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_126),
.B(n_59),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_195),
.B(n_121),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_130),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_197),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_134),
.B(n_32),
.Y(n_197)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_150),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_199),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_124),
.Y(n_199)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_146),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_201),
.Y(n_213)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_116),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_206),
.A2(n_239),
.B1(n_194),
.B2(n_147),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_214),
.A2(n_98),
.B1(n_105),
.B2(n_139),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_160),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_137),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_225),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_222),
.B(n_183),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_155),
.B(n_129),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_155),
.B(n_144),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_226),
.B(n_236),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_161),
.B(n_133),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_181),
.A2(n_139),
.B1(n_105),
.B2(n_98),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_SL g241 ( 
.A(n_222),
.B(n_189),
.C(n_188),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_241),
.Y(n_296)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_242),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_222),
.A2(n_188),
.B(n_182),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_243),
.A2(n_275),
.B(n_234),
.Y(n_289)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_244),
.Y(n_286)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_246),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_248),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_238),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_249),
.A2(n_255),
.B1(n_264),
.B2(n_266),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_233),
.A2(n_182),
.B1(n_157),
.B2(n_106),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_250),
.Y(n_281)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_213),
.Y(n_251)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_251),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_252),
.A2(n_261),
.B1(n_227),
.B2(n_230),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_240),
.B(n_196),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_253),
.B(n_263),
.Y(n_304)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_254),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_239),
.A2(n_164),
.B1(n_163),
.B2(n_97),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_256),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_174),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_257),
.B(n_272),
.C(n_273),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_206),
.A2(n_187),
.B1(n_179),
.B2(n_165),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_258),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_216),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_265),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_193),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_262),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_240),
.B(n_166),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_214),
.A2(n_220),
.B1(n_215),
.B2(n_205),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_238),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_215),
.A2(n_127),
.B1(n_150),
.B2(n_201),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_217),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_267),
.Y(n_291)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_213),
.Y(n_268)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_268),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_223),
.A2(n_146),
.B1(n_127),
.B2(n_198),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_269),
.A2(n_209),
.B1(n_204),
.B2(n_208),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_205),
.B(n_185),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_271),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_203),
.B(n_199),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_203),
.B(n_169),
.C(n_191),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_219),
.B(n_154),
.C(n_124),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_211),
.A2(n_223),
.B1(n_231),
.B2(n_207),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_274),
.A2(n_276),
.B1(n_209),
.B2(n_208),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_210),
.B(n_112),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_211),
.A2(n_83),
.B1(n_71),
.B2(n_72),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_236),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_283),
.B(n_284),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_251),
.B(n_210),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_231),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_287),
.B(n_290),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_289),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_259),
.B(n_230),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_292),
.A2(n_299),
.B1(n_275),
.B2(n_209),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_207),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_294),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_295),
.A2(n_249),
.B1(n_255),
.B2(n_276),
.Y(n_323)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_254),
.Y(n_297)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_297),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_243),
.A2(n_227),
.B1(n_178),
.B2(n_184),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_259),
.B(n_224),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_306),
.C(n_272),
.Y(n_313)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_271),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_303),
.B(n_308),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_305),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_245),
.B(n_218),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_264),
.B(n_208),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_266),
.Y(n_310)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_310),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_245),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_311),
.B(n_315),
.C(n_316),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_289),
.A2(n_285),
.B(n_281),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_312),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_313),
.B(n_329),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_257),
.C(n_273),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_260),
.C(n_252),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_309),
.A2(n_250),
.B(n_258),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_317),
.Y(n_363)
);

OAI32xp33_ASAP7_75t_L g318 ( 
.A1(n_296),
.A2(n_241),
.A3(n_252),
.B1(n_262),
.B2(n_275),
.Y(n_318)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_318),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_320),
.A2(n_297),
.B1(n_288),
.B2(n_32),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_262),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_322),
.B(n_326),
.C(n_331),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_323),
.A2(n_327),
.B1(n_328),
.B2(n_340),
.Y(n_356)
);

NAND2xp33_ASAP7_75t_SL g324 ( 
.A(n_308),
.B(n_248),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_324),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_306),
.B(n_235),
.C(n_256),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_295),
.A2(n_111),
.B1(n_267),
.B2(n_202),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_310),
.A2(n_202),
.B1(n_229),
.B2(n_234),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_282),
.B(n_221),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_282),
.B(n_217),
.C(n_221),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_299),
.A2(n_204),
.B(n_212),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_332),
.B(n_333),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_294),
.A2(n_204),
.B(n_212),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g335 ( 
.A(n_298),
.B(n_192),
.Y(n_335)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_335),
.Y(n_348)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_278),
.Y(n_336)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_336),
.Y(n_372)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_278),
.Y(n_338)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_338),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_304),
.A2(n_237),
.B(n_232),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_339),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_298),
.A2(n_302),
.B1(n_284),
.B2(n_287),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_302),
.A2(n_86),
.B1(n_74),
.B2(n_237),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_341),
.A2(n_291),
.B1(n_286),
.B2(n_293),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_304),
.A2(n_27),
.B(n_156),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_343),
.B(n_344),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_290),
.B(n_200),
.C(n_27),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_337),
.B(n_283),
.Y(n_345)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_345),
.Y(n_383)
);

BUFx8_ASAP7_75t_L g347 ( 
.A(n_317),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_347),
.Y(n_392)
);

FAx1_ASAP7_75t_SL g350 ( 
.A(n_334),
.B(n_300),
.CI(n_280),
.CON(n_350),
.SN(n_350)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_350),
.B(n_376),
.Y(n_386)
);

XOR2x2_ASAP7_75t_L g351 ( 
.A(n_322),
.B(n_280),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_351),
.B(n_323),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_344),
.B(n_279),
.Y(n_353)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_353),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_335),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_355),
.B(n_360),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_337),
.B(n_279),
.Y(n_357)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_357),
.Y(n_395)
);

OA21x2_ASAP7_75t_L g358 ( 
.A1(n_312),
.A2(n_300),
.B(n_292),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_358),
.A2(n_319),
.B(n_320),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_359),
.A2(n_374),
.B1(n_338),
.B2(n_336),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_316),
.B(n_286),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_325),
.A2(n_293),
.B1(n_291),
.B2(n_277),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_361),
.A2(n_364),
.B1(n_369),
.B2(n_368),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_325),
.A2(n_291),
.B1(n_277),
.B2(n_288),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_343),
.B(n_277),
.Y(n_367)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_367),
.Y(n_403)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_335),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_368),
.B(n_314),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_330),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_311),
.B(n_8),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_375),
.B(n_6),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_334),
.B(n_1),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_377),
.A2(n_385),
.B1(n_356),
.B2(n_347),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_366),
.B(n_315),
.C(n_313),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_378),
.B(n_379),
.C(n_381),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_366),
.B(n_326),
.C(n_331),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_363),
.A2(n_321),
.B(n_342),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_380),
.A2(n_397),
.B(n_400),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_373),
.B(n_329),
.C(n_340),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_373),
.B(n_342),
.C(n_339),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_382),
.B(n_389),
.C(n_399),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_365),
.B(n_318),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_387),
.B(n_390),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_388),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_365),
.B(n_333),
.C(n_330),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_351),
.B(n_324),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_391),
.B(n_393),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_346),
.B(n_332),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_357),
.B(n_328),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_396),
.B(n_358),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_363),
.A2(n_314),
.B(n_341),
.Y(n_397)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_398),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_346),
.B(n_327),
.C(n_32),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_354),
.A2(n_9),
.B(n_14),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_354),
.B(n_32),
.C(n_2),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_401),
.B(n_1),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_402),
.B(n_384),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_356),
.A2(n_370),
.B1(n_371),
.B2(n_359),
.Y(n_404)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_404),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_405),
.B(n_390),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_394),
.B(n_350),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_409),
.B(n_411),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_383),
.B(n_350),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_412),
.B(n_416),
.Y(n_435)
);

O2A1O1Ixp33_ASAP7_75t_L g413 ( 
.A1(n_386),
.A2(n_371),
.B(n_348),
.C(n_349),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_413),
.A2(n_420),
.B(n_427),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_386),
.B(n_345),
.Y(n_416)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_395),
.Y(n_419)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_419),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_R g420 ( 
.A(n_392),
.B(n_348),
.C(n_347),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_381),
.B(n_358),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_421),
.B(n_422),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_389),
.B(n_352),
.Y(n_422)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_423),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_424),
.A2(n_396),
.B1(n_400),
.B2(n_362),
.Y(n_437)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_403),
.Y(n_425)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_425),
.Y(n_441)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_380),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_426),
.B(n_393),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_SL g427 ( 
.A(n_387),
.B(n_361),
.C(n_364),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_417),
.A2(n_377),
.B1(n_385),
.B2(n_399),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_428),
.A2(n_433),
.B1(n_418),
.B2(n_6),
.Y(n_458)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_430),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_406),
.B(n_382),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_432),
.B(n_408),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_427),
.A2(n_392),
.B1(n_397),
.B2(n_391),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_434),
.B(n_436),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_415),
.B(n_378),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_437),
.A2(n_442),
.B1(n_413),
.B2(n_410),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_424),
.A2(n_362),
.B1(n_372),
.B2(n_379),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_415),
.B(n_376),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_443),
.B(n_444),
.C(n_445),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_407),
.B(n_401),
.C(n_374),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_407),
.B(n_32),
.C(n_2),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_435),
.B(n_405),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_446),
.B(n_447),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_438),
.B(n_422),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_R g449 ( 
.A(n_440),
.B(n_420),
.Y(n_449)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_449),
.B(n_453),
.Y(n_466)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_450),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_439),
.B(n_408),
.C(n_421),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_452),
.B(n_444),
.C(n_436),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_431),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_442),
.B(n_414),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_454),
.B(n_457),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_440),
.A2(n_410),
.B(n_418),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_455),
.B(n_459),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_458),
.B(n_5),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_437),
.A2(n_6),
.B(n_13),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_429),
.Y(n_460)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_460),
.Y(n_463)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_441),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_461),
.B(n_5),
.Y(n_473)
);

AOI21x1_ASAP7_75t_SL g462 ( 
.A1(n_433),
.A2(n_5),
.B(n_10),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g468 ( 
.A(n_462),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_451),
.A2(n_428),
.B1(n_439),
.B2(n_443),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_464),
.A2(n_448),
.B1(n_462),
.B2(n_457),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_450),
.B(n_445),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_470),
.B(n_474),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_471),
.B(n_472),
.Y(n_486)
);

BUFx24_ASAP7_75t_SL g472 ( 
.A(n_456),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_473),
.B(n_1),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_452),
.B(n_434),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_475),
.B(n_459),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_466),
.A2(n_455),
.B(n_458),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_477),
.A2(n_484),
.B(n_467),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_478),
.B(n_482),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_465),
.A2(n_456),
.B(n_449),
.Y(n_479)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_479),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_480),
.B(n_481),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_476),
.B(n_448),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_467),
.A2(n_5),
.B(n_14),
.Y(n_484)
);

BUFx12f_ASAP7_75t_L g485 ( 
.A(n_468),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_485),
.B(n_469),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_483),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_487),
.B(n_489),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_491),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_490),
.B(n_486),
.C(n_483),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_493),
.Y(n_498)
);

NOR3xp33_ASAP7_75t_L g494 ( 
.A(n_492),
.B(n_485),
.C(n_463),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_494),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_498),
.B(n_496),
.C(n_495),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_499),
.A2(n_488),
.B(n_497),
.Y(n_500)
);

A2O1A1Ixp33_ASAP7_75t_L g501 ( 
.A1(n_500),
.A2(n_473),
.B(n_14),
.C(n_4),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_501),
.A2(n_2),
.B(n_4),
.Y(n_502)
);


endmodule