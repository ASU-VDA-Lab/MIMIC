module fake_ariane_1467_n_2841 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_598, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_587, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_588, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_579, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_616, n_617, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_601, n_565, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_575, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_451, n_613, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_606, n_213, n_110, n_304, n_67, n_509, n_583, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_615, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_618, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_573, n_127, n_531, n_2841);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_587;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_588;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_616;
input n_617;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_601;
input n_565;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_575;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_451;
input n_613;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_583;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_615;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_618;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;

output n_2841;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_2484;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_2818;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_2731;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_737;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_958;
wire n_945;
wire n_2554;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_625;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_2370;
wire n_2233;
wire n_2663;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2782;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_2433;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_661;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_2739;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1021;
wire n_1443;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_2717;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_2527;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_2806;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_1260;
wire n_930;
wire n_1179;
wire n_2703;
wire n_696;
wire n_1442;
wire n_2620;
wire n_798;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_2791;
wire n_2683;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2693;
wire n_2745;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_2628;
wire n_619;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_1139;
wire n_2836;
wire n_2439;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_632;
wire n_650;
wire n_2388;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_712;
wire n_976;
wire n_909;
wire n_1832;
wire n_767;
wire n_1392;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_2467;
wire n_2768;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_1913;
wire n_2495;
wire n_2069;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_760;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_2312;
wire n_670;
wire n_2677;
wire n_1826;
wire n_2834;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_637;
wire n_1592;
wire n_2812;
wire n_2662;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_2811;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_2814;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_1053;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_677;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_2783;
wire n_2599;
wire n_699;
wire n_727;
wire n_1726;
wire n_2075;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2496;
wire n_2031;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_729;
wire n_887;
wire n_2218;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2780;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_957;
wire n_1402;
wire n_1242;
wire n_2754;
wire n_2774;
wire n_2707;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_735;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_888;
wire n_845;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_890;
wire n_842;
wire n_1898;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_2821;
wire n_2690;
wire n_2474;
wire n_2623;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1860;
wire n_1734;
wire n_2785;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_951;
wire n_2772;
wire n_862;
wire n_1700;
wire n_2637;
wire n_659;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_2737;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2576;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_2581;
wire n_1783;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_1191;
wire n_2492;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1856;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_2016;
wire n_2667;
wire n_2725;
wire n_1118;
wire n_943;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_2720;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_1324;
wire n_1429;
wire n_2353;
wire n_2064;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_1154;
wire n_1557;
wire n_1759;
wire n_2325;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2477;
wire n_2314;
wire n_2279;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2203;
wire n_2076;
wire n_2133;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_858;
wire n_2796;
wire n_1185;
wire n_2475;
wire n_2804;
wire n_2173;
wire n_2715;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_825;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_2747;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_644;
wire n_1197;
wire n_2820;
wire n_2613;
wire n_1165;
wire n_1641;
wire n_1517;
wire n_2036;
wire n_843;
wire n_2647;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1603;
wire n_1370;
wire n_728;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2331;
wire n_935;
wire n_2478;
wire n_685;
wire n_911;
wire n_2658;
wire n_623;
wire n_2608;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_2767;
wire n_810;
wire n_1290;
wire n_1959;
wire n_2396;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_2692;
wire n_683;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_1193;
wire n_1345;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_2441;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_692;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1910;
wire n_1816;
wire n_2803;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_621;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_697;
wire n_2828;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_1262;
wire n_792;
wire n_1942;
wire n_2180;
wire n_1579;
wire n_2809;
wire n_2181;
wire n_2014;
wire n_975;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2586;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_1024;
wire n_830;
wire n_2291;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_788;
wire n_908;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_2630;
wire n_2794;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2597;
wire n_1077;
wire n_2321;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_2787;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_2395;
wire n_917;
wire n_2723;
wire n_1271;
wire n_2440;
wire n_2096;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_631;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_898;
wire n_857;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_2583;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_701;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_2775;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2447;
wire n_2538;
wire n_1845;
wire n_2034;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2552;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2105;
wire n_2372;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_2587;
wire n_1347;
wire n_2839;
wire n_860;
wire n_1043;
wire n_1923;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_2644;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_2673;
wire n_664;
wire n_1591;
wire n_2585;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2275;
wire n_2205;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_937;
wire n_1474;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_1211;
wire n_996;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_719;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2798;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2797;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_1308;
wire n_796;
wire n_2823;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_88),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_608),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_263),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_377),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_207),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_17),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_492),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_234),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_576),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_191),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_208),
.Y(n_629)
);

INVxp33_ASAP7_75t_L g630 ( 
.A(n_577),
.Y(n_630)
);

CKINVDCx14_ASAP7_75t_R g631 ( 
.A(n_3),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_164),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_15),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_4),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_307),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_467),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_316),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_491),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_263),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_536),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_403),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_149),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_351),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_447),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_10),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_565),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_421),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_99),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_381),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_24),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_347),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_488),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_247),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_372),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_524),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_298),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_573),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_110),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_453),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_122),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_23),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_474),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_67),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g664 ( 
.A(n_596),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_568),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_288),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_512),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_51),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_20),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_93),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_470),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_322),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_546),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_121),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_223),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_567),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_480),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_152),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_459),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_408),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_489),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_166),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_547),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_449),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_140),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_66),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_583),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_611),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_503),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_45),
.Y(n_690)
);

CKINVDCx14_ASAP7_75t_R g691 ( 
.A(n_588),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_174),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_275),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_158),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_334),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_539),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_483),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_572),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_89),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_444),
.Y(n_700)
);

INVx1_ASAP7_75t_SL g701 ( 
.A(n_257),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_167),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_112),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_469),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_437),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_550),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_535),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_578),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_344),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_348),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_591),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_569),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_349),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_525),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_471),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_300),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_6),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_213),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_500),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_553),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_416),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_158),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_64),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_124),
.Y(n_724)
);

BUFx8_ASAP7_75t_SL g725 ( 
.A(n_243),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_543),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_251),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_586),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_593),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_41),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_236),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_363),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_252),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_229),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_615),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_526),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_490),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_75),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_404),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_109),
.Y(n_740)
);

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_296),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_337),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_413),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_90),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_394),
.Y(n_745)
);

INVxp67_ASAP7_75t_L g746 ( 
.A(n_267),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_528),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_606),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_355),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_135),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_595),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_479),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_463),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_63),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_597),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_222),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_554),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_357),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_249),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_496),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_473),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_241),
.Y(n_762)
);

INVx1_ASAP7_75t_SL g763 ( 
.A(n_21),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_361),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_196),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_272),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_519),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_239),
.Y(n_768)
);

BUFx2_ASAP7_75t_L g769 ( 
.A(n_175),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_97),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_271),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_518),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_378),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_52),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_609),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_545),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_412),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_126),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_188),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_610),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_98),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_84),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_257),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_286),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_465),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_178),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_464),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_113),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_429),
.Y(n_789)
);

CKINVDCx20_ASAP7_75t_R g790 ( 
.A(n_534),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_132),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_506),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_48),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_384),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_443),
.Y(n_795)
);

INVx1_ASAP7_75t_SL g796 ( 
.A(n_352),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_300),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_587),
.Y(n_798)
);

BUFx10_ASAP7_75t_L g799 ( 
.A(n_603),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_78),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_356),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_484),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_57),
.Y(n_803)
);

BUFx10_ASAP7_75t_L g804 ( 
.A(n_387),
.Y(n_804)
);

INVx1_ASAP7_75t_SL g805 ( 
.A(n_49),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_504),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_249),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_194),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_507),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_83),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_589),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_558),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_236),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_40),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_456),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_382),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_425),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_581),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_498),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_555),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_118),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_75),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_618),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_274),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_184),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_225),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_287),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_580),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_302),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_440),
.Y(n_830)
);

BUFx3_ASAP7_75t_L g831 ( 
.A(n_95),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_102),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_538),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_147),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_218),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_269),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_485),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_515),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_15),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_67),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_562),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_303),
.Y(n_842)
);

INVxp67_ASAP7_75t_SL g843 ( 
.A(n_154),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_574),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_154),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_600),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_43),
.Y(n_847)
);

CKINVDCx20_ASAP7_75t_R g848 ( 
.A(n_359),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_139),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_454),
.Y(n_850)
);

BUFx5_ASAP7_75t_L g851 ( 
.A(n_150),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_0),
.Y(n_852)
);

INVx2_ASAP7_75t_SL g853 ( 
.A(n_426),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_319),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_168),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_105),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_157),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_566),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_510),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_190),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_14),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_439),
.Y(n_862)
);

BUFx5_ASAP7_75t_L g863 ( 
.A(n_216),
.Y(n_863)
);

BUFx10_ASAP7_75t_L g864 ( 
.A(n_422),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_297),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_77),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_112),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_159),
.Y(n_868)
);

INVx1_ASAP7_75t_SL g869 ( 
.A(n_182),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_516),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_430),
.Y(n_871)
);

CKINVDCx20_ASAP7_75t_R g872 ( 
.A(n_268),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_271),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_237),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_445),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_151),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_462),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_388),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_278),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_579),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_235),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_476),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_511),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_18),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_187),
.Y(n_885)
);

CKINVDCx14_ASAP7_75t_R g886 ( 
.A(n_301),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_358),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_272),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_448),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_601),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_561),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_282),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_442),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_571),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_22),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_286),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_329),
.Y(n_897)
);

BUFx10_ASAP7_75t_L g898 ( 
.A(n_614),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_594),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_373),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_192),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_451),
.Y(n_902)
);

INVx1_ASAP7_75t_SL g903 ( 
.A(n_208),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_256),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_590),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_446),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_16),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_280),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_441),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_134),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_410),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_478),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_172),
.Y(n_913)
);

CKINVDCx20_ASAP7_75t_R g914 ( 
.A(n_341),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_156),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_530),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_325),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_338),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_152),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_268),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_7),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_436),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_262),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_279),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_450),
.Y(n_925)
);

CKINVDCx20_ASAP7_75t_R g926 ( 
.A(n_43),
.Y(n_926)
);

CKINVDCx16_ASAP7_75t_R g927 ( 
.A(n_402),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_475),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_499),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_607),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_187),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_521),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_548),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_339),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_457),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_612),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_540),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_461),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_460),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_482),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_419),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_513),
.Y(n_942)
);

INVx1_ASAP7_75t_SL g943 ( 
.A(n_477),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_564),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_604),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_505),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_99),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_487),
.Y(n_948)
);

BUFx5_ASAP7_75t_L g949 ( 
.A(n_103),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_105),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_160),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_342),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_256),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_433),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_210),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_103),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_309),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_584),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_585),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_315),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_40),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_232),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_18),
.Y(n_963)
);

INVx1_ASAP7_75t_SL g964 ( 
.A(n_537),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_218),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_551),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_129),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_196),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_360),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_122),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_531),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_549),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_235),
.Y(n_973)
);

INVx1_ASAP7_75t_SL g974 ( 
.A(n_114),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_542),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_582),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_375),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_431),
.Y(n_978)
);

INVxp67_ASAP7_75t_L g979 ( 
.A(n_560),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_552),
.Y(n_980)
);

CKINVDCx11_ASAP7_75t_R g981 ( 
.A(n_230),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_502),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_340),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_486),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_228),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_366),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_186),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_520),
.Y(n_988)
);

BUFx10_ASAP7_75t_L g989 ( 
.A(n_57),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_522),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_165),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_501),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_223),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_270),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_407),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_497),
.Y(n_996)
);

CKINVDCx16_ASAP7_75t_R g997 ( 
.A(n_254),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_157),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_142),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_390),
.Y(n_1000)
);

CKINVDCx20_ASAP7_75t_R g1001 ( 
.A(n_466),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_29),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_262),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_222),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_118),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_284),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_599),
.Y(n_1007)
);

BUFx8_ASAP7_75t_SL g1008 ( 
.A(n_532),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_354),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_523),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_211),
.Y(n_1011)
);

INVx1_ASAP7_75t_SL g1012 ( 
.A(n_613),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_126),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_237),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_136),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_207),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_414),
.Y(n_1017)
);

INVx2_ASAP7_75t_SL g1018 ( 
.A(n_81),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_113),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_179),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_514),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_95),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_598),
.Y(n_1023)
);

CKINVDCx20_ASAP7_75t_R g1024 ( 
.A(n_85),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_213),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_435),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_570),
.Y(n_1027)
);

CKINVDCx20_ASAP7_75t_R g1028 ( 
.A(n_259),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_31),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_209),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_541),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_102),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_495),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_493),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_163),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_452),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_438),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_279),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_275),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_164),
.Y(n_1040)
);

CKINVDCx16_ASAP7_75t_R g1041 ( 
.A(n_557),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_22),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_46),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_0),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_405),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_66),
.Y(n_1046)
);

BUFx5_ASAP7_75t_L g1047 ( 
.A(n_87),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_307),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_323),
.Y(n_1049)
);

CKINVDCx20_ASAP7_75t_R g1050 ( 
.A(n_168),
.Y(n_1050)
);

CKINVDCx20_ASAP7_75t_R g1051 ( 
.A(n_304),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_188),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_517),
.Y(n_1053)
);

CKINVDCx14_ASAP7_75t_R g1054 ( 
.A(n_88),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_79),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_243),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_494),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_56),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_132),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_559),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_617),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_149),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_247),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_455),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_37),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_162),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_137),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_556),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_227),
.Y(n_1069)
);

BUFx8_ASAP7_75t_SL g1070 ( 
.A(n_602),
.Y(n_1070)
);

BUFx5_ASAP7_75t_L g1071 ( 
.A(n_261),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_94),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_527),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_217),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_41),
.Y(n_1075)
);

CKINVDCx14_ASAP7_75t_R g1076 ( 
.A(n_311),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_420),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_468),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_90),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_227),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_108),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_147),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_244),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_201),
.Y(n_1084)
);

CKINVDCx20_ASAP7_75t_R g1085 ( 
.A(n_509),
.Y(n_1085)
);

CKINVDCx20_ASAP7_75t_R g1086 ( 
.A(n_592),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_458),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_385),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_605),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_575),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_544),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_508),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_533),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_380),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_293),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_161),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_529),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_276),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_26),
.Y(n_1099)
);

INVxp67_ASAP7_75t_L g1100 ( 
.A(n_481),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_367),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_472),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_30),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_87),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_53),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_246),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_301),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_269),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_54),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_283),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_24),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_94),
.Y(n_1112)
);

CKINVDCx20_ASAP7_75t_R g1113 ( 
.A(n_48),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_55),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_31),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_178),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_317),
.Y(n_1117)
);

INVx2_ASAP7_75t_SL g1118 ( 
.A(n_255),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_221),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_204),
.Y(n_1120)
);

BUFx10_ASAP7_75t_L g1121 ( 
.A(n_411),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_216),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_616),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_563),
.Y(n_1124)
);

CKINVDCx20_ASAP7_75t_R g1125 ( 
.A(n_252),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_12),
.Y(n_1126)
);

BUFx8_ASAP7_75t_SL g1127 ( 
.A(n_219),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_886),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_886),
.B(n_1),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_953),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_769),
.B(n_1),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_642),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_642),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_642),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_989),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_642),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1054),
.B(n_2),
.Y(n_1137)
);

CKINVDCx11_ASAP7_75t_R g1138 ( 
.A(n_981),
.Y(n_1138)
);

NOR2x1_ASAP7_75t_L g1139 ( 
.A(n_641),
.B(n_310),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_851),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1054),
.B(n_2),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_997),
.B(n_3),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_1004),
.Y(n_1143)
);

BUFx3_ASAP7_75t_L g1144 ( 
.A(n_1023),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_744),
.Y(n_1145)
);

BUFx12f_ASAP7_75t_L g1146 ( 
.A(n_799),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_884),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_680),
.B(n_4),
.Y(n_1148)
);

INVx5_ASAP7_75t_L g1149 ( 
.A(n_799),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_686),
.B(n_5),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_744),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_989),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_725),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_631),
.B(n_691),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_686),
.B(n_5),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_831),
.Y(n_1156)
);

INVx4_ASAP7_75t_L g1157 ( 
.A(n_641),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_743),
.B(n_6),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_831),
.Y(n_1159)
);

NOR2x1_ASAP7_75t_L g1160 ( 
.A(n_698),
.B(n_312),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_744),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_764),
.B(n_7),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_895),
.Y(n_1163)
);

INVx2_ASAP7_75t_SL g1164 ( 
.A(n_895),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_1006),
.B(n_8),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_1112),
.Y(n_1166)
);

BUFx3_ASAP7_75t_L g1167 ( 
.A(n_804),
.Y(n_1167)
);

CKINVDCx20_ASAP7_75t_R g1168 ( 
.A(n_1127),
.Y(n_1168)
);

INVx5_ASAP7_75t_L g1169 ( 
.A(n_804),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_744),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_691),
.B(n_8),
.Y(n_1171)
);

AND2x6_ASAP7_75t_L g1172 ( 
.A(n_698),
.B(n_313),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_781),
.Y(n_1173)
);

HB1xp67_ASAP7_75t_L g1174 ( 
.A(n_1006),
.Y(n_1174)
);

BUFx12f_ASAP7_75t_L g1175 ( 
.A(n_864),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_794),
.B(n_9),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1076),
.B(n_9),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_830),
.B(n_10),
.Y(n_1178)
);

BUFx12f_ASAP7_75t_L g1179 ( 
.A(n_864),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1076),
.B(n_11),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_922),
.B(n_630),
.Y(n_1181)
);

BUFx12f_ASAP7_75t_L g1182 ( 
.A(n_898),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_622),
.B(n_11),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_851),
.B(n_12),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_637),
.B(n_13),
.Y(n_1185)
);

INVx2_ASAP7_75t_SL g1186 ( 
.A(n_898),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_621),
.B(n_13),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1018),
.B(n_14),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_851),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1118),
.B(n_16),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_621),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_719),
.B(n_17),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_851),
.B(n_19),
.Y(n_1193)
);

BUFx8_ASAP7_75t_SL g1194 ( 
.A(n_650),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_927),
.B(n_19),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_647),
.B(n_20),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_719),
.B(n_21),
.Y(n_1197)
);

INVx5_ASAP7_75t_L g1198 ( 
.A(n_1121),
.Y(n_1198)
);

INVx5_ASAP7_75t_L g1199 ( 
.A(n_1121),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_858),
.B(n_23),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_851),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_654),
.B(n_25),
.Y(n_1202)
);

INVx4_ASAP7_75t_L g1203 ( 
.A(n_858),
.Y(n_1203)
);

BUFx6f_ASAP7_75t_L g1204 ( 
.A(n_781),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_781),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_851),
.Y(n_1206)
);

BUFx12f_ASAP7_75t_L g1207 ( 
.A(n_619),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_781),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_813),
.Y(n_1209)
);

INVx2_ASAP7_75t_SL g1210 ( 
.A(n_634),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_958),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_813),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_863),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_958),
.B(n_25),
.Y(n_1214)
);

INVx1_ASAP7_75t_SL g1215 ( 
.A(n_663),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_813),
.Y(n_1216)
);

INVx5_ASAP7_75t_L g1217 ( 
.A(n_1008),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_634),
.B(n_26),
.Y(n_1218)
);

INVx5_ASAP7_75t_L g1219 ( 
.A(n_667),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_657),
.B(n_27),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_675),
.B(n_685),
.Y(n_1221)
);

BUFx8_ASAP7_75t_SL g1222 ( 
.A(n_668),
.Y(n_1222)
);

INVx5_ASAP7_75t_L g1223 ( 
.A(n_667),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_659),
.B(n_27),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_671),
.B(n_28),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_675),
.B(n_28),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_685),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_676),
.B(n_29),
.Y(n_1228)
);

HB1xp67_ASAP7_75t_L g1229 ( 
.A(n_623),
.Y(n_1229)
);

INVx5_ASAP7_75t_L g1230 ( 
.A(n_667),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_863),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_813),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_863),
.B(n_30),
.Y(n_1233)
);

INVx5_ASAP7_75t_L g1234 ( 
.A(n_667),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_863),
.Y(n_1235)
);

INVx5_ASAP7_75t_L g1236 ( 
.A(n_801),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_863),
.Y(n_1237)
);

BUFx8_ASAP7_75t_L g1238 ( 
.A(n_715),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_863),
.Y(n_1239)
);

AND2x6_ASAP7_75t_L g1240 ( 
.A(n_620),
.B(n_640),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_SL g1241 ( 
.A(n_1041),
.B(n_314),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_684),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_731),
.B(n_32),
.Y(n_1243)
);

INVx4_ASAP7_75t_L g1244 ( 
.A(n_801),
.Y(n_1244)
);

CKINVDCx6p67_ASAP7_75t_R g1245 ( 
.A(n_649),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_949),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_949),
.B(n_32),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_688),
.B(n_33),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_829),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_689),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_700),
.B(n_33),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_829),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_731),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_949),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_829),
.Y(n_1255)
);

INVx5_ASAP7_75t_L g1256 ( 
.A(n_1070),
.Y(n_1256)
);

INVx4_ASAP7_75t_L g1257 ( 
.A(n_801),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_651),
.Y(n_1258)
);

BUFx12f_ASAP7_75t_L g1259 ( 
.A(n_626),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_707),
.B(n_34),
.Y(n_1260)
);

INVx4_ASAP7_75t_L g1261 ( 
.A(n_801),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_949),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_710),
.B(n_712),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_720),
.B(n_34),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_733),
.B(n_35),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_949),
.Y(n_1266)
);

INVx4_ASAP7_75t_L g1267 ( 
.A(n_935),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_829),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_733),
.B(n_35),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_840),
.Y(n_1270)
);

AND2x6_ASAP7_75t_L g1271 ( 
.A(n_620),
.B(n_318),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_840),
.B(n_36),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_949),
.B(n_36),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_857),
.B(n_37),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_857),
.B(n_38),
.Y(n_1275)
);

BUFx12f_ASAP7_75t_L g1276 ( 
.A(n_629),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_1002),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_729),
.B(n_38),
.Y(n_1278)
);

BUFx12f_ASAP7_75t_L g1279 ( 
.A(n_633),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1002),
.B(n_1046),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1047),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_737),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1046),
.B(n_39),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_748),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_758),
.B(n_39),
.Y(n_1285)
);

BUFx8_ASAP7_75t_L g1286 ( 
.A(n_721),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1047),
.B(n_42),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_888),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_635),
.Y(n_1289)
);

INVx3_ASAP7_75t_L g1290 ( 
.A(n_1048),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1048),
.Y(n_1291)
);

BUFx8_ASAP7_75t_SL g1292 ( 
.A(n_738),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_761),
.B(n_42),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_888),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_888),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1084),
.B(n_44),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1084),
.B(n_44),
.Y(n_1297)
);

CKINVDCx6p67_ASAP7_75t_R g1298 ( 
.A(n_652),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1047),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1047),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1132),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1189),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1132),
.Y(n_1303)
);

AOI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1181),
.A2(n_1050),
.B1(n_771),
.B2(n_788),
.Y(n_1304)
);

AOI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1171),
.A2(n_1180),
.B1(n_1177),
.B2(n_1137),
.Y(n_1305)
);

OAI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1147),
.A2(n_741),
.B1(n_872),
.B2(n_847),
.Y(n_1306)
);

OR2x6_ASAP7_75t_L g1307 ( 
.A(n_1146),
.B(n_746),
.Y(n_1307)
);

AOI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1171),
.A2(n_1024),
.B1(n_1025),
.B2(n_926),
.Y(n_1308)
);

AOI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1177),
.A2(n_1113),
.B1(n_1051),
.B2(n_1111),
.Y(n_1309)
);

AOI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1180),
.A2(n_1125),
.B1(n_1028),
.B2(n_713),
.Y(n_1310)
);

BUFx10_ASAP7_75t_L g1311 ( 
.A(n_1153),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1128),
.B(n_1116),
.Y(n_1312)
);

OAI22xp33_ASAP7_75t_SL g1313 ( 
.A1(n_1195),
.A2(n_1142),
.B1(n_1162),
.B2(n_1148),
.Y(n_1313)
);

AOI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1129),
.A2(n_726),
.B1(n_790),
.B2(n_755),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1128),
.B(n_1116),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1149),
.B(n_664),
.Y(n_1316)
);

NAND2xp33_ASAP7_75t_SL g1317 ( 
.A(n_1129),
.B(n_888),
.Y(n_1317)
);

AO22x2_ASAP7_75t_L g1318 ( 
.A1(n_1137),
.A2(n_763),
.B1(n_805),
.B2(n_701),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1133),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1147),
.B(n_624),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1154),
.B(n_1122),
.Y(n_1321)
);

BUFx6f_ASAP7_75t_SL g1322 ( 
.A(n_1167),
.Y(n_1322)
);

OAI22xp33_ASAP7_75t_SL g1323 ( 
.A1(n_1176),
.A2(n_1108),
.B1(n_903),
.B2(n_923),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1254),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1133),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_1166),
.B(n_628),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1134),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1134),
.Y(n_1328)
);

AO22x2_ASAP7_75t_L g1329 ( 
.A1(n_1141),
.A2(n_869),
.B1(n_974),
.B2(n_843),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1141),
.A2(n_900),
.B1(n_914),
.B2(n_848),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1266),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1281),
.Y(n_1332)
);

AOI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1241),
.A2(n_939),
.B1(n_944),
.B2(n_929),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1154),
.B(n_901),
.Y(n_1334)
);

INVxp67_ASAP7_75t_SL g1335 ( 
.A(n_1211),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1149),
.B(n_1122),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_SL g1337 ( 
.A1(n_1215),
.A2(n_1085),
.B1(n_1086),
.B2(n_1001),
.Y(n_1337)
);

INVx8_ASAP7_75t_L g1338 ( 
.A(n_1217),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1156),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1136),
.Y(n_1340)
);

AOI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1166),
.A2(n_661),
.B1(n_674),
.B2(n_645),
.Y(n_1341)
);

INVxp67_ASAP7_75t_L g1342 ( 
.A(n_1229),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1136),
.Y(n_1343)
);

AO22x2_ASAP7_75t_L g1344 ( 
.A1(n_1131),
.A2(n_648),
.B1(n_660),
.B2(n_632),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1145),
.Y(n_1345)
);

AO22x2_ASAP7_75t_L g1346 ( 
.A1(n_1188),
.A2(n_666),
.B1(n_692),
.B2(n_682),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1258),
.Y(n_1347)
);

OAI22xp33_ASAP7_75t_SL g1348 ( 
.A1(n_1178),
.A2(n_656),
.B1(n_658),
.B2(n_639),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1145),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1151),
.Y(n_1350)
);

AO22x2_ASAP7_75t_L g1351 ( 
.A1(n_1190),
.A2(n_702),
.B1(n_716),
.B2(n_699),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1159),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1151),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_SL g1354 ( 
.A1(n_1168),
.A2(n_653),
.B1(n_670),
.B2(n_669),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1161),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1149),
.B(n_767),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1161),
.Y(n_1357)
);

AOI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1144),
.A2(n_717),
.B1(n_791),
.B2(n_703),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1163),
.Y(n_1359)
);

AO22x2_ASAP7_75t_L g1360 ( 
.A1(n_1226),
.A2(n_1265),
.B1(n_1275),
.B2(n_1243),
.Y(n_1360)
);

OAI22xp33_ASAP7_75t_SL g1361 ( 
.A1(n_1158),
.A2(n_690),
.B1(n_693),
.B2(n_678),
.Y(n_1361)
);

AOI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1186),
.A2(n_810),
.B1(n_861),
.B2(n_727),
.Y(n_1362)
);

AO22x2_ASAP7_75t_L g1363 ( 
.A1(n_1192),
.A2(n_740),
.B1(n_754),
.B2(n_730),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1169),
.B(n_1047),
.Y(n_1364)
);

AOI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1130),
.A2(n_1143),
.B1(n_1289),
.B2(n_1200),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1174),
.B(n_756),
.Y(n_1366)
);

OAI22xp33_ASAP7_75t_R g1367 ( 
.A1(n_1183),
.A2(n_836),
.B1(n_1042),
.B2(n_783),
.Y(n_1367)
);

AND2x6_ASAP7_75t_L g1368 ( 
.A(n_1197),
.B(n_640),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1169),
.B(n_762),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1214),
.A2(n_694),
.B1(n_722),
.B2(n_718),
.Y(n_1370)
);

AO22x2_ASAP7_75t_L g1371 ( 
.A1(n_1150),
.A2(n_766),
.B1(n_784),
.B2(n_778),
.Y(n_1371)
);

AO22x2_ASAP7_75t_L g1372 ( 
.A1(n_1155),
.A2(n_808),
.B1(n_822),
.B2(n_786),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1135),
.A2(n_797),
.B1(n_832),
.B2(n_782),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1140),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1170),
.Y(n_1375)
);

AOI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1152),
.A2(n_1175),
.B1(n_1182),
.B2(n_1179),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1198),
.B(n_1047),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1198),
.B(n_1071),
.Y(n_1378)
);

OAI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1245),
.A2(n_1119),
.B1(n_1120),
.B2(n_1114),
.Y(n_1379)
);

AO22x2_ASAP7_75t_L g1380 ( 
.A1(n_1165),
.A2(n_826),
.B1(n_827),
.B2(n_824),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_SL g1381 ( 
.A1(n_1207),
.A2(n_724),
.B1(n_734),
.B2(n_723),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1199),
.B(n_1071),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_SL g1383 ( 
.A1(n_1259),
.A2(n_759),
.B1(n_765),
.B2(n_750),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1201),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1199),
.B(n_839),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1170),
.Y(n_1386)
);

AOI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1185),
.A2(n_768),
.B1(n_874),
.B2(n_779),
.Y(n_1387)
);

AOI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1196),
.A2(n_770),
.B1(n_814),
.B2(n_800),
.Y(n_1388)
);

AO22x2_ASAP7_75t_L g1389 ( 
.A1(n_1221),
.A2(n_845),
.B1(n_856),
.B2(n_842),
.Y(n_1389)
);

OAI22xp33_ASAP7_75t_R g1390 ( 
.A1(n_1202),
.A2(n_867),
.B1(n_881),
.B2(n_860),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1206),
.Y(n_1391)
);

OAI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1298),
.A2(n_1104),
.B1(n_1105),
.B2(n_1103),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1173),
.Y(n_1393)
);

AO22x2_ASAP7_75t_L g1394 ( 
.A1(n_1280),
.A2(n_908),
.B1(n_913),
.B2(n_896),
.Y(n_1394)
);

INVx2_ASAP7_75t_SL g1395 ( 
.A(n_1217),
.Y(n_1395)
);

AOI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1220),
.A2(n_849),
.B1(n_865),
.B2(n_803),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1164),
.B(n_1071),
.Y(n_1397)
);

AOI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1224),
.A2(n_852),
.B1(n_892),
.B2(n_834),
.Y(n_1398)
);

BUFx6f_ASAP7_75t_SL g1399 ( 
.A(n_1210),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1256),
.Y(n_1400)
);

AO22x2_ASAP7_75t_L g1401 ( 
.A1(n_1187),
.A2(n_951),
.B1(n_956),
.B2(n_931),
.Y(n_1401)
);

AOI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1225),
.A2(n_873),
.B1(n_910),
.B2(n_835),
.Y(n_1402)
);

AOI22x1_ASAP7_75t_L g1403 ( 
.A1(n_1187),
.A2(n_774),
.B1(n_807),
.B2(n_793),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1157),
.Y(n_1404)
);

OAI22xp33_ASAP7_75t_SL g1405 ( 
.A1(n_1227),
.A2(n_825),
.B1(n_868),
.B2(n_855),
.Y(n_1405)
);

AO22x2_ASAP7_75t_L g1406 ( 
.A1(n_1218),
.A2(n_962),
.B1(n_970),
.B2(n_961),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1173),
.Y(n_1407)
);

INVx4_ASAP7_75t_L g1408 ( 
.A(n_1256),
.Y(n_1408)
);

INVx1_ASAP7_75t_SL g1409 ( 
.A(n_1138),
.Y(n_1409)
);

AO22x2_ASAP7_75t_L g1410 ( 
.A1(n_1218),
.A2(n_985),
.B1(n_991),
.B2(n_973),
.Y(n_1410)
);

OAI22xp33_ASAP7_75t_SL g1411 ( 
.A1(n_1227),
.A2(n_866),
.B1(n_879),
.B2(n_876),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1270),
.B(n_1071),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1213),
.Y(n_1413)
);

AO22x2_ASAP7_75t_L g1414 ( 
.A1(n_1269),
.A2(n_1003),
.B1(n_1011),
.B2(n_998),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1203),
.B(n_979),
.Y(n_1415)
);

AOI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1228),
.A2(n_904),
.B1(n_963),
.B2(n_821),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1263),
.B(n_1100),
.Y(n_1417)
);

OA22x2_ASAP7_75t_L g1418 ( 
.A1(n_1270),
.A2(n_1030),
.B1(n_1035),
.B2(n_1019),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1276),
.Y(n_1419)
);

AO22x2_ASAP7_75t_L g1420 ( 
.A1(n_1269),
.A2(n_1274),
.B1(n_1283),
.B2(n_1272),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1204),
.Y(n_1421)
);

AND2x2_ASAP7_75t_SL g1422 ( 
.A(n_1272),
.B(n_672),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1248),
.A2(n_885),
.B1(n_915),
.B2(n_907),
.Y(n_1423)
);

OAI22xp33_ASAP7_75t_SL g1424 ( 
.A1(n_1291),
.A2(n_920),
.B1(n_924),
.B2(n_919),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1291),
.B(n_1071),
.Y(n_1425)
);

OAI22xp33_ASAP7_75t_SL g1426 ( 
.A1(n_1242),
.A2(n_947),
.B1(n_950),
.B2(n_921),
.Y(n_1426)
);

AOI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1251),
.A2(n_1005),
.B1(n_1016),
.B2(n_967),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1231),
.Y(n_1428)
);

AO22x2_ASAP7_75t_L g1429 ( 
.A1(n_1274),
.A2(n_1043),
.B1(n_1052),
.B2(n_1038),
.Y(n_1429)
);

AOI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1260),
.A2(n_1278),
.B1(n_1285),
.B2(n_1264),
.Y(n_1430)
);

AOI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1293),
.A2(n_1099),
.B1(n_1080),
.B2(n_965),
.Y(n_1431)
);

INVx2_ASAP7_75t_SL g1432 ( 
.A(n_1238),
.Y(n_1432)
);

AO22x2_ASAP7_75t_L g1433 ( 
.A1(n_1283),
.A2(n_1067),
.B1(n_1072),
.B2(n_1066),
.Y(n_1433)
);

OAI22xp33_ASAP7_75t_R g1434 ( 
.A1(n_1194),
.A2(n_1081),
.B1(n_1083),
.B2(n_1079),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1279),
.A2(n_1022),
.B1(n_1055),
.B2(n_993),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1250),
.B(n_1071),
.Y(n_1436)
);

AOI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1286),
.A2(n_1039),
.B1(n_1058),
.B2(n_994),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_1282),
.B(n_1284),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1191),
.B(n_968),
.Y(n_1439)
);

AO22x2_ASAP7_75t_L g1440 ( 
.A1(n_1296),
.A2(n_1115),
.B1(n_1109),
.B2(n_776),
.Y(n_1440)
);

OAI22xp33_ASAP7_75t_SL g1441 ( 
.A1(n_1184),
.A2(n_987),
.B1(n_1013),
.B2(n_999),
.Y(n_1441)
);

AO22x2_ASAP7_75t_L g1442 ( 
.A1(n_1296),
.A2(n_796),
.B1(n_943),
.B2(n_644),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_SL g1443 ( 
.A1(n_1222),
.A2(n_1014),
.B1(n_1015),
.B2(n_955),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1204),
.Y(n_1444)
);

AO22x2_ASAP7_75t_L g1445 ( 
.A1(n_1297),
.A2(n_1012),
.B1(n_964),
.B2(n_681),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1253),
.B(n_1277),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1290),
.B(n_968),
.Y(n_1447)
);

OAI22xp33_ASAP7_75t_R g1448 ( 
.A1(n_1292),
.A2(n_1029),
.B1(n_1032),
.B2(n_1020),
.Y(n_1448)
);

OAI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1297),
.A2(n_1126),
.B1(n_1040),
.B2(n_1056),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1205),
.B(n_1059),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1235),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1205),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1237),
.Y(n_1453)
);

INVx3_ASAP7_75t_L g1454 ( 
.A(n_1208),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1219),
.B(n_1223),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1208),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_SL g1457 ( 
.A1(n_1193),
.A2(n_1044),
.B1(n_1065),
.B2(n_1063),
.Y(n_1457)
);

AO22x2_ASAP7_75t_L g1458 ( 
.A1(n_1233),
.A2(n_681),
.B1(n_714),
.B2(n_672),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1244),
.B(n_773),
.Y(n_1459)
);

AOI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1172),
.A2(n_1074),
.B1(n_1098),
.B2(n_1082),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1209),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1239),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1246),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_1257),
.Y(n_1464)
);

AO22x2_ASAP7_75t_L g1465 ( 
.A1(n_1247),
.A2(n_802),
.B1(n_844),
.B2(n_714),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1209),
.Y(n_1466)
);

INVx3_ASAP7_75t_L g1467 ( 
.A(n_1212),
.Y(n_1467)
);

OAI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1273),
.A2(n_1110),
.B1(n_1107),
.B2(n_1095),
.Y(n_1468)
);

OA22x2_ASAP7_75t_L g1469 ( 
.A1(n_1287),
.A2(n_1096),
.B1(n_1106),
.B2(n_1069),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1212),
.Y(n_1470)
);

INVx3_ASAP7_75t_L g1471 ( 
.A(n_1216),
.Y(n_1471)
);

INVxp33_ASAP7_75t_L g1472 ( 
.A(n_1216),
.Y(n_1472)
);

INVxp33_ASAP7_75t_L g1473 ( 
.A(n_1232),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1219),
.B(n_968),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1232),
.Y(n_1475)
);

AOI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1172),
.A2(n_853),
.B1(n_1033),
.B2(n_850),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1249),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_1261),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1267),
.B(n_775),
.Y(n_1479)
);

OAI22xp33_ASAP7_75t_R g1480 ( 
.A1(n_1262),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_1480)
);

OAI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1139),
.A2(n_1075),
.B1(n_968),
.B2(n_1062),
.Y(n_1481)
);

CKINVDCx20_ASAP7_75t_R g1482 ( 
.A(n_1249),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1172),
.A2(n_1094),
.B1(n_844),
.B2(n_936),
.Y(n_1483)
);

OAI22xp33_ASAP7_75t_SL g1484 ( 
.A1(n_1160),
.A2(n_785),
.B1(n_787),
.B2(n_780),
.Y(n_1484)
);

AO22x2_ASAP7_75t_L g1485 ( 
.A1(n_1300),
.A2(n_936),
.B1(n_952),
.B2(n_802),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1252),
.Y(n_1486)
);

OAI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1252),
.A2(n_1075),
.B1(n_1062),
.B2(n_982),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_SL g1488 ( 
.A1(n_1255),
.A2(n_1075),
.B1(n_1062),
.B2(n_982),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1299),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1255),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1268),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1219),
.B(n_1062),
.Y(n_1492)
);

AO22x2_ASAP7_75t_L g1493 ( 
.A1(n_1240),
.A2(n_1094),
.B1(n_952),
.B2(n_795),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1268),
.Y(n_1494)
);

AND2x2_ASAP7_75t_SL g1495 ( 
.A(n_1288),
.B(n_1075),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1288),
.Y(n_1496)
);

OAI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1294),
.A2(n_798),
.B1(n_811),
.B2(n_792),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1223),
.B(n_1092),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1294),
.B(n_815),
.Y(n_1499)
);

AOI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1240),
.A2(n_838),
.B1(n_859),
.B2(n_833),
.Y(n_1500)
);

OAI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1295),
.A2(n_880),
.B1(n_882),
.B2(n_878),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_SL g1502 ( 
.A1(n_1295),
.A2(n_887),
.B1(n_889),
.B2(n_883),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1223),
.Y(n_1503)
);

AOI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1240),
.A2(n_1271),
.B1(n_917),
.B2(n_928),
.Y(n_1504)
);

AO22x2_ASAP7_75t_L g1505 ( 
.A1(n_1271),
.A2(n_933),
.B1(n_934),
.B2(n_911),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1230),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1230),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1230),
.Y(n_1508)
);

NOR2x1p5_ASAP7_75t_L g1509 ( 
.A(n_1271),
.B(n_1091),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1234),
.Y(n_1510)
);

AOI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1234),
.A2(n_941),
.B1(n_942),
.B2(n_940),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1234),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1236),
.B(n_946),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1236),
.Y(n_1514)
);

OAI22x1_ASAP7_75t_L g1515 ( 
.A1(n_1236),
.A2(n_977),
.B1(n_986),
.B2(n_976),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1132),
.Y(n_1516)
);

AO22x2_ASAP7_75t_L g1517 ( 
.A1(n_1171),
.A2(n_992),
.B1(n_996),
.B2(n_988),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1132),
.Y(n_1518)
);

OAI22xp33_ASAP7_75t_R g1519 ( 
.A1(n_1158),
.A2(n_50),
.B1(n_47),
.B2(n_49),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1128),
.B(n_1087),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1132),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1181),
.A2(n_1078),
.B1(n_1026),
.B2(n_1009),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1181),
.A2(n_1017),
.B1(n_1027),
.B2(n_1007),
.Y(n_1523)
);

INVx2_ASAP7_75t_SL g1524 ( 
.A(n_1149),
.Y(n_1524)
);

INVx3_ASAP7_75t_L g1525 ( 
.A(n_1211),
.Y(n_1525)
);

AOI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1181),
.A2(n_1049),
.B1(n_1068),
.B2(n_1045),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1128),
.B(n_1124),
.Y(n_1527)
);

AOI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1181),
.A2(n_1088),
.B1(n_1097),
.B2(n_1077),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1189),
.Y(n_1529)
);

OAI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1147),
.A2(n_1123),
.B1(n_1101),
.B2(n_627),
.Y(n_1530)
);

AOI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1181),
.A2(n_636),
.B1(n_638),
.B2(n_625),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1189),
.Y(n_1532)
);

INVx8_ASAP7_75t_L g1533 ( 
.A(n_1217),
.Y(n_1533)
);

OAI22xp33_ASAP7_75t_SL g1534 ( 
.A1(n_1195),
.A2(n_646),
.B1(n_655),
.B2(n_643),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1128),
.B(n_662),
.Y(n_1535)
);

AOI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1181),
.A2(n_673),
.B1(n_677),
.B2(n_665),
.Y(n_1536)
);

OAI22xp33_ASAP7_75t_R g1537 ( 
.A1(n_1158),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_1537)
);

OAI22xp33_ASAP7_75t_SL g1538 ( 
.A1(n_1195),
.A2(n_683),
.B1(n_687),
.B2(n_679),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1132),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1132),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1128),
.B(n_935),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1189),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1181),
.A2(n_696),
.B1(n_697),
.B2(n_695),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1128),
.B(n_704),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1181),
.A2(n_706),
.B1(n_708),
.B2(n_705),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_1258),
.Y(n_1546)
);

AND2x2_ASAP7_75t_SL g1547 ( 
.A(n_1241),
.B(n_935),
.Y(n_1547)
);

AO22x2_ASAP7_75t_L g1548 ( 
.A1(n_1171),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1189),
.Y(n_1549)
);

AOI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1181),
.A2(n_711),
.B1(n_728),
.B2(n_709),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1132),
.Y(n_1551)
);

AOI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1181),
.A2(n_735),
.B1(n_736),
.B2(n_732),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1128),
.B(n_935),
.Y(n_1553)
);

OAI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1147),
.A2(n_742),
.B1(n_745),
.B2(n_739),
.Y(n_1554)
);

OA22x2_ASAP7_75t_L g1555 ( 
.A1(n_1130),
.A2(n_749),
.B1(n_751),
.B2(n_747),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1128),
.B(n_752),
.Y(n_1556)
);

AO22x2_ASAP7_75t_L g1557 ( 
.A1(n_1171),
.A2(n_59),
.B1(n_56),
.B2(n_58),
.Y(n_1557)
);

AO22x2_ASAP7_75t_L g1558 ( 
.A1(n_1171),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1189),
.Y(n_1559)
);

AO22x2_ASAP7_75t_L g1560 ( 
.A1(n_1171),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_1560)
);

INVx3_ASAP7_75t_L g1561 ( 
.A(n_1211),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1181),
.A2(n_757),
.B1(n_760),
.B2(n_753),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1258),
.Y(n_1563)
);

OAI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1147),
.A2(n_777),
.B1(n_789),
.B2(n_772),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1189),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1132),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_SL g1567 ( 
.A1(n_1215),
.A2(n_809),
.B1(n_812),
.B2(n_806),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1132),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1181),
.A2(n_817),
.B1(n_818),
.B2(n_816),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_SL g1570 ( 
.A(n_1154),
.B(n_819),
.Y(n_1570)
);

BUFx6f_ASAP7_75t_L g1571 ( 
.A(n_1132),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1189),
.Y(n_1572)
);

OAI22xp33_ASAP7_75t_SL g1573 ( 
.A1(n_1195),
.A2(n_823),
.B1(n_828),
.B2(n_820),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1128),
.B(n_837),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1189),
.Y(n_1575)
);

INVxp67_ASAP7_75t_SL g1576 ( 
.A(n_1211),
.Y(n_1576)
);

OAI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1147),
.A2(n_846),
.B1(n_854),
.B2(n_841),
.Y(n_1577)
);

AOI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1181),
.A2(n_870),
.B1(n_871),
.B2(n_862),
.Y(n_1578)
);

AOI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1181),
.A2(n_877),
.B1(n_890),
.B2(n_875),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1128),
.B(n_891),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_SL g1581 ( 
.A1(n_1215),
.A2(n_894),
.B1(n_897),
.B2(n_893),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1211),
.Y(n_1582)
);

AOI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1181),
.A2(n_902),
.B1(n_905),
.B2(n_899),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1128),
.B(n_906),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1132),
.Y(n_1585)
);

AOI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1181),
.A2(n_912),
.B1(n_916),
.B2(n_909),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1128),
.B(n_918),
.Y(n_1587)
);

AO22x2_ASAP7_75t_L g1588 ( 
.A1(n_1171),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_1588)
);

OR2x6_ASAP7_75t_L g1589 ( 
.A(n_1146),
.B(n_1073),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_1154),
.B(n_925),
.Y(n_1590)
);

OR2x6_ASAP7_75t_L g1591 ( 
.A(n_1146),
.B(n_1073),
.Y(n_1591)
);

AO22x2_ASAP7_75t_L g1592 ( 
.A1(n_1171),
.A2(n_68),
.B1(n_64),
.B2(n_65),
.Y(n_1592)
);

AO22x2_ASAP7_75t_L g1593 ( 
.A1(n_1171),
.A2(n_69),
.B1(n_65),
.B2(n_68),
.Y(n_1593)
);

NAND2xp33_ASAP7_75t_SL g1594 ( 
.A(n_1129),
.B(n_1073),
.Y(n_1594)
);

OA22x2_ASAP7_75t_L g1595 ( 
.A1(n_1130),
.A2(n_932),
.B1(n_937),
.B2(n_930),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_1149),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1132),
.Y(n_1597)
);

AO22x2_ASAP7_75t_L g1598 ( 
.A1(n_1171),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_1598)
);

BUFx10_ASAP7_75t_L g1599 ( 
.A(n_1153),
.Y(n_1599)
);

OAI22xp33_ASAP7_75t_SL g1600 ( 
.A1(n_1195),
.A2(n_945),
.B1(n_948),
.B2(n_938),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1189),
.Y(n_1601)
);

OAI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1147),
.A2(n_957),
.B1(n_959),
.B2(n_954),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1128),
.B(n_1073),
.Y(n_1603)
);

AOI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1181),
.A2(n_966),
.B1(n_969),
.B2(n_960),
.Y(n_1604)
);

OAI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1147),
.A2(n_972),
.B1(n_975),
.B2(n_971),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1128),
.B(n_978),
.Y(n_1606)
);

OAI22xp33_ASAP7_75t_SL g1607 ( 
.A1(n_1195),
.A2(n_983),
.B1(n_984),
.B2(n_980),
.Y(n_1607)
);

AOI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1181),
.A2(n_995),
.B1(n_1000),
.B2(n_990),
.Y(n_1608)
);

BUFx6f_ASAP7_75t_SL g1609 ( 
.A(n_1167),
.Y(n_1609)
);

AO22x2_ASAP7_75t_L g1610 ( 
.A1(n_1171),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_1610)
);

OAI22xp33_ASAP7_75t_SL g1611 ( 
.A1(n_1195),
.A2(n_1021),
.B1(n_1031),
.B2(n_1010),
.Y(n_1611)
);

AND2x4_ASAP7_75t_L g1612 ( 
.A(n_1128),
.B(n_1034),
.Y(n_1612)
);

AND2x2_ASAP7_75t_SL g1613 ( 
.A(n_1241),
.B(n_1036),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1128),
.B(n_1037),
.Y(n_1614)
);

AO22x2_ASAP7_75t_L g1615 ( 
.A1(n_1171),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1181),
.A2(n_1057),
.B1(n_1060),
.B2(n_1053),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1132),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1128),
.B(n_1061),
.Y(n_1618)
);

AOI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1181),
.A2(n_1089),
.B1(n_1090),
.B2(n_1064),
.Y(n_1619)
);

AOI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1181),
.A2(n_1102),
.B1(n_1117),
.B2(n_1093),
.Y(n_1620)
);

INVx4_ASAP7_75t_L g1621 ( 
.A(n_1149),
.Y(n_1621)
);

AO22x2_ASAP7_75t_L g1622 ( 
.A1(n_1171),
.A2(n_76),
.B1(n_73),
.B2(n_74),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1189),
.Y(n_1623)
);

AOI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1181),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_1624)
);

AOI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1181),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_1625)
);

OAI22xp33_ASAP7_75t_SL g1626 ( 
.A1(n_1195),
.A2(n_83),
.B1(n_80),
.B2(n_82),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1147),
.B(n_82),
.Y(n_1627)
);

OAI22xp33_ASAP7_75t_SL g1628 ( 
.A1(n_1195),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1628)
);

OAI22xp33_ASAP7_75t_SL g1629 ( 
.A1(n_1195),
.A2(n_91),
.B1(n_86),
.B2(n_89),
.Y(n_1629)
);

INVx2_ASAP7_75t_SL g1630 ( 
.A(n_1149),
.Y(n_1630)
);

OAI22xp33_ASAP7_75t_SL g1631 ( 
.A1(n_1195),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1215),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1215),
.Y(n_1633)
);

OAI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1147),
.A2(n_97),
.B1(n_92),
.B2(n_96),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1154),
.B(n_96),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1189),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1632),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1404),
.B(n_98),
.Y(n_1638)
);

XOR2xp5_ASAP7_75t_L g1639 ( 
.A(n_1347),
.B(n_100),
.Y(n_1639)
);

INVx1_ASAP7_75t_SL g1640 ( 
.A(n_1633),
.Y(n_1640)
);

XNOR2x2_ASAP7_75t_L g1641 ( 
.A(n_1304),
.B(n_100),
.Y(n_1641)
);

XNOR2x2_ASAP7_75t_L g1642 ( 
.A(n_1442),
.B(n_101),
.Y(n_1642)
);

XNOR2xp5_ASAP7_75t_L g1643 ( 
.A(n_1333),
.B(n_101),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1422),
.B(n_104),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1374),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1339),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1352),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1359),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1302),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1324),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1331),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1541),
.B(n_104),
.Y(n_1652)
);

BUFx6f_ASAP7_75t_L g1653 ( 
.A(n_1444),
.Y(n_1653)
);

CKINVDCx20_ASAP7_75t_R g1654 ( 
.A(n_1546),
.Y(n_1654)
);

NAND2x1p5_ASAP7_75t_L g1655 ( 
.A(n_1525),
.B(n_106),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1332),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1529),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1532),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1542),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1342),
.B(n_106),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1553),
.B(n_107),
.Y(n_1661)
);

BUFx5_ASAP7_75t_L g1662 ( 
.A(n_1384),
.Y(n_1662)
);

BUFx6f_ASAP7_75t_L g1663 ( 
.A(n_1444),
.Y(n_1663)
);

CKINVDCx16_ASAP7_75t_R g1664 ( 
.A(n_1311),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1549),
.Y(n_1665)
);

AOI21x1_ASAP7_75t_L g1666 ( 
.A1(n_1559),
.A2(n_321),
.B(n_320),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1565),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1391),
.Y(n_1668)
);

INVxp33_ASAP7_75t_L g1669 ( 
.A(n_1337),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1430),
.B(n_107),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1572),
.Y(n_1671)
);

INVxp33_ASAP7_75t_L g1672 ( 
.A(n_1438),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1575),
.A2(n_326),
.B(n_324),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1601),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1417),
.B(n_108),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1623),
.Y(n_1676)
);

NOR2xp67_ASAP7_75t_L g1677 ( 
.A(n_1432),
.B(n_327),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1335),
.B(n_109),
.Y(n_1678)
);

OAI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1483),
.A2(n_1636),
.B(n_1476),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1413),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1368),
.B(n_110),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_1563),
.Y(n_1682)
);

XNOR2xp5_ASAP7_75t_L g1683 ( 
.A(n_1306),
.B(n_111),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1368),
.B(n_111),
.Y(n_1684)
);

XNOR2x2_ASAP7_75t_L g1685 ( 
.A(n_1442),
.B(n_114),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1428),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_SL g1687 ( 
.A(n_1547),
.B(n_115),
.Y(n_1687)
);

INVxp67_ASAP7_75t_SL g1688 ( 
.A(n_1561),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1451),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1453),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1462),
.Y(n_1691)
);

INVxp33_ASAP7_75t_L g1692 ( 
.A(n_1446),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1463),
.Y(n_1693)
);

INVxp67_ASAP7_75t_L g1694 ( 
.A(n_1582),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1489),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1301),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1439),
.Y(n_1697)
);

INVxp33_ASAP7_75t_SL g1698 ( 
.A(n_1409),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1303),
.Y(n_1699)
);

INVx2_ASAP7_75t_SL g1700 ( 
.A(n_1612),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1520),
.B(n_115),
.Y(n_1701)
);

INVxp67_ASAP7_75t_SL g1702 ( 
.A(n_1474),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1447),
.Y(n_1703)
);

BUFx2_ASAP7_75t_R g1704 ( 
.A(n_1419),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_SL g1705 ( 
.A(n_1613),
.B(n_116),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1368),
.B(n_116),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1603),
.B(n_117),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1527),
.B(n_117),
.Y(n_1708)
);

BUFx6f_ASAP7_75t_L g1709 ( 
.A(n_1452),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1499),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1535),
.B(n_119),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1544),
.B(n_119),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1556),
.B(n_120),
.Y(n_1713)
);

XNOR2x2_ASAP7_75t_L g1714 ( 
.A(n_1445),
.B(n_120),
.Y(n_1714)
);

OAI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1412),
.A2(n_330),
.B(n_328),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1397),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1319),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1576),
.B(n_121),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1436),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1425),
.Y(n_1720)
);

OAI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1504),
.A2(n_332),
.B(n_331),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_1599),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1492),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1321),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1336),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1364),
.Y(n_1726)
);

XOR2xp5_ASAP7_75t_L g1727 ( 
.A(n_1314),
.B(n_123),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1377),
.Y(n_1728)
);

INVx4_ASAP7_75t_SL g1729 ( 
.A(n_1322),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1378),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1325),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1382),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1503),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_SL g1734 ( 
.A(n_1554),
.B(n_123),
.Y(n_1734)
);

AND2x2_ASAP7_75t_SL g1735 ( 
.A(n_1330),
.B(n_124),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_1609),
.Y(n_1736)
);

CKINVDCx16_ASAP7_75t_R g1737 ( 
.A(n_1589),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_L g1738 ( 
.A(n_1570),
.B(n_125),
.Y(n_1738)
);

OAI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1460),
.A2(n_335),
.B(n_333),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1506),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1512),
.Y(n_1741)
);

XOR2xp5_ASAP7_75t_L g1742 ( 
.A(n_1310),
.B(n_125),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1514),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1450),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1507),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1590),
.B(n_127),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1508),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1510),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1312),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1315),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1327),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1543),
.B(n_127),
.Y(n_1752)
);

INVxp67_ASAP7_75t_SL g1753 ( 
.A(n_1455),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1328),
.Y(n_1754)
);

OAI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1635),
.A2(n_343),
.B(n_336),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1340),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1343),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1498),
.B(n_128),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1345),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1349),
.Y(n_1760)
);

XOR2xp5_ASAP7_75t_L g1761 ( 
.A(n_1308),
.B(n_128),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1350),
.Y(n_1762)
);

CKINVDCx20_ASAP7_75t_R g1763 ( 
.A(n_1482),
.Y(n_1763)
);

XOR2xp5_ASAP7_75t_L g1764 ( 
.A(n_1309),
.B(n_129),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1353),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1355),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1357),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1574),
.B(n_130),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1375),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1386),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1393),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1545),
.B(n_130),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1407),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1421),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1320),
.B(n_131),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1305),
.B(n_131),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1456),
.Y(n_1777)
);

CKINVDCx5p33_ASAP7_75t_R g1778 ( 
.A(n_1338),
.Y(n_1778)
);

INVxp33_ASAP7_75t_L g1779 ( 
.A(n_1341),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1461),
.Y(n_1780)
);

INVxp67_ASAP7_75t_SL g1781 ( 
.A(n_1459),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1562),
.B(n_133),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1466),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1334),
.B(n_133),
.Y(n_1784)
);

CKINVDCx20_ASAP7_75t_R g1785 ( 
.A(n_1567),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1470),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1580),
.B(n_134),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1475),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1477),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1569),
.B(n_135),
.Y(n_1790)
);

XOR2xp5_ASAP7_75t_L g1791 ( 
.A(n_1443),
.B(n_136),
.Y(n_1791)
);

CKINVDCx20_ASAP7_75t_R g1792 ( 
.A(n_1581),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_1338),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1486),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1584),
.B(n_137),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1490),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1491),
.Y(n_1797)
);

XOR2xp5_ASAP7_75t_L g1798 ( 
.A(n_1354),
.B(n_138),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1587),
.B(n_138),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1494),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1496),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1516),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1518),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1606),
.B(n_139),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1521),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1539),
.Y(n_1806)
);

CKINVDCx20_ASAP7_75t_R g1807 ( 
.A(n_1589),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1540),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1551),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1566),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1568),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1585),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1614),
.B(n_140),
.Y(n_1813)
);

XNOR2x2_ASAP7_75t_L g1814 ( 
.A(n_1445),
.B(n_141),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1597),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1420),
.B(n_141),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1420),
.B(n_142),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1617),
.Y(n_1818)
);

INVx2_ASAP7_75t_SL g1819 ( 
.A(n_1591),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1485),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1485),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1454),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1618),
.B(n_143),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1360),
.B(n_143),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1467),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1471),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1478),
.Y(n_1827)
);

NOR2x1p5_ASAP7_75t_L g1828 ( 
.A(n_1627),
.B(n_144),
.Y(n_1828)
);

XNOR2xp5_ASAP7_75t_L g1829 ( 
.A(n_1376),
.B(n_144),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1452),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1513),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1479),
.Y(n_1832)
);

OR2x6_ASAP7_75t_L g1833 ( 
.A(n_1548),
.B(n_1557),
.Y(n_1833)
);

NOR2xp67_ASAP7_75t_L g1834 ( 
.A(n_1395),
.B(n_345),
.Y(n_1834)
);

INVxp33_ASAP7_75t_L g1835 ( 
.A(n_1326),
.Y(n_1835)
);

INVxp33_ASAP7_75t_L g1836 ( 
.A(n_1365),
.Y(n_1836)
);

OAI21xp5_ASAP7_75t_L g1837 ( 
.A1(n_1531),
.A2(n_350),
.B(n_346),
.Y(n_1837)
);

XOR2x2_ASAP7_75t_L g1838 ( 
.A(n_1555),
.B(n_145),
.Y(n_1838)
);

CKINVDCx5p33_ASAP7_75t_R g1839 ( 
.A(n_1533),
.Y(n_1839)
);

XNOR2xp5_ASAP7_75t_L g1840 ( 
.A(n_1318),
.B(n_1329),
.Y(n_1840)
);

OAI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1536),
.A2(n_362),
.B(n_353),
.Y(n_1841)
);

CKINVDCx5p33_ASAP7_75t_R g1842 ( 
.A(n_1533),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1493),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1493),
.Y(n_1844)
);

AND2x2_ASAP7_75t_SL g1845 ( 
.A(n_1495),
.B(n_145),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1360),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1369),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1616),
.B(n_146),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1385),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1571),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1571),
.Y(n_1851)
);

NOR2xp33_ASAP7_75t_SL g1852 ( 
.A(n_1379),
.B(n_146),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1366),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1418),
.Y(n_1854)
);

INVx4_ASAP7_75t_SL g1855 ( 
.A(n_1591),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1356),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1389),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1358),
.B(n_148),
.Y(n_1858)
);

XOR2xp5_ASAP7_75t_L g1859 ( 
.A(n_1435),
.B(n_148),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1389),
.Y(n_1860)
);

NAND2xp33_ASAP7_75t_SL g1861 ( 
.A(n_1457),
.B(n_150),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1394),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1394),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1621),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1401),
.B(n_1406),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1472),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1473),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1401),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1406),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1410),
.B(n_151),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1410),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1550),
.B(n_153),
.Y(n_1872)
);

AND2x6_ASAP7_75t_L g1873 ( 
.A(n_1500),
.B(n_1526),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1414),
.Y(n_1874)
);

INVxp33_ASAP7_75t_L g1875 ( 
.A(n_1423),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1552),
.B(n_153),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1578),
.B(n_155),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1414),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1429),
.Y(n_1879)
);

AND2x4_ASAP7_75t_L g1880 ( 
.A(n_1524),
.B(n_155),
.Y(n_1880)
);

INVx2_ASAP7_75t_SL g1881 ( 
.A(n_1596),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1429),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1433),
.B(n_156),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1509),
.Y(n_1884)
);

BUFx6f_ASAP7_75t_L g1885 ( 
.A(n_1630),
.Y(n_1885)
);

CKINVDCx5p33_ASAP7_75t_R g1886 ( 
.A(n_1399),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1433),
.Y(n_1887)
);

HB1xp67_ASAP7_75t_SL g1888 ( 
.A(n_1318),
.Y(n_1888)
);

INVxp33_ASAP7_75t_L g1889 ( 
.A(n_1316),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1458),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1458),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1307),
.B(n_159),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1464),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1465),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1465),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1346),
.Y(n_1896)
);

NAND2xp33_ASAP7_75t_R g1897 ( 
.A(n_1307),
.B(n_160),
.Y(n_1897)
);

XOR2x2_ASAP7_75t_L g1898 ( 
.A(n_1595),
.B(n_161),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1346),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1403),
.Y(n_1900)
);

HB1xp67_ASAP7_75t_L g1901 ( 
.A(n_1415),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1351),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1579),
.B(n_162),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1351),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1522),
.Y(n_1905)
);

OAI21xp5_ASAP7_75t_L g1906 ( 
.A1(n_1583),
.A2(n_365),
.B(n_364),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1523),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1317),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1528),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1517),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1517),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1371),
.Y(n_1912)
);

BUFx3_ASAP7_75t_L g1913 ( 
.A(n_1400),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1371),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1372),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1515),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1372),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1586),
.B(n_163),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1380),
.Y(n_1919)
);

XOR2xp5_ASAP7_75t_L g1920 ( 
.A(n_1381),
.B(n_1383),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1380),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1363),
.Y(n_1922)
);

AND2x4_ASAP7_75t_L g1923 ( 
.A(n_1373),
.B(n_165),
.Y(n_1923)
);

OR2x2_ASAP7_75t_L g1924 ( 
.A(n_1362),
.B(n_166),
.Y(n_1924)
);

INVxp33_ASAP7_75t_L g1925 ( 
.A(n_1329),
.Y(n_1925)
);

NOR2xp33_ASAP7_75t_L g1926 ( 
.A(n_1604),
.B(n_167),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1363),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1344),
.B(n_169),
.Y(n_1928)
);

OR2x2_ASAP7_75t_SL g1929 ( 
.A(n_1367),
.B(n_169),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1344),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1469),
.Y(n_1931)
);

XOR2xp5_ASAP7_75t_L g1932 ( 
.A(n_1437),
.B(n_170),
.Y(n_1932)
);

INVxp67_ASAP7_75t_SL g1933 ( 
.A(n_1481),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1594),
.Y(n_1934)
);

AND2x4_ASAP7_75t_L g1935 ( 
.A(n_1387),
.B(n_170),
.Y(n_1935)
);

CKINVDCx20_ASAP7_75t_R g1936 ( 
.A(n_1608),
.Y(n_1936)
);

CKINVDCx14_ASAP7_75t_R g1937 ( 
.A(n_1370),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1388),
.B(n_171),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1396),
.B(n_1398),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1505),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1619),
.B(n_171),
.Y(n_1941)
);

BUFx6f_ASAP7_75t_L g1942 ( 
.A(n_1408),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1313),
.Y(n_1943)
);

NOR2xp33_ASAP7_75t_L g1944 ( 
.A(n_1620),
.B(n_172),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1402),
.B(n_173),
.Y(n_1945)
);

CKINVDCx20_ASAP7_75t_R g1946 ( 
.A(n_1416),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1505),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1468),
.B(n_173),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1511),
.Y(n_1949)
);

OAI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1484),
.A2(n_369),
.B(n_368),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1440),
.Y(n_1951)
);

OR2x6_ASAP7_75t_L g1952 ( 
.A(n_1548),
.B(n_1557),
.Y(n_1952)
);

XNOR2x2_ASAP7_75t_L g1953 ( 
.A(n_1558),
.B(n_1560),
.Y(n_1953)
);

INVxp33_ASAP7_75t_L g1954 ( 
.A(n_1427),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1440),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1624),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1625),
.Y(n_1957)
);

BUFx6f_ASAP7_75t_L g1958 ( 
.A(n_1626),
.Y(n_1958)
);

BUFx3_ASAP7_75t_L g1959 ( 
.A(n_1488),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1502),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1628),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1649),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1640),
.B(n_1431),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1650),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1637),
.B(n_1558),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1835),
.B(n_1560),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1781),
.B(n_1449),
.Y(n_1967)
);

BUFx3_ASAP7_75t_L g1968 ( 
.A(n_1763),
.Y(n_1968)
);

INVx2_ASAP7_75t_SL g1969 ( 
.A(n_1700),
.Y(n_1969)
);

INVx8_ASAP7_75t_L g1970 ( 
.A(n_1778),
.Y(n_1970)
);

AND2x4_ASAP7_75t_L g1971 ( 
.A(n_1855),
.B(n_1846),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1853),
.B(n_1588),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1832),
.B(n_1564),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1651),
.Y(n_1974)
);

BUFx3_ASAP7_75t_L g1975 ( 
.A(n_1654),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1656),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1749),
.B(n_1588),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1702),
.B(n_1577),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1657),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1645),
.Y(n_1980)
);

BUFx3_ASAP7_75t_L g1981 ( 
.A(n_1682),
.Y(n_1981)
);

AND2x6_ASAP7_75t_L g1982 ( 
.A(n_1940),
.B(n_1592),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1658),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1750),
.B(n_1592),
.Y(n_1984)
);

AND2x2_ASAP7_75t_SL g1985 ( 
.A(n_1735),
.B(n_1448),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1668),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1659),
.Y(n_1987)
);

INVx3_ASAP7_75t_L g1988 ( 
.A(n_1696),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1665),
.Y(n_1989)
);

OAI21xp5_ASAP7_75t_L g1990 ( 
.A1(n_1900),
.A2(n_1538),
.B(n_1534),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1680),
.Y(n_1991)
);

AND2x4_ASAP7_75t_L g1992 ( 
.A(n_1855),
.B(n_1573),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1686),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1689),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1901),
.B(n_1602),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1672),
.B(n_1593),
.Y(n_1996)
);

OAI21xp5_ASAP7_75t_L g1997 ( 
.A1(n_1716),
.A2(n_1607),
.B(n_1600),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1692),
.B(n_1593),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1690),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1664),
.B(n_1598),
.Y(n_2000)
);

NOR2xp33_ASAP7_75t_L g2001 ( 
.A(n_1954),
.B(n_1611),
.Y(n_2001)
);

HB1xp67_ASAP7_75t_L g2002 ( 
.A(n_1652),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1667),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1710),
.B(n_1598),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1691),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1720),
.B(n_1753),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1671),
.Y(n_2007)
);

INVx3_ASAP7_75t_L g2008 ( 
.A(n_1699),
.Y(n_2008)
);

BUFx4f_ASAP7_75t_L g2009 ( 
.A(n_1845),
.Y(n_2009)
);

BUFx6f_ASAP7_75t_L g2010 ( 
.A(n_1653),
.Y(n_2010)
);

BUFx6f_ASAP7_75t_L g2011 ( 
.A(n_1653),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1693),
.Y(n_2012)
);

BUFx4f_ASAP7_75t_SL g2013 ( 
.A(n_1807),
.Y(n_2013)
);

INVxp67_ASAP7_75t_L g2014 ( 
.A(n_1705),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1724),
.B(n_1610),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1695),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1717),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1731),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1675),
.B(n_1605),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1933),
.B(n_1530),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1808),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1939),
.B(n_1856),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1674),
.Y(n_2023)
);

INVxp67_ASAP7_75t_SL g2024 ( 
.A(n_1652),
.Y(n_2024)
);

INVxp67_ASAP7_75t_L g2025 ( 
.A(n_1704),
.Y(n_2025)
);

INVxp67_ASAP7_75t_SL g2026 ( 
.A(n_1661),
.Y(n_2026)
);

INVx2_ASAP7_75t_SL g2027 ( 
.A(n_1819),
.Y(n_2027)
);

NOR2xp33_ASAP7_75t_SL g2028 ( 
.A(n_1687),
.B(n_1392),
.Y(n_2028)
);

BUFx3_ASAP7_75t_L g2029 ( 
.A(n_1722),
.Y(n_2029)
);

OAI21xp5_ASAP7_75t_L g2030 ( 
.A1(n_1755),
.A2(n_1441),
.B(n_1361),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1676),
.Y(n_2031)
);

NAND2xp33_ASAP7_75t_SL g2032 ( 
.A(n_1875),
.B(n_1480),
.Y(n_2032)
);

HB1xp67_ASAP7_75t_L g2033 ( 
.A(n_1661),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1662),
.Y(n_2034)
);

INVx4_ASAP7_75t_L g2035 ( 
.A(n_1729),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1670),
.B(n_1726),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_SL g2037 ( 
.A(n_1876),
.B(n_1629),
.Y(n_2037)
);

AND2x4_ASAP7_75t_L g2038 ( 
.A(n_1784),
.B(n_174),
.Y(n_2038)
);

BUFx6f_ASAP7_75t_L g2039 ( 
.A(n_1653),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1662),
.Y(n_2040)
);

HB1xp67_ASAP7_75t_L g2041 ( 
.A(n_1698),
.Y(n_2041)
);

BUFx6f_ASAP7_75t_L g2042 ( 
.A(n_1663),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1728),
.B(n_1631),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1836),
.B(n_1610),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1737),
.B(n_1615),
.Y(n_2045)
);

BUFx3_ASAP7_75t_L g2046 ( 
.A(n_1793),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1779),
.B(n_1615),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1733),
.Y(n_2048)
);

CKINVDCx5p33_ASAP7_75t_R g2049 ( 
.A(n_1736),
.Y(n_2049)
);

BUFx6f_ASAP7_75t_L g2050 ( 
.A(n_1663),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1660),
.B(n_1865),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1744),
.B(n_1622),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1662),
.Y(n_2053)
);

INVx4_ASAP7_75t_L g2054 ( 
.A(n_1729),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1824),
.B(n_1622),
.Y(n_2055)
);

INVxp67_ASAP7_75t_L g2056 ( 
.A(n_1877),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1662),
.Y(n_2057)
);

BUFx3_ASAP7_75t_L g2058 ( 
.A(n_1839),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1730),
.B(n_1323),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1732),
.B(n_1348),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1662),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1646),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1740),
.Y(n_2063)
);

INVx3_ASAP7_75t_L g2064 ( 
.A(n_1864),
.Y(n_2064)
);

AND2x4_ASAP7_75t_L g2065 ( 
.A(n_1784),
.B(n_175),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_1909),
.B(n_1390),
.Y(n_2066)
);

INVxp67_ASAP7_75t_SL g2067 ( 
.A(n_1694),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_1886),
.B(n_1842),
.Y(n_2068)
);

BUFx5_ASAP7_75t_L g2069 ( 
.A(n_1843),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1644),
.B(n_1497),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1741),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_1743),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1647),
.Y(n_2073)
);

INVx3_ASAP7_75t_L g2074 ( 
.A(n_1663),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_1913),
.B(n_176),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1751),
.Y(n_2076)
);

NOR2xp33_ASAP7_75t_L g2077 ( 
.A(n_1889),
.B(n_1426),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1648),
.Y(n_2078)
);

OR2x2_ASAP7_75t_L g2079 ( 
.A(n_1775),
.B(n_1634),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1719),
.B(n_1501),
.Y(n_2080)
);

BUFx3_ASAP7_75t_L g2081 ( 
.A(n_1942),
.Y(n_2081)
);

BUFx3_ASAP7_75t_L g2082 ( 
.A(n_1942),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_1935),
.B(n_176),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1873),
.B(n_1405),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1844),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1754),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_1935),
.B(n_177),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_1870),
.B(n_177),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1873),
.B(n_1411),
.Y(n_2089)
);

INVx3_ASAP7_75t_L g2090 ( 
.A(n_1709),
.Y(n_2090)
);

BUFx6f_ASAP7_75t_L g2091 ( 
.A(n_1709),
.Y(n_2091)
);

BUFx6f_ASAP7_75t_L g2092 ( 
.A(n_1709),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1756),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_1873),
.B(n_1424),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_1883),
.B(n_179),
.Y(n_2095)
);

INVx3_ASAP7_75t_L g2096 ( 
.A(n_1745),
.Y(n_2096)
);

OR2x2_ASAP7_75t_L g2097 ( 
.A(n_1905),
.B(n_1487),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_1907),
.B(n_180),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1747),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1873),
.B(n_180),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_1757),
.Y(n_2101)
);

OAI21xp5_ASAP7_75t_L g2102 ( 
.A1(n_1679),
.A2(n_371),
.B(n_370),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_1827),
.B(n_181),
.Y(n_2103)
);

BUFx6f_ASAP7_75t_L g2104 ( 
.A(n_1942),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1748),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1723),
.B(n_181),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1820),
.Y(n_2107)
);

NOR2xp33_ASAP7_75t_L g2108 ( 
.A(n_1943),
.B(n_182),
.Y(n_2108)
);

HB1xp67_ASAP7_75t_L g2109 ( 
.A(n_1833),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1759),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1821),
.Y(n_2111)
);

INVxp67_ASAP7_75t_L g2112 ( 
.A(n_1903),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_1923),
.B(n_183),
.Y(n_2113)
);

NOR2xp33_ASAP7_75t_L g2114 ( 
.A(n_1949),
.B(n_183),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1760),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_1923),
.B(n_184),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1697),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_1703),
.B(n_185),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1762),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_1833),
.B(n_185),
.Y(n_2120)
);

AND2x2_ASAP7_75t_SL g2121 ( 
.A(n_1852),
.B(n_1519),
.Y(n_2121)
);

AND2x2_ASAP7_75t_SL g2122 ( 
.A(n_1926),
.B(n_1537),
.Y(n_2122)
);

NOR2xp33_ASAP7_75t_L g2123 ( 
.A(n_1823),
.B(n_186),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_1952),
.B(n_189),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1765),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_1952),
.B(n_189),
.Y(n_2126)
);

NAND2x1p5_ASAP7_75t_L g2127 ( 
.A(n_1896),
.B(n_1434),
.Y(n_2127)
);

HB1xp67_ASAP7_75t_L g2128 ( 
.A(n_1928),
.Y(n_2128)
);

BUFx2_ASAP7_75t_L g2129 ( 
.A(n_1953),
.Y(n_2129)
);

NOR2xp33_ASAP7_75t_L g2130 ( 
.A(n_1884),
.B(n_190),
.Y(n_2130)
);

INVx1_ASAP7_75t_SL g2131 ( 
.A(n_1701),
.Y(n_2131)
);

OAI21xp5_ASAP7_75t_L g2132 ( 
.A1(n_1715),
.A2(n_376),
.B(n_374),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1766),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1725),
.B(n_191),
.Y(n_2134)
);

INVxp67_ASAP7_75t_SL g2135 ( 
.A(n_1688),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_1937),
.B(n_192),
.Y(n_2136)
);

NOR2xp33_ASAP7_75t_L g2137 ( 
.A(n_1893),
.B(n_193),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1767),
.Y(n_2138)
);

NOR2xp33_ASAP7_75t_L g2139 ( 
.A(n_1956),
.B(n_193),
.Y(n_2139)
);

INVx2_ASAP7_75t_SL g2140 ( 
.A(n_1718),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_1708),
.B(n_194),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1947),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1769),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1770),
.Y(n_2144)
);

BUFx3_ASAP7_75t_L g2145 ( 
.A(n_1866),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1771),
.Y(n_2146)
);

NOR2xp33_ASAP7_75t_R g2147 ( 
.A(n_1936),
.B(n_379),
.Y(n_2147)
);

AND2x2_ASAP7_75t_L g2148 ( 
.A(n_1711),
.B(n_195),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_1712),
.B(n_195),
.Y(n_2149)
);

AND2x4_ASAP7_75t_L g2150 ( 
.A(n_1857),
.B(n_197),
.Y(n_2150)
);

INVx1_ASAP7_75t_SL g2151 ( 
.A(n_1713),
.Y(n_2151)
);

BUFx2_ASAP7_75t_L g2152 ( 
.A(n_1938),
.Y(n_2152)
);

INVx4_ASAP7_75t_L g2153 ( 
.A(n_1885),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1773),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_1774),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_1777),
.Y(n_2156)
);

HB1xp67_ASAP7_75t_L g2157 ( 
.A(n_1768),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1780),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1783),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_1787),
.B(n_197),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_1795),
.B(n_198),
.Y(n_2161)
);

HB1xp67_ASAP7_75t_L g2162 ( 
.A(n_1799),
.Y(n_2162)
);

BUFx8_ASAP7_75t_L g2163 ( 
.A(n_1858),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_L g2164 ( 
.A(n_1804),
.B(n_198),
.Y(n_2164)
);

BUFx6f_ASAP7_75t_L g2165 ( 
.A(n_1885),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1786),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_1788),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1789),
.Y(n_2168)
);

INVxp67_ASAP7_75t_SL g2169 ( 
.A(n_1718),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_1813),
.B(n_199),
.Y(n_2170)
);

BUFx6f_ASAP7_75t_L g2171 ( 
.A(n_1885),
.Y(n_2171)
);

NOR2xp33_ASAP7_75t_L g2172 ( 
.A(n_1957),
.B(n_199),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_1794),
.Y(n_2173)
);

INVx3_ASAP7_75t_L g2174 ( 
.A(n_1796),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_1868),
.B(n_1869),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_1871),
.B(n_1874),
.Y(n_2176)
);

HB1xp67_ASAP7_75t_L g2177 ( 
.A(n_1912),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_1878),
.B(n_1879),
.Y(n_2178)
);

OAI21xp33_ASAP7_75t_L g2179 ( 
.A1(n_1752),
.A2(n_1782),
.B(n_1772),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_1797),
.Y(n_2180)
);

AND2x4_ASAP7_75t_L g2181 ( 
.A(n_1860),
.B(n_200),
.Y(n_2181)
);

BUFx3_ASAP7_75t_L g2182 ( 
.A(n_1867),
.Y(n_2182)
);

BUFx2_ASAP7_75t_L g2183 ( 
.A(n_1945),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_1882),
.B(n_200),
.Y(n_2184)
);

OAI21xp5_ASAP7_75t_L g2185 ( 
.A1(n_1758),
.A2(n_386),
.B(n_383),
.Y(n_2185)
);

INVx4_ASAP7_75t_L g2186 ( 
.A(n_1880),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_1776),
.B(n_201),
.Y(n_2187)
);

BUFx3_ASAP7_75t_L g2188 ( 
.A(n_1830),
.Y(n_2188)
);

OAI21xp5_ASAP7_75t_L g2189 ( 
.A1(n_1934),
.A2(n_1908),
.B(n_1673),
.Y(n_2189)
);

BUFx3_ASAP7_75t_L g2190 ( 
.A(n_1851),
.Y(n_2190)
);

NOR2xp33_ASAP7_75t_L g2191 ( 
.A(n_1961),
.B(n_1914),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_1800),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_1801),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_1887),
.B(n_202),
.Y(n_2194)
);

AND2x4_ASAP7_75t_L g2195 ( 
.A(n_1862),
.B(n_202),
.Y(n_2195)
);

AND2x2_ASAP7_75t_SL g2196 ( 
.A(n_1944),
.B(n_203),
.Y(n_2196)
);

NOR2xp67_ASAP7_75t_L g2197 ( 
.A(n_1837),
.B(n_389),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_1738),
.B(n_203),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_1899),
.B(n_204),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_1902),
.B(n_205),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_1746),
.B(n_205),
.Y(n_2201)
);

BUFx3_ASAP7_75t_L g2202 ( 
.A(n_1850),
.Y(n_2202)
);

INVxp67_ASAP7_75t_L g2203 ( 
.A(n_1790),
.Y(n_2203)
);

AND2x2_ASAP7_75t_SL g2204 ( 
.A(n_1848),
.B(n_206),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_1802),
.Y(n_2205)
);

AND2x4_ASAP7_75t_L g2206 ( 
.A(n_1863),
.B(n_206),
.Y(n_2206)
);

INVx4_ASAP7_75t_L g2207 ( 
.A(n_1880),
.Y(n_2207)
);

BUFx6f_ASAP7_75t_L g2208 ( 
.A(n_1655),
.Y(n_2208)
);

INVxp67_ASAP7_75t_SL g2209 ( 
.A(n_2169),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2022),
.B(n_1961),
.Y(n_2210)
);

BUFx12f_ASAP7_75t_L g2211 ( 
.A(n_2035),
.Y(n_2211)
);

AND2x4_ASAP7_75t_L g2212 ( 
.A(n_1968),
.B(n_1904),
.Y(n_2212)
);

AND2x4_ASAP7_75t_L g2213 ( 
.A(n_2035),
.B(n_1930),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_1963),
.B(n_1946),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_1980),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_1986),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_2048),
.Y(n_2217)
);

CKINVDCx20_ASAP7_75t_R g2218 ( 
.A(n_2041),
.Y(n_2218)
);

AND2x2_ASAP7_75t_SL g2219 ( 
.A(n_2196),
.B(n_1924),
.Y(n_2219)
);

BUFx8_ASAP7_75t_L g2220 ( 
.A(n_1975),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2142),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2066),
.B(n_1910),
.Y(n_2222)
);

BUFx6f_ASAP7_75t_L g2223 ( 
.A(n_2054),
.Y(n_2223)
);

AND2x4_ASAP7_75t_L g2224 ( 
.A(n_2054),
.B(n_1981),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2142),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2019),
.B(n_1958),
.Y(n_2226)
);

BUFx6f_ASAP7_75t_L g2227 ( 
.A(n_2104),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_2056),
.B(n_1958),
.Y(n_2228)
);

AND2x4_ASAP7_75t_L g2229 ( 
.A(n_1971),
.B(n_1915),
.Y(n_2229)
);

NAND2x1p5_ASAP7_75t_L g2230 ( 
.A(n_2081),
.B(n_1917),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_2063),
.Y(n_2231)
);

NOR2xp33_ASAP7_75t_L g2232 ( 
.A(n_2179),
.B(n_1958),
.Y(n_2232)
);

AND2x6_ASAP7_75t_L g2233 ( 
.A(n_2150),
.B(n_1919),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2085),
.Y(n_2234)
);

INVx4_ASAP7_75t_L g2235 ( 
.A(n_1970),
.Y(n_2235)
);

AND2x4_ASAP7_75t_L g2236 ( 
.A(n_1971),
.B(n_1921),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_2112),
.B(n_1911),
.Y(n_2237)
);

BUFx2_ASAP7_75t_L g2238 ( 
.A(n_2013),
.Y(n_2238)
);

CKINVDCx16_ASAP7_75t_R g2239 ( 
.A(n_2029),
.Y(n_2239)
);

NOR2xp33_ASAP7_75t_SL g2240 ( 
.A(n_2028),
.B(n_1785),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_2071),
.Y(n_2241)
);

NAND2x1p5_ASAP7_75t_L g2242 ( 
.A(n_2082),
.B(n_1922),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_2203),
.B(n_1669),
.Y(n_2243)
);

INVx5_ASAP7_75t_L g2244 ( 
.A(n_1970),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2085),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_2191),
.B(n_1927),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2177),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_1973),
.B(n_1816),
.Y(n_2248)
);

OR2x2_ASAP7_75t_L g2249 ( 
.A(n_2032),
.B(n_1929),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2107),
.Y(n_2250)
);

AND2x4_ASAP7_75t_L g2251 ( 
.A(n_2046),
.B(n_1847),
.Y(n_2251)
);

INVx3_ASAP7_75t_L g2252 ( 
.A(n_2058),
.Y(n_2252)
);

NOR2x1_ASAP7_75t_L g2253 ( 
.A(n_2153),
.B(n_1959),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_2072),
.Y(n_2254)
);

BUFx12f_ASAP7_75t_L g2255 ( 
.A(n_2049),
.Y(n_2255)
);

OR2x2_ASAP7_75t_L g2256 ( 
.A(n_2128),
.B(n_1854),
.Y(n_2256)
);

AND2x6_ASAP7_75t_L g2257 ( 
.A(n_2150),
.B(n_1890),
.Y(n_2257)
);

INVx3_ASAP7_75t_L g2258 ( 
.A(n_2104),
.Y(n_2258)
);

BUFx6f_ASAP7_75t_L g2259 ( 
.A(n_2104),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2076),
.Y(n_2260)
);

NOR2xp33_ASAP7_75t_L g2261 ( 
.A(n_2014),
.B(n_1960),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2107),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2111),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2111),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2024),
.B(n_1817),
.Y(n_2265)
);

NOR2xp33_ASAP7_75t_L g2266 ( 
.A(n_1995),
.B(n_1792),
.Y(n_2266)
);

CKINVDCx5p33_ASAP7_75t_R g2267 ( 
.A(n_2068),
.Y(n_2267)
);

OR2x6_ASAP7_75t_L g2268 ( 
.A(n_2109),
.B(n_1892),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2026),
.B(n_1951),
.Y(n_2269)
);

BUFx12f_ASAP7_75t_L g2270 ( 
.A(n_1969),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2204),
.B(n_1916),
.Y(n_2271)
);

BUFx6f_ASAP7_75t_L g2272 ( 
.A(n_2165),
.Y(n_2272)
);

BUFx3_ASAP7_75t_L g2273 ( 
.A(n_2145),
.Y(n_2273)
);

OR2x6_ASAP7_75t_L g2274 ( 
.A(n_2038),
.B(n_1734),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_1962),
.Y(n_2275)
);

NAND2x1p5_ASAP7_75t_L g2276 ( 
.A(n_2153),
.B(n_1828),
.Y(n_2276)
);

OR2x2_ASAP7_75t_L g2277 ( 
.A(n_2079),
.B(n_1931),
.Y(n_2277)
);

INVx5_ASAP7_75t_L g2278 ( 
.A(n_2208),
.Y(n_2278)
);

AND2x4_ASAP7_75t_L g2279 ( 
.A(n_2140),
.B(n_1849),
.Y(n_2279)
);

NOR2xp33_ASAP7_75t_SL g2280 ( 
.A(n_2121),
.B(n_1841),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_1967),
.B(n_1955),
.Y(n_2281)
);

HB1xp67_ASAP7_75t_L g2282 ( 
.A(n_2002),
.Y(n_2282)
);

AND2x6_ASAP7_75t_L g2283 ( 
.A(n_2181),
.B(n_1891),
.Y(n_2283)
);

HB1xp67_ASAP7_75t_L g2284 ( 
.A(n_2033),
.Y(n_2284)
);

BUFx12f_ASAP7_75t_L g2285 ( 
.A(n_2027),
.Y(n_2285)
);

AND2x2_ASAP7_75t_SL g2286 ( 
.A(n_2122),
.B(n_1872),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1962),
.Y(n_2287)
);

BUFx4f_ASAP7_75t_L g2288 ( 
.A(n_2208),
.Y(n_2288)
);

BUFx6f_ASAP7_75t_L g2289 ( 
.A(n_2165),
.Y(n_2289)
);

INVx4_ASAP7_75t_L g2290 ( 
.A(n_2165),
.Y(n_2290)
);

NAND2x1p5_ASAP7_75t_L g2291 ( 
.A(n_2171),
.B(n_1822),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2086),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_2152),
.B(n_1683),
.Y(n_2293)
);

AND2x4_ASAP7_75t_L g2294 ( 
.A(n_2182),
.B(n_1831),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_2093),
.Y(n_2295)
);

OR2x6_ASAP7_75t_L g2296 ( 
.A(n_2038),
.B(n_1906),
.Y(n_2296)
);

NOR2x1_ASAP7_75t_L g2297 ( 
.A(n_2186),
.B(n_1918),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_2101),
.Y(n_2298)
);

OR2x6_ASAP7_75t_L g2299 ( 
.A(n_2065),
.B(n_1894),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_1982),
.B(n_1941),
.Y(n_2300)
);

AND2x4_ASAP7_75t_L g2301 ( 
.A(n_2175),
.B(n_1881),
.Y(n_2301)
);

OR2x2_ASAP7_75t_L g2302 ( 
.A(n_2020),
.B(n_1727),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_1982),
.B(n_1895),
.Y(n_2303)
);

INVxp67_ASAP7_75t_SL g2304 ( 
.A(n_2065),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_2051),
.B(n_1707),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_1964),
.Y(n_2306)
);

AND2x6_ASAP7_75t_L g2307 ( 
.A(n_2181),
.B(n_1681),
.Y(n_2307)
);

OR2x2_ASAP7_75t_L g2308 ( 
.A(n_2036),
.B(n_1742),
.Y(n_2308)
);

CKINVDCx20_ASAP7_75t_R g2309 ( 
.A(n_2147),
.Y(n_2309)
);

NOR2xp67_ASAP7_75t_L g2310 ( 
.A(n_2025),
.B(n_1677),
.Y(n_2310)
);

OR2x6_ASAP7_75t_SL g2311 ( 
.A(n_2100),
.B(n_1948),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_1982),
.B(n_1678),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_1982),
.B(n_1638),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2135),
.B(n_1925),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2110),
.Y(n_2315)
);

BUFx4f_ASAP7_75t_L g2316 ( 
.A(n_2208),
.Y(n_2316)
);

NOR2xp33_ASAP7_75t_L g2317 ( 
.A(n_2037),
.B(n_1643),
.Y(n_2317)
);

INVx4_ASAP7_75t_L g2318 ( 
.A(n_2171),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2098),
.B(n_1684),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_1964),
.Y(n_2320)
);

INVx3_ASAP7_75t_L g2321 ( 
.A(n_2010),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2115),
.Y(n_2322)
);

AND2x4_ASAP7_75t_L g2323 ( 
.A(n_2176),
.B(n_1825),
.Y(n_2323)
);

AND2x4_ASAP7_75t_L g2324 ( 
.A(n_2178),
.B(n_1826),
.Y(n_2324)
);

NOR2xp33_ASAP7_75t_L g2325 ( 
.A(n_2001),
.B(n_1859),
.Y(n_2325)
);

AND2x4_ASAP7_75t_L g2326 ( 
.A(n_2186),
.B(n_1803),
.Y(n_2326)
);

BUFx3_ASAP7_75t_L g2327 ( 
.A(n_2171),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_2131),
.B(n_1706),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_1974),
.Y(n_2329)
);

AND2x4_ASAP7_75t_L g2330 ( 
.A(n_2207),
.B(n_1805),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_2151),
.B(n_1739),
.Y(n_2331)
);

INVx6_ASAP7_75t_L g2332 ( 
.A(n_2163),
.Y(n_2332)
);

AND2x4_ASAP7_75t_L g2333 ( 
.A(n_2207),
.B(n_1806),
.Y(n_2333)
);

BUFx6f_ASAP7_75t_L g2334 ( 
.A(n_2010),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_1974),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_2119),
.Y(n_2336)
);

AND2x2_ASAP7_75t_SL g2337 ( 
.A(n_1985),
.B(n_1714),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_2183),
.B(n_1838),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2006),
.B(n_1950),
.Y(n_2339)
);

BUFx3_ASAP7_75t_L g2340 ( 
.A(n_2010),
.Y(n_2340)
);

AND2x4_ASAP7_75t_L g2341 ( 
.A(n_2129),
.B(n_1809),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2055),
.B(n_1898),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_1976),
.B(n_1810),
.Y(n_2343)
);

HB1xp67_ASAP7_75t_L g2344 ( 
.A(n_2195),
.Y(n_2344)
);

OR2x2_ASAP7_75t_L g2345 ( 
.A(n_2044),
.B(n_1761),
.Y(n_2345)
);

INVx4_ASAP7_75t_L g2346 ( 
.A(n_2011),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_1976),
.B(n_1811),
.Y(n_2347)
);

AND2x4_ASAP7_75t_L g2348 ( 
.A(n_1992),
.B(n_1812),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_1979),
.B(n_1983),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_2125),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_1979),
.Y(n_2351)
);

INVx3_ASAP7_75t_L g2352 ( 
.A(n_2011),
.Y(n_2352)
);

BUFx4_ASAP7_75t_SL g2353 ( 
.A(n_2202),
.Y(n_2353)
);

INVx2_ASAP7_75t_SL g2354 ( 
.A(n_2009),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_1966),
.B(n_1764),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_1983),
.B(n_1815),
.Y(n_2356)
);

INVxp67_ASAP7_75t_L g2357 ( 
.A(n_2157),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_SL g2358 ( 
.A(n_2009),
.B(n_1861),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2047),
.B(n_1840),
.Y(n_2359)
);

INVx1_ASAP7_75t_SL g2360 ( 
.A(n_2120),
.Y(n_2360)
);

OR2x2_ASAP7_75t_L g2361 ( 
.A(n_1996),
.B(n_1641),
.Y(n_2361)
);

INVxp67_ASAP7_75t_SL g2362 ( 
.A(n_2195),
.Y(n_2362)
);

INVx3_ASAP7_75t_L g2363 ( 
.A(n_2011),
.Y(n_2363)
);

OR2x2_ASAP7_75t_L g2364 ( 
.A(n_1972),
.B(n_1814),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_1987),
.B(n_1818),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_1987),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_1989),
.B(n_1834),
.Y(n_2367)
);

OR2x2_ASAP7_75t_L g2368 ( 
.A(n_2084),
.B(n_1642),
.Y(n_2368)
);

NOR2xp33_ASAP7_75t_L g2369 ( 
.A(n_1978),
.B(n_1920),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_1989),
.B(n_1721),
.Y(n_2370)
);

OR2x2_ASAP7_75t_L g2371 ( 
.A(n_2226),
.B(n_2089),
.Y(n_2371)
);

INVx4_ASAP7_75t_L g2372 ( 
.A(n_2244),
.Y(n_2372)
);

INVx5_ASAP7_75t_SL g2373 ( 
.A(n_2224),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_2362),
.B(n_2083),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2234),
.Y(n_2375)
);

BUFx6f_ASAP7_75t_L g2376 ( 
.A(n_2211),
.Y(n_2376)
);

INVx1_ASAP7_75t_SL g2377 ( 
.A(n_2218),
.Y(n_2377)
);

INVx2_ASAP7_75t_SL g2378 ( 
.A(n_2244),
.Y(n_2378)
);

BUFx6f_ASAP7_75t_SL g2379 ( 
.A(n_2235),
.Y(n_2379)
);

BUFx6f_ASAP7_75t_L g2380 ( 
.A(n_2223),
.Y(n_2380)
);

HB1xp67_ASAP7_75t_L g2381 ( 
.A(n_2353),
.Y(n_2381)
);

OR2x2_ASAP7_75t_L g2382 ( 
.A(n_2308),
.B(n_2094),
.Y(n_2382)
);

INVx5_ASAP7_75t_L g2383 ( 
.A(n_2255),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2369),
.B(n_2087),
.Y(n_2384)
);

BUFx3_ASAP7_75t_L g2385 ( 
.A(n_2220),
.Y(n_2385)
);

BUFx6f_ASAP7_75t_L g2386 ( 
.A(n_2223),
.Y(n_2386)
);

AND2x4_ASAP7_75t_L g2387 ( 
.A(n_2278),
.B(n_2124),
.Y(n_2387)
);

AOI22xp5_ASAP7_75t_L g2388 ( 
.A1(n_2280),
.A2(n_2136),
.B1(n_2172),
.B2(n_2139),
.Y(n_2388)
);

INVx1_ASAP7_75t_SL g2389 ( 
.A(n_2273),
.Y(n_2389)
);

BUFx4_ASAP7_75t_SL g2390 ( 
.A(n_2238),
.Y(n_2390)
);

INVx4_ASAP7_75t_L g2391 ( 
.A(n_2278),
.Y(n_2391)
);

INVx2_ASAP7_75t_SL g2392 ( 
.A(n_2288),
.Y(n_2392)
);

BUFx6f_ASAP7_75t_L g2393 ( 
.A(n_2316),
.Y(n_2393)
);

BUFx12f_ASAP7_75t_L g2394 ( 
.A(n_2332),
.Y(n_2394)
);

BUFx8_ASAP7_75t_SL g2395 ( 
.A(n_2270),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2245),
.Y(n_2396)
);

INVxp67_ASAP7_75t_SL g2397 ( 
.A(n_2304),
.Y(n_2397)
);

BUFx2_ASAP7_75t_L g2398 ( 
.A(n_2299),
.Y(n_2398)
);

BUFx2_ASAP7_75t_L g2399 ( 
.A(n_2239),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2250),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2262),
.Y(n_2401)
);

BUFx3_ASAP7_75t_L g2402 ( 
.A(n_2252),
.Y(n_2402)
);

INVx4_ASAP7_75t_L g2403 ( 
.A(n_2332),
.Y(n_2403)
);

INVx1_ASAP7_75t_SL g2404 ( 
.A(n_2214),
.Y(n_2404)
);

INVx4_ASAP7_75t_L g2405 ( 
.A(n_2285),
.Y(n_2405)
);

BUFx4_ASAP7_75t_SL g2406 ( 
.A(n_2267),
.Y(n_2406)
);

INVx4_ASAP7_75t_L g2407 ( 
.A(n_2251),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2261),
.B(n_2088),
.Y(n_2408)
);

BUFx6f_ASAP7_75t_L g2409 ( 
.A(n_2272),
.Y(n_2409)
);

BUFx5_ASAP7_75t_L g2410 ( 
.A(n_2263),
.Y(n_2410)
);

BUFx5_ASAP7_75t_L g2411 ( 
.A(n_2264),
.Y(n_2411)
);

CKINVDCx16_ASAP7_75t_R g2412 ( 
.A(n_2309),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2217),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2275),
.Y(n_2414)
);

CKINVDCx5p33_ASAP7_75t_R g2415 ( 
.A(n_2354),
.Y(n_2415)
);

BUFx6f_ASAP7_75t_L g2416 ( 
.A(n_2272),
.Y(n_2416)
);

BUFx2_ASAP7_75t_L g2417 ( 
.A(n_2299),
.Y(n_2417)
);

BUFx6f_ASAP7_75t_SL g2418 ( 
.A(n_2212),
.Y(n_2418)
);

INVx6_ASAP7_75t_L g2419 ( 
.A(n_2341),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2287),
.Y(n_2420)
);

INVxp67_ASAP7_75t_SL g2421 ( 
.A(n_2209),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2222),
.B(n_2206),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_2266),
.B(n_2095),
.Y(n_2423)
);

INVx5_ASAP7_75t_SL g2424 ( 
.A(n_2274),
.Y(n_2424)
);

BUFx10_ASAP7_75t_L g2425 ( 
.A(n_2294),
.Y(n_2425)
);

INVxp67_ASAP7_75t_SL g2426 ( 
.A(n_2344),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2306),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2320),
.Y(n_2428)
);

CKINVDCx20_ASAP7_75t_R g2429 ( 
.A(n_2282),
.Y(n_2429)
);

INVx1_ASAP7_75t_SL g2430 ( 
.A(n_2360),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_2231),
.Y(n_2431)
);

CKINVDCx20_ASAP7_75t_R g2432 ( 
.A(n_2284),
.Y(n_2432)
);

BUFx2_ASAP7_75t_SL g2433 ( 
.A(n_2233),
.Y(n_2433)
);

BUFx8_ASAP7_75t_L g2434 ( 
.A(n_2249),
.Y(n_2434)
);

BUFx6f_ASAP7_75t_L g2435 ( 
.A(n_2289),
.Y(n_2435)
);

INVx5_ASAP7_75t_L g2436 ( 
.A(n_2233),
.Y(n_2436)
);

INVx4_ASAP7_75t_L g2437 ( 
.A(n_2289),
.Y(n_2437)
);

NAND2x1p5_ASAP7_75t_L g2438 ( 
.A(n_2327),
.B(n_2039),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2241),
.Y(n_2439)
);

INVx1_ASAP7_75t_SL g2440 ( 
.A(n_2243),
.Y(n_2440)
);

INVx2_ASAP7_75t_SL g2441 ( 
.A(n_2213),
.Y(n_2441)
);

AOI22xp33_ASAP7_75t_L g2442 ( 
.A1(n_2219),
.A2(n_2163),
.B1(n_2116),
.B2(n_2113),
.Y(n_2442)
);

BUFx3_ASAP7_75t_L g2443 ( 
.A(n_2229),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2210),
.B(n_2162),
.Y(n_2444)
);

INVx3_ASAP7_75t_L g2445 ( 
.A(n_2227),
.Y(n_2445)
);

INVx2_ASAP7_75t_SL g2446 ( 
.A(n_2301),
.Y(n_2446)
);

BUFx3_ASAP7_75t_L g2447 ( 
.A(n_2236),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2329),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2335),
.Y(n_2449)
);

BUFx2_ASAP7_75t_SL g2450 ( 
.A(n_2233),
.Y(n_2450)
);

NAND2x1p5_ASAP7_75t_L g2451 ( 
.A(n_2290),
.B(n_2039),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2254),
.Y(n_2452)
);

BUFx2_ASAP7_75t_SL g2453 ( 
.A(n_2257),
.Y(n_2453)
);

INVx1_ASAP7_75t_SL g2454 ( 
.A(n_2277),
.Y(n_2454)
);

BUFx12f_ASAP7_75t_L g2455 ( 
.A(n_2268),
.Y(n_2455)
);

BUFx2_ASAP7_75t_L g2456 ( 
.A(n_2268),
.Y(n_2456)
);

BUFx3_ASAP7_75t_L g2457 ( 
.A(n_2348),
.Y(n_2457)
);

BUFx10_ASAP7_75t_L g2458 ( 
.A(n_2323),
.Y(n_2458)
);

BUFx12f_ASAP7_75t_L g2459 ( 
.A(n_2256),
.Y(n_2459)
);

BUFx3_ASAP7_75t_L g2460 ( 
.A(n_2247),
.Y(n_2460)
);

BUFx2_ASAP7_75t_L g2461 ( 
.A(n_2257),
.Y(n_2461)
);

BUFx6f_ASAP7_75t_L g2462 ( 
.A(n_2227),
.Y(n_2462)
);

INVx2_ASAP7_75t_SL g2463 ( 
.A(n_2253),
.Y(n_2463)
);

INVx3_ASAP7_75t_L g2464 ( 
.A(n_2259),
.Y(n_2464)
);

BUFx3_ASAP7_75t_L g2465 ( 
.A(n_2259),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2232),
.B(n_2015),
.Y(n_2466)
);

NAND2x1p5_ASAP7_75t_L g2467 ( 
.A(n_2318),
.B(n_2039),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2271),
.B(n_2206),
.Y(n_2468)
);

BUFx2_ASAP7_75t_L g2469 ( 
.A(n_2274),
.Y(n_2469)
);

NOR2xp33_ASAP7_75t_L g2470 ( 
.A(n_2228),
.B(n_2077),
.Y(n_2470)
);

INVx3_ASAP7_75t_L g2471 ( 
.A(n_2340),
.Y(n_2471)
);

INVx3_ASAP7_75t_L g2472 ( 
.A(n_2334),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2351),
.Y(n_2473)
);

INVx5_ASAP7_75t_L g2474 ( 
.A(n_2257),
.Y(n_2474)
);

BUFx3_ASAP7_75t_L g2475 ( 
.A(n_2324),
.Y(n_2475)
);

BUFx2_ASAP7_75t_R g2476 ( 
.A(n_2311),
.Y(n_2476)
);

BUFx2_ASAP7_75t_L g2477 ( 
.A(n_2429),
.Y(n_2477)
);

INVx3_ASAP7_75t_SL g2478 ( 
.A(n_2383),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2375),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2413),
.Y(n_2480)
);

AOI22xp5_ASAP7_75t_L g2481 ( 
.A1(n_2388),
.A2(n_2325),
.B1(n_2240),
.B2(n_2337),
.Y(n_2481)
);

HB1xp67_ASAP7_75t_L g2482 ( 
.A(n_2460),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2470),
.B(n_2454),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2396),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2400),
.Y(n_2485)
);

INVx6_ASAP7_75t_L g2486 ( 
.A(n_2394),
.Y(n_2486)
);

AOI22xp33_ASAP7_75t_SL g2487 ( 
.A1(n_2423),
.A2(n_1685),
.B1(n_2317),
.B2(n_2338),
.Y(n_2487)
);

AOI22xp33_ASAP7_75t_L g2488 ( 
.A1(n_2384),
.A2(n_2302),
.B1(n_2296),
.B2(n_2293),
.Y(n_2488)
);

OAI22xp5_ASAP7_75t_L g2489 ( 
.A1(n_2408),
.A2(n_2296),
.B1(n_2339),
.B2(n_2349),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2401),
.Y(n_2490)
);

INVx8_ASAP7_75t_L g2491 ( 
.A(n_2379),
.Y(n_2491)
);

INVx4_ASAP7_75t_L g2492 ( 
.A(n_2393),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2414),
.Y(n_2493)
);

BUFx2_ASAP7_75t_L g2494 ( 
.A(n_2432),
.Y(n_2494)
);

BUFx3_ASAP7_75t_L g2495 ( 
.A(n_2393),
.Y(n_2495)
);

AOI22xp33_ASAP7_75t_SL g2496 ( 
.A1(n_2404),
.A2(n_2286),
.B1(n_2342),
.B2(n_2368),
.Y(n_2496)
);

INVx5_ASAP7_75t_L g2497 ( 
.A(n_2436),
.Y(n_2497)
);

AOI22xp5_ASAP7_75t_SL g2498 ( 
.A1(n_2476),
.A2(n_1798),
.B1(n_1791),
.B2(n_1829),
.Y(n_2498)
);

CKINVDCx20_ASAP7_75t_R g2499 ( 
.A(n_2395),
.Y(n_2499)
);

BUFx2_ASAP7_75t_L g2500 ( 
.A(n_2407),
.Y(n_2500)
);

BUFx8_ASAP7_75t_SL g2501 ( 
.A(n_2385),
.Y(n_2501)
);

AOI22xp33_ASAP7_75t_L g2502 ( 
.A1(n_2440),
.A2(n_2342),
.B1(n_2345),
.B2(n_2355),
.Y(n_2502)
);

OAI22xp33_ASAP7_75t_L g2503 ( 
.A1(n_2374),
.A2(n_1897),
.B1(n_2197),
.B2(n_2331),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2420),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_2431),
.Y(n_2505)
);

INVx6_ASAP7_75t_L g2506 ( 
.A(n_2403),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2439),
.Y(n_2507)
);

BUFx2_ASAP7_75t_L g2508 ( 
.A(n_2399),
.Y(n_2508)
);

AOI22xp33_ASAP7_75t_SL g2509 ( 
.A1(n_2459),
.A2(n_2000),
.B1(n_2045),
.B2(n_2364),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2427),
.Y(n_2510)
);

AOI22xp33_ASAP7_75t_SL g2511 ( 
.A1(n_2424),
.A2(n_2030),
.B1(n_2361),
.B2(n_2359),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2452),
.Y(n_2512)
);

BUFx6f_ASAP7_75t_L g2513 ( 
.A(n_2436),
.Y(n_2513)
);

INVxp67_ASAP7_75t_SL g2514 ( 
.A(n_2421),
.Y(n_2514)
);

AOI22xp5_ASAP7_75t_L g2515 ( 
.A1(n_2397),
.A2(n_2197),
.B1(n_1932),
.B2(n_2114),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2428),
.Y(n_2516)
);

AOI22xp33_ASAP7_75t_L g2517 ( 
.A1(n_2382),
.A2(n_2422),
.B1(n_2419),
.B2(n_2468),
.Y(n_2517)
);

AOI22xp33_ASAP7_75t_L g2518 ( 
.A1(n_2382),
.A2(n_2283),
.B1(n_2271),
.B2(n_2108),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2444),
.B(n_2248),
.Y(n_2519)
);

AOI22xp33_ASAP7_75t_SL g2520 ( 
.A1(n_2424),
.A2(n_2283),
.B1(n_1888),
.B2(n_2307),
.Y(n_2520)
);

AOI22xp33_ASAP7_75t_L g2521 ( 
.A1(n_2422),
.A2(n_2283),
.B1(n_2307),
.B2(n_2292),
.Y(n_2521)
);

BUFx3_ASAP7_75t_L g2522 ( 
.A(n_2402),
.Y(n_2522)
);

INVx2_ASAP7_75t_SL g2523 ( 
.A(n_2390),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2448),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2449),
.Y(n_2525)
);

AOI22xp33_ASAP7_75t_L g2526 ( 
.A1(n_2419),
.A2(n_2307),
.B1(n_2295),
.B2(n_2298),
.Y(n_2526)
);

OAI22xp5_ASAP7_75t_L g2527 ( 
.A1(n_2371),
.A2(n_2164),
.B1(n_2170),
.B2(n_2141),
.Y(n_2527)
);

AOI22xp33_ASAP7_75t_L g2528 ( 
.A1(n_2468),
.A2(n_2442),
.B1(n_2371),
.B2(n_2418),
.Y(n_2528)
);

AOI22xp33_ASAP7_75t_SL g2529 ( 
.A1(n_2461),
.A2(n_2126),
.B1(n_1997),
.B2(n_1990),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2473),
.Y(n_2530)
);

INVx4_ASAP7_75t_L g2531 ( 
.A(n_2383),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2426),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2466),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2410),
.Y(n_2534)
);

OAI22xp5_ASAP7_75t_L g2535 ( 
.A1(n_2415),
.A2(n_2149),
.B1(n_2160),
.B2(n_2148),
.Y(n_2535)
);

OAI22xp33_ASAP7_75t_L g2536 ( 
.A1(n_2377),
.A2(n_2198),
.B1(n_2201),
.B2(n_2311),
.Y(n_2536)
);

OAI22xp5_ASAP7_75t_L g2537 ( 
.A1(n_2461),
.A2(n_2161),
.B1(n_2123),
.B2(n_2370),
.Y(n_2537)
);

INVx3_ASAP7_75t_L g2538 ( 
.A(n_2391),
.Y(n_2538)
);

INVxp67_ASAP7_75t_L g2539 ( 
.A(n_2446),
.Y(n_2539)
);

INVx3_ASAP7_75t_L g2540 ( 
.A(n_2474),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2398),
.Y(n_2541)
);

OAI22xp5_ASAP7_75t_L g2542 ( 
.A1(n_2474),
.A2(n_2357),
.B1(n_2366),
.B2(n_2313),
.Y(n_2542)
);

AOI22xp33_ASAP7_75t_L g2543 ( 
.A1(n_2475),
.A2(n_2260),
.B1(n_2322),
.B2(n_2315),
.Y(n_2543)
);

AOI22xp33_ASAP7_75t_L g2544 ( 
.A1(n_2430),
.A2(n_2336),
.B1(n_2350),
.B2(n_1998),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2398),
.Y(n_2545)
);

OAI22xp5_ASAP7_75t_L g2546 ( 
.A1(n_2469),
.A2(n_2312),
.B1(n_2187),
.B2(n_2096),
.Y(n_2546)
);

AOI22xp33_ASAP7_75t_SL g2547 ( 
.A1(n_2433),
.A2(n_1965),
.B1(n_2319),
.B2(n_2137),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_2443),
.B(n_2052),
.Y(n_2548)
);

AOI22xp33_ASAP7_75t_L g2549 ( 
.A1(n_2457),
.A2(n_2215),
.B1(n_2216),
.B2(n_2281),
.Y(n_2549)
);

OAI21xp33_ASAP7_75t_L g2550 ( 
.A1(n_2381),
.A2(n_2130),
.B(n_2106),
.Y(n_2550)
);

BUFx10_ASAP7_75t_L g2551 ( 
.A(n_2376),
.Y(n_2551)
);

AOI22xp33_ASAP7_75t_L g2552 ( 
.A1(n_2434),
.A2(n_2305),
.B1(n_2059),
.B2(n_2117),
.Y(n_2552)
);

CKINVDCx6p67_ASAP7_75t_R g2553 ( 
.A(n_2412),
.Y(n_2553)
);

AOI22xp33_ASAP7_75t_L g2554 ( 
.A1(n_2441),
.A2(n_2305),
.B1(n_2117),
.B2(n_1993),
.Y(n_2554)
);

BUFx12f_ASAP7_75t_L g2555 ( 
.A(n_2376),
.Y(n_2555)
);

CKINVDCx5p33_ASAP7_75t_R g2556 ( 
.A(n_2406),
.Y(n_2556)
);

OAI22xp5_ASAP7_75t_L g2557 ( 
.A1(n_2450),
.A2(n_2096),
.B1(n_2132),
.B2(n_2007),
.Y(n_2557)
);

AND2x4_ASAP7_75t_L g2558 ( 
.A(n_2497),
.B(n_2417),
.Y(n_2558)
);

OR2x2_ASAP7_75t_L g2559 ( 
.A(n_2483),
.B(n_2456),
.Y(n_2559)
);

CKINVDCx8_ASAP7_75t_R g2560 ( 
.A(n_2556),
.Y(n_2560)
);

HB1xp67_ASAP7_75t_L g2561 ( 
.A(n_2482),
.Y(n_2561)
);

AOI22xp33_ASAP7_75t_L g2562 ( 
.A1(n_2487),
.A2(n_2060),
.B1(n_1994),
.B2(n_1999),
.Y(n_2562)
);

AOI22xp33_ASAP7_75t_L g2563 ( 
.A1(n_2511),
.A2(n_2005),
.B1(n_2012),
.B2(n_1991),
.Y(n_2563)
);

AOI22xp5_ASAP7_75t_L g2564 ( 
.A1(n_2481),
.A2(n_1639),
.B1(n_2358),
.B2(n_2075),
.Y(n_2564)
);

OAI22xp5_ASAP7_75t_L g2565 ( 
.A1(n_2515),
.A2(n_2276),
.B1(n_2003),
.B2(n_2023),
.Y(n_2565)
);

OAI22xp5_ASAP7_75t_L g2566 ( 
.A1(n_2536),
.A2(n_2003),
.B1(n_2023),
.B2(n_2007),
.Y(n_2566)
);

AOI22xp33_ASAP7_75t_L g2567 ( 
.A1(n_2496),
.A2(n_2016),
.B1(n_2138),
.B2(n_2133),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2479),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2480),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2519),
.B(n_2533),
.Y(n_2570)
);

AOI22xp33_ASAP7_75t_L g2571 ( 
.A1(n_2529),
.A2(n_2154),
.B1(n_2155),
.B2(n_2146),
.Y(n_2571)
);

AOI22xp33_ASAP7_75t_L g2572 ( 
.A1(n_2502),
.A2(n_2158),
.B1(n_2166),
.B2(n_2156),
.Y(n_2572)
);

AOI22xp33_ASAP7_75t_L g2573 ( 
.A1(n_2509),
.A2(n_2168),
.B1(n_2173),
.B2(n_2167),
.Y(n_2573)
);

AOI222xp33_ASAP7_75t_L g2574 ( 
.A1(n_2535),
.A2(n_2004),
.B1(n_1984),
.B2(n_1977),
.C1(n_2237),
.C2(n_2070),
.Y(n_2574)
);

INVx2_ASAP7_75t_L g2575 ( 
.A(n_2505),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_2514),
.B(n_2517),
.Y(n_2576)
);

BUFx2_ASAP7_75t_L g2577 ( 
.A(n_2508),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_2507),
.Y(n_2578)
);

BUFx4f_ASAP7_75t_L g2579 ( 
.A(n_2486),
.Y(n_2579)
);

AOI22xp33_ASAP7_75t_L g2580 ( 
.A1(n_2518),
.A2(n_2180),
.B1(n_2193),
.B2(n_2192),
.Y(n_2580)
);

BUFx4f_ASAP7_75t_SL g2581 ( 
.A(n_2499),
.Y(n_2581)
);

OAI21xp5_ASAP7_75t_L g2582 ( 
.A1(n_2537),
.A2(n_2489),
.B(n_2527),
.Y(n_2582)
);

NAND2x1p5_ASAP7_75t_L g2583 ( 
.A(n_2497),
.B(n_2417),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2484),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2532),
.B(n_2488),
.Y(n_2585)
);

OAI22xp33_ASAP7_75t_L g2586 ( 
.A1(n_2553),
.A2(n_2265),
.B1(n_2102),
.B2(n_2300),
.Y(n_2586)
);

AOI22xp33_ASAP7_75t_L g2587 ( 
.A1(n_2503),
.A2(n_2205),
.B1(n_2455),
.B2(n_1992),
.Y(n_2587)
);

CKINVDCx5p33_ASAP7_75t_R g2588 ( 
.A(n_2501),
.Y(n_2588)
);

CKINVDCx5p33_ASAP7_75t_R g2589 ( 
.A(n_2555),
.Y(n_2589)
);

BUFx2_ASAP7_75t_L g2590 ( 
.A(n_2500),
.Y(n_2590)
);

NOR2xp33_ASAP7_75t_L g2591 ( 
.A(n_2477),
.B(n_2389),
.Y(n_2591)
);

CKINVDCx8_ASAP7_75t_R g2592 ( 
.A(n_2491),
.Y(n_2592)
);

INVx1_ASAP7_75t_SL g2593 ( 
.A(n_2506),
.Y(n_2593)
);

OAI22xp33_ASAP7_75t_L g2594 ( 
.A1(n_2494),
.A2(n_2328),
.B1(n_2367),
.B2(n_2246),
.Y(n_2594)
);

CKINVDCx5p33_ASAP7_75t_R g2595 ( 
.A(n_2491),
.Y(n_2595)
);

OAI22xp5_ASAP7_75t_L g2596 ( 
.A1(n_2550),
.A2(n_2062),
.B1(n_2073),
.B2(n_2031),
.Y(n_2596)
);

OAI21xp33_ASAP7_75t_L g2597 ( 
.A1(n_2557),
.A2(n_2118),
.B(n_2134),
.Y(n_2597)
);

AND2x2_ASAP7_75t_L g2598 ( 
.A(n_2548),
.B(n_2387),
.Y(n_2598)
);

INVx2_ASAP7_75t_L g2599 ( 
.A(n_2512),
.Y(n_2599)
);

NOR2xp33_ASAP7_75t_L g2600 ( 
.A(n_2486),
.B(n_2458),
.Y(n_2600)
);

INVx5_ASAP7_75t_SL g2601 ( 
.A(n_2513),
.Y(n_2601)
);

AOI22xp33_ASAP7_75t_L g2602 ( 
.A1(n_2552),
.A2(n_2310),
.B1(n_2062),
.B2(n_2073),
.Y(n_2602)
);

AND2x2_ASAP7_75t_L g2603 ( 
.A(n_2541),
.B(n_2465),
.Y(n_2603)
);

NAND3xp33_ASAP7_75t_L g2604 ( 
.A(n_2546),
.B(n_2185),
.C(n_2297),
.Y(n_2604)
);

CKINVDCx20_ASAP7_75t_R g2605 ( 
.A(n_2478),
.Y(n_2605)
);

BUFx2_ASAP7_75t_L g2606 ( 
.A(n_2522),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2485),
.Y(n_2607)
);

CKINVDCx5p33_ASAP7_75t_R g2608 ( 
.A(n_2495),
.Y(n_2608)
);

OAI21xp5_ASAP7_75t_SL g2609 ( 
.A1(n_2547),
.A2(n_2103),
.B(n_2184),
.Y(n_2609)
);

AOI22xp33_ASAP7_75t_L g2610 ( 
.A1(n_2544),
.A2(n_2078),
.B1(n_2031),
.B2(n_2314),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2490),
.Y(n_2611)
);

HB1xp67_ASAP7_75t_L g2612 ( 
.A(n_2545),
.Y(n_2612)
);

AOI22xp33_ASAP7_75t_L g2613 ( 
.A1(n_2528),
.A2(n_2078),
.B1(n_2453),
.B2(n_2144),
.Y(n_2613)
);

OAI22xp5_ASAP7_75t_L g2614 ( 
.A1(n_2554),
.A2(n_2521),
.B1(n_2520),
.B2(n_2542),
.Y(n_2614)
);

OAI222xp33_ASAP7_75t_L g2615 ( 
.A1(n_2498),
.A2(n_2269),
.B1(n_2127),
.B2(n_2303),
.C1(n_2347),
.C2(n_2343),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_2493),
.B(n_2194),
.Y(n_2616)
);

OAI21xp5_ASAP7_75t_SL g2617 ( 
.A1(n_2523),
.A2(n_2200),
.B(n_2199),
.Y(n_2617)
);

AOI22xp5_ASAP7_75t_L g2618 ( 
.A1(n_2506),
.A2(n_2279),
.B1(n_2392),
.B2(n_2447),
.Y(n_2618)
);

AOI22xp33_ASAP7_75t_L g2619 ( 
.A1(n_2549),
.A2(n_2144),
.B1(n_2159),
.B2(n_2143),
.Y(n_2619)
);

AND2x2_ASAP7_75t_SL g2620 ( 
.A(n_2513),
.B(n_2405),
.Y(n_2620)
);

AOI22xp33_ASAP7_75t_L g2621 ( 
.A1(n_2543),
.A2(n_2526),
.B1(n_2159),
.B2(n_2143),
.Y(n_2621)
);

AOI22xp33_ASAP7_75t_L g2622 ( 
.A1(n_2539),
.A2(n_2018),
.B1(n_2021),
.B2(n_2017),
.Y(n_2622)
);

OAI21xp5_ASAP7_75t_SL g2623 ( 
.A1(n_2538),
.A2(n_2378),
.B(n_2189),
.Y(n_2623)
);

AOI22xp33_ASAP7_75t_SL g2624 ( 
.A1(n_2497),
.A2(n_2463),
.B1(n_2410),
.B2(n_2411),
.Y(n_2624)
);

OAI22xp5_ASAP7_75t_L g2625 ( 
.A1(n_2504),
.A2(n_2105),
.B1(n_2099),
.B2(n_2356),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2510),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2516),
.Y(n_2627)
);

CKINVDCx20_ASAP7_75t_R g2628 ( 
.A(n_2551),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2524),
.Y(n_2629)
);

OAI222xp33_ASAP7_75t_L g2630 ( 
.A1(n_2525),
.A2(n_2365),
.B1(n_2221),
.B2(n_2225),
.C1(n_2099),
.C2(n_2105),
.Y(n_2630)
);

BUFx4f_ASAP7_75t_SL g2631 ( 
.A(n_2531),
.Y(n_2631)
);

INVxp67_ASAP7_75t_L g2632 ( 
.A(n_2530),
.Y(n_2632)
);

AOI22xp5_ASAP7_75t_L g2633 ( 
.A1(n_2540),
.A2(n_2326),
.B1(n_2333),
.B2(n_2330),
.Y(n_2633)
);

INVx2_ASAP7_75t_L g2634 ( 
.A(n_2513),
.Y(n_2634)
);

OAI21xp5_ASAP7_75t_L g2635 ( 
.A1(n_2534),
.A2(n_2040),
.B(n_2034),
.Y(n_2635)
);

INVxp67_ASAP7_75t_SL g2636 ( 
.A(n_2540),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_SL g2637 ( 
.A(n_2531),
.B(n_2410),
.Y(n_2637)
);

AOI22xp33_ASAP7_75t_L g2638 ( 
.A1(n_2562),
.A2(n_1988),
.B1(n_2008),
.B2(n_2174),
.Y(n_2638)
);

OAI21xp5_ASAP7_75t_SL g2639 ( 
.A1(n_2582),
.A2(n_2617),
.B(n_2609),
.Y(n_2639)
);

AOI22xp33_ASAP7_75t_L g2640 ( 
.A1(n_2574),
.A2(n_2043),
.B1(n_2174),
.B2(n_2097),
.Y(n_2640)
);

INVx2_ASAP7_75t_L g2641 ( 
.A(n_2607),
.Y(n_2641)
);

AOI22xp33_ASAP7_75t_L g2642 ( 
.A1(n_2563),
.A2(n_1988),
.B1(n_2008),
.B2(n_2188),
.Y(n_2642)
);

AOI22xp33_ASAP7_75t_L g2643 ( 
.A1(n_2573),
.A2(n_2190),
.B1(n_2411),
.B2(n_2410),
.Y(n_2643)
);

AOI22xp33_ASAP7_75t_L g2644 ( 
.A1(n_2614),
.A2(n_2411),
.B1(n_2069),
.B2(n_2425),
.Y(n_2644)
);

OAI211xp5_ASAP7_75t_L g2645 ( 
.A1(n_2617),
.A2(n_2067),
.B(n_2372),
.C(n_2080),
.Y(n_2645)
);

OAI22xp5_ASAP7_75t_L g2646 ( 
.A1(n_2564),
.A2(n_2373),
.B1(n_2034),
.B2(n_2053),
.Y(n_2646)
);

AOI22xp33_ASAP7_75t_L g2647 ( 
.A1(n_2567),
.A2(n_2602),
.B1(n_2566),
.B2(n_2613),
.Y(n_2647)
);

AOI22xp33_ASAP7_75t_L g2648 ( 
.A1(n_2587),
.A2(n_2411),
.B1(n_2069),
.B2(n_2242),
.Y(n_2648)
);

AOI22xp33_ASAP7_75t_L g2649 ( 
.A1(n_2585),
.A2(n_2069),
.B1(n_2230),
.B2(n_2064),
.Y(n_2649)
);

AOI22xp33_ASAP7_75t_L g2650 ( 
.A1(n_2571),
.A2(n_2069),
.B1(n_2064),
.B2(n_2040),
.Y(n_2650)
);

AND2x2_ASAP7_75t_L g2651 ( 
.A(n_2561),
.B(n_2409),
.Y(n_2651)
);

AOI22xp33_ASAP7_75t_L g2652 ( 
.A1(n_2610),
.A2(n_2572),
.B1(n_2586),
.B2(n_2565),
.Y(n_2652)
);

OAI221xp5_ASAP7_75t_L g2653 ( 
.A1(n_2609),
.A2(n_2492),
.B1(n_2291),
.B2(n_2464),
.C(n_2472),
.Y(n_2653)
);

AOI22xp5_ASAP7_75t_L g2654 ( 
.A1(n_2594),
.A2(n_2576),
.B1(n_2596),
.B2(n_2625),
.Y(n_2654)
);

AOI22xp33_ASAP7_75t_L g2655 ( 
.A1(n_2597),
.A2(n_2069),
.B1(n_2057),
.B2(n_2061),
.Y(n_2655)
);

OAI22xp5_ASAP7_75t_L g2656 ( 
.A1(n_2604),
.A2(n_2577),
.B1(n_2623),
.B2(n_2579),
.Y(n_2656)
);

AOI221xp5_ASAP7_75t_L g2657 ( 
.A1(n_2615),
.A2(n_2471),
.B1(n_2445),
.B2(n_2492),
.C(n_2386),
.Y(n_2657)
);

AOI22xp33_ASAP7_75t_L g2658 ( 
.A1(n_2569),
.A2(n_2057),
.B1(n_2061),
.B2(n_2053),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2570),
.B(n_2632),
.Y(n_2659)
);

OAI22xp33_ASAP7_75t_L g2660 ( 
.A1(n_2616),
.A2(n_2416),
.B1(n_2435),
.B2(n_2409),
.Y(n_2660)
);

AOI22xp33_ASAP7_75t_L g2661 ( 
.A1(n_2575),
.A2(n_2258),
.B1(n_2090),
.B2(n_2074),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2629),
.B(n_2373),
.Y(n_2662)
);

AND2x2_ASAP7_75t_SL g2663 ( 
.A(n_2620),
.B(n_2334),
.Y(n_2663)
);

AOI22xp33_ASAP7_75t_SL g2664 ( 
.A1(n_2604),
.A2(n_2603),
.B1(n_2558),
.B2(n_2583),
.Y(n_2664)
);

AOI22xp5_ASAP7_75t_L g2665 ( 
.A1(n_2633),
.A2(n_2090),
.B1(n_2074),
.B2(n_2380),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_2612),
.B(n_2416),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2568),
.B(n_2584),
.Y(n_2667)
);

OAI22xp5_ASAP7_75t_L g2668 ( 
.A1(n_2579),
.A2(n_2352),
.B1(n_2363),
.B2(n_2321),
.Y(n_2668)
);

AOI22xp33_ASAP7_75t_L g2669 ( 
.A1(n_2578),
.A2(n_2042),
.B1(n_2091),
.B2(n_2050),
.Y(n_2669)
);

AOI22xp33_ASAP7_75t_SL g2670 ( 
.A1(n_2558),
.A2(n_2386),
.B1(n_2380),
.B2(n_2435),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_L g2671 ( 
.A(n_2611),
.B(n_2462),
.Y(n_2671)
);

OAI22xp33_ASAP7_75t_L g2672 ( 
.A1(n_2559),
.A2(n_2462),
.B1(n_2437),
.B2(n_2050),
.Y(n_2672)
);

AOI22xp33_ASAP7_75t_L g2673 ( 
.A1(n_2599),
.A2(n_2042),
.B1(n_2091),
.B2(n_2050),
.Y(n_2673)
);

OAI22xp5_ASAP7_75t_L g2674 ( 
.A1(n_2590),
.A2(n_2438),
.B1(n_2467),
.B2(n_2451),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2626),
.B(n_2551),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2627),
.Y(n_2676)
);

AOI22xp33_ASAP7_75t_L g2677 ( 
.A1(n_2621),
.A2(n_2580),
.B1(n_2619),
.B2(n_2622),
.Y(n_2677)
);

NAND3xp33_ASAP7_75t_L g2678 ( 
.A(n_2591),
.B(n_2091),
.C(n_2042),
.Y(n_2678)
);

OAI222xp33_ASAP7_75t_L g2679 ( 
.A1(n_2618),
.A2(n_1666),
.B1(n_2346),
.B2(n_211),
.C1(n_212),
.C2(n_214),
.Y(n_2679)
);

AOI22xp33_ASAP7_75t_L g2680 ( 
.A1(n_2598),
.A2(n_2092),
.B1(n_212),
.B2(n_209),
.Y(n_2680)
);

OAI22xp5_ASAP7_75t_L g2681 ( 
.A1(n_2606),
.A2(n_2636),
.B1(n_2628),
.B2(n_2631),
.Y(n_2681)
);

OAI22xp5_ASAP7_75t_L g2682 ( 
.A1(n_2605),
.A2(n_2092),
.B1(n_215),
.B2(n_210),
.Y(n_2682)
);

AOI221xp5_ASAP7_75t_L g2683 ( 
.A1(n_2630),
.A2(n_2092),
.B1(n_215),
.B2(n_217),
.C(n_219),
.Y(n_2683)
);

AOI22xp33_ASAP7_75t_L g2684 ( 
.A1(n_2634),
.A2(n_221),
.B1(n_214),
.B2(n_220),
.Y(n_2684)
);

AOI22xp33_ASAP7_75t_L g2685 ( 
.A1(n_2600),
.A2(n_225),
.B1(n_220),
.B2(n_224),
.Y(n_2685)
);

AOI22xp33_ASAP7_75t_L g2686 ( 
.A1(n_2593),
.A2(n_228),
.B1(n_224),
.B2(n_226),
.Y(n_2686)
);

OAI222xp33_ASAP7_75t_L g2687 ( 
.A1(n_2583),
.A2(n_226),
.B1(n_229),
.B2(n_230),
.C1(n_231),
.C2(n_232),
.Y(n_2687)
);

AOI22xp33_ASAP7_75t_L g2688 ( 
.A1(n_2608),
.A2(n_234),
.B1(n_231),
.B2(n_233),
.Y(n_2688)
);

OAI222xp33_ASAP7_75t_L g2689 ( 
.A1(n_2592),
.A2(n_233),
.B1(n_238),
.B2(n_239),
.C1(n_240),
.C2(n_241),
.Y(n_2689)
);

AOI22xp33_ASAP7_75t_L g2690 ( 
.A1(n_2635),
.A2(n_242),
.B1(n_238),
.B2(n_240),
.Y(n_2690)
);

OAI22xp33_ASAP7_75t_SL g2691 ( 
.A1(n_2637),
.A2(n_245),
.B1(n_242),
.B2(n_244),
.Y(n_2691)
);

OAI22xp5_ASAP7_75t_L g2692 ( 
.A1(n_2601),
.A2(n_248),
.B1(n_245),
.B2(n_246),
.Y(n_2692)
);

OAI22xp5_ASAP7_75t_L g2693 ( 
.A1(n_2601),
.A2(n_251),
.B1(n_248),
.B2(n_250),
.Y(n_2693)
);

AOI221xp5_ASAP7_75t_L g2694 ( 
.A1(n_2589),
.A2(n_250),
.B1(n_253),
.B2(n_254),
.C(n_255),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2624),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2659),
.B(n_2601),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2676),
.B(n_253),
.Y(n_2697)
);

AND2x2_ASAP7_75t_L g2698 ( 
.A(n_2651),
.B(n_2595),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_L g2699 ( 
.A(n_2667),
.B(n_2654),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_L g2700 ( 
.A(n_2666),
.B(n_2639),
.Y(n_2700)
);

AND2x2_ASAP7_75t_L g2701 ( 
.A(n_2681),
.B(n_2588),
.Y(n_2701)
);

AND2x2_ASAP7_75t_L g2702 ( 
.A(n_2675),
.B(n_2560),
.Y(n_2702)
);

NAND3xp33_ASAP7_75t_L g2703 ( 
.A(n_2694),
.B(n_258),
.C(n_259),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2656),
.B(n_2641),
.Y(n_2704)
);

OAI21xp5_ASAP7_75t_SL g2705 ( 
.A1(n_2689),
.A2(n_2581),
.B(n_258),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2671),
.B(n_260),
.Y(n_2706)
);

OAI21xp33_ASAP7_75t_L g2707 ( 
.A1(n_2688),
.A2(n_260),
.B(n_261),
.Y(n_2707)
);

OAI211xp5_ASAP7_75t_L g2708 ( 
.A1(n_2645),
.A2(n_266),
.B(n_264),
.C(n_265),
.Y(n_2708)
);

NAND3xp33_ASAP7_75t_L g2709 ( 
.A(n_2683),
.B(n_264),
.C(n_265),
.Y(n_2709)
);

OAI22xp5_ASAP7_75t_L g2710 ( 
.A1(n_2652),
.A2(n_270),
.B1(n_266),
.B2(n_267),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2664),
.B(n_273),
.Y(n_2711)
);

AOI21xp5_ASAP7_75t_SL g2712 ( 
.A1(n_2646),
.A2(n_273),
.B(n_274),
.Y(n_2712)
);

AND2x2_ASAP7_75t_L g2713 ( 
.A(n_2662),
.B(n_276),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_SL g2714 ( 
.A(n_2660),
.B(n_277),
.Y(n_2714)
);

AND2x2_ASAP7_75t_L g2715 ( 
.A(n_2663),
.B(n_277),
.Y(n_2715)
);

AND2x2_ASAP7_75t_L g2716 ( 
.A(n_2663),
.B(n_278),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2695),
.B(n_280),
.Y(n_2717)
);

NAND4xp25_ASAP7_75t_L g2718 ( 
.A(n_2685),
.B(n_281),
.C(n_282),
.D(n_283),
.Y(n_2718)
);

AND2x2_ASAP7_75t_L g2719 ( 
.A(n_2670),
.B(n_281),
.Y(n_2719)
);

INVxp67_ASAP7_75t_SL g2720 ( 
.A(n_2678),
.Y(n_2720)
);

OA21x2_ASAP7_75t_L g2721 ( 
.A1(n_2644),
.A2(n_284),
.B(n_285),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2660),
.Y(n_2722)
);

NAND3xp33_ASAP7_75t_L g2723 ( 
.A(n_2690),
.B(n_285),
.C(n_287),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_SL g2724 ( 
.A(n_2672),
.B(n_288),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2672),
.B(n_2640),
.Y(n_2725)
);

OAI221xp5_ASAP7_75t_L g2726 ( 
.A1(n_2682),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.C(n_292),
.Y(n_2726)
);

OAI21xp5_ASAP7_75t_SL g2727 ( 
.A1(n_2687),
.A2(n_289),
.B(n_290),
.Y(n_2727)
);

AND2x2_ASAP7_75t_L g2728 ( 
.A(n_2674),
.B(n_2657),
.Y(n_2728)
);

OAI21xp5_ASAP7_75t_SL g2729 ( 
.A1(n_2692),
.A2(n_2693),
.B(n_2686),
.Y(n_2729)
);

NOR2xp33_ASAP7_75t_L g2730 ( 
.A(n_2653),
.B(n_2691),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2669),
.Y(n_2731)
);

INVx2_ASAP7_75t_L g2732 ( 
.A(n_2665),
.Y(n_2732)
);

OAI221xp5_ASAP7_75t_L g2733 ( 
.A1(n_2680),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.C(n_294),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2704),
.Y(n_2734)
);

NOR2xp33_ASAP7_75t_L g2735 ( 
.A(n_2701),
.B(n_2700),
.Y(n_2735)
);

NAND4xp75_ASAP7_75t_L g2736 ( 
.A(n_2714),
.B(n_2679),
.C(n_2640),
.D(n_2684),
.Y(n_2736)
);

OR2x2_ASAP7_75t_L g2737 ( 
.A(n_2699),
.B(n_2647),
.Y(n_2737)
);

AO21x2_ASAP7_75t_L g2738 ( 
.A1(n_2720),
.A2(n_2668),
.B(n_2673),
.Y(n_2738)
);

AND2x4_ASAP7_75t_L g2739 ( 
.A(n_2720),
.B(n_2643),
.Y(n_2739)
);

AND2x2_ASAP7_75t_L g2740 ( 
.A(n_2698),
.B(n_2655),
.Y(n_2740)
);

NAND3xp33_ASAP7_75t_L g2741 ( 
.A(n_2730),
.B(n_2661),
.C(n_2649),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_L g2742 ( 
.A(n_2696),
.B(n_2658),
.Y(n_2742)
);

NAND4xp75_ASAP7_75t_L g2743 ( 
.A(n_2714),
.B(n_2677),
.C(n_2648),
.D(n_2638),
.Y(n_2743)
);

INVxp67_ASAP7_75t_SL g2744 ( 
.A(n_2722),
.Y(n_2744)
);

NAND3xp33_ASAP7_75t_L g2745 ( 
.A(n_2730),
.B(n_2650),
.C(n_2642),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2697),
.Y(n_2746)
);

AOI22xp5_ASAP7_75t_L g2747 ( 
.A1(n_2727),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_2747)
);

AOI22xp5_ASAP7_75t_L g2748 ( 
.A1(n_2705),
.A2(n_295),
.B1(n_297),
.B2(n_298),
.Y(n_2748)
);

AND2x2_ASAP7_75t_L g2749 ( 
.A(n_2702),
.B(n_299),
.Y(n_2749)
);

AOI221xp5_ASAP7_75t_L g2750 ( 
.A1(n_2726),
.A2(n_299),
.B1(n_302),
.B2(n_303),
.C(n_304),
.Y(n_2750)
);

AOI22xp33_ASAP7_75t_L g2751 ( 
.A1(n_2725),
.A2(n_305),
.B1(n_306),
.B2(n_308),
.Y(n_2751)
);

AND2x2_ASAP7_75t_L g2752 ( 
.A(n_2713),
.B(n_305),
.Y(n_2752)
);

BUFx2_ASAP7_75t_L g2753 ( 
.A(n_2706),
.Y(n_2753)
);

AND2x2_ASAP7_75t_L g2754 ( 
.A(n_2715),
.B(n_306),
.Y(n_2754)
);

NAND3xp33_ASAP7_75t_L g2755 ( 
.A(n_2703),
.B(n_308),
.C(n_391),
.Y(n_2755)
);

AND2x2_ASAP7_75t_L g2756 ( 
.A(n_2716),
.B(n_392),
.Y(n_2756)
);

AOI22xp5_ASAP7_75t_L g2757 ( 
.A1(n_2718),
.A2(n_393),
.B1(n_395),
.B2(n_396),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2744),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_L g2759 ( 
.A(n_2746),
.B(n_2717),
.Y(n_2759)
);

INVx2_ASAP7_75t_L g2760 ( 
.A(n_2734),
.Y(n_2760)
);

AND2x2_ASAP7_75t_L g2761 ( 
.A(n_2753),
.B(n_2728),
.Y(n_2761)
);

NAND4xp75_ASAP7_75t_L g2762 ( 
.A(n_2748),
.B(n_2724),
.C(n_2719),
.D(n_2711),
.Y(n_2762)
);

BUFx3_ASAP7_75t_L g2763 ( 
.A(n_2749),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2739),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_2735),
.B(n_2721),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2739),
.Y(n_2766)
);

AND2x2_ASAP7_75t_L g2767 ( 
.A(n_2740),
.B(n_2721),
.Y(n_2767)
);

AND2x2_ASAP7_75t_L g2768 ( 
.A(n_2754),
.B(n_2721),
.Y(n_2768)
);

AOI211xp5_ASAP7_75t_SL g2769 ( 
.A1(n_2747),
.A2(n_2712),
.B(n_2708),
.C(n_2729),
.Y(n_2769)
);

XOR2x1_ASAP7_75t_L g2770 ( 
.A(n_2737),
.B(n_2732),
.Y(n_2770)
);

XNOR2xp5_ASAP7_75t_L g2771 ( 
.A(n_2752),
.B(n_2724),
.Y(n_2771)
);

INVxp67_ASAP7_75t_L g2772 ( 
.A(n_2761),
.Y(n_2772)
);

XOR2x2_ASAP7_75t_L g2773 ( 
.A(n_2771),
.B(n_2748),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2758),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2759),
.Y(n_2775)
);

INVx2_ASAP7_75t_SL g2776 ( 
.A(n_2763),
.Y(n_2776)
);

INVxp67_ASAP7_75t_L g2777 ( 
.A(n_2768),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2759),
.Y(n_2778)
);

AOI22x1_ASAP7_75t_L g2779 ( 
.A1(n_2776),
.A2(n_2769),
.B1(n_2767),
.B2(n_2756),
.Y(n_2779)
);

OA22x2_ASAP7_75t_L g2780 ( 
.A1(n_2772),
.A2(n_2747),
.B1(n_2765),
.B2(n_2766),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2774),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2775),
.Y(n_2782)
);

INVx1_ASAP7_75t_SL g2783 ( 
.A(n_2773),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2778),
.Y(n_2784)
);

XOR2x2_ASAP7_75t_L g2785 ( 
.A(n_2777),
.B(n_2762),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2781),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2782),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2784),
.Y(n_2788)
);

BUFx2_ASAP7_75t_L g2789 ( 
.A(n_2785),
.Y(n_2789)
);

INVx1_ASAP7_75t_SL g2790 ( 
.A(n_2783),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2786),
.Y(n_2791)
);

AOI22xp5_ASAP7_75t_L g2792 ( 
.A1(n_2789),
.A2(n_2780),
.B1(n_2765),
.B2(n_2736),
.Y(n_2792)
);

INVx1_ASAP7_75t_SL g2793 ( 
.A(n_2790),
.Y(n_2793)
);

AOI22xp33_ASAP7_75t_L g2794 ( 
.A1(n_2792),
.A2(n_2779),
.B1(n_2745),
.B2(n_2741),
.Y(n_2794)
);

OAI211xp5_ASAP7_75t_SL g2795 ( 
.A1(n_2793),
.A2(n_2769),
.B(n_2788),
.C(n_2787),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2791),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2793),
.Y(n_2797)
);

AO22x1_ASAP7_75t_L g2798 ( 
.A1(n_2797),
.A2(n_2763),
.B1(n_2779),
.B2(n_2710),
.Y(n_2798)
);

AOI22xp5_ASAP7_75t_L g2799 ( 
.A1(n_2795),
.A2(n_2757),
.B1(n_2743),
.B2(n_2755),
.Y(n_2799)
);

NOR2x1_ASAP7_75t_L g2800 ( 
.A(n_2796),
.B(n_2723),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2794),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2797),
.Y(n_2802)
);

NOR2x1_ASAP7_75t_L g2803 ( 
.A(n_2795),
.B(n_2709),
.Y(n_2803)
);

AOI221xp5_ASAP7_75t_L g2804 ( 
.A1(n_2795),
.A2(n_2750),
.B1(n_2707),
.B2(n_2751),
.C(n_2733),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2802),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2800),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2801),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2803),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_SL g2809 ( 
.A(n_2799),
.B(n_2757),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2804),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2798),
.Y(n_2811)
);

OR3x2_ASAP7_75t_L g2812 ( 
.A(n_2808),
.B(n_2770),
.C(n_2731),
.Y(n_2812)
);

OAI22xp5_ASAP7_75t_L g2813 ( 
.A1(n_2811),
.A2(n_2764),
.B1(n_2742),
.B2(n_2760),
.Y(n_2813)
);

NAND2x1_ASAP7_75t_L g2814 ( 
.A(n_2806),
.B(n_2805),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2807),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2810),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2809),
.Y(n_2817)
);

INVx2_ASAP7_75t_L g2818 ( 
.A(n_2814),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2817),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2816),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2815),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2813),
.Y(n_2822)
);

OR3x2_ASAP7_75t_L g2823 ( 
.A(n_2812),
.B(n_2770),
.C(n_2738),
.Y(n_2823)
);

OAI22xp33_ASAP7_75t_SL g2824 ( 
.A1(n_2814),
.A2(n_2732),
.B1(n_2738),
.B2(n_399),
.Y(n_2824)
);

AOI22xp5_ASAP7_75t_L g2825 ( 
.A1(n_2820),
.A2(n_2819),
.B1(n_2823),
.B2(n_2818),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2822),
.Y(n_2826)
);

NAND4xp75_ASAP7_75t_L g2827 ( 
.A(n_2821),
.B(n_397),
.C(n_398),
.D(n_400),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2824),
.Y(n_2828)
);

AOI22xp5_ASAP7_75t_L g2829 ( 
.A1(n_2820),
.A2(n_401),
.B1(n_406),
.B2(n_409),
.Y(n_2829)
);

NOR2x1_ASAP7_75t_L g2830 ( 
.A(n_2818),
.B(n_415),
.Y(n_2830)
);

INVx3_ASAP7_75t_L g2831 ( 
.A(n_2826),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2825),
.Y(n_2832)
);

HB1xp67_ASAP7_75t_L g2833 ( 
.A(n_2830),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2828),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2827),
.Y(n_2835)
);

AO22x1_ASAP7_75t_L g2836 ( 
.A1(n_2831),
.A2(n_2829),
.B1(n_418),
.B2(n_423),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2836),
.Y(n_2837)
);

AOI22xp5_ASAP7_75t_L g2838 ( 
.A1(n_2837),
.A2(n_2834),
.B1(n_2832),
.B2(n_2833),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2838),
.Y(n_2839)
);

AOI221xp5_ASAP7_75t_L g2840 ( 
.A1(n_2839),
.A2(n_2835),
.B1(n_424),
.B2(n_427),
.C(n_428),
.Y(n_2840)
);

AOI211xp5_ASAP7_75t_L g2841 ( 
.A1(n_2840),
.A2(n_417),
.B(n_432),
.C(n_434),
.Y(n_2841)
);


endmodule