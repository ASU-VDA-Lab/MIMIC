module fake_ariane_2074_n_2073 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2073);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2073;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_177),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_153),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_188),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_165),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_169),
.Y(n_214)
);

INVxp67_ASAP7_75t_SL g215 ( 
.A(n_137),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_70),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_86),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_75),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_38),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_92),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_192),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_24),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_208),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_4),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_5),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_144),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_126),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_22),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_112),
.Y(n_232)
);

INVxp33_ASAP7_75t_R g233 ( 
.A(n_62),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_131),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_15),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_8),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_22),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_76),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_39),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_111),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_167),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_98),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_207),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_33),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_187),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_34),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_182),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_59),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_107),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_29),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_184),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_82),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_110),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_114),
.Y(n_254)
);

BUFx5_ASAP7_75t_L g255 ( 
.A(n_176),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_163),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_189),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_56),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_19),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_37),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_1),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_23),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_2),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_63),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_62),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_118),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_74),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_119),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_51),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_84),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_66),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_172),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_19),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_18),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_83),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_175),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_6),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_156),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_191),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_20),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_43),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_106),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_34),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_69),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_99),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_97),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_75),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_44),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_206),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_133),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_193),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_142),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_31),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_204),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_17),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_54),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_74),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_17),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_101),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_154),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_139),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_85),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_64),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_94),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_161),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_196),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_51),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_198),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_105),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_53),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_55),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_25),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_128),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_160),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_49),
.Y(n_315)
);

BUFx2_ASAP7_75t_SL g316 ( 
.A(n_26),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_140),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_54),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_42),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_141),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_56),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_23),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_27),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_91),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_43),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_9),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_158),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_159),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_162),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g330 ( 
.A(n_8),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_127),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_49),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_14),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_151),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_152),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_38),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_39),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_4),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_11),
.Y(n_339)
);

BUFx10_ASAP7_75t_L g340 ( 
.A(n_77),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_146),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_18),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_10),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_21),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_179),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_37),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_135),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_35),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_41),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_46),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_73),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_3),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_0),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_120),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_72),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_197),
.Y(n_356)
);

CKINVDCx14_ASAP7_75t_R g357 ( 
.A(n_203),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_40),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_195),
.Y(n_359)
);

BUFx8_ASAP7_75t_SL g360 ( 
.A(n_11),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_80),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_1),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_164),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_178),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_63),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_0),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_66),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_199),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_108),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_113),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_15),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_42),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_28),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_117),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_103),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_89),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_3),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_45),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_35),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_81),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_157),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_136),
.Y(n_382)
);

BUFx10_ASAP7_75t_L g383 ( 
.A(n_64),
.Y(n_383)
);

BUFx10_ASAP7_75t_L g384 ( 
.A(n_104),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_20),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_14),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_155),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_26),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_125),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_205),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_173),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_171),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_73),
.Y(n_393)
);

BUFx10_ASAP7_75t_L g394 ( 
.A(n_45),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_57),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_76),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_132),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_201),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_53),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_109),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_129),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_67),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_33),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_69),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_90),
.Y(n_405)
);

BUFx10_ASAP7_75t_L g406 ( 
.A(n_16),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_190),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_47),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_121),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_12),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_31),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_168),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_57),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_150),
.Y(n_414)
);

INVxp33_ASAP7_75t_R g415 ( 
.A(n_71),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_330),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_360),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_352),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_243),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_234),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_245),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_308),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_352),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_355),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_253),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_257),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_389),
.Y(n_427)
);

INVxp33_ASAP7_75t_SL g428 ( 
.A(n_235),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_363),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_405),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_374),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_355),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_217),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_259),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_225),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_219),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_231),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_238),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_236),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_236),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_331),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_340),
.B(n_383),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_239),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_244),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_236),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_250),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_263),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_267),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_278),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_278),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_280),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_340),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_281),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_283),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_278),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_257),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_293),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_260),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_384),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_315),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_340),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_264),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_384),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_298),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_318),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_348),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_384),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_319),
.Y(n_468)
);

BUFx2_ASAP7_75t_L g469 ( 
.A(n_222),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_305),
.B(n_2),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_209),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_209),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_323),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_316),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_386),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_388),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_396),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_336),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_343),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_349),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_247),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_383),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_213),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_282),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_214),
.B(n_5),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_350),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_213),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_345),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_365),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_216),
.B(n_220),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_223),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_357),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_223),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_383),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_221),
.B(n_6),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_379),
.Y(n_496)
);

INVxp33_ASAP7_75t_L g497 ( 
.A(n_393),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_229),
.B(n_7),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_212),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_212),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_402),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_218),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_403),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_218),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_226),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_232),
.B(n_7),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_271),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_271),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_222),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_287),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_287),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_347),
.Y(n_512)
);

INVxp67_ASAP7_75t_SL g513 ( 
.A(n_236),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_332),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_332),
.Y(n_515)
);

INVxp67_ASAP7_75t_SL g516 ( 
.A(n_236),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_347),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_399),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_226),
.Y(n_519)
);

INVxp67_ASAP7_75t_SL g520 ( 
.A(n_265),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_426),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_439),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_416),
.B(n_394),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_426),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_439),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_440),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_513),
.B(n_399),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_426),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_440),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_516),
.B(n_265),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_520),
.B(n_240),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_442),
.B(n_265),
.Y(n_532)
);

INVx6_ASAP7_75t_L g533 ( 
.A(n_426),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_426),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_456),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_456),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_456),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_445),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_456),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_474),
.B(n_211),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_481),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_456),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_442),
.B(n_490),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_445),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_418),
.B(n_265),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_507),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_434),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_434),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_508),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_469),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_469),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_510),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_511),
.Y(n_553)
);

OA21x2_ASAP7_75t_L g554 ( 
.A1(n_485),
.A2(n_241),
.B(n_224),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_514),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_515),
.Y(n_556)
);

CKINVDCx8_ASAP7_75t_R g557 ( 
.A(n_417),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_449),
.B(n_265),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_423),
.B(n_413),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_497),
.B(n_413),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_518),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_509),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_495),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_433),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_435),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_437),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_509),
.B(n_339),
.Y(n_567)
);

AND2x2_ASAP7_75t_SL g568 ( 
.A(n_470),
.B(n_224),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_438),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_424),
.B(n_249),
.Y(n_570)
);

BUFx8_ASAP7_75t_L g571 ( 
.A(n_432),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_443),
.B(n_252),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_446),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_447),
.B(n_256),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_448),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_451),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_453),
.B(n_268),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_454),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_457),
.B(n_299),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_471),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_460),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_465),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_468),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_473),
.B(n_300),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_478),
.B(n_413),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_436),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_479),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_480),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_486),
.B(n_413),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_489),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_496),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_501),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_503),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_498),
.B(n_302),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_506),
.Y(n_595)
);

AND2x2_ASAP7_75t_SL g596 ( 
.A(n_452),
.B(n_241),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_471),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_472),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_449),
.B(n_450),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_450),
.B(n_304),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_455),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_472),
.Y(n_602)
);

AND2x2_ASAP7_75t_SL g603 ( 
.A(n_461),
.B(n_309),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_541),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_543),
.B(n_455),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_598),
.B(n_420),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_598),
.B(n_420),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_522),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_602),
.B(n_422),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_543),
.B(n_459),
.Y(n_610)
);

OAI22xp33_ASAP7_75t_SL g611 ( 
.A1(n_594),
.A2(n_428),
.B1(n_441),
.B2(n_459),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_601),
.B(n_483),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_543),
.B(n_463),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_522),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_543),
.B(n_482),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_601),
.B(n_483),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_525),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_547),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_601),
.B(n_487),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_530),
.Y(n_620)
);

BUFx10_ASAP7_75t_L g621 ( 
.A(n_601),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_601),
.B(n_487),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_525),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_543),
.B(n_463),
.Y(n_624)
);

INVxp67_ASAP7_75t_SL g625 ( 
.A(n_531),
.Y(n_625)
);

BUFx4f_ASAP7_75t_L g626 ( 
.A(n_601),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_567),
.B(n_494),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_526),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_547),
.Y(n_629)
);

BUFx4f_ASAP7_75t_L g630 ( 
.A(n_601),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_602),
.B(n_422),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_526),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_601),
.B(n_491),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_529),
.Y(n_634)
);

AND3x2_ASAP7_75t_L g635 ( 
.A(n_523),
.B(n_411),
.C(n_385),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_563),
.B(n_532),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_558),
.B(n_427),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_529),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_568),
.A2(n_428),
.B1(n_441),
.B2(n_499),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_538),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_596),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_563),
.B(n_467),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_538),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_530),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_558),
.B(n_427),
.Y(n_645)
);

AO22x2_ASAP7_75t_L g646 ( 
.A1(n_567),
.A2(n_415),
.B1(n_233),
.B2(n_362),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_600),
.B(n_430),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_530),
.Y(n_648)
);

INVx5_ASAP7_75t_L g649 ( 
.A(n_524),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_544),
.Y(n_650)
);

INVxp33_ASAP7_75t_L g651 ( 
.A(n_547),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_564),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_544),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_564),
.Y(n_654)
);

XNOR2xp5_ASAP7_75t_L g655 ( 
.A(n_586),
.B(n_444),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_560),
.B(n_532),
.Y(n_656)
);

OAI22xp33_ASAP7_75t_SL g657 ( 
.A1(n_594),
.A2(n_467),
.B1(n_228),
.B2(n_237),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_596),
.Y(n_658)
);

AO22x2_ASAP7_75t_L g659 ( 
.A1(n_567),
.A2(n_211),
.B1(n_290),
.B2(n_309),
.Y(n_659)
);

INVxp33_ASAP7_75t_L g660 ( 
.A(n_548),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_544),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_600),
.B(n_430),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_532),
.B(n_491),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_586),
.Y(n_664)
);

OR2x6_ASAP7_75t_L g665 ( 
.A(n_570),
.B(n_290),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_596),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_564),
.Y(n_667)
);

INVxp67_ASAP7_75t_SL g668 ( 
.A(n_531),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_560),
.B(n_493),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_596),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_597),
.B(n_493),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_544),
.Y(n_672)
);

INVx5_ASAP7_75t_L g673 ( 
.A(n_524),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_564),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_544),
.Y(n_675)
);

AND3x1_ASAP7_75t_L g676 ( 
.A(n_595),
.B(n_406),
.C(n_394),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_595),
.B(n_505),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_544),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_597),
.B(n_505),
.Y(n_679)
);

INVx6_ASAP7_75t_L g680 ( 
.A(n_530),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_548),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_548),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_544),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_568),
.A2(n_502),
.B1(n_504),
.B2(n_500),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_595),
.B(n_519),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_544),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_530),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_564),
.Y(n_688)
);

AO21x2_ASAP7_75t_L g689 ( 
.A1(n_595),
.A2(n_320),
.B(n_313),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_549),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_565),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_549),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_549),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_549),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_560),
.B(n_519),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_524),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_565),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_565),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_597),
.B(n_603),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_597),
.B(n_484),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_565),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_597),
.B(n_488),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_556),
.Y(n_703)
);

INVx4_ASAP7_75t_L g704 ( 
.A(n_575),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_603),
.B(n_512),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_557),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_542),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_603),
.B(n_517),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_568),
.B(n_492),
.Y(n_709)
);

INVx4_ASAP7_75t_L g710 ( 
.A(n_575),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_565),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_575),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_603),
.B(n_599),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_556),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_566),
.B(n_394),
.Y(n_715)
);

OAI22xp33_ASAP7_75t_L g716 ( 
.A1(n_523),
.A2(n_358),
.B1(n_248),
.B2(n_246),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_575),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_568),
.B(n_210),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_542),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_575),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_557),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_562),
.A2(n_246),
.B1(n_366),
.B2(n_367),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_571),
.Y(n_723)
);

NAND3xp33_ASAP7_75t_L g724 ( 
.A(n_575),
.B(n_413),
.C(n_335),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_556),
.Y(n_725)
);

BUFx4f_ASAP7_75t_L g726 ( 
.A(n_554),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_554),
.A2(n_406),
.B1(n_317),
.B2(n_376),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_556),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_575),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_521),
.Y(n_730)
);

NAND2xp33_ASAP7_75t_L g731 ( 
.A(n_599),
.B(n_230),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_575),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_587),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_599),
.B(n_230),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_540),
.B(n_562),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_587),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_587),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_557),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_580),
.B(n_242),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_580),
.B(n_251),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_551),
.B(n_251),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_521),
.Y(n_742)
);

INVx4_ASAP7_75t_L g743 ( 
.A(n_587),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_587),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_587),
.Y(n_745)
);

INVx4_ASAP7_75t_L g746 ( 
.A(n_587),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_521),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_566),
.B(n_406),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_527),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_527),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_566),
.B(n_227),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_587),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_569),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_569),
.Y(n_754)
);

NOR3xp33_ASAP7_75t_L g755 ( 
.A(n_735),
.B(n_610),
.C(n_605),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_625),
.B(n_527),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_618),
.B(n_551),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_668),
.B(n_527),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_626),
.B(n_551),
.Y(n_759)
);

OAI221xp5_ASAP7_75t_L g760 ( 
.A1(n_639),
.A2(n_576),
.B1(n_592),
.B2(n_591),
.C(n_590),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_679),
.B(n_550),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_713),
.A2(n_550),
.B1(n_576),
.B2(n_573),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_626),
.B(n_571),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_618),
.B(n_541),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_677),
.B(n_571),
.Y(n_765)
);

OAI21xp5_ASAP7_75t_L g766 ( 
.A1(n_726),
.A2(n_554),
.B(n_572),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_685),
.B(n_571),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_715),
.B(n_571),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_715),
.B(n_585),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_690),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_748),
.B(n_585),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_626),
.B(n_593),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_630),
.B(n_593),
.Y(n_773)
);

INVxp67_ASAP7_75t_SL g774 ( 
.A(n_620),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_681),
.B(n_419),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_680),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_642),
.B(n_582),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_748),
.B(n_585),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_630),
.B(n_593),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_692),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_641),
.B(n_582),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_681),
.B(n_421),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_641),
.B(n_590),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_630),
.B(n_569),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_692),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_621),
.B(n_569),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_658),
.B(n_591),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_658),
.B(n_592),
.Y(n_788)
);

NAND2x1p5_ASAP7_75t_L g789 ( 
.A(n_666),
.B(n_588),
.Y(n_789)
);

AND2x2_ASAP7_75t_SL g790 ( 
.A(n_676),
.B(n_554),
.Y(n_790)
);

OR2x6_ASAP7_75t_L g791 ( 
.A(n_615),
.B(n_578),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_621),
.B(n_593),
.Y(n_792)
);

A2O1A1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_718),
.A2(n_588),
.B(n_572),
.C(n_577),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_621),
.B(n_588),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_666),
.B(n_588),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_670),
.B(n_578),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_670),
.B(n_578),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_693),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_680),
.Y(n_799)
);

NOR2xp67_ASAP7_75t_SL g800 ( 
.A(n_612),
.B(n_227),
.Y(n_800)
);

INVxp33_ASAP7_75t_L g801 ( 
.A(n_655),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_620),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_647),
.B(n_581),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_620),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_662),
.B(n_581),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_644),
.B(n_581),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_613),
.B(n_574),
.Y(n_807)
);

NAND2x1p5_ASAP7_75t_L g808 ( 
.A(n_644),
.B(n_583),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_624),
.B(n_574),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_663),
.B(n_570),
.Y(n_810)
);

O2A1O1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_636),
.A2(n_577),
.B(n_584),
.C(n_579),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_694),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_680),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_621),
.B(n_254),
.Y(n_814)
);

AOI221xp5_ASAP7_75t_L g815 ( 
.A1(n_716),
.A2(n_408),
.B1(n_366),
.B2(n_367),
.C(n_353),
.Y(n_815)
);

NAND3x1_ASAP7_75t_L g816 ( 
.A(n_709),
.B(n_462),
.C(n_458),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_656),
.B(n_583),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_604),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_699),
.B(n_671),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_644),
.B(n_583),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_656),
.B(n_751),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_627),
.B(n_425),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_751),
.B(n_579),
.Y(n_823)
);

INVx8_ASAP7_75t_L g824 ( 
.A(n_706),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_726),
.B(n_615),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_629),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_648),
.B(n_584),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_SL g828 ( 
.A(n_706),
.B(n_429),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_637),
.B(n_546),
.Y(n_829)
);

INVxp33_ASAP7_75t_L g830 ( 
.A(n_655),
.Y(n_830)
);

BUFx5_ASAP7_75t_L g831 ( 
.A(n_652),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_SL g832 ( 
.A1(n_664),
.A2(n_466),
.B1(n_464),
.B2(n_475),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_680),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_682),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_648),
.B(n_545),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_648),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_726),
.B(n_254),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_687),
.B(n_545),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_687),
.B(n_749),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_687),
.B(n_545),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_627),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_608),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_608),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_652),
.B(n_654),
.Y(n_844)
);

AND2x2_ASAP7_75t_SL g845 ( 
.A(n_676),
.B(n_554),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_749),
.B(n_545),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_749),
.B(n_545),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_614),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_SL g849 ( 
.A(n_721),
.B(n_431),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_614),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_623),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_750),
.B(n_559),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_750),
.B(n_559),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_651),
.B(n_660),
.Y(n_854)
);

OR2x6_ASAP7_75t_L g855 ( 
.A(n_705),
.B(n_546),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_694),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_654),
.B(n_354),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_623),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_645),
.B(n_552),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_750),
.B(n_559),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_700),
.Y(n_861)
);

NAND2xp33_ASAP7_75t_L g862 ( 
.A(n_720),
.B(n_354),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_632),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_606),
.B(n_356),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_703),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_667),
.B(n_356),
.Y(n_866)
);

BUFx3_ASAP7_75t_L g867 ( 
.A(n_721),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_703),
.Y(n_868)
);

AO22x2_ASAP7_75t_L g869 ( 
.A1(n_708),
.A2(n_555),
.B1(n_552),
.B2(n_553),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_667),
.B(n_361),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_669),
.B(n_559),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_632),
.Y(n_872)
);

INVxp67_ASAP7_75t_L g873 ( 
.A(n_702),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_714),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_669),
.B(n_559),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_738),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_720),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_714),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_634),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_674),
.B(n_361),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_738),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_695),
.B(n_589),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_720),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_695),
.Y(n_884)
);

NAND2xp33_ASAP7_75t_L g885 ( 
.A(n_720),
.B(n_364),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_607),
.B(n_589),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_674),
.B(n_364),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_734),
.B(n_553),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_665),
.A2(n_215),
.B1(n_554),
.B2(n_589),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_634),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_720),
.Y(n_891)
);

INVx4_ASAP7_75t_L g892 ( 
.A(n_635),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_609),
.B(n_589),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_631),
.B(n_555),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_611),
.B(n_368),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_725),
.Y(n_896)
);

OR2x6_ASAP7_75t_L g897 ( 
.A(n_646),
.B(n_589),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_638),
.Y(n_898)
);

NAND2xp33_ASAP7_75t_L g899 ( 
.A(n_688),
.B(n_368),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_638),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_665),
.B(n_561),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_665),
.B(n_561),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_665),
.B(n_561),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_665),
.B(n_369),
.Y(n_904)
);

O2A1O1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_616),
.A2(n_375),
.B(n_324),
.C(n_341),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_725),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_659),
.A2(n_371),
.B1(n_344),
.B2(n_346),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_688),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_691),
.B(n_369),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_739),
.B(n_258),
.Y(n_910)
);

A2O1A1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_691),
.A2(n_390),
.B(n_407),
.C(n_228),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_684),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_L g913 ( 
.A1(n_659),
.A2(n_358),
.B1(n_248),
.B2(n_237),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_697),
.B(n_370),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_722),
.B(n_417),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_728),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_697),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_698),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_698),
.B(n_370),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_701),
.B(n_380),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_728),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_617),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_701),
.B(n_380),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_711),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_842),
.Y(n_925)
);

OAI21xp5_ASAP7_75t_L g926 ( 
.A1(n_766),
.A2(n_711),
.B(n_753),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_818),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_843),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_761),
.A2(n_861),
.B(n_873),
.C(n_821),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_844),
.A2(n_622),
.B(n_619),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_831),
.B(n_704),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_831),
.B(n_790),
.Y(n_932)
);

BUFx4f_ASAP7_75t_L g933 ( 
.A(n_824),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_844),
.A2(n_633),
.B(n_712),
.Y(n_934)
);

CKINVDCx10_ASAP7_75t_R g935 ( 
.A(n_832),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_848),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_810),
.B(n_741),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_831),
.B(n_790),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_810),
.B(n_740),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_772),
.A2(n_729),
.B(n_717),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_772),
.A2(n_732),
.B(n_729),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_894),
.B(n_659),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_773),
.A2(n_784),
.B(n_779),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_755),
.A2(n_657),
.B(n_611),
.C(n_731),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_773),
.A2(n_733),
.B(n_732),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_779),
.A2(n_736),
.B(n_733),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_894),
.B(n_659),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_831),
.B(n_704),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_825),
.B(n_657),
.Y(n_949)
);

AO21x1_ASAP7_75t_L g950 ( 
.A1(n_837),
.A2(n_754),
.B(n_753),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_829),
.B(n_723),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_793),
.A2(n_754),
.B(n_737),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_784),
.A2(n_792),
.B(n_786),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_757),
.B(n_646),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_859),
.B(n_727),
.Y(n_955)
);

INVx11_ASAP7_75t_L g956 ( 
.A(n_824),
.Y(n_956)
);

CKINVDCx10_ASAP7_75t_R g957 ( 
.A(n_801),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_850),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_770),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_786),
.A2(n_737),
.B(n_736),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_825),
.A2(n_689),
.B1(n_640),
.B2(n_617),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_859),
.B(n_689),
.Y(n_962)
);

O2A1O1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_807),
.A2(n_707),
.B(n_719),
.C(n_628),
.Y(n_963)
);

BUFx2_ASAP7_75t_L g964 ( 
.A(n_764),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_823),
.B(n_689),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_824),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_804),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_792),
.A2(n_745),
.B(n_744),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_884),
.B(n_707),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_827),
.B(n_640),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_SL g971 ( 
.A(n_828),
.B(n_849),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_769),
.B(n_628),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_794),
.A2(n_745),
.B(n_744),
.Y(n_973)
);

NAND3xp33_ASAP7_75t_SL g974 ( 
.A(n_815),
.B(n_477),
.C(n_476),
.Y(n_974)
);

AOI21x1_ASAP7_75t_L g975 ( 
.A1(n_794),
.A2(n_837),
.B(n_795),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_791),
.A2(n_704),
.B1(n_746),
.B2(n_743),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_851),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_771),
.B(n_643),
.Y(n_978)
);

O2A1O1Ixp5_ASAP7_75t_L g979 ( 
.A1(n_814),
.A2(n_777),
.B(n_800),
.C(n_809),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_819),
.A2(n_752),
.B(n_710),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_803),
.A2(n_752),
.B(n_672),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_804),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_805),
.A2(n_814),
.B(n_817),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_811),
.A2(n_819),
.B(n_908),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_917),
.A2(n_672),
.B(n_650),
.Y(n_985)
);

BUFx4_ASAP7_75t_SL g986 ( 
.A(n_867),
.Y(n_986)
);

BUFx4f_ASAP7_75t_L g987 ( 
.A(n_826),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_918),
.A2(n_672),
.B(n_650),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_924),
.A2(n_672),
.B(n_650),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_804),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_841),
.B(n_646),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_759),
.A2(n_678),
.B(n_650),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_778),
.B(n_643),
.Y(n_993)
);

INVxp67_ASAP7_75t_L g994 ( 
.A(n_854),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_831),
.B(n_704),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_822),
.B(n_646),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_858),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_863),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_872),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_879),
.A2(n_707),
.B1(n_719),
.B2(n_743),
.Y(n_1000)
);

OAI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_922),
.A2(n_743),
.B(n_710),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_759),
.A2(n_678),
.B(n_710),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_871),
.A2(n_707),
.B(n_719),
.C(n_678),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_875),
.A2(n_719),
.B(n_678),
.C(n_696),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_922),
.A2(n_743),
.B(n_710),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_890),
.A2(n_746),
.B(n_661),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_898),
.A2(n_746),
.B(n_661),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_804),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_900),
.A2(n_746),
.B(n_661),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_780),
.A2(n_675),
.B(n_653),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_886),
.A2(n_675),
.B(n_653),
.Y(n_1011)
);

NOR2x1_ASAP7_75t_L g1012 ( 
.A(n_867),
.B(n_724),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_775),
.B(n_344),
.Y(n_1013)
);

OR2x2_ASAP7_75t_L g1014 ( 
.A(n_782),
.B(n_346),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_791),
.B(n_683),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_876),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_756),
.B(n_683),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_876),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_791),
.B(n_686),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_785),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_758),
.B(n_686),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_893),
.A2(n_696),
.B(n_673),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_909),
.A2(n_696),
.B(n_673),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_914),
.A2(n_673),
.B(n_649),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_806),
.B(n_730),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_774),
.A2(n_381),
.B1(n_414),
.B2(n_412),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_802),
.B(n_730),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_882),
.A2(n_747),
.B(n_742),
.C(n_542),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_806),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_802),
.A2(n_353),
.B1(n_351),
.B2(n_371),
.Y(n_1030)
);

INVx1_ASAP7_75t_SL g1031 ( 
.A(n_834),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_820),
.B(n_742),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_785),
.A2(n_747),
.B(n_724),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_839),
.A2(n_351),
.B1(n_372),
.B2(n_373),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_920),
.A2(n_673),
.B(n_649),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_907),
.A2(n_372),
.B(n_373),
.C(n_377),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_798),
.A2(n_673),
.B(n_649),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_781),
.A2(n_787),
.B1(n_788),
.B2(n_783),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_808),
.A2(n_377),
.B1(n_378),
.B2(n_395),
.Y(n_1039)
);

NOR2x1p5_ASAP7_75t_L g1040 ( 
.A(n_881),
.B(n_378),
.Y(n_1040)
);

O2A1O1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_864),
.A2(n_542),
.B(n_535),
.C(n_539),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_798),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_812),
.A2(n_673),
.B(n_649),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_820),
.B(n_395),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_888),
.B(n_404),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_907),
.A2(n_404),
.B1(n_408),
.B2(n_410),
.Y(n_1046)
);

NAND2x1p5_ASAP7_75t_L g1047 ( 
.A(n_881),
.B(n_649),
.Y(n_1047)
);

NOR2xp67_ASAP7_75t_L g1048 ( 
.A(n_892),
.B(n_381),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_856),
.A2(n_649),
.B(n_542),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_856),
.A2(n_537),
.B(n_535),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_865),
.A2(n_537),
.B(n_535),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_776),
.B(n_410),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_865),
.A2(n_537),
.B(n_535),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_913),
.A2(n_312),
.B(n_261),
.C(n_262),
.Y(n_1054)
);

INVx4_ASAP7_75t_L g1055 ( 
.A(n_808),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_799),
.B(n_269),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_913),
.A2(n_321),
.B1(n_310),
.B2(n_273),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_836),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_835),
.Y(n_1059)
);

AND2x2_ASAP7_75t_SL g1060 ( 
.A(n_845),
.B(n_257),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_868),
.Y(n_1061)
);

NOR2xp67_ASAP7_75t_L g1062 ( 
.A(n_892),
.B(n_382),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_813),
.B(n_274),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_888),
.B(n_277),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_831),
.B(n_382),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_874),
.A2(n_539),
.B(n_537),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_874),
.A2(n_539),
.B(n_387),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_762),
.B(n_284),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_878),
.A2(n_539),
.B(n_528),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_912),
.B(n_288),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_845),
.B(n_387),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_878),
.A2(n_391),
.B(n_392),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_833),
.B(n_295),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_768),
.B(n_296),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_765),
.B(n_391),
.Y(n_1075)
);

OAI21xp33_ASAP7_75t_L g1076 ( 
.A1(n_910),
.A2(n_337),
.B(n_297),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_855),
.B(n_904),
.Y(n_1077)
);

NOR2x1_ASAP7_75t_L g1078 ( 
.A(n_855),
.B(n_528),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_896),
.A2(n_392),
.B(n_397),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_846),
.B(n_303),
.Y(n_1080)
);

INVx5_ASAP7_75t_L g1081 ( 
.A(n_877),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_767),
.B(n_397),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_915),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_896),
.Y(n_1084)
);

O2A1O1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_911),
.A2(n_528),
.B(n_338),
.C(n_333),
.Y(n_1085)
);

INVx3_ASAP7_75t_L g1086 ( 
.A(n_877),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_906),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_847),
.B(n_307),
.Y(n_1088)
);

O2A1O1Ixp5_ASAP7_75t_L g1089 ( 
.A1(n_857),
.A2(n_533),
.B(n_398),
.C(n_400),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_852),
.B(n_311),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_877),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_910),
.A2(n_322),
.B(n_325),
.C(n_326),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_855),
.B(n_342),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_906),
.A2(n_398),
.B(n_400),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_760),
.A2(n_414),
.B(n_412),
.C(n_409),
.Y(n_1095)
);

OAI21xp33_ASAP7_75t_L g1096 ( 
.A1(n_857),
.A2(n_409),
.B(n_266),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_889),
.A2(n_257),
.B(n_359),
.C(n_401),
.Y(n_1097)
);

AOI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_899),
.A2(n_294),
.B1(n_270),
.B2(n_285),
.Y(n_1098)
);

O2A1O1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_866),
.A2(n_9),
.B(n_10),
.C(n_12),
.Y(n_1099)
);

BUFx4f_ASAP7_75t_L g1100 ( 
.A(n_877),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_883),
.B(n_891),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_853),
.B(n_272),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_916),
.A2(n_306),
.B(n_275),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_916),
.A2(n_314),
.B(n_276),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_921),
.A2(n_327),
.B(n_279),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_860),
.B(n_286),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_921),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_883),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_964),
.Y(n_1109)
);

INVx6_ASAP7_75t_L g1110 ( 
.A(n_1018),
.Y(n_1110)
);

BUFx12f_ASAP7_75t_L g1111 ( 
.A(n_1016),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_987),
.B(n_1031),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_987),
.B(n_883),
.Y(n_1113)
);

AOI22xp33_ASAP7_75t_L g1114 ( 
.A1(n_974),
.A2(n_897),
.B1(n_830),
.B2(n_869),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_951),
.A2(n_891),
.B(n_763),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_937),
.B(n_869),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_937),
.B(n_869),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_959),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_939),
.A2(n_895),
.B1(n_838),
.B2(n_840),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_1018),
.B(n_891),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_925),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_962),
.A2(n_970),
.B(n_984),
.Y(n_1122)
);

NOR2x1_ASAP7_75t_L g1123 ( 
.A(n_990),
.B(n_1008),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_929),
.B(n_901),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_983),
.A2(n_763),
.B(n_862),
.Y(n_1125)
);

NAND3xp33_ASAP7_75t_L g1126 ( 
.A(n_939),
.B(n_905),
.C(n_919),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_931),
.A2(n_885),
.B(n_919),
.Y(n_1127)
);

BUFx12f_ASAP7_75t_L g1128 ( 
.A(n_966),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_1070),
.B(n_923),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1045),
.B(n_796),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_1077),
.B(n_994),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1059),
.B(n_797),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_955),
.A2(n_923),
.B1(n_866),
.B2(n_870),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_933),
.B(n_971),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_1100),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_931),
.A2(n_870),
.B(n_887),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_928),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1077),
.B(n_1093),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_933),
.B(n_902),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1064),
.B(n_903),
.Y(n_1140)
);

INVx4_ASAP7_75t_L g1141 ( 
.A(n_956),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_1083),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_948),
.A2(n_887),
.B(n_880),
.Y(n_1143)
);

BUFx3_ASAP7_75t_L g1144 ( 
.A(n_927),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_1100),
.B(n_789),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_1093),
.B(n_880),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1046),
.A2(n_789),
.B1(n_897),
.B2(n_816),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_948),
.A2(n_329),
.B(n_289),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_995),
.A2(n_334),
.B(n_291),
.Y(n_1149)
);

HB1xp67_ASAP7_75t_L g1150 ( 
.A(n_986),
.Y(n_1150)
);

BUFx12f_ASAP7_75t_L g1151 ( 
.A(n_1040),
.Y(n_1151)
);

OR2x2_ASAP7_75t_L g1152 ( 
.A(n_1014),
.B(n_897),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_995),
.A2(n_292),
.B(n_301),
.Y(n_1153)
);

AO21x1_ASAP7_75t_L g1154 ( 
.A1(n_965),
.A2(n_255),
.B(n_401),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_1057),
.B(n_328),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_967),
.Y(n_1156)
);

O2A1O1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_1092),
.A2(n_13),
.B(n_16),
.C(n_21),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_942),
.B(n_13),
.Y(n_1158)
);

NAND3xp33_ASAP7_75t_SL g1159 ( 
.A(n_1046),
.B(n_24),
.C(n_25),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_947),
.B(n_27),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_986),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_967),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_926),
.A2(n_255),
.B(n_533),
.Y(n_1163)
);

INVx2_ASAP7_75t_SL g1164 ( 
.A(n_957),
.Y(n_1164)
);

AO32x2_ASAP7_75t_L g1165 ( 
.A1(n_1038),
.A2(n_28),
.A3(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_949),
.A2(n_401),
.B(n_359),
.C(n_257),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_967),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_936),
.B(n_30),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1057),
.B(n_1081),
.Y(n_1169)
);

NOR2x1_ASAP7_75t_SL g1170 ( 
.A(n_1081),
.B(n_401),
.Y(n_1170)
);

AND2x2_ASAP7_75t_SL g1171 ( 
.A(n_1060),
.B(n_359),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_958),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_977),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1060),
.A2(n_359),
.B1(n_533),
.B2(n_40),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_997),
.B(n_32),
.Y(n_1175)
);

AOI22x1_ASAP7_75t_L g1176 ( 
.A1(n_930),
.A2(n_536),
.B1(n_534),
.B2(n_524),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_949),
.A2(n_536),
.B(n_534),
.C(n_524),
.Y(n_1177)
);

CKINVDCx20_ASAP7_75t_R g1178 ( 
.A(n_1013),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_1029),
.B(n_36),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_967),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_972),
.A2(n_536),
.B(n_534),
.Y(n_1181)
);

NAND2x1p5_ASAP7_75t_L g1182 ( 
.A(n_1055),
.B(n_536),
.Y(n_1182)
);

INVx2_ASAP7_75t_SL g1183 ( 
.A(n_935),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_982),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_954),
.B(n_996),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_998),
.A2(n_533),
.B1(n_41),
.B2(n_44),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_999),
.B(n_36),
.Y(n_1187)
);

OA22x2_ASAP7_75t_L g1188 ( 
.A1(n_991),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_1081),
.B(n_982),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_943),
.A2(n_536),
.B(n_534),
.Y(n_1190)
);

BUFx10_ASAP7_75t_L g1191 ( 
.A(n_1052),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1052),
.B(n_48),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1076),
.B(n_1092),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1058),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_982),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_982),
.Y(n_1196)
);

INVxp67_ASAP7_75t_L g1197 ( 
.A(n_1056),
.Y(n_1197)
);

INVx4_ASAP7_75t_L g1198 ( 
.A(n_1081),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_969),
.B(n_50),
.Y(n_1199)
);

INVx6_ASAP7_75t_L g1200 ( 
.A(n_1055),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_969),
.B(n_50),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_944),
.A2(n_52),
.B(n_55),
.C(n_58),
.Y(n_1202)
);

INVx5_ASAP7_75t_L g1203 ( 
.A(n_1091),
.Y(n_1203)
);

A2O1A1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_1095),
.A2(n_536),
.B(n_534),
.C(n_524),
.Y(n_1204)
);

NAND2x1p5_ASAP7_75t_L g1205 ( 
.A(n_990),
.B(n_536),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_R g1206 ( 
.A(n_1008),
.B(n_1086),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1020),
.Y(n_1207)
);

INVxp33_ASAP7_75t_SL g1208 ( 
.A(n_1026),
.Y(n_1208)
);

AOI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1015),
.A2(n_255),
.B1(n_533),
.B2(n_534),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_981),
.A2(n_536),
.B(n_534),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1095),
.A2(n_534),
.B(n_524),
.C(n_255),
.Y(n_1211)
);

INVxp67_ASAP7_75t_SL g1212 ( 
.A(n_1091),
.Y(n_1212)
);

INVx2_ASAP7_75t_SL g1213 ( 
.A(n_1078),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1054),
.A2(n_524),
.B(n_255),
.C(n_59),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1006),
.A2(n_116),
.B(n_145),
.Y(n_1215)
);

INVx2_ASAP7_75t_SL g1216 ( 
.A(n_1047),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1036),
.A2(n_1054),
.B1(n_978),
.B2(n_993),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1036),
.A2(n_533),
.B1(n_58),
.B2(n_60),
.Y(n_1218)
);

INVx1_ASAP7_75t_SL g1219 ( 
.A(n_1091),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1007),
.A2(n_115),
.B(n_200),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1048),
.B(n_52),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1097),
.A2(n_60),
.B1(n_61),
.B2(n_65),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_1091),
.Y(n_1223)
);

NOR3xp33_ASAP7_75t_SL g1224 ( 
.A(n_1030),
.B(n_61),
.C(n_65),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_953),
.A2(n_255),
.B(n_68),
.Y(n_1225)
);

INVx3_ASAP7_75t_L g1226 ( 
.A(n_1047),
.Y(n_1226)
);

INVx4_ASAP7_75t_L g1227 ( 
.A(n_1086),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1074),
.B(n_67),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_1062),
.B(n_255),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1044),
.B(n_68),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_1012),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1042),
.Y(n_1232)
);

OR2x2_ASAP7_75t_L g1233 ( 
.A(n_1034),
.B(n_70),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_SL g1234 ( 
.A(n_1097),
.B(n_255),
.Y(n_1234)
);

AO32x2_ASAP7_75t_L g1235 ( 
.A1(n_1000),
.A2(n_71),
.A3(n_72),
.B1(n_77),
.B2(n_78),
.Y(n_1235)
);

AOI22x1_ASAP7_75t_L g1236 ( 
.A1(n_1009),
.A2(n_1024),
.B1(n_1035),
.B2(n_934),
.Y(n_1236)
);

AOI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1071),
.A2(n_79),
.B(n_87),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1022),
.A2(n_88),
.B(n_93),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1023),
.A2(n_95),
.B(n_96),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1061),
.Y(n_1240)
);

NOR3xp33_ASAP7_75t_L g1241 ( 
.A(n_1099),
.B(n_1096),
.C(n_1039),
.Y(n_1241)
);

INVxp67_ASAP7_75t_SL g1242 ( 
.A(n_1015),
.Y(n_1242)
);

AOI221xp5_ASAP7_75t_L g1243 ( 
.A1(n_1068),
.A2(n_100),
.B1(n_102),
.B2(n_122),
.C(n_123),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1071),
.A2(n_124),
.B1(n_130),
.B2(n_134),
.Y(n_1244)
);

INVx5_ASAP7_75t_L g1245 ( 
.A(n_1108),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1056),
.B(n_138),
.Y(n_1246)
);

O2A1O1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_1080),
.A2(n_143),
.B(n_147),
.C(n_148),
.Y(n_1247)
);

OR2x2_ASAP7_75t_L g1248 ( 
.A(n_1088),
.B(n_149),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1090),
.B(n_166),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_976),
.A2(n_170),
.B1(n_174),
.B2(n_180),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1063),
.B(n_186),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1063),
.B(n_194),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1073),
.B(n_1075),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1017),
.A2(n_1021),
.B1(n_961),
.B2(n_932),
.Y(n_1254)
);

AND2x4_ASAP7_75t_L g1255 ( 
.A(n_1019),
.B(n_1108),
.Y(n_1255)
);

OAI321xp33_ASAP7_75t_L g1256 ( 
.A1(n_952),
.A2(n_1075),
.A3(n_1082),
.B1(n_1085),
.B2(n_980),
.C(n_1073),
.Y(n_1256)
);

NAND3xp33_ASAP7_75t_SL g1257 ( 
.A(n_1098),
.B(n_979),
.C(n_1082),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1102),
.A2(n_1106),
.B1(n_938),
.B2(n_932),
.Y(n_1258)
);

INVxp67_ASAP7_75t_L g1259 ( 
.A(n_1019),
.Y(n_1259)
);

O2A1O1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1003),
.A2(n_938),
.B(n_1004),
.C(n_1065),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1101),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1065),
.B(n_1087),
.Y(n_1262)
);

INVx3_ASAP7_75t_L g1263 ( 
.A(n_1084),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1107),
.B(n_1025),
.Y(n_1264)
);

AO31x2_ASAP7_75t_L g1265 ( 
.A1(n_1154),
.A2(n_950),
.A3(n_1011),
.B(n_1067),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1121),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1109),
.Y(n_1267)
);

O2A1O1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1197),
.A2(n_1028),
.B(n_963),
.C(n_1089),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1254),
.A2(n_1037),
.A3(n_992),
.B(n_945),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1236),
.A2(n_975),
.B(n_941),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1122),
.A2(n_1043),
.B(n_1101),
.Y(n_1271)
);

OA21x2_ASAP7_75t_L g1272 ( 
.A1(n_1225),
.A2(n_1033),
.B(n_1010),
.Y(n_1272)
);

A2O1A1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1193),
.A2(n_1027),
.B(n_1079),
.C(n_1072),
.Y(n_1273)
);

OAI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1208),
.A2(n_1032),
.B1(n_1027),
.B2(n_1005),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_SL g1275 ( 
.A(n_1171),
.B(n_1001),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1203),
.Y(n_1276)
);

BUFx2_ASAP7_75t_L g1277 ( 
.A(n_1178),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1137),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1190),
.A2(n_1210),
.B(n_1176),
.Y(n_1279)
);

AOI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1138),
.A2(n_1094),
.B1(n_1104),
.B2(n_1103),
.Y(n_1280)
);

OAI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1225),
.A2(n_989),
.B(n_988),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_1203),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1181),
.A2(n_940),
.B(n_946),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1174),
.A2(n_1002),
.B1(n_985),
.B2(n_973),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1172),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1163),
.A2(n_960),
.B(n_968),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1258),
.A2(n_1049),
.B(n_1041),
.Y(n_1287)
);

A2O1A1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1253),
.A2(n_1105),
.B(n_1053),
.C(n_1066),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1142),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1173),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1254),
.A2(n_1050),
.B(n_1051),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1163),
.A2(n_1069),
.B(n_1239),
.Y(n_1292)
);

BUFx3_ASAP7_75t_L g1293 ( 
.A(n_1111),
.Y(n_1293)
);

INVx5_ASAP7_75t_L g1294 ( 
.A(n_1198),
.Y(n_1294)
);

O2A1O1Ixp33_ASAP7_75t_SL g1295 ( 
.A1(n_1246),
.A2(n_1251),
.B(n_1192),
.C(n_1201),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1115),
.A2(n_1237),
.B(n_1238),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_SL g1297 ( 
.A(n_1191),
.B(n_1146),
.Y(n_1297)
);

AOI211x1_ASAP7_75t_L g1298 ( 
.A1(n_1159),
.A2(n_1218),
.B(n_1186),
.C(n_1168),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1260),
.A2(n_1127),
.B(n_1143),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1242),
.B(n_1132),
.Y(n_1300)
);

A2O1A1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1228),
.A2(n_1129),
.B(n_1252),
.C(n_1126),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1134),
.B(n_1191),
.Y(n_1302)
);

OAI221xp5_ASAP7_75t_L g1303 ( 
.A1(n_1224),
.A2(n_1174),
.B1(n_1218),
.B2(n_1233),
.C(n_1202),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1179),
.B(n_1131),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1130),
.B(n_1140),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1118),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1249),
.A2(n_1257),
.B(n_1256),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1198),
.Y(n_1308)
);

OAI22x1_ASAP7_75t_L g1309 ( 
.A1(n_1152),
.A2(n_1179),
.B1(n_1221),
.B2(n_1116),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1136),
.A2(n_1220),
.B(n_1215),
.Y(n_1310)
);

AO31x2_ASAP7_75t_L g1311 ( 
.A1(n_1177),
.A2(n_1166),
.A3(n_1204),
.B(n_1211),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1117),
.B(n_1264),
.Y(n_1312)
);

CKINVDCx6p67_ASAP7_75t_R g1313 ( 
.A(n_1128),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1196),
.Y(n_1314)
);

AO21x2_ASAP7_75t_L g1315 ( 
.A1(n_1256),
.A2(n_1217),
.B(n_1133),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_SL g1316 ( 
.A1(n_1244),
.A2(n_1248),
.B(n_1250),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1194),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1259),
.B(n_1255),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_SL g1319 ( 
.A(n_1234),
.B(n_1147),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1182),
.A2(n_1244),
.B(n_1119),
.Y(n_1320)
);

BUFx2_ASAP7_75t_L g1321 ( 
.A(n_1144),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_L g1322 ( 
.A(n_1112),
.B(n_1110),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1110),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1255),
.B(n_1124),
.Y(n_1324)
);

AOI31xp67_ASAP7_75t_L g1325 ( 
.A1(n_1158),
.A2(n_1160),
.A3(n_1209),
.B(n_1229),
.Y(n_1325)
);

AO21x2_ASAP7_75t_L g1326 ( 
.A1(n_1217),
.A2(n_1262),
.B(n_1119),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1126),
.A2(n_1199),
.B(n_1234),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1120),
.B(n_1203),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1182),
.A2(n_1205),
.B(n_1247),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1250),
.A2(n_1241),
.B(n_1169),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1222),
.A2(n_1145),
.B(n_1212),
.Y(n_1331)
);

O2A1O1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1157),
.A2(n_1214),
.B(n_1186),
.C(n_1230),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1139),
.A2(n_1219),
.B(n_1170),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1205),
.A2(n_1123),
.B(n_1189),
.Y(n_1334)
);

AO32x2_ASAP7_75t_L g1335 ( 
.A1(n_1213),
.A2(n_1165),
.A3(n_1235),
.B1(n_1227),
.B2(n_1216),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1207),
.B(n_1240),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1185),
.B(n_1183),
.Y(n_1337)
);

O2A1O1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1155),
.A2(n_1187),
.B(n_1175),
.C(n_1113),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_1223),
.Y(n_1339)
);

NAND2xp33_ASAP7_75t_L g1340 ( 
.A(n_1135),
.B(n_1223),
.Y(n_1340)
);

AO31x2_ASAP7_75t_L g1341 ( 
.A1(n_1232),
.A2(n_1231),
.A3(n_1184),
.B(n_1195),
.Y(n_1341)
);

CKINVDCx11_ASAP7_75t_R g1342 ( 
.A(n_1151),
.Y(n_1342)
);

NOR2x1_ASAP7_75t_L g1343 ( 
.A(n_1120),
.B(n_1135),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1263),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1263),
.B(n_1219),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1243),
.A2(n_1223),
.B(n_1227),
.Y(n_1346)
);

AO31x2_ASAP7_75t_L g1347 ( 
.A1(n_1148),
.A2(n_1149),
.A3(n_1153),
.B(n_1165),
.Y(n_1347)
);

A2O1A1Ixp33_ASAP7_75t_L g1348 ( 
.A1(n_1221),
.A2(n_1114),
.B(n_1226),
.C(n_1261),
.Y(n_1348)
);

AO31x2_ASAP7_75t_L g1349 ( 
.A1(n_1165),
.A2(n_1235),
.A3(n_1188),
.B(n_1261),
.Y(n_1349)
);

OA21x2_ASAP7_75t_L g1350 ( 
.A1(n_1235),
.A2(n_1261),
.B(n_1188),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1161),
.B(n_1141),
.Y(n_1351)
);

BUFx8_ASAP7_75t_L g1352 ( 
.A(n_1164),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1150),
.B(n_1141),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1200),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1180),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1180),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_SL g1357 ( 
.A(n_1206),
.B(n_1245),
.Y(n_1357)
);

AO22x1_ASAP7_75t_L g1358 ( 
.A1(n_1245),
.A2(n_1226),
.B1(n_1162),
.B2(n_1167),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1200),
.A2(n_1245),
.B1(n_1162),
.B2(n_1167),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_1156),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1167),
.A2(n_1156),
.B(n_1162),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1156),
.A2(n_1225),
.B(n_1122),
.Y(n_1362)
);

INVx5_ASAP7_75t_L g1363 ( 
.A(n_1198),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1111),
.Y(n_1364)
);

INVx1_ASAP7_75t_SL g1365 ( 
.A(n_1109),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1236),
.A2(n_1190),
.B(n_1210),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1109),
.B(n_964),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1138),
.B(n_1070),
.Y(n_1368)
);

AOI211x1_ASAP7_75t_L g1369 ( 
.A1(n_1159),
.A2(n_1218),
.B(n_1192),
.C(n_895),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1134),
.B(n_1018),
.Y(n_1370)
);

CKINVDCx11_ASAP7_75t_R g1371 ( 
.A(n_1111),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1134),
.B(n_1018),
.Y(n_1372)
);

OA21x2_ASAP7_75t_L g1373 ( 
.A1(n_1154),
.A2(n_1122),
.B(n_1225),
.Y(n_1373)
);

OAI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1225),
.A2(n_1122),
.B(n_939),
.Y(n_1374)
);

O2A1O1Ixp33_ASAP7_75t_SL g1375 ( 
.A1(n_1246),
.A2(n_1251),
.B(n_1192),
.C(n_938),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1171),
.A2(n_937),
.B1(n_1046),
.B2(n_1174),
.Y(n_1376)
);

OR2x6_ASAP7_75t_L g1377 ( 
.A(n_1142),
.B(n_824),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1242),
.B(n_1132),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_SL g1379 ( 
.A(n_1197),
.B(n_1138),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1208),
.B(n_861),
.Y(n_1380)
);

INVx2_ASAP7_75t_SL g1381 ( 
.A(n_1110),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_SL g1382 ( 
.A(n_1197),
.B(n_1138),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1242),
.B(n_1132),
.Y(n_1383)
);

O2A1O1Ixp33_ASAP7_75t_SL g1384 ( 
.A1(n_1246),
.A2(n_1251),
.B(n_1192),
.C(n_938),
.Y(n_1384)
);

AO31x2_ASAP7_75t_L g1385 ( 
.A1(n_1154),
.A2(n_950),
.A3(n_1254),
.B(n_1258),
.Y(n_1385)
);

A2O1A1Ixp33_ASAP7_75t_L g1386 ( 
.A1(n_1193),
.A2(n_1253),
.B(n_939),
.C(n_937),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1111),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1118),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1225),
.A2(n_1122),
.B(n_939),
.Y(n_1389)
);

O2A1O1Ixp33_ASAP7_75t_SL g1390 ( 
.A1(n_1246),
.A2(n_1251),
.B(n_1192),
.C(n_938),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1236),
.A2(n_1190),
.B(n_1210),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1121),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1121),
.Y(n_1393)
);

AO31x2_ASAP7_75t_L g1394 ( 
.A1(n_1154),
.A2(n_950),
.A3(n_1254),
.B(n_1258),
.Y(n_1394)
);

AO31x2_ASAP7_75t_L g1395 ( 
.A1(n_1154),
.A2(n_950),
.A3(n_1254),
.B(n_1258),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1122),
.A2(n_630),
.B(n_626),
.Y(n_1396)
);

OAI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1225),
.A2(n_1122),
.B(n_939),
.Y(n_1397)
);

O2A1O1Ixp33_ASAP7_75t_SL g1398 ( 
.A1(n_1246),
.A2(n_1251),
.B(n_1192),
.C(n_938),
.Y(n_1398)
);

AO31x2_ASAP7_75t_L g1399 ( 
.A1(n_1154),
.A2(n_950),
.A3(n_1254),
.B(n_1258),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1122),
.A2(n_630),
.B(n_626),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1171),
.A2(n_937),
.B1(n_1046),
.B2(n_1174),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1236),
.A2(n_1190),
.B(n_1210),
.Y(n_1402)
);

INVxp67_ASAP7_75t_L g1403 ( 
.A(n_1109),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1118),
.Y(n_1404)
);

AO31x2_ASAP7_75t_L g1405 ( 
.A1(n_1154),
.A2(n_950),
.A3(n_1254),
.B(n_1258),
.Y(n_1405)
);

A2O1A1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1193),
.A2(n_1253),
.B(n_939),
.C(n_937),
.Y(n_1406)
);

O2A1O1Ixp33_ASAP7_75t_SL g1407 ( 
.A1(n_1246),
.A2(n_1251),
.B(n_1192),
.C(n_938),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1122),
.A2(n_630),
.B(n_626),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1138),
.B(n_1070),
.Y(n_1409)
);

INVx4_ASAP7_75t_L g1410 ( 
.A(n_1141),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1242),
.B(n_1132),
.Y(n_1411)
);

BUFx2_ASAP7_75t_L g1412 ( 
.A(n_1109),
.Y(n_1412)
);

INVx3_ASAP7_75t_L g1413 ( 
.A(n_1198),
.Y(n_1413)
);

NAND2x1p5_ASAP7_75t_L g1414 ( 
.A(n_1203),
.B(n_1081),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1225),
.A2(n_1122),
.B(n_939),
.Y(n_1415)
);

INVx5_ASAP7_75t_L g1416 ( 
.A(n_1198),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1236),
.A2(n_1190),
.B(n_1210),
.Y(n_1417)
);

NAND3xp33_ASAP7_75t_L g1418 ( 
.A(n_1193),
.B(n_1251),
.C(n_1246),
.Y(n_1418)
);

OA21x2_ASAP7_75t_L g1419 ( 
.A1(n_1154),
.A2(n_1122),
.B(n_1225),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1138),
.B(n_1070),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1121),
.Y(n_1421)
);

AO21x2_ASAP7_75t_L g1422 ( 
.A1(n_1154),
.A2(n_1122),
.B(n_1071),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1242),
.B(n_1132),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1122),
.A2(n_630),
.B(n_626),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_SL g1425 ( 
.A(n_1197),
.B(n_1138),
.Y(n_1425)
);

AOI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1122),
.A2(n_1125),
.B(n_1154),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1236),
.A2(n_1190),
.B(n_1210),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1134),
.B(n_1018),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1236),
.A2(n_1190),
.B(n_1210),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_1111),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_SL g1431 ( 
.A1(n_1225),
.A2(n_1143),
.B(n_1136),
.Y(n_1431)
);

INVx4_ASAP7_75t_L g1432 ( 
.A(n_1276),
.Y(n_1432)
);

OAI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1376),
.A2(n_1401),
.B1(n_1319),
.B2(n_1303),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1376),
.A2(n_1401),
.B1(n_1418),
.B2(n_1303),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1266),
.Y(n_1435)
);

CKINVDCx11_ASAP7_75t_R g1436 ( 
.A(n_1342),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1276),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1278),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1276),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1377),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1418),
.A2(n_1386),
.B1(n_1406),
.B2(n_1301),
.Y(n_1441)
);

OAI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1319),
.A2(n_1275),
.B1(n_1305),
.B2(n_1330),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1285),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1380),
.A2(n_1316),
.B1(n_1425),
.B2(n_1382),
.Y(n_1444)
);

BUFx3_ASAP7_75t_L g1445 ( 
.A(n_1354),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1300),
.B(n_1378),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1377),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1290),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1317),
.Y(n_1449)
);

CKINVDCx11_ASAP7_75t_R g1450 ( 
.A(n_1371),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1368),
.A2(n_1409),
.B1(n_1420),
.B2(n_1315),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1315),
.A2(n_1350),
.B1(n_1326),
.B2(n_1305),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_SL g1453 ( 
.A1(n_1377),
.A2(n_1302),
.B1(n_1298),
.B2(n_1277),
.Y(n_1453)
);

CKINVDCx20_ASAP7_75t_R g1454 ( 
.A(n_1352),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1304),
.B(n_1337),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1350),
.A2(n_1326),
.B1(n_1330),
.B2(n_1397),
.Y(n_1456)
);

OAI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1275),
.A2(n_1415),
.B1(n_1389),
.B2(n_1397),
.Y(n_1457)
);

BUFx4f_ASAP7_75t_SL g1458 ( 
.A(n_1352),
.Y(n_1458)
);

AOI22xp5_ASAP7_75t_SL g1459 ( 
.A1(n_1370),
.A2(n_1372),
.B1(n_1428),
.B2(n_1309),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1282),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1374),
.A2(n_1415),
.B1(n_1389),
.B2(n_1378),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1374),
.A2(n_1300),
.B1(n_1383),
.B2(n_1423),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1383),
.B(n_1411),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_SL g1464 ( 
.A1(n_1307),
.A2(n_1411),
.B1(n_1423),
.B2(n_1327),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1379),
.A2(n_1365),
.B1(n_1369),
.B2(n_1403),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1392),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1393),
.Y(n_1467)
);

BUFx8_ASAP7_75t_SL g1468 ( 
.A(n_1430),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1295),
.A2(n_1407),
.B(n_1375),
.Y(n_1469)
);

OAI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1274),
.A2(n_1324),
.B1(n_1327),
.B2(n_1367),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1365),
.B(n_1318),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_1313),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1421),
.Y(n_1473)
);

CKINVDCx8_ASAP7_75t_R g1474 ( 
.A(n_1351),
.Y(n_1474)
);

CKINVDCx11_ASAP7_75t_R g1475 ( 
.A(n_1293),
.Y(n_1475)
);

OAI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1297),
.A2(n_1267),
.B1(n_1412),
.B2(n_1332),
.Y(n_1476)
);

BUFx3_ASAP7_75t_L g1477 ( 
.A(n_1321),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1336),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1289),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1388),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1336),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1318),
.B(n_1312),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1414),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1312),
.B(n_1370),
.Y(n_1484)
);

OAI22xp33_ASAP7_75t_R g1485 ( 
.A1(n_1322),
.A2(n_1314),
.B1(n_1381),
.B2(n_1323),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1324),
.A2(n_1280),
.B1(n_1273),
.B2(n_1351),
.Y(n_1486)
);

AOI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1372),
.A2(n_1428),
.B1(n_1384),
.B2(n_1390),
.Y(n_1487)
);

OAI22x1_ASAP7_75t_L g1488 ( 
.A1(n_1344),
.A2(n_1343),
.B1(n_1355),
.B2(n_1356),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1404),
.A2(n_1272),
.B1(n_1320),
.B2(n_1431),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1272),
.A2(n_1373),
.B1(n_1419),
.B2(n_1331),
.Y(n_1490)
);

OAI21xp5_ASAP7_75t_SL g1491 ( 
.A1(n_1338),
.A2(n_1353),
.B(n_1362),
.Y(n_1491)
);

INVx4_ASAP7_75t_L g1492 ( 
.A(n_1410),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1373),
.A2(n_1419),
.B1(n_1331),
.B2(n_1362),
.Y(n_1493)
);

OAI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1287),
.A2(n_1335),
.B1(n_1346),
.B2(n_1345),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1345),
.B(n_1348),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1287),
.A2(n_1387),
.B1(n_1364),
.B2(n_1422),
.Y(n_1496)
);

BUFx2_ASAP7_75t_L g1497 ( 
.A(n_1339),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1357),
.B(n_1349),
.Y(n_1498)
);

OAI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1335),
.A2(n_1346),
.B1(n_1294),
.B2(n_1363),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1422),
.A2(n_1281),
.B1(n_1284),
.B2(n_1291),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1410),
.A2(n_1284),
.B1(n_1281),
.B2(n_1308),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1349),
.B(n_1341),
.Y(n_1502)
);

OAI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1335),
.A2(n_1363),
.B1(n_1294),
.B2(n_1416),
.Y(n_1503)
);

INVx3_ASAP7_75t_SL g1504 ( 
.A(n_1339),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_SL g1505 ( 
.A1(n_1349),
.A2(n_1359),
.B1(n_1398),
.B2(n_1340),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1360),
.B(n_1341),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1291),
.A2(n_1328),
.B1(n_1359),
.B2(n_1271),
.Y(n_1507)
);

INVx1_ASAP7_75t_SL g1508 ( 
.A(n_1360),
.Y(n_1508)
);

AOI21xp33_ASAP7_75t_SL g1509 ( 
.A1(n_1308),
.A2(n_1413),
.B(n_1268),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1333),
.A2(n_1299),
.B1(n_1292),
.B2(n_1286),
.Y(n_1510)
);

INVx1_ASAP7_75t_SL g1511 ( 
.A(n_1358),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1413),
.A2(n_1363),
.B1(n_1294),
.B2(n_1416),
.Y(n_1512)
);

AOI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1363),
.A2(n_1416),
.B1(n_1361),
.B2(n_1334),
.Y(n_1513)
);

INVx4_ASAP7_75t_L g1514 ( 
.A(n_1361),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_1396),
.Y(n_1515)
);

BUFx6f_ASAP7_75t_L g1516 ( 
.A(n_1329),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1325),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1396),
.A2(n_1310),
.B1(n_1408),
.B2(n_1424),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_SL g1519 ( 
.A1(n_1296),
.A2(n_1405),
.B1(n_1394),
.B2(n_1385),
.Y(n_1519)
);

OAI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1400),
.A2(n_1426),
.B1(n_1395),
.B2(n_1385),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1288),
.A2(n_1347),
.B1(n_1395),
.B2(n_1385),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1394),
.B(n_1395),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1283),
.A2(n_1405),
.B1(n_1399),
.B2(n_1394),
.Y(n_1523)
);

BUFx8_ASAP7_75t_SL g1524 ( 
.A(n_1347),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_SL g1525 ( 
.A1(n_1399),
.A2(n_1405),
.B1(n_1311),
.B2(n_1279),
.Y(n_1525)
);

BUFx12f_ASAP7_75t_L g1526 ( 
.A(n_1269),
.Y(n_1526)
);

BUFx4f_ASAP7_75t_SL g1527 ( 
.A(n_1269),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1399),
.A2(n_1270),
.B1(n_1429),
.B2(n_1391),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1366),
.A2(n_1402),
.B1(n_1417),
.B2(n_1427),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1269),
.B(n_1311),
.Y(n_1530)
);

CKINVDCx11_ASAP7_75t_R g1531 ( 
.A(n_1265),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_SL g1532 ( 
.A1(n_1311),
.A2(n_1319),
.B1(n_1401),
.B2(n_1376),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1265),
.A2(n_1401),
.B1(n_1376),
.B2(n_1418),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1418),
.A2(n_1386),
.B1(n_1406),
.B2(n_1301),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1418),
.A2(n_1386),
.B1(n_1406),
.B2(n_1301),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1266),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1266),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1306),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_SL g1539 ( 
.A1(n_1319),
.A2(n_1401),
.B1(n_1376),
.B2(n_1147),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_SL g1540 ( 
.A1(n_1319),
.A2(n_1401),
.B1(n_1376),
.B2(n_1147),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1376),
.A2(n_1401),
.B1(n_1418),
.B2(n_897),
.Y(n_1541)
);

INVx2_ASAP7_75t_SL g1542 ( 
.A(n_1354),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1376),
.A2(n_1401),
.B1(n_1418),
.B2(n_897),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1377),
.Y(n_1544)
);

OAI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1376),
.A2(n_1401),
.B1(n_1319),
.B2(n_1303),
.Y(n_1545)
);

CKINVDCx6p67_ASAP7_75t_R g1546 ( 
.A(n_1342),
.Y(n_1546)
);

CKINVDCx6p67_ASAP7_75t_R g1547 ( 
.A(n_1342),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1376),
.A2(n_1401),
.B1(n_1418),
.B2(n_897),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1376),
.A2(n_1401),
.B1(n_1418),
.B2(n_897),
.Y(n_1549)
);

CKINVDCx11_ASAP7_75t_R g1550 ( 
.A(n_1342),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1266),
.Y(n_1551)
);

INVx3_ASAP7_75t_L g1552 ( 
.A(n_1276),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_SL g1553 ( 
.A1(n_1319),
.A2(n_1401),
.B1(n_1376),
.B2(n_1147),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1418),
.A2(n_1386),
.B1(n_1406),
.B2(n_1301),
.Y(n_1554)
);

INVxp67_ASAP7_75t_SL g1555 ( 
.A(n_1345),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1266),
.Y(n_1556)
);

BUFx2_ASAP7_75t_L g1557 ( 
.A(n_1377),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1266),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1266),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1418),
.A2(n_1386),
.B1(n_1406),
.B2(n_1301),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_SL g1561 ( 
.A1(n_1319),
.A2(n_1401),
.B1(n_1376),
.B2(n_1147),
.Y(n_1561)
);

CKINVDCx16_ASAP7_75t_R g1562 ( 
.A(n_1293),
.Y(n_1562)
);

INVx2_ASAP7_75t_SL g1563 ( 
.A(n_1354),
.Y(n_1563)
);

BUFx12f_ASAP7_75t_L g1564 ( 
.A(n_1342),
.Y(n_1564)
);

BUFx10_ASAP7_75t_L g1565 ( 
.A(n_1380),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1266),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1266),
.Y(n_1567)
);

INVx4_ASAP7_75t_L g1568 ( 
.A(n_1276),
.Y(n_1568)
);

BUFx3_ASAP7_75t_L g1569 ( 
.A(n_1354),
.Y(n_1569)
);

BUFx4f_ASAP7_75t_SL g1570 ( 
.A(n_1352),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1376),
.A2(n_1401),
.B1(n_1418),
.B2(n_897),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1376),
.A2(n_1401),
.B1(n_1418),
.B2(n_897),
.Y(n_1572)
);

BUFx2_ASAP7_75t_L g1573 ( 
.A(n_1377),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_SL g1574 ( 
.A1(n_1319),
.A2(n_1401),
.B1(n_1376),
.B2(n_1147),
.Y(n_1574)
);

INVx2_ASAP7_75t_SL g1575 ( 
.A(n_1354),
.Y(n_1575)
);

INVx6_ASAP7_75t_L g1576 ( 
.A(n_1276),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_SL g1577 ( 
.A1(n_1319),
.A2(n_1401),
.B1(n_1376),
.B2(n_1147),
.Y(n_1577)
);

BUFx4f_ASAP7_75t_SL g1578 ( 
.A(n_1352),
.Y(n_1578)
);

AOI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1376),
.A2(n_1401),
.B1(n_1208),
.B2(n_1418),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1266),
.Y(n_1580)
);

OAI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1376),
.A2(n_1401),
.B1(n_1319),
.B2(n_1303),
.Y(n_1581)
);

INVx2_ASAP7_75t_SL g1582 ( 
.A(n_1506),
.Y(n_1582)
);

OAI21x1_ASAP7_75t_L g1583 ( 
.A1(n_1529),
.A2(n_1528),
.B(n_1518),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1446),
.B(n_1463),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1555),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1530),
.B(n_1532),
.Y(n_1586)
);

INVx3_ASAP7_75t_L g1587 ( 
.A(n_1516),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1471),
.Y(n_1588)
);

AOI21x1_ASAP7_75t_L g1589 ( 
.A1(n_1469),
.A2(n_1517),
.B(n_1521),
.Y(n_1589)
);

AOI21x1_ASAP7_75t_L g1590 ( 
.A1(n_1522),
.A2(n_1534),
.B(n_1441),
.Y(n_1590)
);

AO21x2_ASAP7_75t_L g1591 ( 
.A1(n_1520),
.A2(n_1494),
.B(n_1433),
.Y(n_1591)
);

OAI21x1_ASAP7_75t_L g1592 ( 
.A1(n_1529),
.A2(n_1528),
.B(n_1518),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1479),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1498),
.Y(n_1594)
);

BUFx2_ASAP7_75t_L g1595 ( 
.A(n_1515),
.Y(n_1595)
);

AOI21xp5_ASAP7_75t_L g1596 ( 
.A1(n_1433),
.A2(n_1581),
.B(n_1545),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1482),
.B(n_1462),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1502),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_SL g1599 ( 
.A1(n_1535),
.A2(n_1560),
.B1(n_1554),
.B2(n_1459),
.Y(n_1599)
);

OAI21x1_ASAP7_75t_L g1600 ( 
.A1(n_1510),
.A2(n_1490),
.B(n_1500),
.Y(n_1600)
);

INVx5_ASAP7_75t_L g1601 ( 
.A(n_1526),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1435),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1451),
.B(n_1533),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1514),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1438),
.Y(n_1605)
);

INVx4_ASAP7_75t_SL g1606 ( 
.A(n_1527),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1539),
.A2(n_1574),
.B1(n_1561),
.B2(n_1553),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1527),
.Y(n_1608)
);

AOI21x1_ASAP7_75t_L g1609 ( 
.A1(n_1501),
.A2(n_1486),
.B(n_1488),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1451),
.B(n_1533),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1443),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1565),
.B(n_1444),
.Y(n_1612)
);

INVx2_ASAP7_75t_SL g1613 ( 
.A(n_1477),
.Y(n_1613)
);

OAI21x1_ASAP7_75t_L g1614 ( 
.A1(n_1510),
.A2(n_1490),
.B(n_1500),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1448),
.Y(n_1615)
);

OAI21x1_ASAP7_75t_L g1616 ( 
.A1(n_1493),
.A2(n_1489),
.B(n_1523),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1449),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1466),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1467),
.Y(n_1619)
);

OAI21x1_ASAP7_75t_L g1620 ( 
.A1(n_1493),
.A2(n_1489),
.B(n_1523),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1462),
.B(n_1478),
.Y(n_1621)
);

OAI21x1_ASAP7_75t_L g1622 ( 
.A1(n_1507),
.A2(n_1456),
.B(n_1513),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1473),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1536),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1537),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1456),
.B(n_1540),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1551),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1556),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1558),
.Y(n_1629)
);

OAI21x1_ASAP7_75t_L g1630 ( 
.A1(n_1507),
.A2(n_1496),
.B(n_1461),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1559),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1566),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1567),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1580),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1434),
.A2(n_1579),
.B1(n_1581),
.B2(n_1545),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1481),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1452),
.Y(n_1637)
);

BUFx12f_ASAP7_75t_L g1638 ( 
.A(n_1436),
.Y(n_1638)
);

AOI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1577),
.A2(n_1434),
.B1(n_1541),
.B2(n_1548),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1461),
.B(n_1452),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1464),
.B(n_1541),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1457),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1484),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1457),
.Y(n_1644)
);

OA21x2_ASAP7_75t_L g1645 ( 
.A1(n_1543),
.A2(n_1549),
.B(n_1571),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1494),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1524),
.Y(n_1647)
);

OAI21x1_ASAP7_75t_L g1648 ( 
.A1(n_1496),
.A2(n_1487),
.B(n_1512),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1519),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1440),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1531),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1525),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1520),
.Y(n_1653)
);

OR2x6_ASAP7_75t_L g1654 ( 
.A(n_1495),
.B(n_1491),
.Y(n_1654)
);

AOI21x1_ASAP7_75t_L g1655 ( 
.A1(n_1465),
.A2(n_1476),
.B(n_1557),
.Y(n_1655)
);

BUFx5_ASAP7_75t_L g1656 ( 
.A(n_1503),
.Y(n_1656)
);

OAI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1572),
.A2(n_1442),
.B1(n_1453),
.B2(n_1470),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1477),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1442),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1447),
.Y(n_1660)
);

OA21x2_ASAP7_75t_L g1661 ( 
.A1(n_1572),
.A2(n_1480),
.B(n_1538),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1544),
.Y(n_1662)
);

OAI21x1_ASAP7_75t_L g1663 ( 
.A1(n_1512),
.A2(n_1483),
.B(n_1552),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1573),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1470),
.B(n_1499),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1499),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1455),
.B(n_1503),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1505),
.B(n_1497),
.Y(n_1668)
);

AO21x1_ASAP7_75t_SL g1669 ( 
.A1(n_1509),
.A2(n_1485),
.B(n_1504),
.Y(n_1669)
);

BUFx3_ASAP7_75t_L g1670 ( 
.A(n_1437),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1437),
.Y(n_1671)
);

INVx3_ASAP7_75t_L g1672 ( 
.A(n_1437),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1439),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1439),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1508),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1565),
.B(n_1460),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1460),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1432),
.B(n_1568),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1511),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1576),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1576),
.Y(n_1681)
);

INVx2_ASAP7_75t_SL g1682 ( 
.A(n_1445),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1474),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_1468),
.Y(n_1684)
);

OAI21x1_ASAP7_75t_L g1685 ( 
.A1(n_1492),
.A2(n_1445),
.B(n_1569),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1492),
.Y(n_1686)
);

HB1xp67_ASAP7_75t_L g1687 ( 
.A(n_1569),
.Y(n_1687)
);

OAI21x1_ASAP7_75t_L g1688 ( 
.A1(n_1458),
.A2(n_1578),
.B(n_1570),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1542),
.Y(n_1689)
);

BUFx2_ASAP7_75t_L g1690 ( 
.A(n_1563),
.Y(n_1690)
);

BUFx4f_ASAP7_75t_L g1691 ( 
.A(n_1575),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1562),
.Y(n_1692)
);

AOI221xp5_ASAP7_75t_L g1693 ( 
.A1(n_1635),
.A2(n_1472),
.B1(n_1454),
.B2(n_1550),
.C(n_1450),
.Y(n_1693)
);

OAI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1596),
.A2(n_1458),
.B(n_1570),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1595),
.B(n_1578),
.Y(n_1695)
);

BUFx2_ASAP7_75t_L g1696 ( 
.A(n_1595),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1658),
.B(n_1613),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1602),
.B(n_1546),
.Y(n_1698)
);

OA21x2_ASAP7_75t_L g1699 ( 
.A1(n_1583),
.A2(n_1475),
.B(n_1547),
.Y(n_1699)
);

NOR2x1_ASAP7_75t_SL g1700 ( 
.A(n_1669),
.B(n_1564),
.Y(n_1700)
);

O2A1O1Ixp33_ASAP7_75t_SL g1701 ( 
.A1(n_1692),
.A2(n_1613),
.B(n_1687),
.C(n_1593),
.Y(n_1701)
);

OAI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1599),
.A2(n_1607),
.B(n_1657),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1682),
.B(n_1690),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1650),
.B(n_1660),
.Y(n_1704)
);

OR2x6_ASAP7_75t_L g1705 ( 
.A(n_1665),
.B(n_1648),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1650),
.B(n_1662),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1664),
.B(n_1690),
.Y(n_1707)
);

AO32x2_ASAP7_75t_L g1708 ( 
.A1(n_1582),
.A2(n_1682),
.A3(n_1588),
.B1(n_1643),
.B2(n_1590),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1639),
.A2(n_1654),
.B1(n_1665),
.B2(n_1644),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1642),
.B(n_1644),
.Y(n_1710)
);

BUFx6f_ASAP7_75t_L g1711 ( 
.A(n_1691),
.Y(n_1711)
);

A2O1A1Ixp33_ASAP7_75t_L g1712 ( 
.A1(n_1626),
.A2(n_1612),
.B(n_1641),
.C(n_1639),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1676),
.Y(n_1713)
);

OAI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1630),
.A2(n_1642),
.B(n_1590),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1606),
.B(n_1601),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1625),
.B(n_1627),
.Y(n_1716)
);

BUFx2_ASAP7_75t_L g1717 ( 
.A(n_1689),
.Y(n_1717)
);

AO21x2_ASAP7_75t_L g1718 ( 
.A1(n_1646),
.A2(n_1637),
.B(n_1591),
.Y(n_1718)
);

O2A1O1Ixp33_ASAP7_75t_SL g1719 ( 
.A1(n_1686),
.A2(n_1632),
.B(n_1638),
.C(n_1597),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1654),
.Y(n_1720)
);

AOI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1591),
.A2(n_1630),
.B(n_1654),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1685),
.Y(n_1722)
);

OAI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1659),
.A2(n_1654),
.B(n_1609),
.Y(n_1723)
);

AOI221xp5_ASAP7_75t_L g1724 ( 
.A1(n_1646),
.A2(n_1640),
.B1(n_1649),
.B2(n_1653),
.C(n_1652),
.Y(n_1724)
);

BUFx12f_ASAP7_75t_L g1725 ( 
.A(n_1638),
.Y(n_1725)
);

NOR2x1_ASAP7_75t_SL g1726 ( 
.A(n_1669),
.B(n_1654),
.Y(n_1726)
);

OAI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1659),
.A2(n_1603),
.B1(n_1610),
.B2(n_1609),
.C(n_1653),
.Y(n_1727)
);

NOR2x1_ASAP7_75t_SL g1728 ( 
.A(n_1667),
.B(n_1591),
.Y(n_1728)
);

OA21x2_ASAP7_75t_L g1729 ( 
.A1(n_1583),
.A2(n_1592),
.B(n_1622),
.Y(n_1729)
);

AO21x1_ASAP7_75t_L g1730 ( 
.A1(n_1621),
.A2(n_1640),
.B(n_1655),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1689),
.B(n_1647),
.Y(n_1731)
);

CKINVDCx20_ASAP7_75t_R g1732 ( 
.A(n_1684),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1585),
.Y(n_1733)
);

INVxp33_ASAP7_75t_SL g1734 ( 
.A(n_1688),
.Y(n_1734)
);

AOI221xp5_ASAP7_75t_L g1735 ( 
.A1(n_1666),
.A2(n_1586),
.B1(n_1637),
.B2(n_1594),
.C(n_1610),
.Y(n_1735)
);

OA21x2_ASAP7_75t_L g1736 ( 
.A1(n_1592),
.A2(n_1614),
.B(n_1600),
.Y(n_1736)
);

OAI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1655),
.A2(n_1614),
.B(n_1600),
.Y(n_1737)
);

OA21x2_ASAP7_75t_L g1738 ( 
.A1(n_1616),
.A2(n_1620),
.B(n_1666),
.Y(n_1738)
);

AOI221xp5_ASAP7_75t_L g1739 ( 
.A1(n_1603),
.A2(n_1586),
.B1(n_1605),
.B2(n_1611),
.C(n_1617),
.Y(n_1739)
);

A2O1A1Ixp33_ASAP7_75t_L g1740 ( 
.A1(n_1616),
.A2(n_1620),
.B(n_1651),
.C(n_1679),
.Y(n_1740)
);

NAND3xp33_ASAP7_75t_L g1741 ( 
.A(n_1585),
.B(n_1675),
.C(n_1686),
.Y(n_1741)
);

AO21x1_ASAP7_75t_L g1742 ( 
.A1(n_1605),
.A2(n_1634),
.B(n_1633),
.Y(n_1742)
);

A2O1A1Ixp33_ASAP7_75t_L g1743 ( 
.A1(n_1679),
.A2(n_1668),
.B(n_1691),
.C(n_1683),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1673),
.B(n_1674),
.Y(n_1744)
);

A2O1A1Ixp33_ASAP7_75t_L g1745 ( 
.A1(n_1679),
.A2(n_1668),
.B(n_1691),
.C(n_1683),
.Y(n_1745)
);

A2O1A1Ixp33_ASAP7_75t_L g1746 ( 
.A1(n_1691),
.A2(n_1584),
.B(n_1608),
.C(n_1685),
.Y(n_1746)
);

AND2x4_ASAP7_75t_L g1747 ( 
.A(n_1606),
.B(n_1601),
.Y(n_1747)
);

AND2x4_ASAP7_75t_L g1748 ( 
.A(n_1606),
.B(n_1601),
.Y(n_1748)
);

AOI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1604),
.A2(n_1645),
.B(n_1587),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1678),
.B(n_1681),
.Y(n_1750)
);

OAI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1645),
.A2(n_1611),
.B1(n_1617),
.B2(n_1634),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_1606),
.B(n_1601),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1636),
.B(n_1615),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1677),
.B(n_1670),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1680),
.B(n_1619),
.Y(n_1755)
);

BUFx2_ASAP7_75t_L g1756 ( 
.A(n_1681),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1680),
.B(n_1619),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_L g1758 ( 
.A(n_1672),
.B(n_1680),
.Y(n_1758)
);

OAI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1645),
.A2(n_1589),
.B(n_1663),
.Y(n_1759)
);

AOI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1645),
.A2(n_1656),
.B1(n_1633),
.B2(n_1629),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1672),
.B(n_1629),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1636),
.B(n_1628),
.Y(n_1762)
);

OAI222xp33_ASAP7_75t_L g1763 ( 
.A1(n_1727),
.A2(n_1709),
.B1(n_1760),
.B2(n_1705),
.C1(n_1721),
.C2(n_1751),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1736),
.B(n_1729),
.Y(n_1764)
);

AND2x2_ASAP7_75t_SL g1765 ( 
.A(n_1739),
.B(n_1656),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1751),
.B(n_1624),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1742),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1736),
.B(n_1656),
.Y(n_1768)
);

NOR2x1_ASAP7_75t_L g1769 ( 
.A(n_1741),
.B(n_1671),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1729),
.B(n_1656),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1738),
.B(n_1755),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1733),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1753),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1716),
.B(n_1624),
.Y(n_1774)
);

INVxp67_ASAP7_75t_L g1775 ( 
.A(n_1717),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1738),
.B(n_1656),
.Y(n_1776)
);

INVxp67_ASAP7_75t_L g1777 ( 
.A(n_1756),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1753),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1762),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1757),
.B(n_1656),
.Y(n_1780)
);

INVx4_ASAP7_75t_L g1781 ( 
.A(n_1715),
.Y(n_1781)
);

INVxp67_ASAP7_75t_L g1782 ( 
.A(n_1741),
.Y(n_1782)
);

AOI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1702),
.A2(n_1656),
.B1(n_1598),
.B2(n_1661),
.Y(n_1783)
);

INVx3_ASAP7_75t_L g1784 ( 
.A(n_1722),
.Y(n_1784)
);

AOI22xp33_ASAP7_75t_L g1785 ( 
.A1(n_1702),
.A2(n_1656),
.B1(n_1598),
.B2(n_1661),
.Y(n_1785)
);

INVxp67_ASAP7_75t_L g1786 ( 
.A(n_1696),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1713),
.B(n_1628),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1730),
.B(n_1631),
.Y(n_1788)
);

NOR2x1_ASAP7_75t_L g1789 ( 
.A(n_1746),
.B(n_1671),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_L g1790 ( 
.A(n_1704),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_SL g1791 ( 
.A1(n_1709),
.A2(n_1661),
.B1(n_1623),
.B2(n_1631),
.Y(n_1791)
);

BUFx3_ASAP7_75t_L g1792 ( 
.A(n_1725),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1706),
.Y(n_1793)
);

INVx4_ASAP7_75t_L g1794 ( 
.A(n_1747),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1718),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1710),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1710),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1708),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1708),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1708),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1728),
.Y(n_1801)
);

INVx3_ASAP7_75t_L g1802 ( 
.A(n_1722),
.Y(n_1802)
);

AOI31xp33_ASAP7_75t_L g1803 ( 
.A1(n_1782),
.A2(n_1693),
.A3(n_1694),
.B(n_1712),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1782),
.B(n_1707),
.Y(n_1804)
);

CKINVDCx14_ASAP7_75t_R g1805 ( 
.A(n_1792),
.Y(n_1805)
);

INVx4_ASAP7_75t_L g1806 ( 
.A(n_1792),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1790),
.B(n_1697),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1775),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1764),
.Y(n_1809)
);

NOR2x1_ASAP7_75t_L g1810 ( 
.A(n_1769),
.B(n_1699),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_1792),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1796),
.B(n_1720),
.Y(n_1812)
);

AND2x2_ASAP7_75t_SL g1813 ( 
.A(n_1765),
.B(n_1739),
.Y(n_1813)
);

AOI221xp5_ASAP7_75t_L g1814 ( 
.A1(n_1763),
.A2(n_1724),
.B1(n_1714),
.B2(n_1735),
.C(n_1737),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1790),
.B(n_1713),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1793),
.B(n_1731),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1765),
.A2(n_1785),
.B1(n_1783),
.B2(n_1791),
.Y(n_1817)
);

INVxp67_ASAP7_75t_SL g1818 ( 
.A(n_1769),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1773),
.Y(n_1819)
);

OA21x2_ASAP7_75t_L g1820 ( 
.A1(n_1795),
.A2(n_1737),
.B(n_1759),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1764),
.Y(n_1821)
);

AOI22xp33_ASAP7_75t_L g1822 ( 
.A1(n_1765),
.A2(n_1791),
.B1(n_1723),
.B2(n_1776),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1773),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1778),
.Y(n_1824)
);

NAND3xp33_ASAP7_75t_L g1825 ( 
.A(n_1767),
.B(n_1693),
.C(n_1723),
.Y(n_1825)
);

INVx1_ASAP7_75t_SL g1826 ( 
.A(n_1774),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1764),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1793),
.B(n_1786),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1778),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1780),
.B(n_1699),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1796),
.B(n_1703),
.Y(n_1831)
);

AOI22xp33_ASAP7_75t_L g1832 ( 
.A1(n_1776),
.A2(n_1661),
.B1(n_1759),
.B2(n_1734),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1780),
.B(n_1754),
.Y(n_1833)
);

OAI322xp33_ASAP7_75t_L g1834 ( 
.A1(n_1767),
.A2(n_1698),
.A3(n_1695),
.B1(n_1761),
.B2(n_1749),
.C1(n_1618),
.C2(n_1623),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1780),
.B(n_1777),
.Y(n_1835)
);

AOI221xp5_ASAP7_75t_L g1836 ( 
.A1(n_1763),
.A2(n_1740),
.B1(n_1743),
.B2(n_1745),
.C(n_1701),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1774),
.B(n_1744),
.Y(n_1837)
);

CKINVDCx16_ASAP7_75t_R g1838 ( 
.A(n_1781),
.Y(n_1838)
);

INVx2_ASAP7_75t_SL g1839 ( 
.A(n_1787),
.Y(n_1839)
);

INVxp67_ASAP7_75t_SL g1840 ( 
.A(n_1766),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1771),
.B(n_1750),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1771),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1797),
.B(n_1758),
.Y(n_1843)
);

NOR2x1p5_ASAP7_75t_L g1844 ( 
.A(n_1781),
.B(n_1711),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1779),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1771),
.B(n_1726),
.Y(n_1846)
);

AOI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1776),
.A2(n_1694),
.B1(n_1748),
.B2(n_1752),
.Y(n_1847)
);

INVx2_ASAP7_75t_SL g1848 ( 
.A(n_1838),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1842),
.B(n_1768),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1842),
.B(n_1768),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1842),
.Y(n_1851)
);

AOI22xp33_ASAP7_75t_L g1852 ( 
.A1(n_1813),
.A2(n_1799),
.B1(n_1800),
.B2(n_1798),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1830),
.B(n_1768),
.Y(n_1853)
);

NAND2x1_ASAP7_75t_L g1854 ( 
.A(n_1810),
.B(n_1781),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1830),
.B(n_1770),
.Y(n_1855)
);

OR2x2_ASAP7_75t_L g1856 ( 
.A(n_1840),
.B(n_1766),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1819),
.Y(n_1857)
);

INVx2_ASAP7_75t_SL g1858 ( 
.A(n_1838),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1819),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1823),
.Y(n_1860)
);

INVx1_ASAP7_75t_SL g1861 ( 
.A(n_1808),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1809),
.Y(n_1862)
);

NOR2x1_ASAP7_75t_L g1863 ( 
.A(n_1806),
.B(n_1801),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1824),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1829),
.B(n_1772),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1809),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1809),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1841),
.B(n_1770),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1846),
.B(n_1835),
.Y(n_1869)
);

INVx4_ASAP7_75t_L g1870 ( 
.A(n_1806),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1826),
.B(n_1798),
.Y(n_1871)
);

NAND2x1_ASAP7_75t_L g1872 ( 
.A(n_1810),
.B(n_1781),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1818),
.B(n_1784),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1815),
.B(n_1833),
.Y(n_1874)
);

INVx3_ASAP7_75t_L g1875 ( 
.A(n_1821),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1845),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1821),
.Y(n_1877)
);

AND2x4_ASAP7_75t_SL g1878 ( 
.A(n_1847),
.B(n_1794),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1821),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1828),
.B(n_1802),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1826),
.B(n_1799),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1839),
.B(n_1800),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1861),
.B(n_1825),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1857),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1857),
.Y(n_1885)
);

INVxp33_ASAP7_75t_L g1886 ( 
.A(n_1854),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1874),
.B(n_1828),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1875),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1856),
.B(n_1812),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1856),
.B(n_1839),
.Y(n_1890)
);

AOI22xp33_ASAP7_75t_L g1891 ( 
.A1(n_1852),
.A2(n_1813),
.B1(n_1817),
.B2(n_1814),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1874),
.B(n_1806),
.Y(n_1892)
);

NOR2x1p5_ASAP7_75t_L g1893 ( 
.A(n_1854),
.B(n_1806),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1875),
.Y(n_1894)
);

OR2x2_ASAP7_75t_L g1895 ( 
.A(n_1856),
.B(n_1843),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1859),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1874),
.B(n_1816),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1875),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1859),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1860),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1875),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1860),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1875),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1861),
.B(n_1825),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1852),
.B(n_1804),
.Y(n_1905)
);

AND2x4_ASAP7_75t_L g1906 ( 
.A(n_1878),
.B(n_1870),
.Y(n_1906)
);

AND2x4_ASAP7_75t_L g1907 ( 
.A(n_1878),
.B(n_1844),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1849),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1864),
.Y(n_1909)
);

INVxp67_ASAP7_75t_L g1910 ( 
.A(n_1848),
.Y(n_1910)
);

OR2x2_ASAP7_75t_L g1911 ( 
.A(n_1871),
.B(n_1827),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1865),
.B(n_1831),
.Y(n_1912)
);

NAND2x1_ASAP7_75t_L g1913 ( 
.A(n_1863),
.B(n_1827),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1865),
.B(n_1803),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1849),
.Y(n_1915)
);

OR2x2_ASAP7_75t_L g1916 ( 
.A(n_1871),
.B(n_1827),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1878),
.B(n_1816),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1849),
.Y(n_1918)
);

OR2x2_ASAP7_75t_L g1919 ( 
.A(n_1871),
.B(n_1837),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1850),
.Y(n_1920)
);

AND3x2_ASAP7_75t_L g1921 ( 
.A(n_1873),
.B(n_1836),
.C(n_1700),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1864),
.Y(n_1922)
);

OR2x2_ASAP7_75t_L g1923 ( 
.A(n_1881),
.B(n_1837),
.Y(n_1923)
);

NOR2x1p5_ASAP7_75t_SL g1924 ( 
.A(n_1862),
.B(n_1801),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1878),
.B(n_1807),
.Y(n_1925)
);

OAI22xp33_ASAP7_75t_L g1926 ( 
.A1(n_1854),
.A2(n_1803),
.B1(n_1847),
.B2(n_1813),
.Y(n_1926)
);

AOI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1872),
.A2(n_1834),
.B(n_1822),
.Y(n_1927)
);

INVx4_ASAP7_75t_L g1928 ( 
.A(n_1870),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1851),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_L g1930 ( 
.A(n_1914),
.B(n_1805),
.Y(n_1930)
);

INVx2_ASAP7_75t_SL g1931 ( 
.A(n_1906),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1883),
.B(n_1869),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1884),
.Y(n_1933)
);

OR2x2_ASAP7_75t_L g1934 ( 
.A(n_1895),
.B(n_1881),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1884),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1908),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1895),
.B(n_1881),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1885),
.Y(n_1938)
);

BUFx2_ASAP7_75t_L g1939 ( 
.A(n_1910),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_L g1940 ( 
.A(n_1904),
.B(n_1811),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1885),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1908),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1926),
.B(n_1732),
.Y(n_1943)
);

AND2x4_ASAP7_75t_L g1944 ( 
.A(n_1906),
.B(n_1870),
.Y(n_1944)
);

OR2x2_ASAP7_75t_L g1945 ( 
.A(n_1912),
.B(n_1882),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1891),
.B(n_1869),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_SL g1947 ( 
.A(n_1907),
.B(n_1848),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1896),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1896),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1897),
.B(n_1869),
.Y(n_1950)
);

NOR2xp33_ASAP7_75t_L g1951 ( 
.A(n_1928),
.B(n_1870),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1899),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1905),
.B(n_1887),
.Y(n_1953)
);

INVx2_ASAP7_75t_SL g1954 ( 
.A(n_1906),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1899),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1887),
.B(n_1853),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1897),
.B(n_1853),
.Y(n_1957)
);

OR2x2_ASAP7_75t_L g1958 ( 
.A(n_1889),
.B(n_1882),
.Y(n_1958)
);

INVx3_ASAP7_75t_L g1959 ( 
.A(n_1907),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1892),
.B(n_1848),
.Y(n_1960)
);

INVx4_ASAP7_75t_L g1961 ( 
.A(n_1928),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1889),
.B(n_1853),
.Y(n_1962)
);

OAI21xp5_ASAP7_75t_SL g1963 ( 
.A1(n_1921),
.A2(n_1863),
.B(n_1858),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1892),
.B(n_1858),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1900),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1907),
.B(n_1858),
.Y(n_1966)
);

AOI221xp5_ASAP7_75t_L g1967 ( 
.A1(n_1946),
.A2(n_1927),
.B1(n_1953),
.B2(n_1932),
.C(n_1939),
.Y(n_1967)
);

AOI21xp5_ASAP7_75t_L g1968 ( 
.A1(n_1963),
.A2(n_1872),
.B(n_1886),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1933),
.Y(n_1969)
);

INVxp67_ASAP7_75t_L g1970 ( 
.A(n_1940),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1933),
.Y(n_1971)
);

OAI21xp33_ASAP7_75t_L g1972 ( 
.A1(n_1960),
.A2(n_1890),
.B(n_1915),
.Y(n_1972)
);

AOI21xp5_ASAP7_75t_L g1973 ( 
.A1(n_1943),
.A2(n_1872),
.B(n_1913),
.Y(n_1973)
);

AOI22xp5_ASAP7_75t_L g1974 ( 
.A1(n_1930),
.A2(n_1832),
.B1(n_1820),
.B2(n_1788),
.Y(n_1974)
);

OR2x2_ASAP7_75t_L g1975 ( 
.A(n_1934),
.B(n_1890),
.Y(n_1975)
);

A2O1A1Ixp33_ASAP7_75t_L g1976 ( 
.A1(n_1934),
.A2(n_1924),
.B(n_1923),
.C(n_1919),
.Y(n_1976)
);

AOI22xp5_ASAP7_75t_L g1977 ( 
.A1(n_1936),
.A2(n_1942),
.B1(n_1966),
.B2(n_1959),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1948),
.Y(n_1978)
);

INVx1_ASAP7_75t_SL g1979 ( 
.A(n_1939),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1948),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1936),
.B(n_1900),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1955),
.Y(n_1982)
);

AOI31xp33_ASAP7_75t_L g1983 ( 
.A1(n_1931),
.A2(n_1906),
.A3(n_1907),
.B(n_1925),
.Y(n_1983)
);

OAI21xp5_ASAP7_75t_SL g1984 ( 
.A1(n_1959),
.A2(n_1925),
.B(n_1917),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1942),
.B(n_1902),
.Y(n_1985)
);

OAI21xp33_ASAP7_75t_L g1986 ( 
.A1(n_1960),
.A2(n_1918),
.B(n_1915),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1955),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1935),
.Y(n_1988)
);

OAI21xp33_ASAP7_75t_L g1989 ( 
.A1(n_1964),
.A2(n_1920),
.B(n_1918),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1938),
.Y(n_1990)
);

OAI221xp5_ASAP7_75t_L g1991 ( 
.A1(n_1937),
.A2(n_1919),
.B1(n_1923),
.B2(n_1916),
.C(n_1911),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1941),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1949),
.Y(n_1993)
);

AOI22xp5_ASAP7_75t_L g1994 ( 
.A1(n_1966),
.A2(n_1820),
.B1(n_1788),
.B2(n_1855),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1979),
.B(n_1950),
.Y(n_1995)
);

NAND4xp25_ASAP7_75t_L g1996 ( 
.A(n_1967),
.B(n_1951),
.C(n_1959),
.D(n_1961),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1975),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1970),
.B(n_1931),
.Y(n_1998)
);

AOI22xp5_ASAP7_75t_L g1999 ( 
.A1(n_1974),
.A2(n_1954),
.B1(n_1937),
.B2(n_1947),
.Y(n_1999)
);

OAI21xp33_ASAP7_75t_L g2000 ( 
.A1(n_1972),
.A2(n_1984),
.B(n_1986),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1969),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1971),
.Y(n_2002)
);

NOR4xp25_ASAP7_75t_SL g2003 ( 
.A(n_1976),
.B(n_1965),
.C(n_1952),
.D(n_1954),
.Y(n_2003)
);

NOR2xp33_ASAP7_75t_L g2004 ( 
.A(n_1983),
.B(n_1944),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1977),
.B(n_1950),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1989),
.B(n_1962),
.Y(n_2006)
);

AOI31xp33_ASAP7_75t_L g2007 ( 
.A1(n_1968),
.A2(n_1944),
.A3(n_1964),
.B(n_1958),
.Y(n_2007)
);

HB1xp67_ASAP7_75t_L g2008 ( 
.A(n_1978),
.Y(n_2008)
);

OAI22xp5_ASAP7_75t_L g2009 ( 
.A1(n_1994),
.A2(n_1956),
.B1(n_1957),
.B2(n_1958),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1988),
.B(n_1944),
.Y(n_2010)
);

OAI22xp33_ASAP7_75t_L g2011 ( 
.A1(n_1991),
.A2(n_1945),
.B1(n_1911),
.B2(n_1916),
.Y(n_2011)
);

INVx1_ASAP7_75t_SL g2012 ( 
.A(n_1981),
.Y(n_2012)
);

AOI22xp33_ASAP7_75t_L g2013 ( 
.A1(n_1981),
.A2(n_1929),
.B1(n_1945),
.B2(n_1820),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1980),
.Y(n_2014)
);

OAI22xp33_ASAP7_75t_L g2015 ( 
.A1(n_1999),
.A2(n_1985),
.B1(n_1987),
.B2(n_1982),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_2008),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_2008),
.Y(n_2017)
);

INVxp67_ASAP7_75t_L g2018 ( 
.A(n_1998),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_2003),
.B(n_1961),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1997),
.Y(n_2020)
);

NOR2xp67_ASAP7_75t_L g2021 ( 
.A(n_1996),
.B(n_1961),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1995),
.Y(n_2022)
);

OAI21xp5_ASAP7_75t_SL g2023 ( 
.A1(n_2007),
.A2(n_1973),
.B(n_1990),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_2001),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_2002),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_2014),
.Y(n_2026)
);

OAI22xp5_ASAP7_75t_L g2027 ( 
.A1(n_2015),
.A2(n_2005),
.B1(n_2013),
.B2(n_2006),
.Y(n_2027)
);

INVx1_ASAP7_75t_SL g2028 ( 
.A(n_2019),
.Y(n_2028)
);

AOI22xp33_ASAP7_75t_L g2029 ( 
.A1(n_2015),
.A2(n_2013),
.B1(n_2012),
.B2(n_2009),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_2018),
.B(n_2010),
.Y(n_2030)
);

AOI22xp5_ASAP7_75t_L g2031 ( 
.A1(n_2019),
.A2(n_2011),
.B1(n_2000),
.B2(n_2004),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_2016),
.Y(n_2032)
);

NAND4xp25_ASAP7_75t_L g2033 ( 
.A(n_2021),
.B(n_1993),
.C(n_1992),
.D(n_1928),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_2016),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_2022),
.B(n_2020),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_SL g2036 ( 
.A(n_2017),
.B(n_2011),
.Y(n_2036)
);

OAI211xp5_ASAP7_75t_L g2037 ( 
.A1(n_2023),
.A2(n_1928),
.B(n_1985),
.C(n_1870),
.Y(n_2037)
);

AOI31xp33_ASAP7_75t_L g2038 ( 
.A1(n_2028),
.A2(n_2026),
.A3(n_2025),
.B(n_2024),
.Y(n_2038)
);

AOI211xp5_ASAP7_75t_L g2039 ( 
.A1(n_2027),
.A2(n_1834),
.B(n_1920),
.C(n_1855),
.Y(n_2039)
);

AOI31xp33_ASAP7_75t_L g2040 ( 
.A1(n_2030),
.A2(n_1917),
.A3(n_1901),
.B(n_1898),
.Y(n_2040)
);

NOR2xp33_ASAP7_75t_L g2041 ( 
.A(n_2037),
.B(n_2033),
.Y(n_2041)
);

AOI321xp33_ASAP7_75t_L g2042 ( 
.A1(n_2029),
.A2(n_2036),
.A3(n_2031),
.B1(n_2034),
.B2(n_2032),
.C(n_2035),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_2028),
.B(n_1902),
.Y(n_2043)
);

NOR3xp33_ASAP7_75t_L g2044 ( 
.A(n_2038),
.B(n_1929),
.C(n_1894),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_2043),
.Y(n_2045)
);

AOI222xp33_ASAP7_75t_L g2046 ( 
.A1(n_2042),
.A2(n_1924),
.B1(n_1929),
.B2(n_1888),
.C1(n_1901),
.C2(n_1898),
.Y(n_2046)
);

AOI22xp5_ASAP7_75t_L g2047 ( 
.A1(n_2039),
.A2(n_1855),
.B1(n_1922),
.B2(n_1909),
.Y(n_2047)
);

AOI222xp33_ASAP7_75t_L g2048 ( 
.A1(n_2041),
.A2(n_1888),
.B1(n_1894),
.B2(n_1898),
.C1(n_1901),
.C2(n_1922),
.Y(n_2048)
);

AOI22xp5_ASAP7_75t_L g2049 ( 
.A1(n_2040),
.A2(n_1909),
.B1(n_1862),
.B2(n_1867),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_2041),
.B(n_1880),
.Y(n_2050)
);

NAND4xp75_ASAP7_75t_L g2051 ( 
.A(n_2045),
.B(n_1873),
.C(n_1888),
.D(n_1894),
.Y(n_2051)
);

NAND4xp75_ASAP7_75t_L g2052 ( 
.A(n_2050),
.B(n_1873),
.C(n_1789),
.D(n_1903),
.Y(n_2052)
);

XNOR2xp5_ASAP7_75t_L g2053 ( 
.A(n_2044),
.B(n_1893),
.Y(n_2053)
);

INVx2_ASAP7_75t_SL g2054 ( 
.A(n_2049),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2046),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_2047),
.Y(n_2056)
);

NOR3xp33_ASAP7_75t_L g2057 ( 
.A(n_2055),
.B(n_2048),
.C(n_1903),
.Y(n_2057)
);

NOR2x1p5_ASAP7_75t_L g2058 ( 
.A(n_2056),
.B(n_1913),
.Y(n_2058)
);

NAND3xp33_ASAP7_75t_L g2059 ( 
.A(n_2054),
.B(n_1882),
.C(n_1866),
.Y(n_2059)
);

NOR4xp75_ASAP7_75t_SL g2060 ( 
.A(n_2057),
.B(n_2053),
.C(n_2051),
.D(n_2054),
.Y(n_2060)
);

HB1xp67_ASAP7_75t_L g2061 ( 
.A(n_2060),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_2061),
.Y(n_2062)
);

AOI21xp33_ASAP7_75t_L g2063 ( 
.A1(n_2061),
.A2(n_2059),
.B(n_2058),
.Y(n_2063)
);

HB1xp67_ASAP7_75t_L g2064 ( 
.A(n_2062),
.Y(n_2064)
);

OAI22xp5_ASAP7_75t_L g2065 ( 
.A1(n_2063),
.A2(n_2052),
.B1(n_1893),
.B2(n_1862),
.Y(n_2065)
);

OAI21xp5_ASAP7_75t_SL g2066 ( 
.A1(n_2064),
.A2(n_2065),
.B(n_1868),
.Y(n_2066)
);

OAI21xp5_ASAP7_75t_L g2067 ( 
.A1(n_2064),
.A2(n_1866),
.B(n_1862),
.Y(n_2067)
);

AOI22xp33_ASAP7_75t_SL g2068 ( 
.A1(n_2067),
.A2(n_1867),
.B1(n_1879),
.B2(n_1877),
.Y(n_2068)
);

OAI21xp5_ASAP7_75t_L g2069 ( 
.A1(n_2066),
.A2(n_1867),
.B(n_1866),
.Y(n_2069)
);

OAI21xp33_ASAP7_75t_L g2070 ( 
.A1(n_2069),
.A2(n_1880),
.B(n_1867),
.Y(n_2070)
);

OAI22xp33_ASAP7_75t_L g2071 ( 
.A1(n_2070),
.A2(n_2068),
.B1(n_1866),
.B2(n_1879),
.Y(n_2071)
);

AOI221xp5_ASAP7_75t_L g2072 ( 
.A1(n_2071),
.A2(n_1879),
.B1(n_1877),
.B2(n_1851),
.C(n_1876),
.Y(n_2072)
);

AOI211xp5_ASAP7_75t_L g2073 ( 
.A1(n_2072),
.A2(n_1719),
.B(n_1879),
.C(n_1877),
.Y(n_2073)
);


endmodule