module fake_jpeg_14112_n_138 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_138);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_138;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_27),
.B(n_26),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

OR2x2_ASAP7_75t_SL g53 ( 
.A(n_16),
.B(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_63),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_47),
.Y(n_70)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_64),
.A2(n_56),
.B1(n_45),
.B2(n_48),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_73),
.B1(n_48),
.B2(n_46),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_49),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_43),
.B1(n_52),
.B2(n_45),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_53),
.B(n_54),
.C(n_51),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_2),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_79),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_66),
.Y(n_80)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

AND2x6_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_81),
.B(n_86),
.Y(n_104)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_78),
.A2(n_42),
.B(n_54),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_96),
.B1(n_20),
.B2(n_33),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_88),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_80),
.A2(n_44),
.B(n_2),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_94),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_72),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_1),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_22),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_90),
.B(n_6),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_75),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_96),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_77),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_23),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_71),
.A2(n_21),
.B1(n_38),
.B2(n_34),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_3),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_105),
.Y(n_115)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_101),
.A2(n_102),
.B1(n_106),
.B2(n_8),
.Y(n_120)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_96),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_83),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_108),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_109),
.A2(n_110),
.B(n_114),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_7),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_8),
.Y(n_118)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_112),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_18),
.C(n_10),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_118),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_120),
.A2(n_106),
.B1(n_102),
.B2(n_101),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_104),
.B(n_11),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_121),
.A2(n_124),
.B(n_123),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_13),
.C(n_15),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_127),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_116),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_128),
.A2(n_113),
.B1(n_119),
.B2(n_103),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_115),
.C(n_121),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_131),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_129),
.B(n_115),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_126),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_SL g136 ( 
.A1(n_135),
.A2(n_122),
.B(n_107),
.C(n_30),
.Y(n_136)
);

FAx1_ASAP7_75t_SL g137 ( 
.A(n_136),
.B(n_28),
.CI(n_29),
.CON(n_137),
.SN(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_31),
.Y(n_138)
);


endmodule