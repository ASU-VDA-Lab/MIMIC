module fake_netlist_5_2205_n_1820 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1820);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1820;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_1809;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_336;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_88),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_64),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_43),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_70),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_31),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_167),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_152),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_49),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_92),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_80),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_13),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_45),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_63),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_19),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_55),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_18),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_57),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_97),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_55),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_98),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_37),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_49),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_131),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_84),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_158),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_144),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_69),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_128),
.Y(n_200)
);

BUFx2_ASAP7_75t_SL g201 ( 
.A(n_114),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_74),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_109),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_40),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_134),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_66),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_48),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_73),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_36),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_96),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_156),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_37),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_62),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_155),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_138),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_6),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_75),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_43),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_124),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_5),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_76),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_87),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_135),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_1),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_23),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_38),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_125),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_56),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_53),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_10),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_46),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_0),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_129),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_107),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_81),
.Y(n_235)
);

BUFx10_ASAP7_75t_L g236 ( 
.A(n_13),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_4),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_65),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_19),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_146),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_12),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_50),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_104),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_149),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_168),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_119),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_48),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_24),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_45),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_91),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_118),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_154),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_44),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_4),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_117),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_62),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_54),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_102),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_126),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_169),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_115),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_160),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_40),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_12),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_110),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_36),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_22),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_95),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_50),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_17),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_139),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_162),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_41),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_111),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_120),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_22),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_116),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_16),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_39),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_58),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_133),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_5),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_42),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_136),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_148),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_44),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_27),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_68),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_61),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_105),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_113),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_6),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_8),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_147),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_132),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_143),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_8),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_141),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_26),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_72),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_59),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_14),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_52),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_7),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_163),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_2),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_79),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_33),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_99),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_170),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_153),
.Y(n_311)
);

BUFx10_ASAP7_75t_L g312 ( 
.A(n_23),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_60),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_58),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_157),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_42),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_32),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_11),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_20),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_31),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_56),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_93),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_54),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_166),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_145),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_32),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_16),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_1),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_15),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_94),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_123),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_51),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_27),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_30),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_150),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_30),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_130),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_15),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_100),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_25),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_173),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_237),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_237),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_308),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_308),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_175),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_282),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_217),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_213),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_213),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_213),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_304),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_248),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_171),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_248),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_248),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_302),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_178),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_180),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_181),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_302),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_246),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_302),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_183),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_304),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_210),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_272),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_183),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_243),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_184),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_207),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_195),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_207),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_265),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_209),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_196),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_192),
.B(n_0),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_197),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_209),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_192),
.B(n_2),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_198),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_216),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_199),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_177),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_200),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_202),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_205),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_216),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_206),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_218),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_316),
.Y(n_391)
);

NOR2xp67_ASAP7_75t_L g392 ( 
.A(n_218),
.B(n_3),
.Y(n_392)
);

NOR2xp67_ASAP7_75t_L g393 ( 
.A(n_225),
.B(n_3),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_225),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_229),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_316),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_335),
.B(n_7),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_208),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_214),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_215),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_222),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_229),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_233),
.Y(n_403)
);

NOR2xp67_ASAP7_75t_L g404 ( 
.A(n_230),
.B(n_9),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_240),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_230),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_232),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_244),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_232),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_242),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_242),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_247),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_247),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_245),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_250),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_176),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_254),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_254),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_257),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_257),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_270),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_251),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_255),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_369),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_380),
.B(n_335),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_369),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_369),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_369),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_377),
.B(n_190),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_369),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_350),
.B(n_210),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_369),
.Y(n_432)
);

AND2x6_ASAP7_75t_L g433 ( 
.A(n_384),
.B(n_243),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_384),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_364),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_364),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_371),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_391),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_342),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_342),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_343),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_343),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_347),
.B(n_231),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_350),
.B(n_210),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_344),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_344),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_345),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_349),
.B(n_177),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_345),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_371),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_373),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_349),
.B(n_259),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_351),
.B(n_260),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_373),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_366),
.Y(n_455)
);

AND2x6_ASAP7_75t_L g456 ( 
.A(n_397),
.B(n_243),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_375),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_375),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_351),
.B(n_261),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_379),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_379),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_353),
.B(n_185),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_348),
.A2(n_182),
.B1(n_226),
.B2(n_313),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_353),
.B(n_271),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_382),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_382),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_388),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_388),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_390),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_355),
.B(n_185),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_374),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_390),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_355),
.B(n_172),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_394),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_356),
.B(n_274),
.Y(n_475)
);

NAND2xp33_ASAP7_75t_R g476 ( 
.A(n_365),
.B(n_179),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_394),
.Y(n_477)
);

AND2x6_ASAP7_75t_L g478 ( 
.A(n_366),
.B(n_243),
.Y(n_478)
);

CKINVDCx8_ASAP7_75t_R g479 ( 
.A(n_347),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_395),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_395),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_396),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_402),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_402),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_406),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_406),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_409),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_409),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_410),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_356),
.B(n_172),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_410),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_392),
.B(n_231),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_411),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_357),
.B(n_221),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_411),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_412),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_412),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_413),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_413),
.Y(n_499)
);

NAND2xp33_ASAP7_75t_R g500 ( 
.A(n_429),
.B(n_365),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_435),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_461),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_429),
.B(n_341),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_454),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_428),
.Y(n_505)
);

AND3x2_ASAP7_75t_L g506 ( 
.A(n_443),
.B(n_352),
.C(n_235),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_455),
.B(n_346),
.Y(n_507)
);

INVxp67_ASAP7_75t_SL g508 ( 
.A(n_455),
.Y(n_508)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_438),
.B(n_416),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_454),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_455),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_425),
.A2(n_389),
.B1(n_399),
.B2(n_398),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_425),
.B(n_358),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_461),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_455),
.B(n_359),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_454),
.Y(n_516)
);

NOR2x1p5_ASAP7_75t_L g517 ( 
.A(n_452),
.B(n_354),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_461),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_461),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_458),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_461),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_461),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_461),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_479),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_456),
.B(n_360),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_461),
.Y(n_526)
);

NAND3xp33_ASAP7_75t_L g527 ( 
.A(n_476),
.B(n_453),
.C(n_452),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_456),
.A2(n_393),
.B1(n_404),
.B2(n_287),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_458),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_453),
.B(n_370),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_458),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_448),
.B(n_357),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_456),
.B(n_372),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_460),
.Y(n_534)
);

NAND3xp33_ASAP7_75t_L g535 ( 
.A(n_476),
.B(n_378),
.C(n_376),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_460),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_466),
.Y(n_537)
);

NAND2xp33_ASAP7_75t_L g538 ( 
.A(n_456),
.B(n_243),
.Y(n_538)
);

AND2x6_ASAP7_75t_L g539 ( 
.A(n_448),
.B(n_243),
.Y(n_539)
);

INVxp67_ASAP7_75t_SL g540 ( 
.A(n_432),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_478),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_456),
.B(n_381),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_466),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_460),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_466),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_435),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_443),
.B(n_383),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_428),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_456),
.B(n_385),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_436),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_466),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_466),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_479),
.B(n_386),
.Y(n_553)
);

OAI22xp33_ASAP7_75t_L g554 ( 
.A1(n_459),
.A2(n_194),
.B1(n_249),
.B2(n_174),
.Y(n_554)
);

INVxp67_ASAP7_75t_SL g555 ( 
.A(n_432),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_466),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_479),
.B(n_387),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_474),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_466),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_474),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_466),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_487),
.Y(n_562)
);

OAI22xp33_ASAP7_75t_SL g563 ( 
.A1(n_492),
.A2(n_252),
.B1(n_296),
.B2(n_298),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_436),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_459),
.B(n_400),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_487),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_478),
.Y(n_567)
);

NAND3xp33_ASAP7_75t_L g568 ( 
.A(n_464),
.B(n_403),
.C(n_401),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_474),
.Y(n_569)
);

INVxp67_ASAP7_75t_SL g570 ( 
.A(n_432),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_448),
.B(n_361),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_487),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_488),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_428),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_464),
.B(n_405),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_431),
.B(n_361),
.Y(n_576)
);

NAND2xp33_ASAP7_75t_L g577 ( 
.A(n_456),
.B(n_311),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_488),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_456),
.B(n_415),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_456),
.B(n_423),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_475),
.B(n_408),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_437),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_475),
.B(n_422),
.Y(n_583)
);

NAND2xp33_ASAP7_75t_SL g584 ( 
.A(n_492),
.B(n_186),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_431),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_428),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_487),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_437),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_471),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_467),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_431),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_467),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_456),
.A2(n_279),
.B1(n_270),
.B2(n_278),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_488),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_438),
.B(n_414),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_491),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_491),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_491),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_482),
.B(n_363),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_493),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_444),
.B(n_281),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_463),
.B(n_362),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_456),
.B(n_363),
.Y(n_603)
);

AND3x2_ASAP7_75t_L g604 ( 
.A(n_482),
.B(n_235),
.C(n_221),
.Y(n_604)
);

AND2x6_ASAP7_75t_L g605 ( 
.A(n_462),
.B(n_311),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_444),
.B(n_284),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_444),
.B(n_285),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_473),
.B(n_288),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_473),
.B(n_291),
.Y(n_609)
);

INVx5_ASAP7_75t_L g610 ( 
.A(n_433),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_469),
.A2(n_188),
.B1(n_189),
.B2(n_187),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_462),
.B(n_294),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_473),
.A2(n_292),
.B1(n_329),
.B2(n_278),
.Y(n_613)
);

INVx4_ASAP7_75t_L g614 ( 
.A(n_478),
.Y(n_614)
);

INVx1_ASAP7_75t_SL g615 ( 
.A(n_471),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_493),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_493),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_428),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_462),
.B(n_300),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_495),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_472),
.B(n_367),
.Y(n_621)
);

XOR2xp5_ASAP7_75t_L g622 ( 
.A(n_463),
.B(n_293),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_470),
.Y(n_623)
);

AND3x2_ASAP7_75t_L g624 ( 
.A(n_470),
.B(n_295),
.C(n_277),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_487),
.Y(n_625)
);

BUFx4f_ASAP7_75t_L g626 ( 
.A(n_478),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_470),
.B(n_309),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_473),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_473),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_473),
.B(n_315),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_490),
.B(n_322),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_469),
.A2(n_266),
.B1(n_264),
.B2(n_267),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_495),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_487),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_428),
.Y(n_635)
);

INVxp33_ASAP7_75t_L g636 ( 
.A(n_483),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_478),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_487),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_483),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_487),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_472),
.B(n_368),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_495),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_490),
.B(n_417),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_490),
.B(n_417),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_472),
.B(n_407),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_472),
.B(n_324),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_497),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_490),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_485),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_490),
.A2(n_314),
.B1(n_330),
.B2(n_339),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_490),
.B(n_203),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_485),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_504),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_503),
.B(n_331),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_513),
.B(n_337),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_629),
.Y(n_656)
);

NAND2xp33_ASAP7_75t_L g657 ( 
.A(n_528),
.B(n_311),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_629),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_585),
.B(n_472),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_510),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_585),
.B(n_477),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_516),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_516),
.Y(n_663)
);

AOI221xp5_ASAP7_75t_L g664 ( 
.A1(n_554),
.A2(n_584),
.B1(n_622),
.B2(n_292),
.C(n_329),
.Y(n_664)
);

NAND2xp33_ASAP7_75t_L g665 ( 
.A(n_539),
.B(n_311),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_520),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_591),
.B(n_477),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_591),
.B(n_530),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_520),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_529),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_565),
.B(n_575),
.Y(n_671)
);

NAND2x1_ASAP7_75t_L g672 ( 
.A(n_541),
.B(n_567),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_641),
.B(n_477),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_527),
.B(n_477),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_535),
.B(n_494),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_623),
.B(n_477),
.Y(n_676)
);

BUFx6f_ASAP7_75t_SL g677 ( 
.A(n_576),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_532),
.B(n_486),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_576),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_615),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_529),
.B(n_486),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_531),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_636),
.B(n_494),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_531),
.B(n_486),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_534),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_534),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_536),
.B(n_486),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_618),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_536),
.Y(n_689)
);

NAND3xp33_ASAP7_75t_L g690 ( 
.A(n_500),
.B(n_193),
.C(n_191),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_544),
.B(n_486),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_544),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_621),
.B(n_494),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_SL g694 ( 
.A(n_524),
.B(n_231),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_558),
.B(n_494),
.Y(n_695)
);

OR2x6_ASAP7_75t_L g696 ( 
.A(n_507),
.B(n_201),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_558),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_501),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_R g699 ( 
.A(n_524),
.B(n_204),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_576),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_560),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_546),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_568),
.B(n_494),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_550),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_618),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_560),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_515),
.B(n_494),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_628),
.A2(n_201),
.B1(n_258),
.B2(n_262),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_650),
.B(n_489),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_569),
.B(n_489),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_569),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_573),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_573),
.B(n_489),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_581),
.B(n_489),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_578),
.Y(n_715)
);

OAI221xp5_ASAP7_75t_L g716 ( 
.A1(n_613),
.A2(n_340),
.B1(n_279),
.B2(n_287),
.C(n_334),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_578),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_594),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_594),
.B(n_489),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_651),
.A2(n_277),
.B1(n_295),
.B2(n_305),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_596),
.B(n_489),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_564),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_SL g723 ( 
.A(n_595),
.B(n_231),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_651),
.A2(n_593),
.B1(n_644),
.B2(n_643),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_596),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_582),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_588),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_597),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_597),
.Y(n_729)
);

NAND2xp33_ASAP7_75t_L g730 ( 
.A(n_539),
.B(n_311),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_598),
.Y(n_731)
);

NAND2x1_ASAP7_75t_L g732 ( 
.A(n_541),
.B(n_567),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_598),
.B(n_489),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_600),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_600),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_616),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_583),
.B(n_489),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_589),
.Y(n_738)
);

NAND2xp33_ASAP7_75t_L g739 ( 
.A(n_539),
.B(n_311),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_511),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_628),
.B(n_203),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_599),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_616),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_617),
.Y(n_744)
);

NAND3xp33_ASAP7_75t_L g745 ( 
.A(n_584),
.B(n_220),
.C(n_212),
.Y(n_745)
);

INVx4_ASAP7_75t_L g746 ( 
.A(n_626),
.Y(n_746)
);

OR2x2_ASAP7_75t_SL g747 ( 
.A(n_509),
.B(n_334),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_617),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_620),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_620),
.B(n_450),
.Y(n_750)
);

NAND2x1_ASAP7_75t_L g751 ( 
.A(n_541),
.B(n_432),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_626),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_626),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_547),
.B(n_224),
.Y(n_754)
);

INVx3_ASAP7_75t_L g755 ( 
.A(n_618),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_633),
.B(n_450),
.Y(n_756)
);

INVxp67_ASAP7_75t_L g757 ( 
.A(n_509),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_R g758 ( 
.A(n_589),
.B(n_228),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_633),
.B(n_450),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_642),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_642),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_639),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_647),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_647),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_643),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_648),
.B(n_211),
.Y(n_766)
);

INVxp67_ASAP7_75t_L g767 ( 
.A(n_611),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_532),
.B(n_450),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_553),
.B(n_557),
.Y(n_769)
);

AND2x6_ASAP7_75t_SL g770 ( 
.A(n_622),
.B(n_340),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_512),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_571),
.B(n_451),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_506),
.B(n_239),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_SL g774 ( 
.A(n_639),
.B(n_236),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_571),
.B(n_451),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_648),
.B(n_211),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_645),
.B(n_241),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_511),
.B(n_451),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_645),
.B(n_253),
.Y(n_779)
);

INVx8_ASAP7_75t_L g780 ( 
.A(n_539),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_590),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_606),
.B(n_219),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_592),
.B(n_451),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_649),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_652),
.B(n_457),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_644),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_508),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_612),
.B(n_457),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_601),
.B(n_256),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_502),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_619),
.B(n_457),
.Y(n_791)
);

NAND2xp33_ASAP7_75t_SL g792 ( 
.A(n_517),
.B(n_219),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_651),
.Y(n_793)
);

AND2x6_ASAP7_75t_SL g794 ( 
.A(n_602),
.B(n_418),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_607),
.B(n_269),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_627),
.B(n_457),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_502),
.Y(n_797)
);

OR2x6_ASAP7_75t_L g798 ( 
.A(n_603),
.B(n_223),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_540),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_514),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_555),
.B(n_465),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_514),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_570),
.B(n_465),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_563),
.B(n_223),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_646),
.B(n_465),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_525),
.B(n_533),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_632),
.B(n_497),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_542),
.A2(n_305),
.B1(n_296),
.B2(n_290),
.Y(n_808)
);

INVx2_ASAP7_75t_SL g809 ( 
.A(n_624),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_518),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_549),
.B(n_273),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_604),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_518),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_519),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_579),
.B(n_497),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_519),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_580),
.B(n_276),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_608),
.B(n_280),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_567),
.B(n_227),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_539),
.A2(n_227),
.B1(n_234),
.B2(n_238),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_609),
.B(n_234),
.Y(n_821)
);

BUFx2_ASAP7_75t_L g822 ( 
.A(n_539),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_614),
.B(n_238),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_672),
.A2(n_732),
.B(n_746),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_671),
.B(n_668),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_752),
.B(n_614),
.Y(n_826)
);

OR2x2_ASAP7_75t_L g827 ( 
.A(n_757),
.B(n_602),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_777),
.B(n_505),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_653),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_672),
.A2(n_637),
.B(n_614),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_779),
.B(n_505),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_752),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_680),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_752),
.B(n_637),
.Y(n_834)
);

O2A1O1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_767),
.A2(n_674),
.B(n_676),
.C(n_742),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_754),
.A2(n_538),
.B(n_577),
.C(n_630),
.Y(n_836)
);

AOI21x1_ASAP7_75t_L g837 ( 
.A1(n_675),
.A2(n_631),
.B(n_522),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_678),
.B(n_740),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_656),
.B(n_505),
.Y(n_839)
);

NOR2xp67_ASAP7_75t_L g840 ( 
.A(n_738),
.B(n_521),
.Y(n_840)
);

O2A1O1Ixp33_ASAP7_75t_SL g841 ( 
.A1(n_709),
.A2(n_298),
.B(n_252),
.C(n_307),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_740),
.Y(n_842)
);

CKINVDCx14_ASAP7_75t_R g843 ( 
.A(n_699),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_732),
.A2(n_637),
.B(n_577),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_678),
.B(n_548),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_746),
.A2(n_538),
.B(n_618),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_818),
.A2(n_258),
.B(n_262),
.C(n_268),
.Y(n_847)
);

AOI21x1_ASAP7_75t_L g848 ( 
.A1(n_707),
.A2(n_522),
.B(n_521),
.Y(n_848)
);

NOR2xp67_ASAP7_75t_L g849 ( 
.A(n_690),
.B(n_745),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_815),
.A2(n_526),
.B(n_523),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_762),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_815),
.A2(n_526),
.B(n_523),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_746),
.A2(n_618),
.B(n_574),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_799),
.B(n_548),
.Y(n_854)
);

A2O1A1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_765),
.A2(n_310),
.B(n_325),
.C(n_307),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_673),
.A2(n_543),
.B(n_537),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_781),
.B(n_548),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_752),
.B(n_537),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_752),
.B(n_543),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_812),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_792),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_806),
.A2(n_586),
.B(n_574),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_781),
.B(n_784),
.Y(n_863)
);

NAND2xp33_ASAP7_75t_SL g864 ( 
.A(n_677),
.B(n_758),
.Y(n_864)
);

BUFx2_ASAP7_75t_L g865 ( 
.A(n_747),
.Y(n_865)
);

AOI21x1_ASAP7_75t_L g866 ( 
.A1(n_703),
.A2(n_551),
.B(n_545),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_666),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_753),
.A2(n_586),
.B(n_574),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_753),
.A2(n_635),
.B(n_586),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_L g870 ( 
.A1(n_659),
.A2(n_640),
.B(n_638),
.Y(n_870)
);

NOR3xp33_ASAP7_75t_L g871 ( 
.A(n_664),
.B(n_771),
.C(n_773),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_658),
.B(n_723),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_753),
.A2(n_635),
.B(n_638),
.Y(n_873)
);

O2A1O1Ixp5_ASAP7_75t_L g874 ( 
.A1(n_782),
.A2(n_640),
.B(n_545),
.C(n_634),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_679),
.B(n_418),
.Y(n_875)
);

A2O1A1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_765),
.A2(n_268),
.B(n_310),
.C(n_290),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_753),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_769),
.A2(n_679),
.B1(n_700),
.B2(n_786),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_753),
.A2(n_635),
.B(n_634),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_788),
.A2(n_796),
.B(n_791),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_812),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_724),
.A2(n_275),
.B1(n_325),
.B2(n_572),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_784),
.B(n_551),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_700),
.B(n_552),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_694),
.B(n_283),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_805),
.A2(n_625),
.B(n_552),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_786),
.B(n_556),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_789),
.A2(n_795),
.B(n_792),
.C(n_821),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_807),
.B(n_236),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_693),
.A2(n_625),
.B(n_556),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_787),
.B(n_559),
.Y(n_891)
);

OAI22xp5_ASAP7_75t_L g892 ( 
.A1(n_793),
.A2(n_275),
.B1(n_587),
.B2(n_572),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_661),
.A2(n_559),
.B(n_561),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_807),
.B(n_236),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_669),
.B(n_670),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_768),
.A2(n_587),
.B(n_566),
.Y(n_896)
);

O2A1O1Ixp33_ASAP7_75t_SL g897 ( 
.A1(n_819),
.A2(n_561),
.B(n_566),
.C(n_562),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_793),
.A2(n_562),
.B1(n_498),
.B2(n_333),
.Y(n_898)
);

INVxp67_ASAP7_75t_L g899 ( 
.A(n_683),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_772),
.A2(n_610),
.B(n_428),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_670),
.B(n_605),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_780),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_775),
.A2(n_610),
.B(n_428),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_771),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_778),
.A2(n_610),
.B(n_432),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_667),
.A2(n_605),
.B(n_426),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_682),
.A2(n_498),
.B1(n_289),
.B2(n_303),
.Y(n_907)
);

AND2x4_ASAP7_75t_SL g908 ( 
.A(n_696),
.B(n_236),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_682),
.B(n_605),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_685),
.B(n_605),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_801),
.A2(n_803),
.B(n_823),
.Y(n_911)
);

NOR3xp33_ASAP7_75t_L g912 ( 
.A(n_654),
.B(n_498),
.C(n_336),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_695),
.A2(n_610),
.B(n_434),
.Y(n_913)
);

A2O1A1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_821),
.A2(n_439),
.B(n_440),
.C(n_442),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_747),
.B(n_286),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_681),
.A2(n_605),
.B(n_427),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_751),
.A2(n_657),
.B(n_780),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_677),
.Y(n_918)
);

O2A1O1Ixp33_ASAP7_75t_SL g919 ( 
.A1(n_684),
.A2(n_440),
.B(n_449),
.C(n_442),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_751),
.A2(n_610),
.B(n_434),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_698),
.B(n_297),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_657),
.A2(n_434),
.B(n_430),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_660),
.B(n_434),
.Y(n_923)
);

NAND3xp33_ASAP7_75t_L g924 ( 
.A(n_655),
.B(n_306),
.C(n_320),
.Y(n_924)
);

AOI22xp5_ASAP7_75t_L g925 ( 
.A1(n_714),
.A2(n_737),
.B1(n_811),
.B2(n_817),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_685),
.A2(n_299),
.B1(n_332),
.B2(n_338),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_702),
.B(n_301),
.Y(n_927)
);

OAI321xp33_ASAP7_75t_L g928 ( 
.A1(n_716),
.A2(n_421),
.A3(n_420),
.B1(n_419),
.B2(n_442),
.C(n_439),
.Y(n_928)
);

AOI21xp33_ASAP7_75t_L g929 ( 
.A1(n_696),
.A2(n_317),
.B(n_318),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_687),
.A2(n_605),
.B(n_430),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_809),
.B(n_419),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_662),
.B(n_434),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_780),
.A2(n_434),
.B(n_430),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_704),
.B(n_319),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_686),
.B(n_465),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_662),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_821),
.B(n_468),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_691),
.A2(n_430),
.B(n_427),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_710),
.A2(n_719),
.B(n_713),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_686),
.B(n_468),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_689),
.B(n_468),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_774),
.B(n_468),
.Y(n_942)
);

AO21x1_ASAP7_75t_L g943 ( 
.A1(n_689),
.A2(n_441),
.B(n_439),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_712),
.B(n_729),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_712),
.B(n_480),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_780),
.A2(n_434),
.B(n_424),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_663),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_721),
.A2(n_424),
.B(n_426),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_722),
.A2(n_441),
.B(n_440),
.C(n_449),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_726),
.B(n_263),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_729),
.B(n_480),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_731),
.B(n_480),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_688),
.A2(n_434),
.B(n_424),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_731),
.B(n_480),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_809),
.B(n_420),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_688),
.A2(n_755),
.B(n_705),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_688),
.A2(n_424),
.B(n_426),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_734),
.B(n_481),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_705),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_734),
.A2(n_321),
.B1(n_323),
.B2(n_326),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_736),
.B(n_481),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_727),
.B(n_481),
.Y(n_962)
);

O2A1O1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_741),
.A2(n_499),
.B(n_496),
.C(n_484),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_733),
.A2(n_426),
.B(n_427),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_705),
.A2(n_427),
.B(n_496),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_736),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_755),
.A2(n_499),
.B(n_496),
.Y(n_967)
);

AOI33xp33_ASAP7_75t_L g968 ( 
.A1(n_708),
.A2(n_421),
.A3(n_449),
.B1(n_441),
.B2(n_481),
.B3(n_496),
.Y(n_968)
);

NAND2x1p5_ASAP7_75t_L g969 ( 
.A(n_822),
.B(n_499),
.Y(n_969)
);

O2A1O1Ixp33_ASAP7_75t_SL g970 ( 
.A1(n_804),
.A2(n_499),
.B(n_484),
.C(n_447),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_794),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_743),
.B(n_484),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_743),
.B(n_484),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_761),
.B(n_447),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_696),
.A2(n_478),
.B1(n_447),
.B2(n_446),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_766),
.B(n_327),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_755),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_783),
.A2(n_447),
.B(n_446),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_761),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_696),
.B(n_263),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_822),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_692),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_776),
.B(n_445),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_692),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_697),
.B(n_445),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_697),
.B(n_446),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_785),
.A2(n_446),
.B(n_445),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_750),
.A2(n_478),
.B(n_433),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_756),
.A2(n_445),
.B(n_478),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_759),
.A2(n_445),
.B(n_478),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_790),
.A2(n_445),
.B(n_478),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_677),
.B(n_328),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_701),
.A2(n_263),
.B(n_312),
.C(n_11),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_701),
.B(n_445),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_790),
.A2(n_445),
.B(n_478),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_706),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_706),
.B(n_9),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_711),
.Y(n_998)
);

BUFx3_ASAP7_75t_L g999 ( 
.A(n_798),
.Y(n_999)
);

AND3x1_ASAP7_75t_L g1000 ( 
.A(n_770),
.B(n_263),
.C(n_312),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_711),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_797),
.A2(n_433),
.B(n_67),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_798),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_715),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_797),
.A2(n_433),
.B(n_108),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_800),
.A2(n_433),
.B(n_106),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_715),
.B(n_433),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_829),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_984),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_825),
.B(n_717),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_984),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_843),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_888),
.A2(n_749),
.B1(n_717),
.B2(n_718),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_917),
.A2(n_730),
.B(n_739),
.Y(n_1014)
);

AO22x1_ASAP7_75t_L g1015 ( 
.A1(n_904),
.A2(n_760),
.B1(n_763),
.B2(n_718),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_880),
.A2(n_730),
.B(n_739),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_999),
.B(n_918),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_872),
.B(n_725),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_861),
.A2(n_763),
.B(n_725),
.C(n_728),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_826),
.A2(n_665),
.B(n_744),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_861),
.B(n_728),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_832),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_872),
.B(n_735),
.Y(n_1023)
);

INVx5_ASAP7_75t_L g1024 ( 
.A(n_832),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_835),
.A2(n_764),
.B(n_748),
.C(n_749),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_981),
.Y(n_1026)
);

AOI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_871),
.A2(n_798),
.B1(n_764),
.B2(n_735),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_899),
.B(n_744),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_851),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_871),
.A2(n_760),
.B(n_748),
.C(n_816),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_976),
.A2(n_810),
.B(n_808),
.C(n_813),
.Y(n_1031)
);

AND2x2_ASAP7_75t_SL g1032 ( 
.A(n_912),
.B(n_665),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_976),
.A2(n_810),
.B(n_814),
.C(n_813),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_838),
.B(n_814),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_826),
.A2(n_802),
.B(n_800),
.Y(n_1035)
);

O2A1O1Ixp5_ASAP7_75t_L g1036 ( 
.A1(n_943),
.A2(n_802),
.B(n_798),
.C(n_720),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_847),
.A2(n_820),
.B(n_312),
.C(n_17),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_925),
.A2(n_103),
.B1(n_165),
.B2(n_164),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_834),
.A2(n_433),
.B(n_161),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_834),
.A2(n_433),
.B(n_151),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_833),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_889),
.B(n_894),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_824),
.A2(n_911),
.B(n_846),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_899),
.B(n_312),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_878),
.A2(n_142),
.B1(n_137),
.B2(n_127),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_844),
.A2(n_831),
.B(n_828),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_875),
.B(n_10),
.Y(n_1047)
);

OAI22x1_ASAP7_75t_L g1048 ( 
.A1(n_885),
.A2(n_14),
.B1(n_18),
.B2(n_20),
.Y(n_1048)
);

AO21x1_ASAP7_75t_L g1049 ( 
.A1(n_997),
.A2(n_21),
.B(n_24),
.Y(n_1049)
);

NOR3xp33_ASAP7_75t_SL g1050 ( 
.A(n_1003),
.B(n_21),
.C(n_25),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_875),
.B(n_26),
.Y(n_1051)
);

NOR2x1_ASAP7_75t_L g1052 ( 
.A(n_924),
.B(n_849),
.Y(n_1052)
);

INVxp67_ASAP7_75t_L g1053 ( 
.A(n_865),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_842),
.B(n_28),
.Y(n_1054)
);

BUFx8_ASAP7_75t_L g1055 ( 
.A(n_860),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_830),
.A2(n_852),
.B(n_850),
.Y(n_1056)
);

INVxp67_ASAP7_75t_L g1057 ( 
.A(n_833),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_SL g1058 ( 
.A1(n_912),
.A2(n_433),
.B(n_122),
.C(n_121),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_853),
.A2(n_433),
.B(n_112),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_845),
.A2(n_433),
.B(n_101),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_827),
.B(n_28),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_929),
.A2(n_29),
.B(n_33),
.C(n_34),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_881),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_862),
.A2(n_939),
.B(n_869),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_915),
.B(n_29),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_918),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_842),
.B(n_867),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_936),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_947),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_885),
.A2(n_34),
.B(n_35),
.C(n_38),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_915),
.A2(n_35),
.B(n_39),
.C(n_41),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_981),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_966),
.B(n_46),
.Y(n_1073)
);

AOI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_882),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_832),
.B(n_77),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_979),
.B(n_47),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_840),
.B(n_53),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_981),
.B(n_82),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_981),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_895),
.B(n_57),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_832),
.B(n_83),
.Y(n_1081)
);

BUFx2_ASAP7_75t_L g1082 ( 
.A(n_931),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_950),
.B(n_59),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_868),
.A2(n_85),
.B(n_89),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_877),
.B(n_71),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_944),
.A2(n_78),
.B1(n_86),
.B2(n_90),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_982),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_931),
.B(n_60),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_955),
.B(n_61),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_955),
.B(n_921),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_863),
.A2(n_836),
.B(n_873),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_877),
.B(n_996),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_921),
.B(n_927),
.Y(n_1093)
);

BUFx3_ASAP7_75t_L g1094 ( 
.A(n_992),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_927),
.B(n_934),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_934),
.B(n_997),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_998),
.A2(n_1004),
.B1(n_1001),
.B2(n_937),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_887),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_980),
.A2(n_864),
.B1(n_942),
.B2(n_992),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_839),
.B(n_968),
.Y(n_1100)
);

INVx4_ASAP7_75t_L g1101 ( 
.A(n_877),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_877),
.B(n_908),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_879),
.A2(n_856),
.B(n_858),
.Y(n_1103)
);

O2A1O1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_855),
.A2(n_876),
.B(n_993),
.C(n_914),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_971),
.B(n_839),
.Y(n_1105)
);

O2A1O1Ixp5_ASAP7_75t_L g1106 ( 
.A1(n_858),
.A2(n_859),
.B(n_837),
.C(n_870),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_891),
.B(n_935),
.Y(n_1107)
);

AO21x1_ASAP7_75t_L g1108 ( 
.A1(n_859),
.A2(n_961),
.B(n_941),
.Y(n_1108)
);

INVx5_ASAP7_75t_L g1109 ( 
.A(n_902),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_883),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_893),
.A2(n_890),
.B(n_857),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_986),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_940),
.B(n_945),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_906),
.A2(n_956),
.B(n_909),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1000),
.B(n_926),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_951),
.B(n_952),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_949),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_969),
.A2(n_902),
.B1(n_901),
.B2(n_910),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_954),
.B(n_972),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_959),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_960),
.B(n_907),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_958),
.B(n_973),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_898),
.A2(n_962),
.B(n_919),
.C(n_892),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_900),
.A2(n_903),
.B(n_854),
.Y(n_1124)
);

INVx1_ASAP7_75t_SL g1125 ( 
.A(n_983),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_959),
.Y(n_1126)
);

OR2x6_ASAP7_75t_L g1127 ( 
.A(n_902),
.B(n_969),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_896),
.A2(n_874),
.B(n_886),
.C(n_930),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_884),
.B(n_977),
.Y(n_1129)
);

AOI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_884),
.A2(n_975),
.B1(n_1007),
.B2(n_977),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_916),
.A2(n_974),
.B(n_985),
.Y(n_1131)
);

OR2x2_ASAP7_75t_L g1132 ( 
.A(n_985),
.B(n_932),
.Y(n_1132)
);

NOR2xp67_ASAP7_75t_SL g1133 ( 
.A(n_902),
.B(n_928),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_959),
.B(n_977),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_959),
.B(n_977),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_994),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_841),
.A2(n_970),
.B(n_932),
.C(n_923),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_866),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_938),
.A2(n_964),
.B(n_948),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_933),
.A2(n_946),
.B(n_913),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_897),
.A2(n_920),
.B(n_905),
.Y(n_1141)
);

O2A1O1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_963),
.A2(n_967),
.B(n_988),
.C(n_965),
.Y(n_1142)
);

INVx4_ASAP7_75t_L g1143 ( 
.A(n_848),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_989),
.B(n_990),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_978),
.B(n_987),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_957),
.A2(n_922),
.B(n_953),
.C(n_991),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_995),
.B(n_1002),
.Y(n_1147)
);

A2O1A1Ixp33_ASAP7_75t_SL g1148 ( 
.A1(n_1005),
.A2(n_671),
.B(n_817),
.C(n_811),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1006),
.B(n_671),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_825),
.B(n_671),
.Y(n_1150)
);

AOI21xp33_ASAP7_75t_L g1151 ( 
.A1(n_976),
.A2(n_671),
.B(n_500),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_888),
.B(n_671),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_984),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_832),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_843),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_889),
.B(n_894),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_889),
.B(n_894),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_917),
.A2(n_753),
.B(n_752),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1008),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_1022),
.Y(n_1160)
);

CKINVDCx12_ASAP7_75t_R g1161 ( 
.A(n_1088),
.Y(n_1161)
);

AO31x2_ASAP7_75t_L g1162 ( 
.A1(n_1128),
.A2(n_1013),
.A3(n_1056),
.B(n_1108),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1150),
.B(n_1093),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1087),
.Y(n_1164)
);

INVx4_ASAP7_75t_L g1165 ( 
.A(n_1024),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1042),
.B(n_1156),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1158),
.A2(n_1152),
.B(n_1149),
.Y(n_1167)
);

INVx3_ASAP7_75t_SL g1168 ( 
.A(n_1012),
.Y(n_1168)
);

AOI21xp33_ASAP7_75t_L g1169 ( 
.A1(n_1096),
.A2(n_1095),
.B(n_1151),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1046),
.A2(n_1043),
.B(n_1139),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1036),
.A2(n_1091),
.B(n_1150),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1140),
.A2(n_1141),
.B(n_1124),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1016),
.A2(n_1148),
.B(n_1014),
.Y(n_1173)
);

AOI21xp33_ASAP7_75t_L g1174 ( 
.A1(n_1065),
.A2(n_1121),
.B(n_1032),
.Y(n_1174)
);

OA21x2_ASAP7_75t_L g1175 ( 
.A1(n_1106),
.A2(n_1036),
.B(n_1064),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_SL g1176 ( 
.A(n_1065),
.B(n_1121),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_1090),
.A2(n_1061),
.B1(n_1157),
.B2(n_1115),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_1063),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1148),
.A2(n_1111),
.B(n_1107),
.Y(n_1179)
);

NOR2xp67_ASAP7_75t_SL g1180 ( 
.A(n_1024),
.B(n_1109),
.Y(n_1180)
);

AND2x6_ASAP7_75t_L g1181 ( 
.A(n_1022),
.B(n_1154),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_1022),
.Y(n_1182)
);

O2A1O1Ixp33_ASAP7_75t_SL g1183 ( 
.A1(n_1075),
.A2(n_1085),
.B(n_1058),
.C(n_1030),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_1155),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1103),
.A2(n_1116),
.B(n_1113),
.Y(n_1185)
);

NOR3xp33_ASAP7_75t_L g1186 ( 
.A(n_1061),
.B(n_1052),
.C(n_1071),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1119),
.A2(n_1122),
.B(n_1020),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1068),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1069),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1105),
.B(n_1094),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1105),
.B(n_1057),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1098),
.B(n_1021),
.Y(n_1192)
);

OA22x2_ASAP7_75t_L g1193 ( 
.A1(n_1048),
.A2(n_1053),
.B1(n_1082),
.B2(n_1057),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1041),
.Y(n_1194)
);

INVx6_ASAP7_75t_L g1195 ( 
.A(n_1055),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1114),
.A2(n_1147),
.B(n_1131),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1144),
.A2(n_1145),
.B(n_1031),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1106),
.A2(n_1025),
.B(n_1033),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1104),
.A2(n_1099),
.B(n_1027),
.C(n_1044),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1044),
.A2(n_1021),
.B(n_1028),
.C(n_1032),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_1029),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1035),
.A2(n_1144),
.B(n_1118),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1010),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1009),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1083),
.B(n_1053),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1019),
.A2(n_1034),
.B(n_1142),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1028),
.B(n_1110),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_SL g1208 ( 
.A1(n_1127),
.A2(n_1038),
.B(n_1045),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1067),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_1055),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1011),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_1127),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1074),
.A2(n_1100),
.B1(n_1080),
.B2(n_1073),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1017),
.B(n_1089),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1066),
.B(n_1051),
.Y(n_1215)
);

INVx1_ASAP7_75t_SL g1216 ( 
.A(n_1054),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1137),
.A2(n_1092),
.B(n_1123),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_R g1218 ( 
.A(n_1026),
.B(n_1072),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_1017),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1112),
.B(n_1136),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1018),
.A2(n_1023),
.B(n_1146),
.Y(n_1221)
);

A2O1A1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1062),
.A2(n_1037),
.B(n_1073),
.C(n_1129),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1047),
.B(n_1102),
.Y(n_1223)
);

INVx2_ASAP7_75t_SL g1224 ( 
.A(n_1026),
.Y(n_1224)
);

AO31x2_ASAP7_75t_L g1225 ( 
.A1(n_1143),
.A2(n_1049),
.A3(n_1117),
.B(n_1129),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1022),
.Y(n_1226)
);

OAI21xp33_ASAP7_75t_L g1227 ( 
.A1(n_1074),
.A2(n_1070),
.B(n_1076),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1077),
.A2(n_1133),
.B(n_1130),
.C(n_1086),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1153),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1024),
.A2(n_1127),
.B(n_1092),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_SL g1231 ( 
.A1(n_1078),
.A2(n_1125),
.B(n_1075),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1024),
.A2(n_1109),
.B(n_1015),
.Y(n_1232)
);

AOI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1134),
.A2(n_1135),
.B(n_1085),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1109),
.A2(n_1138),
.B(n_1084),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1109),
.A2(n_1138),
.B(n_1143),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1081),
.A2(n_1079),
.B1(n_1072),
.B2(n_1097),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1097),
.A2(n_1079),
.B1(n_1132),
.B2(n_1050),
.Y(n_1237)
);

OR2x2_ASAP7_75t_L g1238 ( 
.A(n_1126),
.B(n_1120),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1050),
.A2(n_1058),
.B(n_1039),
.C(n_1040),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1154),
.A2(n_1101),
.B1(n_1120),
.B2(n_1138),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1059),
.A2(n_1060),
.B(n_1138),
.Y(n_1241)
);

INVx1_ASAP7_75t_SL g1242 ( 
.A(n_1154),
.Y(n_1242)
);

O2A1O1Ixp33_ASAP7_75t_SL g1243 ( 
.A1(n_1154),
.A2(n_888),
.B(n_1095),
.C(n_1093),
.Y(n_1243)
);

AOI21xp33_ASAP7_75t_L g1244 ( 
.A1(n_1101),
.A2(n_1096),
.B(n_1095),
.Y(n_1244)
);

AO22x2_ASAP7_75t_L g1245 ( 
.A1(n_1093),
.A2(n_1095),
.B1(n_1096),
.B2(n_1152),
.Y(n_1245)
);

AOI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1152),
.A2(n_1158),
.B(n_1013),
.Y(n_1246)
);

AO31x2_ASAP7_75t_L g1247 ( 
.A1(n_1128),
.A2(n_943),
.A3(n_1013),
.B(n_1056),
.Y(n_1247)
);

NOR3xp33_ASAP7_75t_L g1248 ( 
.A(n_1093),
.B(n_671),
.C(n_1095),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1017),
.B(n_1082),
.Y(n_1249)
);

BUFx12f_ASAP7_75t_L g1250 ( 
.A(n_1012),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1158),
.A2(n_671),
.B(n_752),
.Y(n_1251)
);

BUFx4f_ASAP7_75t_SL g1252 ( 
.A(n_1055),
.Y(n_1252)
);

A2O1A1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1093),
.A2(n_671),
.B(n_1095),
.C(n_1151),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1093),
.A2(n_671),
.B1(n_1095),
.B2(n_1096),
.Y(n_1254)
);

A2O1A1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1093),
.A2(n_671),
.B(n_1095),
.C(n_1151),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1042),
.B(n_1156),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1008),
.Y(n_1257)
);

O2A1O1Ixp33_ASAP7_75t_SL g1258 ( 
.A1(n_1093),
.A2(n_888),
.B(n_1095),
.C(n_1096),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1150),
.B(n_671),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1158),
.A2(n_1140),
.B(n_1043),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_1041),
.Y(n_1261)
);

OA21x2_ASAP7_75t_L g1262 ( 
.A1(n_1106),
.A2(n_1056),
.B(n_1036),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_1042),
.B(n_827),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1008),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1008),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1093),
.A2(n_871),
.B1(n_1095),
.B2(n_671),
.Y(n_1266)
);

NOR2x1_ASAP7_75t_R g1267 ( 
.A(n_1012),
.B(n_524),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1158),
.A2(n_671),
.B(n_752),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1158),
.A2(n_671),
.B(n_752),
.Y(n_1269)
);

AOI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1093),
.A2(n_671),
.B1(n_1095),
.B2(n_871),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1158),
.A2(n_1140),
.B(n_1043),
.Y(n_1271)
);

CKINVDCx20_ASAP7_75t_R g1272 ( 
.A(n_1012),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1008),
.Y(n_1273)
);

A2O1A1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1093),
.A2(n_671),
.B(n_1095),
.C(n_1151),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1093),
.A2(n_1095),
.B(n_671),
.C(n_1151),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1152),
.A2(n_671),
.B(n_1036),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_1127),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1152),
.A2(n_671),
.B(n_1036),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1093),
.B(n_671),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1008),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1150),
.B(n_671),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1008),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1152),
.A2(n_671),
.B(n_1036),
.Y(n_1283)
);

A2O1A1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1093),
.A2(n_671),
.B(n_1095),
.C(n_1151),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1150),
.B(n_671),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1093),
.B(n_671),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1093),
.A2(n_671),
.B1(n_1095),
.B2(n_1096),
.Y(n_1287)
);

O2A1O1Ixp5_ASAP7_75t_SL g1288 ( 
.A1(n_1152),
.A2(n_1144),
.B(n_1151),
.C(n_1145),
.Y(n_1288)
);

OAI21xp33_ASAP7_75t_SL g1289 ( 
.A1(n_1093),
.A2(n_671),
.B(n_1095),
.Y(n_1289)
);

INVx2_ASAP7_75t_SL g1290 ( 
.A(n_1055),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1158),
.A2(n_671),
.B(n_752),
.Y(n_1291)
);

NAND2x1p5_ASAP7_75t_L g1292 ( 
.A(n_1024),
.B(n_1109),
.Y(n_1292)
);

BUFx3_ASAP7_75t_L g1293 ( 
.A(n_1063),
.Y(n_1293)
);

NOR2xp67_ASAP7_75t_L g1294 ( 
.A(n_1012),
.B(n_680),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_SL g1295 ( 
.A(n_1093),
.B(n_1095),
.Y(n_1295)
);

AO32x2_ASAP7_75t_L g1296 ( 
.A1(n_1013),
.A2(n_1143),
.A3(n_882),
.B1(n_1038),
.B2(n_898),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_SL g1297 ( 
.A1(n_1049),
.A2(n_943),
.B(n_1104),
.Y(n_1297)
);

O2A1O1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1093),
.A2(n_1095),
.B(n_671),
.C(n_1151),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1158),
.A2(n_671),
.B(n_752),
.Y(n_1299)
);

AO22x2_ASAP7_75t_L g1300 ( 
.A1(n_1093),
.A2(n_1095),
.B1(n_1096),
.B2(n_1152),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1158),
.A2(n_1140),
.B(n_1043),
.Y(n_1301)
);

AO31x2_ASAP7_75t_L g1302 ( 
.A1(n_1128),
.A2(n_943),
.A3(n_1013),
.B(n_1056),
.Y(n_1302)
);

A2O1A1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_1093),
.A2(n_671),
.B(n_1095),
.C(n_1151),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1008),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1158),
.A2(n_1140),
.B(n_1043),
.Y(n_1305)
);

INVx8_ASAP7_75t_L g1306 ( 
.A(n_1024),
.Y(n_1306)
);

INVx4_ASAP7_75t_L g1307 ( 
.A(n_1024),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1150),
.B(n_671),
.Y(n_1308)
);

INVxp67_ASAP7_75t_L g1309 ( 
.A(n_1041),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_1178),
.Y(n_1310)
);

BUFx10_ASAP7_75t_L g1311 ( 
.A(n_1190),
.Y(n_1311)
);

BUFx8_ASAP7_75t_L g1312 ( 
.A(n_1250),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_1225),
.Y(n_1313)
);

INVx6_ASAP7_75t_L g1314 ( 
.A(n_1306),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1293),
.Y(n_1315)
);

CKINVDCx11_ASAP7_75t_R g1316 ( 
.A(n_1272),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1176),
.A2(n_1174),
.B1(n_1248),
.B2(n_1287),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1306),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1266),
.A2(n_1270),
.B1(n_1285),
.B2(n_1281),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1177),
.A2(n_1191),
.B1(n_1163),
.B2(n_1308),
.Y(n_1320)
);

OAI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1254),
.A2(n_1287),
.B1(n_1259),
.B2(n_1308),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1186),
.A2(n_1223),
.B1(n_1254),
.B2(n_1256),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1174),
.A2(n_1227),
.B1(n_1213),
.B2(n_1169),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_SL g1324 ( 
.A1(n_1213),
.A2(n_1193),
.B1(n_1259),
.B2(n_1289),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1169),
.A2(n_1295),
.B1(n_1263),
.B2(n_1166),
.Y(n_1325)
);

CKINVDCx6p67_ASAP7_75t_R g1326 ( 
.A(n_1168),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1184),
.Y(n_1327)
);

INVx2_ASAP7_75t_SL g1328 ( 
.A(n_1201),
.Y(n_1328)
);

BUFx4_ASAP7_75t_R g1329 ( 
.A(n_1210),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1245),
.A2(n_1300),
.B1(n_1171),
.B2(n_1297),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1245),
.A2(n_1300),
.B1(n_1216),
.B2(n_1276),
.Y(n_1331)
);

OAI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1192),
.A2(n_1207),
.B1(n_1216),
.B2(n_1220),
.Y(n_1332)
);

BUFx12f_ASAP7_75t_L g1333 ( 
.A(n_1195),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_SL g1334 ( 
.A1(n_1171),
.A2(n_1278),
.B1(n_1283),
.B2(n_1276),
.Y(n_1334)
);

CKINVDCx8_ASAP7_75t_R g1335 ( 
.A(n_1249),
.Y(n_1335)
);

BUFx8_ASAP7_75t_L g1336 ( 
.A(n_1261),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1200),
.A2(n_1199),
.B1(n_1192),
.B2(n_1303),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1159),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1253),
.A2(n_1284),
.B1(n_1274),
.B2(n_1255),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1207),
.A2(n_1215),
.B1(n_1222),
.B2(n_1309),
.Y(n_1340)
);

CKINVDCx11_ASAP7_75t_R g1341 ( 
.A(n_1252),
.Y(n_1341)
);

BUFx12f_ASAP7_75t_L g1342 ( 
.A(n_1195),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1275),
.B(n_1298),
.Y(n_1343)
);

BUFx10_ASAP7_75t_L g1344 ( 
.A(n_1290),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1278),
.A2(n_1283),
.B1(n_1244),
.B2(n_1209),
.Y(n_1345)
);

INVx2_ASAP7_75t_SL g1346 ( 
.A(n_1194),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1228),
.A2(n_1220),
.B1(n_1236),
.B2(n_1231),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1203),
.B(n_1214),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1244),
.A2(n_1205),
.B1(n_1237),
.B2(n_1164),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_SL g1350 ( 
.A1(n_1237),
.A2(n_1198),
.B1(n_1273),
.B2(n_1264),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1288),
.A2(n_1258),
.B(n_1221),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1257),
.Y(n_1352)
);

CKINVDCx11_ASAP7_75t_R g1353 ( 
.A(n_1267),
.Y(n_1353)
);

OAI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1265),
.A2(n_1304),
.B1(n_1282),
.B2(n_1280),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1188),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1306),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1219),
.B(n_1204),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1294),
.B(n_1189),
.Y(n_1358)
);

INVx5_ASAP7_75t_L g1359 ( 
.A(n_1181),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_SL g1360 ( 
.A1(n_1198),
.A2(n_1217),
.B1(n_1262),
.B2(n_1175),
.Y(n_1360)
);

CKINVDCx11_ASAP7_75t_R g1361 ( 
.A(n_1160),
.Y(n_1361)
);

CKINVDCx11_ASAP7_75t_R g1362 ( 
.A(n_1160),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1206),
.A2(n_1211),
.B1(n_1229),
.B2(n_1185),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1262),
.A2(n_1212),
.B1(n_1277),
.B2(n_1197),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1238),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_SL g1366 ( 
.A1(n_1175),
.A2(n_1277),
.B1(n_1232),
.B2(n_1167),
.Y(n_1366)
);

INVx6_ASAP7_75t_L g1367 ( 
.A(n_1165),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1187),
.A2(n_1179),
.B1(n_1196),
.B2(n_1173),
.Y(n_1368)
);

BUFx8_ASAP7_75t_SL g1369 ( 
.A(n_1160),
.Y(n_1369)
);

OAI21xp33_ASAP7_75t_L g1370 ( 
.A1(n_1231),
.A2(n_1239),
.B(n_1208),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1251),
.A2(n_1291),
.B1(n_1269),
.B2(n_1268),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_SL g1372 ( 
.A1(n_1165),
.A2(n_1307),
.B1(n_1240),
.B2(n_1299),
.Y(n_1372)
);

BUFx12f_ASAP7_75t_L g1373 ( 
.A(n_1182),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1224),
.Y(n_1374)
);

OAI21xp5_ASAP7_75t_SL g1375 ( 
.A1(n_1246),
.A2(n_1170),
.B(n_1230),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1218),
.A2(n_1202),
.B1(n_1240),
.B2(n_1234),
.Y(n_1376)
);

OAI22xp33_ASAP7_75t_SL g1377 ( 
.A1(n_1233),
.A2(n_1292),
.B1(n_1242),
.B2(n_1243),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1292),
.A2(n_1242),
.B1(n_1235),
.B2(n_1226),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1226),
.A2(n_1180),
.B1(n_1305),
.B2(n_1271),
.Y(n_1379)
);

AOI22xp5_ASAP7_75t_SL g1380 ( 
.A1(n_1161),
.A2(n_1181),
.B1(n_1183),
.B2(n_1296),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_1181),
.Y(n_1381)
);

BUFx12f_ASAP7_75t_L g1382 ( 
.A(n_1241),
.Y(n_1382)
);

INVx3_ASAP7_75t_L g1383 ( 
.A(n_1247),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1260),
.A2(n_1301),
.B1(n_1172),
.B2(n_1296),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1296),
.A2(n_1162),
.B1(n_1247),
.B2(n_1302),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1247),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1302),
.Y(n_1387)
);

INVx6_ASAP7_75t_L g1388 ( 
.A(n_1162),
.Y(n_1388)
);

CKINVDCx20_ASAP7_75t_R g1389 ( 
.A(n_1162),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1279),
.A2(n_671),
.B1(n_1095),
.B2(n_1093),
.Y(n_1390)
);

BUFx8_ASAP7_75t_L g1391 ( 
.A(n_1250),
.Y(n_1391)
);

INVxp67_ASAP7_75t_SL g1392 ( 
.A(n_1180),
.Y(n_1392)
);

INVx3_ASAP7_75t_L g1393 ( 
.A(n_1306),
.Y(n_1393)
);

BUFx3_ASAP7_75t_L g1394 ( 
.A(n_1178),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1306),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1176),
.A2(n_1065),
.B1(n_1095),
.B2(n_1093),
.Y(n_1396)
);

OAI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1176),
.A2(n_671),
.B1(n_1095),
.B2(n_1093),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1184),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1279),
.A2(n_671),
.B1(n_1095),
.B2(n_1093),
.Y(n_1399)
);

CKINVDCx11_ASAP7_75t_R g1400 ( 
.A(n_1272),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1176),
.A2(n_1065),
.B1(n_1095),
.B2(n_1093),
.Y(n_1401)
);

BUFx10_ASAP7_75t_L g1402 ( 
.A(n_1190),
.Y(n_1402)
);

OAI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1176),
.A2(n_671),
.B1(n_1095),
.B2(n_1093),
.Y(n_1403)
);

OAI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1176),
.A2(n_671),
.B1(n_1095),
.B2(n_1093),
.Y(n_1404)
);

INVx2_ASAP7_75t_SL g1405 ( 
.A(n_1178),
.Y(n_1405)
);

INVx6_ASAP7_75t_L g1406 ( 
.A(n_1306),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_1261),
.Y(n_1407)
);

BUFx12f_ASAP7_75t_L g1408 ( 
.A(n_1250),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_SL g1409 ( 
.A1(n_1176),
.A2(n_723),
.B1(n_1095),
.B2(n_1093),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1261),
.Y(n_1410)
);

BUFx4f_ASAP7_75t_SL g1411 ( 
.A(n_1250),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1184),
.Y(n_1412)
);

CKINVDCx11_ASAP7_75t_R g1413 ( 
.A(n_1272),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1279),
.B(n_1286),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1176),
.A2(n_1065),
.B1(n_1095),
.B2(n_1093),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1176),
.A2(n_723),
.B1(n_1095),
.B2(n_1093),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1279),
.B(n_1286),
.Y(n_1417)
);

INVx4_ASAP7_75t_SL g1418 ( 
.A(n_1181),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1176),
.A2(n_1065),
.B1(n_1095),
.B2(n_1093),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1178),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1176),
.A2(n_671),
.B1(n_1065),
.B2(n_1186),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1306),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1176),
.A2(n_671),
.B1(n_1065),
.B2(n_1186),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1263),
.B(n_1163),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_SL g1425 ( 
.A1(n_1176),
.A2(n_723),
.B1(n_1095),
.B2(n_1093),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_SL g1426 ( 
.A1(n_1270),
.A2(n_602),
.B(n_671),
.Y(n_1426)
);

INVx1_ASAP7_75t_SL g1427 ( 
.A(n_1407),
.Y(n_1427)
);

AOI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1343),
.A2(n_1339),
.B(n_1337),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1387),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1383),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1368),
.A2(n_1384),
.B(n_1371),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1386),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1388),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1381),
.Y(n_1434)
);

AO21x2_ASAP7_75t_L g1435 ( 
.A1(n_1351),
.A2(n_1375),
.B(n_1321),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1334),
.B(n_1389),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1313),
.Y(n_1437)
);

INVx3_ASAP7_75t_L g1438 ( 
.A(n_1382),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1385),
.B(n_1331),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1331),
.B(n_1349),
.Y(n_1440)
);

BUFx4f_ASAP7_75t_SL g1441 ( 
.A(n_1408),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1321),
.B(n_1332),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1334),
.B(n_1350),
.Y(n_1443)
);

INVx2_ASAP7_75t_SL g1444 ( 
.A(n_1359),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1338),
.Y(n_1445)
);

AOI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1347),
.A2(n_1319),
.B(n_1320),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1350),
.B(n_1330),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1352),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1330),
.B(n_1323),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1360),
.B(n_1364),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1355),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1354),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1409),
.A2(n_1416),
.B1(n_1425),
.B2(n_1423),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1360),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1323),
.B(n_1349),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1377),
.Y(n_1456)
);

CKINVDCx6p67_ASAP7_75t_R g1457 ( 
.A(n_1333),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1336),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_SL g1459 ( 
.A(n_1335),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1316),
.Y(n_1460)
);

AOI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1397),
.A2(n_1403),
.B(n_1404),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1379),
.A2(n_1363),
.B(n_1376),
.Y(n_1462)
);

OA21x2_ASAP7_75t_L g1463 ( 
.A1(n_1345),
.A2(n_1370),
.B(n_1317),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1380),
.B(n_1418),
.Y(n_1464)
);

INVxp67_ASAP7_75t_L g1465 ( 
.A(n_1340),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1317),
.B(n_1324),
.Y(n_1466)
);

OR2x6_ASAP7_75t_L g1467 ( 
.A(n_1378),
.B(n_1314),
.Y(n_1467)
);

BUFx6f_ASAP7_75t_L g1468 ( 
.A(n_1395),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1365),
.Y(n_1469)
);

O2A1O1Ixp5_ASAP7_75t_L g1470 ( 
.A1(n_1397),
.A2(n_1404),
.B(n_1403),
.C(n_1399),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1324),
.B(n_1345),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1421),
.A2(n_1356),
.B(n_1393),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1366),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1322),
.B(n_1325),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1348),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1366),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1318),
.A2(n_1356),
.B(n_1393),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1372),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1372),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1390),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1357),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1374),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1424),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_1336),
.Y(n_1484)
);

INVx4_ASAP7_75t_L g1485 ( 
.A(n_1422),
.Y(n_1485)
);

CKINVDCx20_ASAP7_75t_R g1486 ( 
.A(n_1400),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1318),
.A2(n_1396),
.B(n_1419),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1392),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1392),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1396),
.A2(n_1415),
.B(n_1401),
.Y(n_1490)
);

INVxp67_ASAP7_75t_R g1491 ( 
.A(n_1329),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1358),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1409),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1401),
.B(n_1415),
.Y(n_1494)
);

OAI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1470),
.A2(n_1419),
.B(n_1425),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1453),
.A2(n_1416),
.B1(n_1417),
.B2(n_1414),
.Y(n_1496)
);

O2A1O1Ixp33_ASAP7_75t_SL g1497 ( 
.A1(n_1465),
.A2(n_1426),
.B(n_1346),
.C(n_1328),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1477),
.B(n_1422),
.Y(n_1498)
);

NAND2xp33_ASAP7_75t_R g1499 ( 
.A(n_1464),
.B(n_1410),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1436),
.B(n_1454),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1486),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1445),
.Y(n_1502)
);

OAI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1470),
.A2(n_1310),
.B(n_1405),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1445),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1483),
.B(n_1311),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1475),
.B(n_1402),
.Y(n_1506)
);

A2O1A1Ixp33_ASAP7_75t_L g1507 ( 
.A1(n_1461),
.A2(n_1422),
.B(n_1315),
.C(n_1420),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1481),
.B(n_1362),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1436),
.B(n_1361),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1436),
.B(n_1454),
.Y(n_1510)
);

OA21x2_ASAP7_75t_L g1511 ( 
.A1(n_1431),
.A2(n_1367),
.B(n_1314),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1450),
.B(n_1367),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1450),
.B(n_1344),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1450),
.B(n_1344),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1469),
.B(n_1326),
.Y(n_1515)
);

OAI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1465),
.A2(n_1398),
.B(n_1327),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1477),
.B(n_1394),
.Y(n_1517)
);

O2A1O1Ixp33_ASAP7_75t_L g1518 ( 
.A1(n_1442),
.A2(n_1342),
.B(n_1411),
.C(n_1369),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1477),
.B(n_1412),
.Y(n_1519)
);

AOI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1474),
.A2(n_1411),
.B1(n_1353),
.B2(n_1391),
.Y(n_1520)
);

AO21x1_ASAP7_75t_L g1521 ( 
.A1(n_1493),
.A2(n_1373),
.B(n_1406),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1469),
.B(n_1413),
.Y(n_1522)
);

OAI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1446),
.A2(n_1312),
.B(n_1391),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1443),
.B(n_1341),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1475),
.B(n_1312),
.Y(n_1525)
);

AOI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1474),
.A2(n_1466),
.B1(n_1455),
.B2(n_1494),
.Y(n_1526)
);

AO32x2_ASAP7_75t_L g1527 ( 
.A1(n_1444),
.A2(n_1439),
.A3(n_1437),
.B1(n_1485),
.B2(n_1432),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_1428),
.B(n_1446),
.Y(n_1528)
);

OAI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1428),
.A2(n_1490),
.B(n_1442),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1448),
.B(n_1492),
.Y(n_1530)
);

O2A1O1Ixp33_ASAP7_75t_L g1531 ( 
.A1(n_1480),
.A2(n_1466),
.B(n_1471),
.C(n_1456),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1443),
.B(n_1473),
.Y(n_1532)
);

INVx3_ASAP7_75t_L g1533 ( 
.A(n_1438),
.Y(n_1533)
);

A2O1A1Ixp33_ASAP7_75t_L g1534 ( 
.A1(n_1443),
.A2(n_1471),
.B(n_1447),
.C(n_1490),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1478),
.B(n_1479),
.Y(n_1535)
);

OR2x6_ASAP7_75t_L g1536 ( 
.A(n_1467),
.B(n_1462),
.Y(n_1536)
);

O2A1O1Ixp33_ASAP7_75t_L g1537 ( 
.A1(n_1471),
.A2(n_1456),
.B(n_1449),
.C(n_1455),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_1460),
.Y(n_1538)
);

A2O1A1Ixp33_ASAP7_75t_L g1539 ( 
.A1(n_1447),
.A2(n_1490),
.B(n_1449),
.C(n_1494),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1434),
.B(n_1451),
.Y(n_1540)
);

INVx4_ASAP7_75t_SL g1541 ( 
.A(n_1467),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1473),
.B(n_1476),
.Y(n_1542)
);

AO21x1_ASAP7_75t_L g1543 ( 
.A1(n_1488),
.A2(n_1489),
.B(n_1464),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1476),
.B(n_1451),
.Y(n_1544)
);

OR2x6_ASAP7_75t_L g1545 ( 
.A(n_1467),
.B(n_1462),
.Y(n_1545)
);

OAI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1487),
.A2(n_1472),
.B(n_1462),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1451),
.B(n_1435),
.Y(n_1547)
);

OAI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1487),
.A2(n_1472),
.B(n_1463),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1429),
.Y(n_1549)
);

INVx2_ASAP7_75t_SL g1550 ( 
.A(n_1517),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1500),
.B(n_1429),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1547),
.B(n_1439),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1502),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1502),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1500),
.B(n_1429),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1547),
.B(n_1432),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1549),
.Y(n_1557)
);

INVxp67_ASAP7_75t_L g1558 ( 
.A(n_1505),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1540),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1515),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1548),
.B(n_1437),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_1498),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1510),
.B(n_1536),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1495),
.A2(n_1463),
.B1(n_1440),
.B2(n_1464),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1504),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1504),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1536),
.B(n_1545),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1544),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1536),
.B(n_1430),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1496),
.A2(n_1463),
.B1(n_1440),
.B2(n_1464),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1498),
.B(n_1433),
.Y(n_1571)
);

INVx1_ASAP7_75t_SL g1572 ( 
.A(n_1506),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1542),
.B(n_1452),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1542),
.B(n_1452),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1498),
.B(n_1519),
.Y(n_1575)
);

NOR2xp67_ASAP7_75t_L g1576 ( 
.A(n_1533),
.B(n_1438),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1530),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1543),
.Y(n_1578)
);

BUFx5_ASAP7_75t_L g1579 ( 
.A(n_1519),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1527),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1527),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1552),
.B(n_1545),
.Y(n_1582)
);

AOI222xp33_ASAP7_75t_L g1583 ( 
.A1(n_1570),
.A2(n_1534),
.B1(n_1539),
.B2(n_1529),
.C1(n_1532),
.C2(n_1535),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1552),
.B(n_1546),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1553),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1567),
.B(n_1519),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1556),
.B(n_1511),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1553),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1572),
.B(n_1539),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1567),
.B(n_1541),
.Y(n_1590)
);

INVx1_ASAP7_75t_SL g1591 ( 
.A(n_1560),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1554),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1565),
.Y(n_1593)
);

AOI221xp5_ASAP7_75t_L g1594 ( 
.A1(n_1578),
.A2(n_1537),
.B1(n_1531),
.B2(n_1534),
.C(n_1497),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1563),
.B(n_1527),
.Y(n_1595)
);

INVxp67_ASAP7_75t_SL g1596 ( 
.A(n_1578),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1556),
.B(n_1511),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1559),
.B(n_1513),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1566),
.Y(n_1599)
);

BUFx2_ASAP7_75t_L g1600 ( 
.A(n_1562),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1568),
.B(n_1511),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1562),
.B(n_1541),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1550),
.B(n_1513),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1557),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1575),
.B(n_1541),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1575),
.B(n_1514),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1575),
.B(n_1514),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1564),
.A2(n_1463),
.B1(n_1525),
.B2(n_1435),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1566),
.Y(n_1609)
);

NAND2x1_ASAP7_75t_L g1610 ( 
.A(n_1576),
.B(n_1571),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1560),
.A2(n_1435),
.B1(n_1524),
.B2(n_1512),
.Y(n_1611)
);

INVxp67_ASAP7_75t_L g1612 ( 
.A(n_1577),
.Y(n_1612)
);

OAI211xp5_ASAP7_75t_L g1613 ( 
.A1(n_1558),
.A2(n_1526),
.B(n_1497),
.C(n_1503),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1585),
.Y(n_1614)
);

NOR2xp67_ASAP7_75t_L g1615 ( 
.A(n_1601),
.B(n_1580),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1585),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1594),
.A2(n_1435),
.B1(n_1528),
.B2(n_1535),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1588),
.Y(n_1618)
);

INVx2_ASAP7_75t_SL g1619 ( 
.A(n_1610),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1589),
.B(n_1524),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1596),
.B(n_1581),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1601),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1587),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1588),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1587),
.B(n_1580),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1595),
.B(n_1569),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1597),
.B(n_1561),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1600),
.B(n_1551),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1603),
.B(n_1555),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1597),
.B(n_1561),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_SL g1631 ( 
.A(n_1583),
.B(n_1579),
.Y(n_1631)
);

BUFx2_ASAP7_75t_L g1632 ( 
.A(n_1590),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1612),
.B(n_1573),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1592),
.B(n_1574),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1606),
.B(n_1579),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1604),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1606),
.B(n_1579),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1607),
.B(n_1579),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1593),
.Y(n_1639)
);

INVx1_ASAP7_75t_SL g1640 ( 
.A(n_1591),
.Y(n_1640)
);

INVx5_ASAP7_75t_SL g1641 ( 
.A(n_1602),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1622),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1622),
.Y(n_1643)
);

INVx1_ASAP7_75t_SL g1644 ( 
.A(n_1640),
.Y(n_1644)
);

INVx1_ASAP7_75t_SL g1645 ( 
.A(n_1640),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1618),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1622),
.Y(n_1647)
);

NOR2x1_ASAP7_75t_L g1648 ( 
.A(n_1631),
.B(n_1610),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1633),
.B(n_1584),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1633),
.B(n_1584),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1622),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1618),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1641),
.B(n_1586),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1641),
.B(n_1586),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1624),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1641),
.B(n_1586),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1623),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1623),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1624),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1639),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1641),
.B(n_1586),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1627),
.B(n_1582),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1639),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1614),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1628),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1614),
.Y(n_1666)
);

INVxp67_ASAP7_75t_L g1667 ( 
.A(n_1620),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1623),
.Y(n_1668)
);

NOR2xp67_ASAP7_75t_SL g1669 ( 
.A(n_1631),
.B(n_1458),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1617),
.B(n_1598),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1617),
.A2(n_1613),
.B1(n_1608),
.B2(n_1611),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1616),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1623),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1620),
.B(n_1441),
.Y(n_1674)
);

AND2x4_ASAP7_75t_L g1675 ( 
.A(n_1632),
.B(n_1605),
.Y(n_1675)
);

INVxp67_ASAP7_75t_L g1676 ( 
.A(n_1632),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1616),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1621),
.B(n_1599),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1621),
.B(n_1599),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1634),
.B(n_1609),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1628),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1634),
.B(n_1609),
.Y(n_1682)
);

INVx2_ASAP7_75t_SL g1683 ( 
.A(n_1632),
.Y(n_1683)
);

OAI32xp33_ASAP7_75t_L g1684 ( 
.A1(n_1627),
.A2(n_1499),
.A3(n_1509),
.B1(n_1528),
.B2(n_1522),
.Y(n_1684)
);

INVx1_ASAP7_75t_SL g1685 ( 
.A(n_1644),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1648),
.B(n_1641),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1655),
.Y(n_1687)
);

AOI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1671),
.A2(n_1641),
.B1(n_1590),
.B2(n_1499),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1664),
.Y(n_1689)
);

XNOR2xp5_ASAP7_75t_L g1690 ( 
.A(n_1671),
.B(n_1520),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1648),
.B(n_1635),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1644),
.B(n_1645),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1649),
.B(n_1627),
.Y(n_1693)
);

AND2x2_ASAP7_75t_SL g1694 ( 
.A(n_1674),
.B(n_1509),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1664),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1667),
.B(n_1501),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1649),
.B(n_1630),
.Y(n_1697)
);

OAI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1669),
.A2(n_1619),
.B1(n_1523),
.B2(n_1630),
.C(n_1516),
.Y(n_1698)
);

OAI31xp33_ASAP7_75t_L g1699 ( 
.A1(n_1670),
.A2(n_1619),
.A3(n_1507),
.B(n_1630),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1653),
.B(n_1635),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1645),
.B(n_1629),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1669),
.B(n_1629),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1653),
.B(n_1635),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1650),
.B(n_1625),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1650),
.B(n_1629),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1666),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1654),
.B(n_1637),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1665),
.B(n_1625),
.Y(n_1708)
);

AND2x4_ASAP7_75t_L g1709 ( 
.A(n_1675),
.B(n_1619),
.Y(n_1709)
);

NAND2x1p5_ASAP7_75t_L g1710 ( 
.A(n_1683),
.B(n_1602),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1675),
.B(n_1637),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1666),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1672),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1654),
.B(n_1656),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1656),
.B(n_1637),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1676),
.B(n_1628),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1672),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1677),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1661),
.B(n_1638),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1681),
.B(n_1625),
.Y(n_1720)
);

NAND3xp33_ASAP7_75t_L g1721 ( 
.A(n_1699),
.B(n_1683),
.C(n_1652),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1710),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1694),
.B(n_1501),
.Y(n_1723)
);

INVxp67_ASAP7_75t_L g1724 ( 
.A(n_1692),
.Y(n_1724)
);

INVx1_ASAP7_75t_SL g1725 ( 
.A(n_1685),
.Y(n_1725)
);

OAI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1690),
.A2(n_1675),
.B1(n_1661),
.B2(n_1662),
.Y(n_1726)
);

INVx1_ASAP7_75t_SL g1727 ( 
.A(n_1694),
.Y(n_1727)
);

AOI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1690),
.A2(n_1675),
.B1(n_1602),
.B2(n_1590),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1687),
.B(n_1626),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1689),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1695),
.Y(n_1731)
);

AOI221xp5_ASAP7_75t_L g1732 ( 
.A1(n_1688),
.A2(n_1684),
.B1(n_1646),
.B2(n_1652),
.C(n_1663),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1710),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1714),
.B(n_1638),
.Y(n_1734)
);

INVx1_ASAP7_75t_SL g1735 ( 
.A(n_1714),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1709),
.Y(n_1736)
);

AOI32xp33_ASAP7_75t_L g1737 ( 
.A1(n_1691),
.A2(n_1686),
.A3(n_1702),
.B1(n_1698),
.B2(n_1701),
.Y(n_1737)
);

NOR4xp25_ASAP7_75t_L g1738 ( 
.A(n_1696),
.B(n_1659),
.C(n_1646),
.D(n_1660),
.Y(n_1738)
);

O2A1O1Ixp33_ASAP7_75t_L g1739 ( 
.A1(n_1686),
.A2(n_1684),
.B(n_1659),
.C(n_1660),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1706),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1709),
.Y(n_1741)
);

INVxp67_ASAP7_75t_L g1742 ( 
.A(n_1716),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1709),
.B(n_1638),
.Y(n_1743)
);

NOR3xp33_ASAP7_75t_L g1744 ( 
.A(n_1712),
.B(n_1518),
.C(n_1663),
.Y(n_1744)
);

AOI221x1_ASAP7_75t_L g1745 ( 
.A1(n_1713),
.A2(n_1677),
.B1(n_1643),
.B2(n_1642),
.C(n_1647),
.Y(n_1745)
);

OAI32xp33_ASAP7_75t_L g1746 ( 
.A1(n_1691),
.A2(n_1662),
.A3(n_1678),
.B1(n_1679),
.B2(n_1643),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1731),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1736),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1725),
.B(n_1705),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1735),
.B(n_1700),
.Y(n_1750)
);

NAND2xp33_ASAP7_75t_R g1751 ( 
.A(n_1738),
.B(n_1538),
.Y(n_1751)
);

OAI22xp33_ASAP7_75t_L g1752 ( 
.A1(n_1721),
.A2(n_1491),
.B1(n_1693),
.B2(n_1697),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_L g1753 ( 
.A(n_1723),
.B(n_1538),
.Y(n_1753)
);

AOI32xp33_ASAP7_75t_L g1754 ( 
.A1(n_1732),
.A2(n_1703),
.A3(n_1719),
.B1(n_1707),
.B2(n_1700),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1727),
.B(n_1703),
.Y(n_1755)
);

OAI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1739),
.A2(n_1715),
.B(n_1707),
.Y(n_1756)
);

OAI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1728),
.A2(n_1711),
.B1(n_1693),
.B2(n_1697),
.Y(n_1757)
);

AOI21xp33_ASAP7_75t_SL g1758 ( 
.A1(n_1726),
.A2(n_1720),
.B(n_1708),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1724),
.B(n_1715),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1731),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1744),
.A2(n_1718),
.B1(n_1717),
.B2(n_1719),
.Y(n_1761)
);

OAI21xp5_ASAP7_75t_L g1762 ( 
.A1(n_1742),
.A2(n_1711),
.B(n_1708),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1736),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1740),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1740),
.Y(n_1765)
);

INVxp67_ASAP7_75t_L g1766 ( 
.A(n_1741),
.Y(n_1766)
);

AOI21xp33_ASAP7_75t_L g1767 ( 
.A1(n_1751),
.A2(n_1737),
.B(n_1746),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1766),
.B(n_1730),
.Y(n_1768)
);

NOR2x1_ASAP7_75t_L g1769 ( 
.A(n_1752),
.B(n_1741),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1750),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1761),
.B(n_1722),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1748),
.Y(n_1772)
);

OR2x2_ASAP7_75t_L g1773 ( 
.A(n_1755),
.B(n_1729),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1763),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1747),
.Y(n_1775)
);

OAI221xp5_ASAP7_75t_L g1776 ( 
.A1(n_1751),
.A2(n_1722),
.B1(n_1733),
.B2(n_1704),
.C(n_1720),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1752),
.A2(n_1756),
.B(n_1761),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1762),
.Y(n_1778)
);

NAND3xp33_ASAP7_75t_SL g1779 ( 
.A(n_1777),
.B(n_1776),
.C(n_1778),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1770),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1769),
.B(n_1753),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1768),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1768),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_SL g1784 ( 
.A(n_1767),
.B(n_1758),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1771),
.B(n_1759),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1767),
.B(n_1754),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_L g1787 ( 
.A(n_1773),
.B(n_1753),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_SL g1788 ( 
.A(n_1772),
.B(n_1733),
.Y(n_1788)
);

OAI321xp33_ASAP7_75t_L g1789 ( 
.A1(n_1784),
.A2(n_1757),
.A3(n_1774),
.B1(n_1775),
.B2(n_1749),
.C(n_1765),
.Y(n_1789)
);

NAND2xp33_ASAP7_75t_SL g1790 ( 
.A(n_1781),
.B(n_1760),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1779),
.A2(n_1734),
.B1(n_1743),
.B2(n_1711),
.Y(n_1791)
);

NAND5xp2_ASAP7_75t_L g1792 ( 
.A(n_1787),
.B(n_1764),
.C(n_1734),
.D(n_1743),
.E(n_1746),
.Y(n_1792)
);

AOI221xp5_ASAP7_75t_L g1793 ( 
.A1(n_1779),
.A2(n_1704),
.B1(n_1642),
.B2(n_1643),
.C(n_1647),
.Y(n_1793)
);

AOI221x1_ASAP7_75t_L g1794 ( 
.A1(n_1790),
.A2(n_1780),
.B1(n_1783),
.B2(n_1782),
.C(n_1786),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1791),
.Y(n_1795)
);

A2O1A1Ixp33_ASAP7_75t_L g1796 ( 
.A1(n_1789),
.A2(n_1785),
.B(n_1788),
.C(n_1458),
.Y(n_1796)
);

NAND4xp25_ASAP7_75t_L g1797 ( 
.A(n_1792),
.B(n_1745),
.C(n_1484),
.D(n_1458),
.Y(n_1797)
);

NOR3xp33_ASAP7_75t_L g1798 ( 
.A(n_1793),
.B(n_1484),
.C(n_1427),
.Y(n_1798)
);

AOI32xp33_ASAP7_75t_L g1799 ( 
.A1(n_1789),
.A2(n_1745),
.A3(n_1484),
.B1(n_1651),
.B2(n_1647),
.Y(n_1799)
);

NOR3xp33_ASAP7_75t_L g1800 ( 
.A(n_1795),
.B(n_1457),
.C(n_1427),
.Y(n_1800)
);

AND2x4_ASAP7_75t_L g1801 ( 
.A(n_1794),
.B(n_1678),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1797),
.Y(n_1802)
);

NAND4xp75_ASAP7_75t_L g1803 ( 
.A(n_1796),
.B(n_1457),
.C(n_1642),
.D(n_1651),
.Y(n_1803)
);

NOR2x1_ASAP7_75t_L g1804 ( 
.A(n_1799),
.B(n_1651),
.Y(n_1804)
);

OAI221xp5_ASAP7_75t_SL g1805 ( 
.A1(n_1802),
.A2(n_1798),
.B1(n_1800),
.B2(n_1803),
.C(n_1801),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1804),
.A2(n_1658),
.B(n_1657),
.Y(n_1806)
);

NAND2x1p5_ASAP7_75t_L g1807 ( 
.A(n_1804),
.B(n_1457),
.Y(n_1807)
);

NAND4xp75_ASAP7_75t_L g1808 ( 
.A(n_1806),
.B(n_1658),
.C(n_1657),
.D(n_1673),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1808),
.Y(n_1809)
);

XOR2xp5_ASAP7_75t_L g1810 ( 
.A(n_1809),
.B(n_1807),
.Y(n_1810)
);

AOI22x1_ASAP7_75t_L g1811 ( 
.A1(n_1809),
.A2(n_1805),
.B1(n_1491),
.B2(n_1668),
.Y(n_1811)
);

AND2x4_ASAP7_75t_SL g1812 ( 
.A(n_1810),
.B(n_1657),
.Y(n_1812)
);

AOI22x1_ASAP7_75t_L g1813 ( 
.A1(n_1811),
.A2(n_1673),
.B1(n_1668),
.B2(n_1658),
.Y(n_1813)
);

OAI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1813),
.A2(n_1668),
.B1(n_1673),
.B2(n_1679),
.Y(n_1814)
);

OAI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1812),
.A2(n_1682),
.B1(n_1680),
.B2(n_1459),
.Y(n_1815)
);

AOI21xp33_ASAP7_75t_L g1816 ( 
.A1(n_1815),
.A2(n_1682),
.B(n_1680),
.Y(n_1816)
);

AOI21xp5_ASAP7_75t_L g1817 ( 
.A1(n_1816),
.A2(n_1814),
.B(n_1508),
.Y(n_1817)
);

XNOR2xp5_ASAP7_75t_L g1818 ( 
.A(n_1817),
.B(n_1459),
.Y(n_1818)
);

AOI22xp33_ASAP7_75t_L g1819 ( 
.A1(n_1818),
.A2(n_1615),
.B1(n_1482),
.B2(n_1636),
.Y(n_1819)
);

AOI211xp5_ASAP7_75t_L g1820 ( 
.A1(n_1819),
.A2(n_1521),
.B(n_1615),
.C(n_1468),
.Y(n_1820)
);


endmodule