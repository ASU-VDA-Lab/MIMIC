module real_jpeg_31826_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_0),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_0),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_0),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_0),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_1),
.A2(n_29),
.B1(n_34),
.B2(n_35),
.Y(n_28)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_1),
.A2(n_34),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g245 ( 
.A1(n_1),
.A2(n_34),
.B1(n_246),
.B2(n_249),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_1),
.A2(n_34),
.B1(n_299),
.B2(n_302),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_3),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_4),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_4),
.Y(n_118)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_4),
.Y(n_153)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_4),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_5),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_5),
.Y(n_96)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_5),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_5),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

AO22x2_ASAP7_75t_L g60 ( 
.A1(n_7),
.A2(n_61),
.B1(n_65),
.B2(n_66),
.Y(n_60)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_7),
.A2(n_65),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_7),
.A2(n_65),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_7),
.A2(n_65),
.B1(n_232),
.B2(n_234),
.Y(n_231)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_8),
.Y(n_110)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_8),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_9),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_9),
.A2(n_42),
.B1(n_134),
.B2(n_137),
.Y(n_133)
);

AO22x1_ASAP7_75t_SL g143 ( 
.A1(n_9),
.A2(n_42),
.B1(n_144),
.B2(n_146),
.Y(n_143)
);

AOI22x1_ASAP7_75t_SL g215 ( 
.A1(n_9),
.A2(n_42),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

NAND2xp33_ASAP7_75t_SL g268 ( 
.A(n_9),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_9),
.B(n_102),
.Y(n_291)
);

OAI32xp33_ASAP7_75t_L g313 ( 
.A1(n_9),
.A2(n_179),
.A3(n_314),
.B1(n_318),
.B2(n_325),
.Y(n_313)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_10),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_11),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_11),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_11),
.A2(n_178),
.B1(n_375),
.B2(n_379),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_365),
.Y(n_12)
);

AO21x1_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_237),
.B(n_363),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_199),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_15),
.B(n_199),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_141),
.C(n_172),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_16),
.B(n_361),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_57),
.Y(n_16)
);

MAJx2_ASAP7_75t_L g236 ( 
.A(n_17),
.B(n_58),
.C(n_105),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_37),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_18),
.B(n_387),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_28),
.Y(n_18)
);

NOR2x1p5_ASAP7_75t_L g48 ( 
.A(n_19),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_19),
.Y(n_167)
);

AO22x2_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_22),
.B1(n_24),
.B2(n_26),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_20),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_22),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_25),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_25),
.Y(n_264)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_28),
.B(n_48),
.Y(n_206)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_36),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_48),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_42),
.B(n_43),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_42),
.B(n_167),
.Y(n_166)
);

AOI32xp33_ASAP7_75t_L g260 ( 
.A1(n_42),
.A2(n_261),
.A3(n_265),
.B1(n_267),
.B2(n_268),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_42),
.B(n_326),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_R g337 ( 
.A(n_42),
.B(n_107),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_42),
.B(n_344),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_43),
.Y(n_189)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_44),
.Y(n_210)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_45),
.Y(n_192)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_48),
.B(n_208),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_53),
.B2(n_55),
.Y(n_49)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_52),
.Y(n_186)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_104),
.B1(n_105),
.B2(n_140),
.Y(n_57)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_58),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_97),
.Y(n_58)
);

NAND2x1_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_69),
.Y(n_59)
);

AND2x4_ASAP7_75t_L g170 ( 
.A(n_60),
.B(n_102),
.Y(n_170)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_63),
.Y(n_217)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_69),
.B(n_98),
.Y(n_171)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2x1_ASAP7_75t_L g256 ( 
.A(n_70),
.B(n_215),
.Y(n_256)
);

AOI21x1_ASAP7_75t_L g384 ( 
.A1(n_70),
.A2(n_215),
.B(n_385),
.Y(n_384)
);

AO21x2_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_79),
.B(n_86),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g267 ( 
.A(n_79),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_89),
.B1(n_92),
.B2(n_95),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_88),
.Y(n_251)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_96),
.Y(n_271)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_96),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_97),
.B(n_255),
.Y(n_254)
);

NAND2xp33_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_102),
.Y(n_97)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_102),
.B(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_102),
.Y(n_385)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_105),
.Y(n_104)
);

OA21x2_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_119),
.B(n_133),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_106),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_106),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_106),
.B(n_133),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_106),
.B(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_120),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_111),
.B1(n_114),
.B2(n_117),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_109),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_112),
.Y(n_342)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_118),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_119),
.B(n_133),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_119),
.B(n_231),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_119),
.B(n_245),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_123),
.B1(n_126),
.B2(n_131),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_130),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_130),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx5_ASAP7_75t_L g321 ( 
.A(n_135),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_141),
.B(n_172),
.Y(n_361)
);

MAJx2_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_165),
.C(n_168),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_142),
.A2(n_165),
.B1(n_166),
.B2(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_142),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_148),
.B(n_154),
.Y(n_142)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_143),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_143),
.B(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_148),
.B(n_160),
.Y(n_181)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_148),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_148),
.B(n_298),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.Y(n_148)
);

AO21x2_ASAP7_75t_L g272 ( 
.A1(n_149),
.A2(n_226),
.B(n_273),
.Y(n_272)
);

INVx4_ASAP7_75t_SL g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_155),
.A2(n_176),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_155),
.B(n_297),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_160),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx2_ASAP7_75t_SL g303 ( 
.A(n_162),
.Y(n_303)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_167),
.Y(n_211)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_168),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_182),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_173),
.A2(n_202),
.B(n_203),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_176),
.B(n_181),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_180),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_181),
.B(n_348),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_181),
.B(n_294),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_190),
.Y(n_182)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_187),
.B(n_189),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

NAND3xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.C(n_195),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_SL g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_223),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_200),
.B(n_224),
.C(n_236),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_201),
.B(n_205),
.C(n_222),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_212),
.B1(n_221),
.B2(n_222),
.Y(n_204)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_212),
.Y(n_222)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVxp67_ASAP7_75t_SL g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_236),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_225),
.B(n_228),
.Y(n_388)
);

OAI21xp33_ASAP7_75t_L g347 ( 
.A1(n_226),
.A2(n_273),
.B(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_229),
.B(n_244),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_230),
.B(n_279),
.Y(n_289)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_233),
.Y(n_235)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

AO21x1_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_358),
.B(n_362),
.Y(n_238)
);

OAI21x1_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_285),
.B(n_357),
.Y(n_239)
);

NOR2x1_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_275),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_241),
.B(n_275),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_253),
.C(n_257),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_243),
.B(n_254),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_252),
.Y(n_243)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_252),
.B(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_305),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_272),
.B2(n_274),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

NOR2x1_ASAP7_75t_SL g280 ( 
.A(n_260),
.B(n_272),
.Y(n_280)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_271),
.Y(n_380)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_272),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_281),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_280),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_277),
.B(n_280),
.C(n_281),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

XOR2x2_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

AOI21x1_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_306),
.B(n_356),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_304),
.Y(n_286)
);

NOR2xp67_ASAP7_75t_SL g356 ( 
.A(n_287),
.B(n_304),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_290),
.C(n_292),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_289),
.A2(n_290),
.B1(n_291),
.B2(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_289),
.Y(n_310)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_309),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_297),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_298),
.B(n_345),
.Y(n_348)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_333),
.B(n_355),
.Y(n_306)
);

NOR2xp67_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_311),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_308),
.B(n_311),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_331),
.Y(n_311)
);

NAND2xp33_ASAP7_75t_SL g352 ( 
.A(n_312),
.B(n_332),
.Y(n_352)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_313),
.B(n_331),
.Y(n_353)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_322),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

AOI21x1_ASAP7_75t_SL g333 ( 
.A1(n_334),
.A2(n_350),
.B(n_354),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_338),
.B(n_349),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_336),
.B(n_337),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_347),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_343),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

BUFx4f_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

NAND3xp33_ASAP7_75t_SL g350 ( 
.A(n_351),
.B(n_352),
.C(n_353),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_351),
.A2(n_352),
.B(n_353),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

NOR2xp67_ASAP7_75t_L g362 ( 
.A(n_359),
.B(n_360),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_390),
.Y(n_365)
);

INVxp33_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

NAND2x1_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_389),
.Y(n_367)
);

OR2x2_ASAP7_75t_L g391 ( 
.A(n_368),
.B(n_389),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_382),
.Y(n_370)
);

XNOR2x2_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_381),
.Y(n_371)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx3_ASAP7_75t_SL g377 ( 
.A(n_378),
.Y(n_377)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_388),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_386),
.Y(n_383)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);


endmodule