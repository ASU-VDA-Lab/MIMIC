module fake_jpeg_27950_n_45 (n_3, n_2, n_1, n_0, n_4, n_5, n_45);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_45;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx4_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

BUFx2_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx8_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_1),
.B(n_5),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_10),
.B(n_3),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_18),
.A2(n_23),
.B1(n_13),
.B2(n_12),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_3),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_19),
.A2(n_21),
.B(n_22),
.Y(n_27)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

OAI22xp33_ASAP7_75t_L g28 ( 
.A1(n_20),
.A2(n_6),
.B1(n_8),
.B2(n_11),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_11),
.A2(n_4),
.B1(n_0),
.B2(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_15),
.A2(n_14),
.B(n_22),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_30),
.B(n_17),
.C(n_13),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_29),
.B1(n_20),
.B2(n_23),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_6),
.C(n_8),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_32),
.B1(n_33),
.B2(n_21),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_18),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_24),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_25),
.C(n_27),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_38),
.Y(n_40)
);

MAJx2_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_31),
.C(n_28),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_9),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_37),
.B(n_4),
.Y(n_42)
);

AO21x1_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_41),
.B(n_39),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);


endmodule