module real_jpeg_10406_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_215;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_187;
wire n_75;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_2),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_2),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_2),
.A2(n_51),
.B1(n_52),
.B2(n_69),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_3),
.A2(n_51),
.B1(n_52),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_3),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_80),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_3),
.A2(n_65),
.B1(n_66),
.B2(n_80),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_4),
.A2(n_65),
.B1(n_66),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_4),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_5),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_5),
.B(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_5),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_5),
.A2(n_183),
.B(n_207),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_7),
.A2(n_65),
.B1(n_66),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_7),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_8),
.A2(n_37),
.B1(n_51),
.B2(n_52),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_8),
.A2(n_37),
.B1(n_65),
.B2(n_66),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_9),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_9),
.A2(n_29),
.B1(n_51),
.B2(n_52),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_9),
.A2(n_29),
.B1(n_65),
.B2(n_66),
.Y(n_173)
);

BUFx6f_ASAP7_75t_SL g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g84 ( 
.A(n_12),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_44),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_13),
.A2(n_44),
.B1(n_65),
.B2(n_66),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_13),
.A2(n_44),
.B1(n_51),
.B2(n_52),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_15),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_15),
.A2(n_31),
.B(n_33),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_61),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_15),
.B(n_99),
.Y(n_138)
);

A2O1A1O1Ixp25_ASAP7_75t_L g150 ( 
.A1(n_15),
.A2(n_52),
.B(n_82),
.C(n_151),
.D(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_15),
.B(n_52),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_15),
.B(n_50),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_L g185 ( 
.A1(n_15),
.A2(n_70),
.B(n_166),
.Y(n_185)
);

A2O1A1O1Ixp25_ASAP7_75t_L g198 ( 
.A1(n_15),
.A2(n_32),
.B(n_46),
.C(n_54),
.D(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_15),
.B(n_32),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_16),
.A2(n_65),
.B1(n_66),
.B2(n_73),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_16),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_16),
.A2(n_51),
.B1(n_52),
.B2(n_73),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_127),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_126),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_103),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_21),
.B(n_103),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_74),
.C(n_89),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_22),
.B(n_143),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_58),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_41),
.B1(n_42),
.B2(n_57),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_24),
.Y(n_57)
);

OAI21xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B(n_35),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_25),
.A2(n_30),
.B1(n_39),
.B2(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_30),
.B(n_34),
.C(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_34),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_27),
.A2(n_34),
.B(n_61),
.C(n_62),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_30),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_47),
.B(n_49),
.C(n_50),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_47),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_36),
.B(n_99),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_38),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_41),
.B(n_57),
.C(n_58),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_45),
.B(n_53),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_43),
.A2(n_45),
.B1(n_56),
.B2(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_46),
.B(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_48),
.B(n_51),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_49),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_50),
.Y(n_56)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

O2A1O1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_51),
.A2(n_83),
.B(n_85),
.C(n_86),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_83),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_52),
.A2(n_199),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_55),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_56),
.A2(n_116),
.B(n_118),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_56),
.A2(n_102),
.B(n_118),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_61),
.B(n_88),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_61),
.B(n_71),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_63),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_64),
.A2(n_70),
.B1(n_71),
.B2(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_66),
.B1(n_83),
.B2(n_84),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_65),
.B(n_83),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_65),
.B(n_187),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_66),
.A2(n_85),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

BUFx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_70),
.A2(n_71),
.B1(n_76),
.B2(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_70),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_70),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_70),
.B(n_168),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_71),
.A2(n_173),
.B(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_74),
.B(n_89),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_78),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_81),
.B1(n_87),
.B2(n_88),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_88),
.B(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_87),
.B1(n_88),
.B2(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_81),
.A2(n_88),
.B1(n_163),
.B2(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_81),
.A2(n_197),
.B(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_82),
.B(n_93),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_86),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_88),
.B(n_94),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_88),
.A2(n_92),
.B(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_95),
.C(n_100),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_90),
.A2(n_91),
.B1(n_100),
.B2(n_101),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_124),
.B2(n_125),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_112),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_120),
.B1(n_121),
.B2(n_123),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_115),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_124),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_144),
.B(n_228),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_142),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_129),
.B(n_142),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.C(n_134),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_130),
.B(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_132),
.A2(n_134),
.B1(n_135),
.B2(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_132),
.Y(n_226)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.C(n_139),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_136),
.A2(n_137),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_138),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_141),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_222),
.B(n_227),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_210),
.B(n_221),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_191),
.B(n_209),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_169),
.B(n_190),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_157),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_149),
.B(n_157),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_150),
.A2(n_153),
.B1(n_154),
.B2(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_150),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_151),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_152),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_164),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_162),
.C(n_164),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_165),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_178),
.B(n_189),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_176),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_171),
.B(n_176),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_184),
.B(n_188),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_180),
.B(n_181),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_192),
.B(n_193),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_202),
.B2(n_208),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_198),
.B1(n_200),
.B2(n_201),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_196),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_198),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_201),
.C(n_208),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_202),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_206),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_211),
.B(n_212),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_218),
.C(n_219),
.Y(n_223)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_214),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_223),
.B(n_224),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);


endmodule