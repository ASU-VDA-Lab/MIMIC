module fake_netlist_1_12020_n_662 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_662);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_662;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g89 ( .A(n_12), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_77), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_16), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_63), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_54), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_52), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_40), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_81), .Y(n_96) );
CKINVDCx14_ASAP7_75t_R g97 ( .A(n_22), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_76), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_73), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_38), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_18), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_62), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_7), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_61), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_67), .Y(n_105) );
INVxp67_ASAP7_75t_SL g106 ( .A(n_72), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_15), .Y(n_107) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_17), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_36), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_26), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_83), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_69), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_24), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_14), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_46), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_33), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_28), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_5), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_25), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_6), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_29), .Y(n_121) );
INVxp33_ASAP7_75t_L g122 ( .A(n_84), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_20), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_3), .Y(n_124) );
INVxp67_ASAP7_75t_SL g125 ( .A(n_68), .Y(n_125) );
INVx1_ASAP7_75t_SL g126 ( .A(n_45), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_0), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_15), .Y(n_128) );
OR2x2_ASAP7_75t_L g129 ( .A(n_70), .B(n_35), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_104), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_90), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_90), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_104), .Y(n_133) );
AND2x4_ASAP7_75t_L g134 ( .A(n_117), .B(n_0), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_97), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_92), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_92), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_104), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_112), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_112), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_94), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_94), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_117), .B(n_1), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_96), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_96), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g146 ( .A(n_122), .B(n_1), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_108), .B(n_2), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_112), .B(n_2), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_116), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_98), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_116), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_116), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_98), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_99), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_99), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_113), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_100), .B(n_3), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_131), .B(n_100), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_149), .Y(n_159) );
OAI22xp5_ASAP7_75t_L g160 ( .A1(n_134), .A2(n_89), .B1(n_114), .B2(n_127), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_135), .B(n_93), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_149), .Y(n_162) );
INVx5_ASAP7_75t_L g163 ( .A(n_149), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_131), .B(n_102), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_149), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_156), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_130), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_147), .B(n_89), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_130), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_130), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_135), .B(n_102), .Y(n_171) );
BUFx3_ASAP7_75t_L g172 ( .A(n_148), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_130), .Y(n_173) );
AND2x6_ASAP7_75t_L g174 ( .A(n_134), .B(n_105), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_134), .B(n_95), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_156), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_134), .A2(n_124), .B1(n_128), .B2(n_127), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_138), .Y(n_178) );
INVx2_ASAP7_75t_SL g179 ( .A(n_134), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_147), .Y(n_180) );
INVxp33_ASAP7_75t_L g181 ( .A(n_147), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_149), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_138), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_138), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_149), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_132), .B(n_105), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_132), .B(n_109), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_138), .Y(n_188) );
INVx3_ASAP7_75t_L g189 ( .A(n_148), .Y(n_189) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_146), .Y(n_190) );
OAI22xp33_ASAP7_75t_L g191 ( .A1(n_136), .A2(n_114), .B1(n_101), .B2(n_103), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_168), .B(n_136), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_180), .A2(n_143), .B1(n_146), .B2(n_148), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_181), .B(n_143), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_172), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_179), .B(n_148), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_168), .B(n_137), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_167), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_174), .B(n_137), .Y(n_199) );
INVx2_ASAP7_75t_SL g200 ( .A(n_174), .Y(n_200) );
NOR2x1_ASAP7_75t_R g201 ( .A(n_176), .B(n_157), .Y(n_201) );
OAI22xp5_ASAP7_75t_SL g202 ( .A1(n_166), .A2(n_91), .B1(n_101), .B2(n_103), .Y(n_202) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_160), .Y(n_203) );
INVx2_ASAP7_75t_SL g204 ( .A(n_174), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_178), .Y(n_205) );
AOI22xp33_ASAP7_75t_L g206 ( .A1(n_174), .A2(n_148), .B1(n_145), .B2(n_150), .Y(n_206) );
AOI211xp5_ASAP7_75t_L g207 ( .A1(n_191), .A2(n_160), .B(n_177), .C(n_171), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_178), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g209 ( .A1(n_177), .A2(n_157), .B1(n_141), .B2(n_142), .Y(n_209) );
OAI21xp33_ASAP7_75t_L g210 ( .A1(n_172), .A2(n_142), .B(n_144), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_174), .B(n_141), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_179), .B(n_154), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_167), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_172), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_174), .B(n_144), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_174), .A2(n_145), .B1(n_150), .B2(n_154), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_174), .B(n_154), .Y(n_217) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_162), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_190), .A2(n_154), .B1(n_155), .B2(n_153), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_189), .A2(n_154), .B1(n_155), .B2(n_153), .Y(n_220) );
NAND2xp33_ASAP7_75t_SL g221 ( .A(n_189), .B(n_129), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_162), .Y(n_222) );
NAND2x1p5_ASAP7_75t_L g223 ( .A(n_189), .B(n_91), .Y(n_223) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_158), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_183), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_189), .B(n_153), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_175), .B(n_155), .Y(n_227) );
NOR2x2_ASAP7_75t_L g228 ( .A(n_161), .B(n_133), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_183), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_158), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_184), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_186), .A2(n_123), .B1(n_107), .B2(n_118), .Y(n_232) );
INVx2_ASAP7_75t_SL g233 ( .A(n_164), .Y(n_233) );
INVx8_ASAP7_75t_L g234 ( .A(n_163), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_164), .B(n_138), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_169), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_198), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_230), .B(n_169), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_234), .Y(n_239) );
BUFx2_ASAP7_75t_L g240 ( .A(n_215), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_203), .A2(n_187), .B1(n_188), .B2(n_184), .Y(n_241) );
AOI21xp5_ASAP7_75t_SL g242 ( .A1(n_215), .A2(n_129), .B(n_170), .Y(n_242) );
INVx4_ASAP7_75t_L g243 ( .A(n_234), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_230), .B(n_188), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_233), .B(n_170), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_212), .A2(n_173), .B(n_182), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_198), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_233), .A2(n_173), .B(n_139), .C(n_151), .Y(n_248) );
INVx6_ASAP7_75t_L g249 ( .A(n_195), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_213), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_213), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_224), .B(n_139), .Y(n_252) );
BUFx2_ASAP7_75t_L g253 ( .A(n_215), .Y(n_253) );
OAI22xp5_ASAP7_75t_SL g254 ( .A1(n_202), .A2(n_120), .B1(n_107), .B2(n_118), .Y(n_254) );
AO21x2_ASAP7_75t_L g255 ( .A1(n_196), .A2(n_110), .B(n_121), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_L g256 ( .A1(n_207), .A2(n_123), .B(n_120), .C(n_140), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_236), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_236), .Y(n_258) );
INVx2_ASAP7_75t_SL g259 ( .A(n_223), .Y(n_259) );
BUFx12f_ASAP7_75t_L g260 ( .A(n_223), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_192), .B(n_139), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_194), .B(n_193), .Y(n_262) );
OR2x2_ASAP7_75t_L g263 ( .A(n_197), .B(n_139), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_205), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_235), .Y(n_265) );
OR2x2_ASAP7_75t_L g266 ( .A(n_209), .B(n_139), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_208), .Y(n_267) );
BUFx4_ASAP7_75t_SL g268 ( .A(n_225), .Y(n_268) );
INVx2_ASAP7_75t_SL g269 ( .A(n_195), .Y(n_269) );
OR2x2_ASAP7_75t_L g270 ( .A(n_221), .B(n_133), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_219), .B(n_133), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_206), .B(n_140), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_229), .Y(n_273) );
INVx2_ASAP7_75t_SL g274 ( .A(n_195), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_231), .Y(n_275) );
O2A1O1Ixp33_ASAP7_75t_L g276 ( .A1(n_196), .A2(n_152), .B(n_151), .C(n_140), .Y(n_276) );
BUFx2_ASAP7_75t_L g277 ( .A(n_200), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_227), .Y(n_278) );
INVxp67_ASAP7_75t_L g279 ( .A(n_221), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_226), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_247), .Y(n_281) );
OR2x2_ASAP7_75t_L g282 ( .A(n_238), .B(n_199), .Y(n_282) );
BUFx2_ASAP7_75t_R g283 ( .A(n_268), .Y(n_283) );
OAI21x1_ASAP7_75t_L g284 ( .A1(n_242), .A2(n_182), .B(n_159), .Y(n_284) );
AO21x2_ASAP7_75t_L g285 ( .A1(n_242), .A2(n_152), .B(n_151), .Y(n_285) );
AND2x4_ASAP7_75t_L g286 ( .A(n_243), .B(n_200), .Y(n_286) );
OA21x2_ASAP7_75t_L g287 ( .A1(n_248), .A2(n_121), .B(n_111), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_246), .A2(n_212), .B(n_226), .Y(n_288) );
A2O1A1Ixp33_ASAP7_75t_L g289 ( .A1(n_256), .A2(n_210), .B(n_216), .C(n_152), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_237), .Y(n_290) );
OAI21x1_ASAP7_75t_L g291 ( .A1(n_271), .A2(n_159), .B(n_165), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_237), .Y(n_292) );
OAI21x1_ASAP7_75t_L g293 ( .A1(n_270), .A2(n_159), .B(n_165), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_250), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_250), .Y(n_295) );
OAI21x1_ASAP7_75t_SL g296 ( .A1(n_259), .A2(n_204), .B(n_217), .Y(n_296) );
OAI21x1_ASAP7_75t_L g297 ( .A1(n_270), .A2(n_165), .B(n_182), .Y(n_297) );
NAND3xp33_ASAP7_75t_L g298 ( .A(n_262), .B(n_232), .C(n_149), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_247), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_243), .B(n_204), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_279), .B(n_201), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_251), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_260), .Y(n_303) );
BUFx12f_ASAP7_75t_L g304 ( .A(n_260), .Y(n_304) );
OAI21x1_ASAP7_75t_L g305 ( .A1(n_276), .A2(n_185), .B(n_211), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_254), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_251), .Y(n_307) );
OA21x2_ASAP7_75t_L g308 ( .A1(n_264), .A2(n_110), .B(n_111), .Y(n_308) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_239), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_245), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_238), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_245), .Y(n_312) );
OAI21x1_ASAP7_75t_L g313 ( .A1(n_266), .A2(n_185), .B(n_109), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_265), .B(n_220), .Y(n_314) );
OAI21x1_ASAP7_75t_L g315 ( .A1(n_266), .A2(n_185), .B(n_214), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_243), .Y(n_316) );
AOI21xp33_ASAP7_75t_L g317 ( .A1(n_298), .A2(n_255), .B(n_244), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_281), .Y(n_318) );
AOI22xp33_ASAP7_75t_SL g319 ( .A1(n_311), .A2(n_259), .B1(n_245), .B2(n_252), .Y(n_319) );
NAND2xp33_ASAP7_75t_SL g320 ( .A(n_316), .B(n_239), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g321 ( .A1(n_288), .A2(n_264), .B(n_257), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_307), .Y(n_322) );
OAI22xp33_ASAP7_75t_L g323 ( .A1(n_304), .A2(n_263), .B1(n_267), .B2(n_275), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_314), .A2(n_252), .B1(n_241), .B2(n_273), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_288), .A2(n_258), .B(n_272), .Y(n_325) );
OAI211xp5_ASAP7_75t_L g326 ( .A1(n_301), .A2(n_261), .B(n_263), .C(n_278), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_290), .B(n_240), .Y(n_327) );
OA21x2_ASAP7_75t_L g328 ( .A1(n_284), .A2(n_280), .B(n_106), .Y(n_328) );
AND2x4_ASAP7_75t_L g329 ( .A(n_290), .B(n_239), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_307), .Y(n_330) );
A2O1A1Ixp33_ASAP7_75t_L g331 ( .A1(n_298), .A2(n_214), .B(n_274), .C(n_269), .Y(n_331) );
AOI21xp5_ASAP7_75t_SL g332 ( .A1(n_285), .A2(n_239), .B(n_274), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_281), .Y(n_333) );
INVx4_ASAP7_75t_L g334 ( .A(n_309), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_281), .A2(n_255), .B(n_269), .Y(n_335) );
OA21x2_ASAP7_75t_L g336 ( .A1(n_284), .A2(n_125), .B(n_255), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_292), .B(n_294), .Y(n_337) );
OAI22xp33_ASAP7_75t_L g338 ( .A1(n_304), .A2(n_253), .B1(n_240), .B2(n_239), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_310), .A2(n_253), .B1(n_249), .B2(n_195), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_304), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_314), .B(n_214), .Y(n_341) );
AO22x2_ASAP7_75t_L g342 ( .A1(n_310), .A2(n_228), .B1(n_126), .B2(n_249), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_314), .A2(n_249), .B1(n_277), .B2(n_228), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_310), .A2(n_249), .B1(n_277), .B2(n_115), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_292), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_345), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_345), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_322), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_318), .B(n_281), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_318), .B(n_299), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_324), .A2(n_285), .B1(n_312), .B2(n_310), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_318), .B(n_299), .Y(n_352) );
BUFx3_ASAP7_75t_L g353 ( .A(n_334), .Y(n_353) );
OAI21xp5_ASAP7_75t_L g354 ( .A1(n_325), .A2(n_289), .B(n_313), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_333), .Y(n_355) );
AND2x4_ASAP7_75t_L g356 ( .A(n_334), .B(n_315), .Y(n_356) );
INVx3_ASAP7_75t_L g357 ( .A(n_334), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_322), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_333), .B(n_299), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_337), .B(n_294), .Y(n_360) );
INVx4_ASAP7_75t_L g361 ( .A(n_334), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_330), .B(n_295), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_333), .Y(n_363) );
BUFx2_ASAP7_75t_L g364 ( .A(n_342), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_330), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_328), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_328), .Y(n_367) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_337), .Y(n_368) );
INVx4_ASAP7_75t_L g369 ( .A(n_329), .Y(n_369) );
BUFx5_ASAP7_75t_L g370 ( .A(n_329), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_341), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_327), .B(n_295), .Y(n_372) );
AOI221xp5_ASAP7_75t_L g373 ( .A1(n_323), .A2(n_306), .B1(n_301), .B2(n_289), .C(n_312), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_355), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_346), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_368), .B(n_308), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_368), .B(n_308), .Y(n_377) );
NAND2xp33_ASAP7_75t_SL g378 ( .A(n_361), .B(n_283), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_372), .B(n_343), .Y(n_379) );
OAI222xp33_ASAP7_75t_L g380 ( .A1(n_364), .A2(n_319), .B1(n_338), .B2(n_344), .C1(n_342), .C2(n_339), .Y(n_380) );
OAI21xp5_ASAP7_75t_L g381 ( .A1(n_351), .A2(n_326), .B(n_317), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_355), .B(n_308), .Y(n_382) );
AOI21xp5_ASAP7_75t_L g383 ( .A1(n_355), .A2(n_332), .B(n_317), .Y(n_383) );
AO21x2_ASAP7_75t_L g384 ( .A1(n_354), .A2(n_332), .B(n_284), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_372), .B(n_327), .Y(n_385) );
NAND5xp2_ASAP7_75t_L g386 ( .A(n_373), .B(n_283), .C(n_321), .D(n_342), .E(n_335), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_346), .B(n_303), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_347), .B(n_303), .Y(n_388) );
NOR2xp67_ASAP7_75t_L g389 ( .A(n_361), .B(n_344), .Y(n_389) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_353), .Y(n_390) );
NAND2x1_ASAP7_75t_L g391 ( .A(n_361), .B(n_328), .Y(n_391) );
OAI21xp5_ASAP7_75t_L g392 ( .A1(n_373), .A2(n_313), .B(n_308), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_349), .B(n_308), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_349), .B(n_308), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_347), .B(n_329), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_356), .B(n_285), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_348), .B(n_329), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_349), .B(n_328), .Y(n_398) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_364), .A2(n_342), .B1(n_340), .B2(n_339), .C(n_285), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_350), .B(n_285), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_355), .B(n_363), .Y(n_401) );
BUFx3_ASAP7_75t_L g402 ( .A(n_353), .Y(n_402) );
BUFx3_ASAP7_75t_L g403 ( .A(n_353), .Y(n_403) );
INVx4_ASAP7_75t_L g404 ( .A(n_361), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_348), .B(n_342), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_358), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_364), .A2(n_371), .B1(n_369), .B2(n_370), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_358), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_400), .B(n_356), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_376), .B(n_363), .Y(n_410) );
OAI33xp33_ASAP7_75t_L g411 ( .A1(n_387), .A2(n_365), .A3(n_360), .B1(n_371), .B2(n_362), .B3(n_366), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_376), .B(n_363), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_400), .B(n_398), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_398), .B(n_356), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_377), .B(n_363), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_396), .B(n_356), .Y(n_416) );
NOR3xp33_ASAP7_75t_L g417 ( .A(n_388), .B(n_320), .C(n_357), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_375), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_377), .B(n_365), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_396), .B(n_356), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_401), .B(n_366), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_401), .B(n_366), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_402), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_385), .B(n_360), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_375), .Y(n_425) );
BUFx3_ASAP7_75t_L g426 ( .A(n_402), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_405), .B(n_366), .Y(n_427) );
INVx1_ASAP7_75t_SL g428 ( .A(n_402), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_406), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_396), .B(n_367), .Y(n_430) );
INVx1_ASAP7_75t_SL g431 ( .A(n_403), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_404), .B(n_361), .Y(n_432) );
NOR3xp33_ASAP7_75t_L g433 ( .A(n_380), .B(n_357), .C(n_369), .Y(n_433) );
NAND3xp33_ASAP7_75t_L g434 ( .A(n_399), .B(n_351), .C(n_354), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_379), .B(n_4), .Y(n_435) );
INVx2_ASAP7_75t_SL g436 ( .A(n_404), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_406), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_396), .B(n_367), .Y(n_438) );
NAND4xp25_ASAP7_75t_L g439 ( .A(n_386), .B(n_369), .C(n_362), .D(n_353), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_408), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_393), .B(n_367), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_393), .B(n_362), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_408), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_394), .B(n_367), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_394), .B(n_350), .Y(n_445) );
INVxp67_ASAP7_75t_L g446 ( .A(n_403), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_374), .B(n_357), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_395), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_374), .B(n_357), .Y(n_449) );
OR2x6_ASAP7_75t_L g450 ( .A(n_404), .B(n_357), .Y(n_450) );
NAND2x1_ASAP7_75t_SL g451 ( .A(n_404), .B(n_369), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_397), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_403), .Y(n_453) );
INVx1_ASAP7_75t_SL g454 ( .A(n_390), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_390), .B(n_350), .Y(n_455) );
AND2x4_ASAP7_75t_L g456 ( .A(n_390), .B(n_369), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_382), .Y(n_457) );
OAI33xp33_ASAP7_75t_L g458 ( .A1(n_382), .A2(n_282), .A3(n_5), .B1(n_6), .B2(n_7), .B3(n_8), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_391), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_418), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_413), .B(n_384), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_425), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_441), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_413), .B(n_390), .Y(n_464) );
INVx1_ASAP7_75t_SL g465 ( .A(n_428), .Y(n_465) );
NAND2x1_ASAP7_75t_L g466 ( .A(n_450), .B(n_389), .Y(n_466) );
INVx1_ASAP7_75t_SL g467 ( .A(n_431), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_414), .B(n_384), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_414), .B(n_384), .Y(n_469) );
OAI221xp5_ASAP7_75t_L g470 ( .A1(n_435), .A2(n_378), .B1(n_381), .B2(n_407), .C(n_392), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_429), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_409), .B(n_383), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_437), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_409), .B(n_390), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_430), .B(n_391), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_445), .B(n_381), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_448), .B(n_370), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_452), .B(n_370), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_440), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_436), .B(n_389), .Y(n_480) );
NAND3xp33_ASAP7_75t_L g481 ( .A(n_434), .B(n_287), .C(n_336), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_442), .B(n_352), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_424), .B(n_370), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_410), .B(n_352), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_410), .B(n_352), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_430), .B(n_370), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_443), .B(n_370), .Y(n_487) );
BUFx3_ASAP7_75t_L g488 ( .A(n_426), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_419), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_438), .B(n_370), .Y(n_490) );
O2A1O1Ixp5_ASAP7_75t_L g491 ( .A1(n_432), .A2(n_458), .B(n_411), .C(n_459), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_441), .B(n_370), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_444), .B(n_370), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_412), .B(n_359), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_444), .B(n_370), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_419), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_421), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_412), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_433), .A2(n_370), .B1(n_287), .B2(n_336), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_457), .B(n_370), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_457), .B(n_359), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_415), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_415), .Y(n_503) );
INVx1_ASAP7_75t_SL g504 ( .A(n_426), .Y(n_504) );
NAND2xp33_ASAP7_75t_SL g505 ( .A(n_451), .B(n_359), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_450), .B(n_315), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_438), .B(n_336), .Y(n_507) );
INVx1_ASAP7_75t_SL g508 ( .A(n_451), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_432), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_423), .B(n_287), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_453), .Y(n_511) );
OAI221xp5_ASAP7_75t_L g512 ( .A1(n_417), .A2(n_282), .B1(n_287), .B2(n_331), .C(n_336), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_SL g513 ( .A1(n_446), .A2(n_299), .B(n_302), .C(n_9), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_421), .Y(n_514) );
NOR2x1_ASAP7_75t_L g515 ( .A(n_450), .B(n_287), .Y(n_515) );
OAI21x1_ASAP7_75t_L g516 ( .A1(n_439), .A2(n_291), .B(n_305), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_427), .B(n_287), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_416), .B(n_315), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_422), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_463), .B(n_427), .Y(n_520) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_511), .Y(n_521) );
INVx1_ASAP7_75t_SL g522 ( .A(n_465), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_467), .B(n_436), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_476), .B(n_422), .Y(n_524) );
OAI221xp5_ASAP7_75t_L g525 ( .A1(n_470), .A2(n_450), .B1(n_454), .B2(n_420), .C(n_416), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_476), .B(n_420), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_474), .B(n_455), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_460), .Y(n_528) );
AOI221xp5_ASAP7_75t_L g529 ( .A1(n_491), .A2(n_449), .B1(n_447), .B2(n_455), .C(n_456), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_463), .B(n_447), .Y(n_530) );
OAI32xp33_ASAP7_75t_L g531 ( .A1(n_505), .A2(n_449), .A3(n_302), .B1(n_456), .B2(n_282), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_489), .B(n_496), .Y(n_532) );
O2A1O1Ixp5_ASAP7_75t_SL g533 ( .A1(n_509), .A2(n_4), .B(n_8), .C(n_9), .Y(n_533) );
AOI211xp5_ASAP7_75t_L g534 ( .A1(n_505), .A2(n_456), .B(n_313), .C(n_309), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_498), .B(n_10), .Y(n_535) );
INVx1_ASAP7_75t_SL g536 ( .A(n_504), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_472), .A2(n_309), .B1(n_296), .B2(n_302), .Y(n_537) );
OAI221xp5_ASAP7_75t_L g538 ( .A1(n_499), .A2(n_119), .B1(n_302), .B2(n_162), .C(n_309), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_508), .B(n_309), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_472), .A2(n_309), .B1(n_296), .B2(n_305), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_484), .B(n_10), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_462), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_471), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_473), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_479), .Y(n_545) );
OAI21xp33_ASAP7_75t_L g546 ( .A1(n_461), .A2(n_468), .B(n_469), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_502), .Y(n_547) );
OAI21xp33_ASAP7_75t_L g548 ( .A1(n_461), .A2(n_162), .B(n_309), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_484), .B(n_485), .Y(n_549) );
INVxp67_ASAP7_75t_L g550 ( .A(n_488), .Y(n_550) );
OAI22xp33_ASAP7_75t_L g551 ( .A1(n_466), .A2(n_309), .B1(n_300), .B2(n_286), .Y(n_551) );
NAND2x1_ASAP7_75t_L g552 ( .A(n_506), .B(n_296), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_503), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_464), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_485), .B(n_11), .Y(n_555) );
AOI221xp5_ASAP7_75t_L g556 ( .A1(n_468), .A2(n_162), .B1(n_12), .B2(n_13), .C(n_14), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_497), .Y(n_557) );
OAI22xp33_ASAP7_75t_L g558 ( .A1(n_488), .A2(n_286), .B1(n_300), .B2(n_16), .Y(n_558) );
OAI22xp33_ASAP7_75t_L g559 ( .A1(n_515), .A2(n_286), .B1(n_300), .B2(n_17), .Y(n_559) );
AND2x2_ASAP7_75t_SL g560 ( .A(n_506), .B(n_286), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_497), .B(n_11), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_464), .Y(n_562) );
INVx1_ASAP7_75t_SL g563 ( .A(n_494), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_513), .A2(n_293), .B(n_297), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_514), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_512), .A2(n_286), .B1(n_300), .B2(n_19), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_514), .B(n_13), .Y(n_567) );
OAI32xp33_ASAP7_75t_L g568 ( .A1(n_517), .A2(n_18), .A3(n_19), .B1(n_20), .B2(n_21), .Y(n_568) );
OAI22xp33_ASAP7_75t_SL g569 ( .A1(n_480), .A2(n_21), .B1(n_22), .B2(n_23), .Y(n_569) );
OAI21xp33_ASAP7_75t_SL g570 ( .A1(n_480), .A2(n_297), .B(n_293), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_519), .Y(n_571) );
NOR3xp33_ASAP7_75t_L g572 ( .A(n_513), .B(n_305), .C(n_297), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_531), .A2(n_506), .B(n_481), .Y(n_573) );
INVx1_ASAP7_75t_SL g574 ( .A(n_536), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_524), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_560), .A2(n_482), .B1(n_483), .B2(n_492), .Y(n_576) );
NOR2x1_ASAP7_75t_L g577 ( .A(n_525), .B(n_517), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_524), .B(n_469), .Y(n_578) );
AOI221xp5_ASAP7_75t_L g579 ( .A1(n_525), .A2(n_519), .B1(n_475), .B2(n_477), .C(n_478), .Y(n_579) );
AOI211xp5_ASAP7_75t_L g580 ( .A1(n_529), .A2(n_475), .B(n_474), .C(n_507), .Y(n_580) );
NAND3xp33_ASAP7_75t_L g581 ( .A(n_521), .B(n_510), .C(n_487), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_526), .B(n_507), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_528), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_563), .B(n_482), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_542), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_549), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_543), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_522), .B(n_493), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_532), .B(n_495), .Y(n_589) );
OA21x2_ASAP7_75t_L g590 ( .A1(n_546), .A2(n_516), .B(n_500), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_547), .B(n_490), .Y(n_591) );
OAI21xp33_ASAP7_75t_SL g592 ( .A1(n_523), .A2(n_490), .B(n_486), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_544), .Y(n_593) );
AOI322xp5_ASAP7_75t_L g594 ( .A1(n_535), .A2(n_486), .A3(n_518), .B1(n_501), .B2(n_494), .C1(n_516), .C2(n_23), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_545), .Y(n_595) );
AOI211xp5_ASAP7_75t_L g596 ( .A1(n_569), .A2(n_518), .B(n_162), .C(n_24), .Y(n_596) );
XOR2x2_ASAP7_75t_L g597 ( .A(n_541), .B(n_27), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_532), .Y(n_598) );
XNOR2xp5_ASAP7_75t_L g599 ( .A(n_527), .B(n_30), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_553), .Y(n_600) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_534), .A2(n_291), .B(n_293), .Y(n_601) );
INVx1_ASAP7_75t_SL g602 ( .A(n_555), .Y(n_602) );
OAI21xp5_ASAP7_75t_L g603 ( .A1(n_559), .A2(n_291), .B(n_300), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_520), .Y(n_604) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_557), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_565), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_571), .Y(n_607) );
AOI322xp5_ASAP7_75t_L g608 ( .A1(n_535), .A2(n_163), .A3(n_32), .B1(n_34), .B2(n_37), .C1(n_39), .C2(n_41), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_575), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g610 ( .A1(n_592), .A2(n_580), .B1(n_579), .B2(n_602), .C(n_589), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_589), .A2(n_566), .B1(n_568), .B2(n_556), .C(n_567), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_605), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_577), .A2(n_566), .B1(n_550), .B2(n_558), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_574), .A2(n_554), .B1(n_562), .B2(n_561), .Y(n_614) );
OAI321xp33_ASAP7_75t_L g615 ( .A1(n_596), .A2(n_561), .A3(n_551), .B1(n_537), .B2(n_548), .C(n_538), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_598), .B(n_530), .Y(n_616) );
CKINVDCx20_ASAP7_75t_R g617 ( .A(n_599), .Y(n_617) );
OAI21xp33_ASAP7_75t_L g618 ( .A1(n_594), .A2(n_570), .B(n_552), .Y(n_618) );
CKINVDCx5p33_ASAP7_75t_R g619 ( .A(n_597), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g620 ( .A1(n_573), .A2(n_539), .B(n_564), .Y(n_620) );
NAND3xp33_ASAP7_75t_L g621 ( .A(n_590), .B(n_533), .C(n_572), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_576), .A2(n_540), .B1(n_163), .B2(n_218), .C(n_222), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_605), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_588), .A2(n_163), .B1(n_222), .B2(n_218), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_588), .B(n_31), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_582), .A2(n_586), .B1(n_584), .B2(n_578), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_573), .A2(n_163), .B1(n_234), .B2(n_44), .Y(n_627) );
OAI21xp33_ASAP7_75t_L g628 ( .A1(n_591), .A2(n_42), .B(n_43), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_583), .Y(n_629) );
AOI322xp5_ASAP7_75t_L g630 ( .A1(n_604), .A2(n_163), .A3(n_48), .B1(n_49), .B2(n_50), .C1(n_51), .C2(n_53), .Y(n_630) );
OA22x2_ASAP7_75t_L g631 ( .A1(n_613), .A2(n_595), .B1(n_593), .B2(n_587), .Y(n_631) );
AOI221x1_ASAP7_75t_L g632 ( .A1(n_618), .A2(n_585), .B1(n_600), .B2(n_606), .C(n_607), .Y(n_632) );
A2O1A1Ixp33_ASAP7_75t_SL g633 ( .A1(n_625), .A2(n_603), .B(n_601), .C(n_608), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_619), .B(n_581), .Y(n_634) );
BUFx2_ASAP7_75t_L g635 ( .A(n_612), .Y(n_635) );
OAI21xp33_ASAP7_75t_L g636 ( .A1(n_610), .A2(n_601), .B(n_590), .Y(n_636) );
AOI211x1_ASAP7_75t_L g637 ( .A1(n_620), .A2(n_47), .B(n_55), .C(n_56), .Y(n_637) );
CKINVDCx5p33_ASAP7_75t_R g638 ( .A(n_617), .Y(n_638) );
OAI211xp5_ASAP7_75t_L g639 ( .A1(n_611), .A2(n_163), .B(n_234), .C(n_59), .Y(n_639) );
OA22x2_ASAP7_75t_L g640 ( .A1(n_614), .A2(n_57), .B1(n_58), .B2(n_60), .Y(n_640) );
NAND3xp33_ASAP7_75t_L g641 ( .A(n_621), .B(n_222), .C(n_218), .Y(n_641) );
OAI221xp5_ASAP7_75t_L g642 ( .A1(n_626), .A2(n_64), .B1(n_65), .B2(n_66), .C(n_71), .Y(n_642) );
AOI211xp5_ASAP7_75t_L g643 ( .A1(n_636), .A2(n_615), .B(n_627), .C(n_622), .Y(n_643) );
OAI211xp5_ASAP7_75t_SL g644 ( .A1(n_636), .A2(n_634), .B(n_633), .C(n_639), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_631), .A2(n_623), .B1(n_616), .B2(n_609), .Y(n_645) );
NOR3x2_ASAP7_75t_L g646 ( .A(n_637), .B(n_615), .C(n_630), .Y(n_646) );
NOR3xp33_ASAP7_75t_SL g647 ( .A(n_638), .B(n_628), .C(n_629), .Y(n_647) );
OAI211xp5_ASAP7_75t_SL g648 ( .A1(n_641), .A2(n_624), .B(n_75), .C(n_78), .Y(n_648) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_635), .Y(n_649) );
OAI221xp5_ASAP7_75t_L g650 ( .A1(n_644), .A2(n_642), .B1(n_640), .B2(n_632), .C(n_82), .Y(n_650) );
AND3x4_ASAP7_75t_L g651 ( .A(n_647), .B(n_74), .C(n_79), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_649), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_645), .B(n_80), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_652), .B(n_643), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_653), .Y(n_655) );
BUFx2_ASAP7_75t_L g656 ( .A(n_651), .Y(n_656) );
NAND3xp33_ASAP7_75t_L g657 ( .A(n_654), .B(n_650), .C(n_646), .Y(n_657) );
AOI22x1_ASAP7_75t_L g658 ( .A1(n_656), .A2(n_648), .B1(n_86), .B2(n_87), .Y(n_658) );
OAI22x1_ASAP7_75t_L g659 ( .A1(n_657), .A2(n_656), .B1(n_655), .B2(n_88), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_659), .A2(n_658), .B1(n_218), .B2(n_222), .Y(n_660) );
INVxp67_ASAP7_75t_L g661 ( .A(n_660), .Y(n_661) );
AOI22xp33_ASAP7_75t_SL g662 ( .A1(n_661), .A2(n_218), .B1(n_222), .B2(n_85), .Y(n_662) );
endmodule