module fake_netlist_5_2088_n_2360 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_226, n_235, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_229, n_108, n_231, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_46, n_233, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_234, n_17, n_92, n_19, n_149, n_120, n_232, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_225, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_223, n_188, n_190, n_8, n_201, n_158, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_230, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2360);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_235;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_46;
input n_233;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_234;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_232;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2360;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_2323;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_291;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_2249;
wire n_344;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2276;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_2300;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_283;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_310;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2324;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_832;
wire n_857;
wire n_2305;
wire n_561;
wire n_1319;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_1194;
wire n_431;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_604;
wire n_433;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2320;
wire n_2339;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_2299;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_1609;
wire n_374;
wire n_1989;
wire n_2359;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_2346;
wire n_662;
wire n_459;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_1574;
wire n_473;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_2277;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_860;
wire n_441;
wire n_450;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1205;
wire n_1044;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_2198;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_2266;
wire n_389;
wire n_418;
wire n_248;
wire n_968;
wire n_912;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_2333;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_2289;
wire n_302;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_321;
wire n_2294;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_2269;
wire n_2309;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_2310;
wire n_323;
wire n_2287;
wire n_356;
wire n_2291;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2318;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_2282;
wire n_510;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2340;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_770;
wire n_458;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2148;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1543;
wire n_1399;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_2286;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_2136;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_2332;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2284;
wire n_2187;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_994;
wire n_386;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_328;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_1321;
wire n_362;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_2278;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_1654;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1956;
wire n_1936;
wire n_437;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_2273;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;
wire n_2268;

INVx1_ASAP7_75t_L g236 ( 
.A(n_46),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_146),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_159),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_69),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_116),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_226),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_169),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_160),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_76),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_183),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_230),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_179),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_24),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_128),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_109),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_86),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_84),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_218),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_201),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_177),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_108),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_148),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_18),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_127),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_187),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_93),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_43),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_7),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_141),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_57),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_82),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_39),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_118),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_197),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_66),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_214),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_176),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_135),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_143),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_6),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_85),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_149),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_36),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_20),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_32),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_203),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_74),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_34),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_3),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_24),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_126),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_4),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_29),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_50),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_138),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_171),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_157),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_97),
.Y(n_293)
);

BUFx10_ASAP7_75t_L g294 ( 
.A(n_99),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_47),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_35),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_73),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_63),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_154),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_167),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_37),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_12),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_14),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_27),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_153),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_119),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_202),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_90),
.Y(n_308)
);

INVxp33_ASAP7_75t_SL g309 ( 
.A(n_58),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_114),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_49),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_88),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_66),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_156),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_120),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_44),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_235),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_170),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_199),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_74),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_38),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_76),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_211),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_189),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_209),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_104),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_98),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_200),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_155),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_172),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_233),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_65),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_158),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_18),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_92),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_168),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_212),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_21),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_38),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_87),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_178),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_32),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_58),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_29),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_140),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_182),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_48),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_101),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_147),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_47),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_31),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_191),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_186),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_121),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_231),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_190),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_224),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_68),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_181),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_56),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_163),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_82),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_11),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_184),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_43),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_87),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_94),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_27),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_112),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_90),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_28),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_62),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_207),
.Y(n_373)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_61),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_7),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_204),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_232),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_215),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_213),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_196),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_49),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_11),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_96),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_193),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_134),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_223),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_192),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_180),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_107),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_220),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_206),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_95),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_5),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_61),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_46),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_194),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_133),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_42),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_106),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_91),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_91),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_161),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_73),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_42),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_110),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_185),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g407 ( 
.A(n_41),
.Y(n_407)
);

INVxp33_ASAP7_75t_R g408 ( 
.A(n_102),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_83),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_139),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_4),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_69),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_142),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_17),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_132),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_103),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_124),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_93),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_5),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_45),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_60),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_80),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_62),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_174),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_0),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_44),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_75),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_34),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_13),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_208),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_198),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_229),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_217),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_57),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_162),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_221),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_166),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_2),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_216),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_75),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_45),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_48),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_10),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_35),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_173),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_85),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_86),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_71),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_23),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_8),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_115),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_137),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_9),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_165),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_130),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_234),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_195),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_79),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_79),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_68),
.Y(n_460)
);

BUFx5_ASAP7_75t_L g461 ( 
.A(n_14),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_80),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_461),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_353),
.B(n_0),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_460),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_461),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_244),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_250),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_461),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_260),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_461),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_461),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_353),
.B(n_1),
.Y(n_473)
);

INVxp67_ASAP7_75t_SL g474 ( 
.A(n_318),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_271),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_251),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_412),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_461),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_461),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_261),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_461),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_262),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_265),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_238),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_238),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_246),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_246),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_412),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_239),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_239),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_318),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_292),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_395),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_303),
.Y(n_494)
);

NOR2xp67_ASAP7_75t_L g495 ( 
.A(n_429),
.B(n_1),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_345),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_402),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_276),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_416),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_273),
.B(n_2),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_445),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_239),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_309),
.B(n_247),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_239),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_278),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_279),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_284),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_247),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_329),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_285),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_255),
.Y(n_511)
);

INVxp67_ASAP7_75t_SL g512 ( 
.A(n_329),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_336),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_289),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_240),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_254),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g517 ( 
.A(n_290),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_295),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_308),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_324),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_255),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_257),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_257),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_311),
.Y(n_524)
);

NOR2xp67_ASAP7_75t_L g525 ( 
.A(n_296),
.B(n_3),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_312),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_269),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_263),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_397),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_269),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_274),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_263),
.Y(n_532)
);

BUFx6f_ASAP7_75t_SL g533 ( 
.A(n_256),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_316),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_259),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_320),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_274),
.B(n_6),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_277),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_277),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_239),
.Y(n_540)
);

INVxp67_ASAP7_75t_SL g541 ( 
.A(n_439),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_281),
.B(n_8),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_281),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_321),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_310),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_310),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_322),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_338),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_339),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_342),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_350),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_360),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_319),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_319),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_325),
.Y(n_555)
);

INVxp33_ASAP7_75t_SL g556 ( 
.A(n_363),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_325),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_314),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_366),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_297),
.Y(n_560)
);

BUFx2_ASAP7_75t_L g561 ( 
.A(n_303),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_336),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_297),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_372),
.Y(n_564)
);

INVxp67_ASAP7_75t_SL g565 ( 
.A(n_439),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_297),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_297),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_382),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_393),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_297),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_400),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_263),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_341),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_237),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_241),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_341),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_243),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_348),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_245),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_348),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_249),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_361),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_401),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_358),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_358),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_358),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_404),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_253),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_474),
.B(n_334),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_566),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_489),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_513),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_512),
.B(n_273),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_489),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_490),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_490),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_502),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_502),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_513),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_504),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_504),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_488),
.A2(n_368),
.B1(n_381),
.B2(n_258),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_566),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_540),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_513),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_465),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_540),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_574),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_513),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_465),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_560),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_513),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_541),
.B(n_305),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_562),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_565),
.B(n_305),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_560),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_467),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_563),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_491),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_562),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_562),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_562),
.Y(n_622)
);

NAND2xp33_ASAP7_75t_SL g623 ( 
.A(n_464),
.B(n_296),
.Y(n_623)
);

BUFx8_ASAP7_75t_L g624 ( 
.A(n_533),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_562),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_563),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_503),
.B(n_417),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_567),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_567),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_570),
.Y(n_630)
);

BUFx2_ASAP7_75t_L g631 ( 
.A(n_467),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_466),
.Y(n_632)
);

BUFx2_ASAP7_75t_L g633 ( 
.A(n_476),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_570),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_584),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_584),
.B(n_417),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_472),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_491),
.B(n_436),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_505),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_478),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_575),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_476),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_585),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_509),
.B(n_436),
.Y(n_644)
);

HB1xp67_ASAP7_75t_L g645 ( 
.A(n_480),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_556),
.B(n_242),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_479),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_481),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_463),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_463),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_469),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_585),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_586),
.Y(n_653)
);

NAND2xp33_ASAP7_75t_L g654 ( 
.A(n_480),
.B(n_358),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_586),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_469),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_471),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_471),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_484),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_509),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_485),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_473),
.B(n_286),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_486),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_487),
.Y(n_664)
);

BUFx2_ASAP7_75t_L g665 ( 
.A(n_482),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_508),
.B(n_437),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_511),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_517),
.B(n_256),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_510),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_521),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_522),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_523),
.B(n_437),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_527),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_529),
.B(n_535),
.Y(n_674)
);

AND2x6_ASAP7_75t_L g675 ( 
.A(n_537),
.B(n_336),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_558),
.B(n_256),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_530),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_531),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_542),
.A2(n_449),
.B1(n_448),
.B2(n_495),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_538),
.Y(n_680)
);

AND2x6_ASAP7_75t_L g681 ( 
.A(n_500),
.B(n_336),
.Y(n_681)
);

AND2x6_ASAP7_75t_L g682 ( 
.A(n_539),
.B(n_336),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_543),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_577),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_545),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_546),
.Y(n_686)
);

INVx1_ASAP7_75t_SL g687 ( 
.A(n_631),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_627),
.A2(n_477),
.B1(n_370),
.B2(n_358),
.Y(n_688)
);

AND3x2_ASAP7_75t_L g689 ( 
.A(n_662),
.B(n_302),
.C(n_283),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_660),
.B(n_553),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_590),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_L g692 ( 
.A(n_675),
.B(n_482),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_619),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_590),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_590),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_589),
.B(n_660),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_675),
.A2(n_370),
.B1(n_407),
.B2(n_374),
.Y(n_697)
);

AND3x1_ASAP7_75t_L g698 ( 
.A(n_679),
.B(n_407),
.C(n_374),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_603),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_656),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_658),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_656),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_646),
.B(n_579),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_603),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_603),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_608),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_619),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_675),
.A2(n_370),
.B1(n_555),
.B2(n_554),
.Y(n_708)
);

INVx4_ASAP7_75t_L g709 ( 
.A(n_658),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_657),
.B(n_675),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_657),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_619),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_658),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_675),
.B(n_557),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_679),
.A2(n_248),
.B1(n_398),
.B2(n_394),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_639),
.B(n_581),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_669),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_666),
.B(n_361),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_675),
.A2(n_370),
.B1(n_576),
.B2(n_573),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_666),
.B(n_369),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_649),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_649),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_675),
.B(n_578),
.Y(n_723)
);

AND2x4_ASAP7_75t_L g724 ( 
.A(n_666),
.B(n_369),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_658),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_649),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_624),
.B(n_483),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_632),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_624),
.B(n_483),
.Y(n_729)
);

AO21x2_ASAP7_75t_L g730 ( 
.A1(n_593),
.A2(n_415),
.B(n_413),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_650),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_632),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_624),
.B(n_498),
.Y(n_733)
);

INVx4_ASAP7_75t_L g734 ( 
.A(n_658),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_632),
.Y(n_735)
);

CKINVDCx20_ASAP7_75t_R g736 ( 
.A(n_641),
.Y(n_736)
);

INVx4_ASAP7_75t_L g737 ( 
.A(n_658),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_589),
.B(n_588),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_613),
.B(n_498),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_650),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_650),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_650),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_651),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_647),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_675),
.A2(n_681),
.B1(n_615),
.B2(n_672),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_647),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_651),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_651),
.Y(n_748)
);

OR2x6_ASAP7_75t_L g749 ( 
.A(n_638),
.B(n_644),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_647),
.Y(n_750)
);

NOR2x1p5_ASAP7_75t_L g751 ( 
.A(n_684),
.B(n_334),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_648),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_651),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_654),
.B(n_506),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_661),
.B(n_580),
.Y(n_755)
);

INVx4_ASAP7_75t_L g756 ( 
.A(n_637),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_592),
.Y(n_757)
);

INVx4_ASAP7_75t_L g758 ( 
.A(n_637),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_661),
.B(n_582),
.Y(n_759)
);

NAND2xp33_ASAP7_75t_SL g760 ( 
.A(n_668),
.B(n_515),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_617),
.B(n_506),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_606),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_592),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_610),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_624),
.B(n_507),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_666),
.B(n_373),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_642),
.B(n_507),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_592),
.Y(n_768)
);

NAND3xp33_ASAP7_75t_L g769 ( 
.A(n_670),
.B(n_525),
.C(n_385),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_648),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_648),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_667),
.Y(n_772)
);

AND2x6_ASAP7_75t_L g773 ( 
.A(n_636),
.B(n_356),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_591),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_667),
.B(n_514),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_645),
.B(n_514),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_591),
.Y(n_777)
);

INVxp67_ASAP7_75t_L g778 ( 
.A(n_631),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_594),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_633),
.B(n_518),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_594),
.Y(n_781)
);

BUFx4f_ASAP7_75t_L g782 ( 
.A(n_637),
.Y(n_782)
);

NAND3xp33_ASAP7_75t_L g783 ( 
.A(n_670),
.B(n_385),
.C(n_373),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_681),
.A2(n_370),
.B1(n_302),
.B2(n_283),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_633),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_637),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_667),
.B(n_673),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_667),
.B(n_518),
.Y(n_788)
);

CKINVDCx6p67_ASAP7_75t_R g789 ( 
.A(n_674),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_673),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_673),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_673),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_L g793 ( 
.A(n_681),
.B(n_519),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_677),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_677),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_680),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_672),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_680),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_685),
.B(n_494),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_592),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_665),
.B(n_519),
.Y(n_801)
);

OAI21xp33_ASAP7_75t_SL g802 ( 
.A1(n_676),
.A2(n_252),
.B(n_236),
.Y(n_802)
);

INVx5_ASAP7_75t_L g803 ( 
.A(n_682),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_685),
.B(n_494),
.Y(n_804)
);

OR2x6_ASAP7_75t_L g805 ( 
.A(n_665),
.B(n_388),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_637),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_595),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_595),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_623),
.B(n_524),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_637),
.B(n_524),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_640),
.B(n_681),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_596),
.Y(n_812)
);

INVx6_ASAP7_75t_L g813 ( 
.A(n_640),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_596),
.Y(n_814)
);

OR2x2_ASAP7_75t_L g815 ( 
.A(n_602),
.B(n_547),
.Y(n_815)
);

BUFx2_ASAP7_75t_L g816 ( 
.A(n_602),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_672),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_681),
.A2(n_375),
.B1(n_493),
.B2(n_252),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_672),
.B(n_388),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_597),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_592),
.Y(n_821)
);

XOR2xp5_ASAP7_75t_L g822 ( 
.A(n_664),
.B(n_468),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_664),
.B(n_526),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_664),
.B(n_561),
.Y(n_824)
);

OR2x6_ASAP7_75t_L g825 ( 
.A(n_636),
.B(n_389),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_597),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_598),
.Y(n_827)
);

AND2x6_ASAP7_75t_L g828 ( 
.A(n_636),
.B(n_356),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_681),
.A2(n_375),
.B1(n_266),
.B2(n_267),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_598),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_592),
.Y(n_831)
);

AND2x2_ASAP7_75t_SL g832 ( 
.A(n_636),
.B(n_356),
.Y(n_832)
);

INVxp67_ASAP7_75t_SL g833 ( 
.A(n_599),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_600),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_612),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_659),
.B(n_526),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_612),
.Y(n_837)
);

BUFx2_ASAP7_75t_L g838 ( 
.A(n_659),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_659),
.B(n_534),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_600),
.Y(n_840)
);

INVx6_ASAP7_75t_L g841 ( 
.A(n_640),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_612),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_671),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_671),
.Y(n_844)
);

AND2x6_ASAP7_75t_L g845 ( 
.A(n_640),
.B(n_356),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_671),
.B(n_561),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_601),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_640),
.B(n_534),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_681),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_681),
.A2(n_266),
.B1(n_267),
.B2(n_236),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_696),
.B(n_640),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_843),
.Y(n_852)
);

OAI22xp33_ASAP7_75t_L g853 ( 
.A1(n_715),
.A2(n_275),
.B1(n_280),
.B2(n_270),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_794),
.Y(n_854)
);

OR2x2_ASAP7_75t_L g855 ( 
.A(n_687),
.B(n_785),
.Y(n_855)
);

INVx5_ASAP7_75t_L g856 ( 
.A(n_845),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_696),
.B(n_659),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_794),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_824),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_739),
.B(n_659),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_797),
.B(n_659),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_730),
.A2(n_275),
.B1(n_280),
.B2(n_270),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_730),
.A2(n_287),
.B1(n_288),
.B2(n_282),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_745),
.A2(n_520),
.B1(n_516),
.B2(n_475),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_754),
.B(n_536),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_795),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_795),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_832),
.B(n_356),
.Y(n_868)
);

AND2x2_ASAP7_75t_SL g869 ( 
.A(n_698),
.B(n_389),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_691),
.Y(n_870)
);

INVxp67_ASAP7_75t_L g871 ( 
.A(n_801),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_797),
.B(n_663),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_844),
.B(n_536),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_817),
.B(n_663),
.Y(n_874)
);

INVx4_ASAP7_75t_L g875 ( 
.A(n_707),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_823),
.B(n_544),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_691),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_817),
.B(n_663),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_775),
.A2(n_492),
.B1(n_496),
.B2(n_470),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_832),
.B(n_380),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_694),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_730),
.A2(n_287),
.B1(n_288),
.B2(n_282),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_788),
.B(n_544),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_796),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_796),
.Y(n_885)
);

NAND2xp33_ASAP7_75t_L g886 ( 
.A(n_810),
.B(n_264),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_SL g887 ( 
.A1(n_816),
.A2(n_499),
.B1(n_501),
.B2(n_497),
.Y(n_887)
);

NAND2xp33_ASAP7_75t_R g888 ( 
.A(n_816),
.B(n_548),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_700),
.B(n_663),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_707),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_848),
.B(n_548),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_700),
.B(n_663),
.Y(n_892)
);

OAI221xp5_ASAP7_75t_L g893 ( 
.A1(n_688),
.A2(n_421),
.B1(n_298),
.B2(n_403),
.C(n_304),
.Y(n_893)
);

BUFx6f_ASAP7_75t_SL g894 ( 
.A(n_762),
.Y(n_894)
);

BUFx5_ASAP7_75t_L g895 ( 
.A(n_731),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_695),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_702),
.B(n_711),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_798),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_702),
.B(n_663),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_707),
.B(n_396),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_798),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_755),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_711),
.B(n_678),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_755),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_832),
.B(n_678),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_759),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_710),
.B(n_380),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_712),
.B(n_678),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_712),
.B(n_807),
.Y(n_909)
);

NOR3xp33_ASAP7_75t_L g910 ( 
.A(n_703),
.B(n_551),
.C(n_550),
.Y(n_910)
);

NAND3xp33_ASAP7_75t_L g911 ( 
.A(n_738),
.B(n_551),
.C(n_550),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_807),
.B(n_678),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_757),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_812),
.B(n_678),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_759),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_699),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_772),
.B(n_380),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_812),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_772),
.B(n_380),
.Y(n_919)
);

O2A1O1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_692),
.A2(n_301),
.B(n_304),
.C(n_298),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_749),
.A2(n_559),
.B1(n_569),
.B2(n_552),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_799),
.B(n_549),
.Y(n_922)
);

NOR2xp67_ASAP7_75t_SL g923 ( 
.A(n_803),
.B(n_849),
.Y(n_923)
);

OR2x6_ASAP7_75t_L g924 ( 
.A(n_762),
.B(n_528),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_699),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_693),
.B(n_552),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_790),
.B(n_380),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_820),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_693),
.B(n_559),
.Y(n_929)
);

INVx8_ASAP7_75t_L g930 ( 
.A(n_805),
.Y(n_930)
);

NOR2xp67_ASAP7_75t_L g931 ( 
.A(n_778),
.B(n_569),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_820),
.B(n_678),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_802),
.B(n_571),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_802),
.B(n_571),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_799),
.B(n_564),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_R g936 ( 
.A(n_706),
.B(n_583),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_704),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_826),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_704),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_826),
.B(n_683),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_790),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_731),
.B(n_683),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_791),
.B(n_683),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_705),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_804),
.B(n_583),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_740),
.B(n_683),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_791),
.B(n_683),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_740),
.B(n_741),
.Y(n_948)
);

AND2x2_ASAP7_75t_SL g949 ( 
.A(n_698),
.B(n_396),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_804),
.B(n_587),
.Y(n_950)
);

INVxp67_ASAP7_75t_L g951 ( 
.A(n_717),
.Y(n_951)
);

OAI22xp33_ASAP7_75t_L g952 ( 
.A1(n_715),
.A2(n_313),
.B1(n_332),
.B2(n_301),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_705),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_749),
.A2(n_587),
.B1(n_272),
.B2(n_291),
.Y(n_954)
);

INVx2_ASAP7_75t_SL g955 ( 
.A(n_824),
.Y(n_955)
);

AND2x4_ASAP7_75t_SL g956 ( 
.A(n_736),
.B(n_568),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_792),
.B(n_683),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_R g958 ( 
.A(n_760),
.B(n_268),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_749),
.A2(n_299),
.B1(n_300),
.B2(n_293),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_741),
.B(n_686),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_742),
.B(n_686),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_742),
.B(n_686),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_815),
.B(n_532),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_743),
.B(n_686),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_743),
.B(n_686),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_846),
.B(n_399),
.Y(n_966)
);

INVx8_ASAP7_75t_L g967 ( 
.A(n_805),
.Y(n_967)
);

OR2x2_ASAP7_75t_L g968 ( 
.A(n_815),
.B(n_572),
.Y(n_968)
);

AOI22xp33_ASAP7_75t_L g969 ( 
.A1(n_697),
.A2(n_850),
.B1(n_829),
.B2(n_784),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_792),
.Y(n_970)
);

INVxp67_ASAP7_75t_L g971 ( 
.A(n_716),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_774),
.Y(n_972)
);

INVxp67_ASAP7_75t_L g973 ( 
.A(n_761),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_744),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_747),
.B(n_686),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_846),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_714),
.B(n_306),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_836),
.B(n_408),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_774),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_744),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_723),
.B(n_307),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_787),
.B(n_315),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_718),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_764),
.B(n_409),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_839),
.B(n_533),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_777),
.Y(n_986)
);

AOI22xp33_ASAP7_75t_L g987 ( 
.A1(n_718),
.A2(n_351),
.B1(n_313),
.B2(n_332),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_747),
.B(n_748),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_749),
.A2(n_352),
.B1(n_317),
.B2(n_323),
.Y(n_989)
);

OR2x6_ASAP7_75t_L g990 ( 
.A(n_764),
.B(n_335),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_L g991 ( 
.A1(n_749),
.A2(n_354),
.B1(n_326),
.B2(n_327),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_811),
.B(n_328),
.Y(n_992)
);

NAND3xp33_ASAP7_75t_L g993 ( 
.A(n_767),
.B(n_418),
.C(n_414),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_748),
.B(n_330),
.Y(n_994)
);

AOI22xp33_ASAP7_75t_L g995 ( 
.A1(n_718),
.A2(n_724),
.B1(n_766),
.B2(n_720),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_753),
.B(n_833),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_690),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_757),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_744),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_753),
.B(n_331),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_838),
.B(n_601),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_779),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_776),
.B(n_333),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_718),
.B(n_337),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_779),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_781),
.Y(n_1006)
);

OR2x6_ASAP7_75t_L g1007 ( 
.A(n_805),
.B(n_335),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_805),
.B(n_419),
.Y(n_1008)
);

NAND2xp33_ASAP7_75t_L g1009 ( 
.A(n_849),
.B(n_708),
.Y(n_1009)
);

INVx2_ASAP7_75t_SL g1010 ( 
.A(n_751),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_781),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_809),
.B(n_533),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_806),
.B(n_346),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_806),
.B(n_349),
.Y(n_1014)
);

AND2x2_ASAP7_75t_SL g1015 ( 
.A(n_818),
.B(n_399),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_805),
.B(n_420),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_806),
.B(n_355),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_719),
.B(n_357),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_780),
.B(n_422),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_808),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_808),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_720),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_922),
.B(n_751),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_976),
.B(n_720),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_891),
.B(n_720),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_891),
.A2(n_793),
.B1(n_838),
.B2(n_766),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_995),
.B(n_701),
.Y(n_1027)
);

INVxp67_ASAP7_75t_L g1028 ( 
.A(n_855),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_941),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_854),
.B(n_724),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_860),
.A2(n_782),
.B(n_734),
.Y(n_1031)
);

OAI21xp33_ASAP7_75t_L g1032 ( 
.A1(n_945),
.A2(n_729),
.B(n_727),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_858),
.B(n_724),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_866),
.B(n_867),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_970),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_976),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_972),
.Y(n_1037)
);

NOR2xp67_ASAP7_75t_L g1038 ( 
.A(n_971),
.B(n_769),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_851),
.A2(n_782),
.B(n_734),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_857),
.A2(n_782),
.B(n_734),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_905),
.A2(n_734),
.B(n_709),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_861),
.A2(n_737),
.B(n_709),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_872),
.A2(n_737),
.B(n_709),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_884),
.B(n_724),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_885),
.B(n_766),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_898),
.B(n_766),
.Y(n_1046)
);

O2A1O1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_853),
.A2(n_847),
.B(n_814),
.C(n_830),
.Y(n_1047)
);

INVx1_ASAP7_75t_SL g1048 ( 
.A(n_956),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_901),
.B(n_819),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_871),
.B(n_789),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_973),
.B(n_789),
.Y(n_1051)
);

INVxp67_ASAP7_75t_L g1052 ( 
.A(n_935),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_995),
.B(n_701),
.Y(n_1053)
);

NOR2x2_ASAP7_75t_L g1054 ( 
.A(n_1007),
.B(n_825),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_979),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_874),
.A2(n_737),
.B(n_709),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_945),
.B(n_822),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_895),
.B(n_701),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_883),
.B(n_918),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_883),
.B(n_819),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_878),
.A2(n_737),
.B(n_756),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_936),
.Y(n_1062)
);

NOR2x1_ASAP7_75t_L g1063 ( 
.A(n_911),
.B(n_931),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_986),
.Y(n_1064)
);

BUFx4f_ASAP7_75t_L g1065 ( 
.A(n_930),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_1002),
.Y(n_1066)
);

AO21x1_ASAP7_75t_L g1067 ( 
.A1(n_868),
.A2(n_435),
.B(n_405),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_950),
.B(n_822),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_1005),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_969),
.A2(n_825),
.B1(n_769),
.B2(n_819),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_890),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_928),
.B(n_819),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_950),
.B(n_733),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_1006),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_963),
.B(n_765),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_938),
.B(n_814),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1009),
.A2(n_758),
.B(n_756),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_997),
.B(n_827),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_908),
.A2(n_758),
.B(n_756),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_948),
.A2(n_722),
.B(n_721),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_895),
.B(n_701),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_890),
.A2(n_758),
.B(n_756),
.Y(n_1082)
);

OAI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_988),
.A2(n_722),
.B(n_721),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_897),
.B(n_827),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_992),
.A2(n_758),
.B(n_786),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_968),
.B(n_830),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_L g1087 ( 
.A(n_859),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_955),
.B(n_909),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_902),
.B(n_834),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_992),
.A2(n_786),
.B(n_763),
.Y(n_1090)
);

OR2x6_ASAP7_75t_L g1091 ( 
.A(n_930),
.B(n_825),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1011),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_996),
.A2(n_786),
.B(n_763),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_913),
.A2(n_763),
.B(n_757),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1020),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_1021),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_984),
.B(n_689),
.Y(n_1097)
);

INVx4_ASAP7_75t_L g1098 ( 
.A(n_983),
.Y(n_1098)
);

CKINVDCx20_ASAP7_75t_R g1099 ( 
.A(n_936),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_904),
.B(n_834),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_913),
.A2(n_998),
.B(n_1001),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_913),
.A2(n_763),
.B(n_757),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_895),
.B(n_713),
.Y(n_1103)
);

CKINVDCx8_ASAP7_75t_R g1104 ( 
.A(n_924),
.Y(n_1104)
);

INVx5_ASAP7_75t_L g1105 ( 
.A(n_913),
.Y(n_1105)
);

OR2x6_ASAP7_75t_L g1106 ( 
.A(n_930),
.B(n_825),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_983),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_906),
.B(n_840),
.Y(n_1108)
);

O2A1O1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_853),
.A2(n_847),
.B(n_840),
.C(n_825),
.Y(n_1109)
);

O2A1O1Ixp5_ASAP7_75t_L g1110 ( 
.A1(n_868),
.A2(n_725),
.B(n_713),
.C(n_728),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_966),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_998),
.A2(n_763),
.B(n_757),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_915),
.B(n_713),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_895),
.B(n_713),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_880),
.A2(n_726),
.B(n_770),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_998),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_952),
.A2(n_783),
.B(n_770),
.C(n_771),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_969),
.B(n_966),
.Y(n_1118)
);

OAI21xp33_ASAP7_75t_L g1119 ( 
.A1(n_1019),
.A2(n_426),
.B(n_423),
.Y(n_1119)
);

HB1xp67_ASAP7_75t_L g1120 ( 
.A(n_1022),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_870),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_900),
.B(n_725),
.Y(n_1122)
);

INVx2_ASAP7_75t_SL g1123 ( 
.A(n_990),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_998),
.A2(n_981),
.B(n_977),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_1022),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_977),
.A2(n_725),
.B(n_803),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_900),
.B(n_725),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1015),
.B(n_726),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_1019),
.A2(n_783),
.B(n_403),
.C(n_371),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_877),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_978),
.A2(n_841),
.B1(n_813),
.B2(n_771),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_881),
.Y(n_1132)
);

NOR2xp67_ASAP7_75t_L g1133 ( 
.A(n_951),
.B(n_728),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_981),
.A2(n_803),
.B(n_800),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_926),
.B(n_732),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_852),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_880),
.A2(n_750),
.B(n_746),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_1010),
.B(n_405),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_889),
.A2(n_803),
.B(n_800),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1015),
.B(n_732),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_896),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_895),
.B(n_803),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_892),
.A2(n_803),
.B(n_800),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_926),
.B(n_735),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_916),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_899),
.A2(n_800),
.B(n_768),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_862),
.B(n_863),
.Y(n_1147)
);

INVxp67_ASAP7_75t_L g1148 ( 
.A(n_924),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_925),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_907),
.A2(n_750),
.B(n_746),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_907),
.A2(n_750),
.B(n_746),
.Y(n_1151)
);

CKINVDCx10_ASAP7_75t_R g1152 ( 
.A(n_894),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_895),
.B(n_752),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_862),
.B(n_735),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_863),
.A2(n_451),
.B1(n_455),
.B2(n_452),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_882),
.B(n_752),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_856),
.B(n_752),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_876),
.B(n_813),
.Y(n_1158)
);

A2O1A1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_882),
.A2(n_365),
.B(n_371),
.C(n_362),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_856),
.B(n_768),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_942),
.A2(n_821),
.B(n_768),
.Y(n_1161)
);

BUFx4f_ASAP7_75t_L g1162 ( 
.A(n_967),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_903),
.A2(n_914),
.B(n_912),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_875),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_875),
.B(n_768),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_865),
.B(n_821),
.Y(n_1166)
);

NAND2xp33_ASAP7_75t_L g1167 ( 
.A(n_967),
.B(n_856),
.Y(n_1167)
);

OAI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_888),
.A2(n_451),
.B1(n_452),
.B2(n_455),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_937),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_932),
.A2(n_831),
.B(n_821),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_978),
.B(n_813),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_856),
.B(n_821),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_987),
.A2(n_442),
.B(n_344),
.C(n_343),
.Y(n_1173)
);

AOI33xp33_ASAP7_75t_L g1174 ( 
.A1(n_952),
.A2(n_411),
.A3(n_421),
.B1(n_425),
.B2(n_427),
.B3(n_453),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_893),
.A2(n_435),
.B(n_457),
.C(n_604),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_994),
.B(n_831),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_994),
.B(n_831),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_939),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_864),
.B(n_831),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1000),
.B(n_835),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_924),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_967),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_944),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_940),
.B(n_835),
.Y(n_1184)
);

NOR2x1p5_ASAP7_75t_L g1185 ( 
.A(n_993),
.B(n_428),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_959),
.B(n_835),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_946),
.A2(n_837),
.B(n_835),
.Y(n_1187)
);

AOI21x1_ASAP7_75t_L g1188 ( 
.A1(n_943),
.A2(n_609),
.B(n_605),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_953),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_960),
.A2(n_842),
.B(n_837),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_974),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_873),
.B(n_434),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1000),
.B(n_837),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_985),
.B(n_837),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_1007),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_980),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_929),
.B(n_813),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_999),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_989),
.A2(n_457),
.B1(n_841),
.B2(n_842),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_985),
.B(n_982),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_961),
.A2(n_842),
.B(n_621),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_962),
.A2(n_842),
.B(n_621),
.Y(n_1202)
);

OAI21xp33_ASAP7_75t_L g1203 ( 
.A1(n_921),
.A2(n_441),
.B(n_440),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_964),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_965),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_879),
.B(n_841),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_888),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_990),
.B(n_841),
.Y(n_1208)
);

BUFx4f_ASAP7_75t_L g1209 ( 
.A(n_990),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_982),
.B(n_604),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_975),
.A2(n_621),
.B(n_612),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_894),
.Y(n_1212)
);

AO21x1_ASAP7_75t_L g1213 ( 
.A1(n_920),
.A2(n_343),
.B(n_340),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_R g1214 ( 
.A(n_1099),
.B(n_1012),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1095),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1059),
.B(n_887),
.Y(n_1216)
);

O2A1O1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1168),
.A2(n_934),
.B(n_933),
.C(n_1003),
.Y(n_1217)
);

O2A1O1Ixp5_ASAP7_75t_L g1218 ( 
.A1(n_1200),
.A2(n_1017),
.B(n_1014),
.C(n_1013),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_1036),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_R g1220 ( 
.A(n_1207),
.B(n_1012),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1105),
.A2(n_886),
.B(n_1004),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1095),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_1073),
.B(n_954),
.Y(n_1223)
);

INVx1_ASAP7_75t_SL g1224 ( 
.A(n_1048),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1147),
.A2(n_991),
.B1(n_987),
.B2(n_869),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1076),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1135),
.B(n_1008),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1105),
.A2(n_1014),
.B(n_1013),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1135),
.B(n_1086),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1086),
.B(n_1016),
.Y(n_1230)
);

AND2x4_ASAP7_75t_L g1231 ( 
.A(n_1036),
.B(n_910),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1168),
.A2(n_1017),
.B(n_919),
.C(n_917),
.Y(n_1232)
);

INVxp67_ASAP7_75t_SL g1233 ( 
.A(n_1116),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1024),
.B(n_869),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_1120),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1055),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_SL g1237 ( 
.A(n_1024),
.B(n_949),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1144),
.B(n_949),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_SL g1239 ( 
.A(n_1075),
.B(n_958),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1052),
.B(n_1028),
.Y(n_1240)
);

O2A1O1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1075),
.A2(n_927),
.B(n_919),
.C(n_917),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_1116),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1116),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1118),
.A2(n_1018),
.B1(n_957),
.B2(n_947),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_1111),
.B(n_1182),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_R g1246 ( 
.A(n_1212),
.B(n_359),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1105),
.A2(n_947),
.B(n_943),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1188),
.A2(n_957),
.B(n_927),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1060),
.A2(n_1018),
.B1(n_364),
.B2(n_391),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1025),
.A2(n_383),
.B1(n_387),
.B2(n_390),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1109),
.A2(n_923),
.B(n_453),
.C(n_340),
.Y(n_1251)
);

AO21x2_ASAP7_75t_L g1252 ( 
.A1(n_1194),
.A2(n_958),
.B(n_611),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1105),
.A2(n_621),
.B(n_612),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1198),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1057),
.B(n_443),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1125),
.B(n_367),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1077),
.A2(n_621),
.B(n_612),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1031),
.A2(n_621),
.B(n_599),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1057),
.B(n_446),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1026),
.A2(n_454),
.B1(n_376),
.B2(n_377),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1079),
.A2(n_609),
.B(n_605),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1088),
.B(n_607),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1125),
.B(n_378),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1068),
.B(n_447),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1120),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1041),
.A2(n_599),
.B(n_605),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1198),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1191),
.Y(n_1268)
);

BUFx2_ASAP7_75t_L g1269 ( 
.A(n_1148),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_1116),
.Y(n_1270)
);

NOR3xp33_ASAP7_75t_SL g1271 ( 
.A(n_1068),
.B(n_450),
.C(n_458),
.Y(n_1271)
);

INVx1_ASAP7_75t_SL g1272 ( 
.A(n_1181),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1078),
.B(n_607),
.Y(n_1273)
);

BUFx12f_ASAP7_75t_L g1274 ( 
.A(n_1138),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1082),
.A2(n_599),
.B(n_620),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1034),
.B(n_611),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1050),
.B(n_459),
.Y(n_1277)
);

OAI22x1_ASAP7_75t_L g1278 ( 
.A1(n_1050),
.A2(n_462),
.B1(n_425),
.B2(n_347),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1051),
.B(n_379),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1039),
.A2(n_622),
.B(n_609),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1195),
.Y(n_1281)
);

OAI21xp33_ASAP7_75t_SL g1282 ( 
.A1(n_1027),
.A2(n_347),
.B(n_344),
.Y(n_1282)
);

NOR3xp33_ASAP7_75t_SL g1283 ( 
.A(n_1203),
.B(n_406),
.C(n_392),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1087),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1092),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_1152),
.Y(n_1286)
);

O2A1O1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1129),
.A2(n_427),
.B(n_411),
.C(n_365),
.Y(n_1287)
);

A2O1A1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1032),
.A2(n_444),
.B(n_442),
.C(n_438),
.Y(n_1288)
);

NAND2xp33_ASAP7_75t_SL g1289 ( 
.A(n_1182),
.B(n_384),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1051),
.B(n_386),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1040),
.A2(n_622),
.B(n_614),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1128),
.A2(n_828),
.B(n_773),
.Y(n_1292)
);

AND2x2_ASAP7_75t_SL g1293 ( 
.A(n_1167),
.B(n_351),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1163),
.A2(n_622),
.B(n_614),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1087),
.B(n_410),
.Y(n_1295)
);

AOI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1206),
.A2(n_430),
.B1(n_433),
.B2(n_432),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1029),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1062),
.B(n_424),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1035),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1037),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1125),
.Y(n_1301)
);

INVx1_ASAP7_75t_SL g1302 ( 
.A(n_1136),
.Y(n_1302)
);

INVxp67_ASAP7_75t_L g1303 ( 
.A(n_1023),
.Y(n_1303)
);

O2A1O1Ixp33_ASAP7_75t_L g1304 ( 
.A1(n_1129),
.A2(n_444),
.B(n_362),
.C(n_438),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1084),
.B(n_616),
.Y(n_1305)
);

NAND2x1p5_ASAP7_75t_L g1306 ( 
.A(n_1164),
.B(n_616),
.Y(n_1306)
);

INVxp67_ASAP7_75t_SL g1307 ( 
.A(n_1164),
.Y(n_1307)
);

O2A1O1Ixp5_ASAP7_75t_L g1308 ( 
.A1(n_1186),
.A2(n_629),
.B(n_626),
.C(n_618),
.Y(n_1308)
);

O2A1O1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1155),
.A2(n_629),
.B(n_653),
.C(n_618),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1089),
.Y(n_1310)
);

INVx1_ASAP7_75t_SL g1311 ( 
.A(n_1192),
.Y(n_1311)
);

OAI21xp33_ASAP7_75t_L g1312 ( 
.A1(n_1119),
.A2(n_431),
.B(n_456),
.Y(n_1312)
);

INVxp67_ASAP7_75t_L g1313 ( 
.A(n_1206),
.Y(n_1313)
);

OR2x6_ASAP7_75t_L g1314 ( 
.A(n_1091),
.B(n_626),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1123),
.B(n_9),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1027),
.A2(n_294),
.B1(n_828),
.B2(n_773),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_1212),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_1125),
.B(n_294),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1124),
.A2(n_614),
.B(n_620),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1071),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1061),
.A2(n_620),
.B(n_625),
.Y(n_1321)
);

AND2x4_ASAP7_75t_SL g1322 ( 
.A(n_1182),
.B(n_294),
.Y(n_1322)
);

NOR2xp67_ASAP7_75t_SL g1323 ( 
.A(n_1164),
.B(n_628),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1205),
.B(n_628),
.Y(n_1324)
);

NAND3xp33_ASAP7_75t_SL g1325 ( 
.A(n_1104),
.B(n_655),
.C(n_653),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1038),
.B(n_630),
.Y(n_1326)
);

O2A1O1Ixp5_ASAP7_75t_L g1327 ( 
.A1(n_1186),
.A2(n_655),
.B(n_635),
.C(n_643),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1030),
.A2(n_643),
.B1(n_634),
.B2(n_635),
.Y(n_1328)
);

BUFx12f_ASAP7_75t_L g1329 ( 
.A(n_1138),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1100),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1042),
.A2(n_625),
.B(n_652),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1204),
.B(n_634),
.Y(n_1332)
);

BUFx4f_ASAP7_75t_SL g1333 ( 
.A(n_1182),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1108),
.B(n_773),
.Y(n_1334)
);

O2A1O1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1179),
.A2(n_1159),
.B(n_1173),
.C(n_1044),
.Y(n_1335)
);

INVx2_ASAP7_75t_SL g1336 ( 
.A(n_1185),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1033),
.A2(n_625),
.B1(n_828),
.B2(n_773),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1064),
.Y(n_1338)
);

A2O1A1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1171),
.A2(n_828),
.B(n_773),
.C(n_13),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1066),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1045),
.A2(n_828),
.B1(n_773),
.B2(n_845),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1043),
.A2(n_828),
.B(n_773),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1069),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_1209),
.B(n_828),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1056),
.A2(n_845),
.B(n_682),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_SL g1346 ( 
.A(n_1209),
.B(n_845),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1164),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1156),
.A2(n_845),
.B(n_682),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1091),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1142),
.A2(n_845),
.B(n_682),
.Y(n_1350)
);

AOI221xp5_ASAP7_75t_L g1351 ( 
.A1(n_1159),
.A2(n_10),
.B1(n_12),
.B2(n_15),
.C(n_16),
.Y(n_1351)
);

OAI21xp33_ASAP7_75t_SL g1352 ( 
.A1(n_1053),
.A2(n_15),
.B(n_16),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1053),
.A2(n_845),
.B1(n_682),
.B2(n_20),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1195),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1142),
.A2(n_682),
.B(n_228),
.Y(n_1355)
);

OR2x6_ASAP7_75t_SL g1356 ( 
.A(n_1166),
.B(n_17),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1171),
.B(n_682),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1074),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_R g1359 ( 
.A(n_1065),
.B(n_100),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1097),
.B(n_1063),
.Y(n_1360)
);

NAND3xp33_ASAP7_75t_SL g1361 ( 
.A(n_1174),
.B(n_1197),
.C(n_1175),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1133),
.B(n_682),
.Y(n_1362)
);

OAI22x1_ASAP7_75t_L g1363 ( 
.A1(n_1208),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1096),
.Y(n_1364)
);

A2O1A1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1197),
.A2(n_19),
.B(n_22),
.C(n_23),
.Y(n_1365)
);

OAI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1140),
.A2(n_227),
.B(n_225),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1154),
.A2(n_222),
.B(n_219),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1085),
.A2(n_210),
.B(n_205),
.Y(n_1368)
);

A2O1A1Ixp33_ASAP7_75t_L g1369 ( 
.A1(n_1158),
.A2(n_25),
.B(n_26),
.C(n_28),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1098),
.B(n_188),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1141),
.Y(n_1371)
);

O2A1O1Ixp33_ASAP7_75t_L g1372 ( 
.A1(n_1173),
.A2(n_25),
.B(n_26),
.C(n_30),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1208),
.B(n_30),
.Y(n_1373)
);

INVx3_ASAP7_75t_SL g1374 ( 
.A(n_1054),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1058),
.A2(n_175),
.B(n_164),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1046),
.A2(n_152),
.B1(n_151),
.B2(n_150),
.Y(n_1376)
);

O2A1O1Ixp33_ASAP7_75t_L g1377 ( 
.A1(n_1049),
.A2(n_31),
.B(n_33),
.C(n_36),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_SL g1378 ( 
.A(n_1098),
.B(n_145),
.Y(n_1378)
);

BUFx8_ASAP7_75t_L g1379 ( 
.A(n_1281),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1261),
.A2(n_1090),
.B(n_1146),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1229),
.B(n_1107),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1215),
.Y(n_1382)
);

AND2x4_ASAP7_75t_L g1383 ( 
.A(n_1245),
.B(n_1107),
.Y(n_1383)
);

NOR2xp67_ASAP7_75t_SL g1384 ( 
.A(n_1274),
.B(n_1071),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1222),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_L g1386 ( 
.A(n_1349),
.Y(n_1386)
);

INVx3_ASAP7_75t_L g1387 ( 
.A(n_1347),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1236),
.Y(n_1388)
);

O2A1O1Ixp5_ASAP7_75t_L g1389 ( 
.A1(n_1239),
.A2(n_1067),
.B(n_1213),
.C(n_1199),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_SL g1390 ( 
.A1(n_1255),
.A2(n_1070),
.B(n_1158),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1307),
.A2(n_1080),
.B(n_1083),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1294),
.A2(n_1170),
.B(n_1187),
.Y(n_1392)
);

AO31x2_ASAP7_75t_L g1393 ( 
.A1(n_1251),
.A2(n_1093),
.A3(n_1101),
.B(n_1180),
.Y(n_1393)
);

O2A1O1Ixp33_ASAP7_75t_L g1394 ( 
.A1(n_1216),
.A2(n_1047),
.B(n_1072),
.C(n_1210),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1313),
.B(n_1145),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1285),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1332),
.Y(n_1397)
);

AO21x1_ASAP7_75t_L g1398 ( 
.A1(n_1217),
.A2(n_1176),
.B(n_1177),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1319),
.A2(n_1161),
.B(n_1190),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1307),
.A2(n_1153),
.B(n_1058),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1280),
.A2(n_1150),
.B(n_1151),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1349),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1313),
.B(n_1169),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1216),
.B(n_1174),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1227),
.A2(n_1153),
.B(n_1081),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1221),
.A2(n_1103),
.B(n_1114),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_1240),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1324),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1291),
.A2(n_1257),
.B(n_1321),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1230),
.B(n_1183),
.Y(n_1410)
);

NAND4xp25_ASAP7_75t_SL g1411 ( 
.A(n_1351),
.B(n_1117),
.C(n_1131),
.D(n_1113),
.Y(n_1411)
);

INVxp67_ASAP7_75t_SL g1412 ( 
.A(n_1235),
.Y(n_1412)
);

O2A1O1Ixp33_ASAP7_75t_SL g1413 ( 
.A1(n_1346),
.A2(n_1193),
.B(n_1122),
.C(n_1127),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1310),
.B(n_1121),
.Y(n_1414)
);

AO31x2_ASAP7_75t_L g1415 ( 
.A1(n_1244),
.A2(n_1202),
.A3(n_1201),
.B(n_1211),
.Y(n_1415)
);

AOI221x1_ASAP7_75t_L g1416 ( 
.A1(n_1225),
.A2(n_1115),
.B1(n_1137),
.B2(n_1126),
.C(n_1165),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1228),
.A2(n_1103),
.B(n_1081),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1357),
.A2(n_1114),
.B(n_1184),
.Y(n_1418)
);

A2O1A1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1255),
.A2(n_1065),
.B(n_1162),
.C(n_1110),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1245),
.B(n_1091),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1311),
.B(n_1132),
.Y(n_1421)
);

AO31x2_ASAP7_75t_L g1422 ( 
.A1(n_1288),
.A2(n_1094),
.A3(n_1102),
.B(n_1112),
.Y(n_1422)
);

NOR2xp67_ASAP7_75t_L g1423 ( 
.A(n_1303),
.B(n_1360),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1218),
.A2(n_1184),
.B(n_1134),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1335),
.A2(n_1162),
.B(n_1139),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1305),
.A2(n_1143),
.B(n_1160),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1258),
.A2(n_1196),
.B(n_1189),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1330),
.B(n_1149),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1268),
.Y(n_1429)
);

OR2x6_ASAP7_75t_L g1430 ( 
.A(n_1329),
.B(n_1106),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1226),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1371),
.Y(n_1432)
);

AO31x2_ASAP7_75t_L g1433 ( 
.A1(n_1331),
.A2(n_1178),
.A3(n_1130),
.B(n_1157),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1286),
.Y(n_1434)
);

OAI21xp5_ASAP7_75t_SL g1435 ( 
.A1(n_1259),
.A2(n_1172),
.B(n_1160),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1266),
.A2(n_1157),
.B(n_1172),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1302),
.B(n_1272),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1223),
.A2(n_1106),
.B(n_144),
.Y(n_1438)
);

OAI22x1_ASAP7_75t_L g1439 ( 
.A1(n_1259),
.A2(n_1106),
.B1(n_37),
.B2(n_39),
.Y(n_1439)
);

AO31x2_ASAP7_75t_L g1440 ( 
.A1(n_1348),
.A2(n_33),
.A3(n_40),
.B(n_41),
.Y(n_1440)
);

O2A1O1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1264),
.A2(n_40),
.B(n_50),
.C(n_51),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1284),
.B(n_51),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1238),
.A2(n_136),
.B(n_131),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1297),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1214),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1349),
.B(n_129),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1264),
.B(n_52),
.Y(n_1447)
);

OAI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1232),
.A2(n_125),
.B(n_123),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1293),
.A2(n_122),
.B(n_117),
.Y(n_1449)
);

AOI221xp5_ASAP7_75t_L g1450 ( 
.A1(n_1278),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.C(n_55),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1248),
.A2(n_113),
.B(n_111),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1299),
.Y(n_1452)
);

O2A1O1Ixp33_ASAP7_75t_L g1453 ( 
.A1(n_1277),
.A2(n_53),
.B(n_54),
.C(n_55),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1293),
.A2(n_105),
.B(n_59),
.Y(n_1454)
);

O2A1O1Ixp33_ASAP7_75t_SL g1455 ( 
.A1(n_1344),
.A2(n_1366),
.B(n_1369),
.C(n_1365),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1303),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_1456)
);

NAND2x1_ASAP7_75t_L g1457 ( 
.A(n_1347),
.B(n_63),
.Y(n_1457)
);

INVx3_ASAP7_75t_L g1458 ( 
.A(n_1242),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1234),
.A2(n_1237),
.B1(n_1279),
.B2(n_1290),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1279),
.B(n_64),
.Y(n_1460)
);

CKINVDCx11_ASAP7_75t_R g1461 ( 
.A(n_1356),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1342),
.A2(n_67),
.B(n_70),
.Y(n_1462)
);

A2O1A1Ixp33_ASAP7_75t_L g1463 ( 
.A1(n_1290),
.A2(n_67),
.B(n_70),
.C(n_71),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1340),
.Y(n_1464)
);

AO31x2_ASAP7_75t_L g1465 ( 
.A1(n_1339),
.A2(n_72),
.A3(n_77),
.B(n_78),
.Y(n_1465)
);

NAND2x1p5_ASAP7_75t_L g1466 ( 
.A(n_1317),
.B(n_72),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1343),
.Y(n_1467)
);

OA21x2_ASAP7_75t_L g1468 ( 
.A1(n_1308),
.A2(n_77),
.B(n_78),
.Y(n_1468)
);

A2O1A1Ixp33_ASAP7_75t_L g1469 ( 
.A1(n_1283),
.A2(n_81),
.B(n_83),
.C(n_84),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1300),
.Y(n_1470)
);

O2A1O1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1373),
.A2(n_81),
.B(n_88),
.C(n_89),
.Y(n_1471)
);

INVx1_ASAP7_75t_SL g1472 ( 
.A(n_1224),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1275),
.A2(n_89),
.B(n_92),
.Y(n_1473)
);

AO31x2_ASAP7_75t_L g1474 ( 
.A1(n_1345),
.A2(n_1328),
.A3(n_1249),
.B(n_1368),
.Y(n_1474)
);

AO31x2_ASAP7_75t_L g1475 ( 
.A1(n_1337),
.A2(n_1341),
.A3(n_1247),
.B(n_1367),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1262),
.B(n_1276),
.Y(n_1476)
);

AOI221xp5_ASAP7_75t_SL g1477 ( 
.A1(n_1363),
.A2(n_1372),
.B1(n_1377),
.B2(n_1352),
.C(n_1315),
.Y(n_1477)
);

NOR2xp67_ASAP7_75t_L g1478 ( 
.A(n_1336),
.B(n_1298),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1295),
.B(n_1284),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1273),
.B(n_1265),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1233),
.A2(n_1349),
.B1(n_1338),
.B2(n_1358),
.Y(n_1481)
);

OAI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1241),
.A2(n_1334),
.B(n_1282),
.Y(n_1482)
);

BUFx4f_ASAP7_75t_L g1483 ( 
.A(n_1231),
.Y(n_1483)
);

AO32x2_ASAP7_75t_L g1484 ( 
.A1(n_1260),
.A2(n_1376),
.A3(n_1250),
.B1(n_1361),
.B2(n_1252),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1364),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1235),
.B(n_1265),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1295),
.B(n_1231),
.Y(n_1487)
);

AOI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1233),
.A2(n_1292),
.B(n_1252),
.Y(n_1488)
);

A2O1A1Ixp33_ASAP7_75t_L g1489 ( 
.A1(n_1283),
.A2(n_1312),
.B(n_1326),
.C(n_1287),
.Y(n_1489)
);

AO31x2_ASAP7_75t_L g1490 ( 
.A1(n_1350),
.A2(n_1375),
.A3(n_1355),
.B(n_1362),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1219),
.B(n_1271),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_L g1492 ( 
.A(n_1242),
.Y(n_1492)
);

OAI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1316),
.A2(n_1327),
.B(n_1353),
.Y(n_1493)
);

AOI211x1_ASAP7_75t_L g1494 ( 
.A1(n_1378),
.A2(n_1325),
.B(n_1318),
.C(n_1263),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1320),
.Y(n_1495)
);

BUFx2_ASAP7_75t_L g1496 ( 
.A(n_1219),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_SL g1497 ( 
.A(n_1220),
.B(n_1269),
.Y(n_1497)
);

NAND3x1_ASAP7_75t_L g1498 ( 
.A(n_1315),
.B(n_1296),
.C(n_1374),
.Y(n_1498)
);

AOI221x1_ASAP7_75t_L g1499 ( 
.A1(n_1289),
.A2(n_1370),
.B1(n_1253),
.B2(n_1254),
.C(n_1267),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1301),
.B(n_1320),
.Y(n_1500)
);

NOR2xp67_ASAP7_75t_L g1501 ( 
.A(n_1354),
.B(n_1301),
.Y(n_1501)
);

INVxp33_ASAP7_75t_L g1502 ( 
.A(n_1246),
.Y(n_1502)
);

CKINVDCx20_ASAP7_75t_R g1503 ( 
.A(n_1333),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1306),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1309),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1306),
.A2(n_1256),
.B(n_1304),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1370),
.B(n_1322),
.Y(n_1507)
);

INVx2_ASAP7_75t_SL g1508 ( 
.A(n_1333),
.Y(n_1508)
);

AOI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1271),
.A2(n_1314),
.B1(n_1323),
.B2(n_1353),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1316),
.A2(n_1314),
.B(n_1243),
.Y(n_1510)
);

AOI221x1_ASAP7_75t_L g1511 ( 
.A1(n_1242),
.A2(n_1243),
.B1(n_1270),
.B2(n_1314),
.C(n_1359),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1242),
.Y(n_1512)
);

OAI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1243),
.A2(n_1270),
.B(n_1261),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1243),
.B(n_1270),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1270),
.A2(n_1229),
.B1(n_1227),
.B2(n_1313),
.Y(n_1515)
);

BUFx2_ASAP7_75t_L g1516 ( 
.A(n_1219),
.Y(n_1516)
);

INVx2_ASAP7_75t_SL g1517 ( 
.A(n_1317),
.Y(n_1517)
);

OA21x2_ASAP7_75t_L g1518 ( 
.A1(n_1218),
.A2(n_1327),
.B(n_1308),
.Y(n_1518)
);

BUFx10_ASAP7_75t_L g1519 ( 
.A(n_1286),
.Y(n_1519)
);

A2O1A1Ixp33_ASAP7_75t_L g1520 ( 
.A1(n_1216),
.A2(n_1217),
.B(n_1075),
.C(n_1032),
.Y(n_1520)
);

BUFx6f_ASAP7_75t_L g1521 ( 
.A(n_1349),
.Y(n_1521)
);

A2O1A1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1216),
.A2(n_1217),
.B(n_1075),
.C(n_1032),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1313),
.B(n_855),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1215),
.Y(n_1524)
);

AO32x2_ASAP7_75t_L g1525 ( 
.A1(n_1225),
.A2(n_1155),
.A3(n_1244),
.B1(n_1070),
.B2(n_1249),
.Y(n_1525)
);

AOI221xp5_ASAP7_75t_L g1526 ( 
.A1(n_1255),
.A2(n_1264),
.B1(n_1259),
.B2(n_1216),
.C(n_816),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1261),
.A2(n_1294),
.B(n_1319),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1216),
.A2(n_1259),
.B1(n_1264),
.B2(n_1255),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1229),
.B(n_1230),
.Y(n_1529)
);

AO21x1_ASAP7_75t_L g1530 ( 
.A1(n_1217),
.A2(n_1200),
.B(n_1366),
.Y(n_1530)
);

OAI22x1_ASAP7_75t_L g1531 ( 
.A1(n_1216),
.A2(n_1313),
.B1(n_1068),
.B2(n_1057),
.Y(n_1531)
);

OA21x2_ASAP7_75t_L g1532 ( 
.A1(n_1218),
.A2(n_1327),
.B(n_1308),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1215),
.Y(n_1533)
);

AOI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1229),
.A2(n_1025),
.B(n_1105),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1236),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1229),
.A2(n_1025),
.B(n_1105),
.Y(n_1536)
);

O2A1O1Ixp33_ASAP7_75t_SL g1537 ( 
.A1(n_1346),
.A2(n_1147),
.B(n_1159),
.C(n_1118),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1261),
.A2(n_1294),
.B(n_1319),
.Y(n_1538)
);

CKINVDCx6p67_ASAP7_75t_R g1539 ( 
.A(n_1274),
.Y(n_1539)
);

OAI21x1_ASAP7_75t_L g1540 ( 
.A1(n_1261),
.A2(n_1294),
.B(n_1319),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1215),
.Y(n_1541)
);

AOI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1229),
.A2(n_1025),
.B(n_1105),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1229),
.A2(n_1025),
.B(n_1105),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1215),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1215),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1245),
.B(n_1349),
.Y(n_1546)
);

AO32x2_ASAP7_75t_L g1547 ( 
.A1(n_1225),
.A2(n_1155),
.A3(n_1244),
.B1(n_1070),
.B2(n_1249),
.Y(n_1547)
);

AO31x2_ASAP7_75t_L g1548 ( 
.A1(n_1251),
.A2(n_1213),
.A3(n_1244),
.B(n_1067),
.Y(n_1548)
);

AO32x2_ASAP7_75t_L g1549 ( 
.A1(n_1225),
.A2(n_1155),
.A3(n_1244),
.B1(n_1070),
.B2(n_1249),
.Y(n_1549)
);

AO31x2_ASAP7_75t_L g1550 ( 
.A1(n_1251),
.A2(n_1213),
.A3(n_1244),
.B(n_1067),
.Y(n_1550)
);

AO31x2_ASAP7_75t_L g1551 ( 
.A1(n_1251),
.A2(n_1213),
.A3(n_1244),
.B(n_1067),
.Y(n_1551)
);

BUFx6f_ASAP7_75t_L g1552 ( 
.A(n_1349),
.Y(n_1552)
);

AOI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1229),
.A2(n_1025),
.B(n_1105),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1229),
.B(n_1230),
.Y(n_1554)
);

AOI21xp5_ASAP7_75t_L g1555 ( 
.A1(n_1229),
.A2(n_1025),
.B(n_1105),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1215),
.Y(n_1556)
);

OAI22x1_ASAP7_75t_L g1557 ( 
.A1(n_1216),
.A2(n_1313),
.B1(n_1068),
.B2(n_1057),
.Y(n_1557)
);

AOI221x1_ASAP7_75t_L g1558 ( 
.A1(n_1225),
.A2(n_1366),
.B1(n_1278),
.B2(n_1255),
.C(n_1264),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1529),
.B(n_1554),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1528),
.A2(n_1526),
.B1(n_1447),
.B2(n_1404),
.Y(n_1560)
);

INVxp67_ASAP7_75t_SL g1561 ( 
.A(n_1486),
.Y(n_1561)
);

BUFx10_ASAP7_75t_L g1562 ( 
.A(n_1434),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1437),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1460),
.A2(n_1459),
.B1(n_1557),
.B2(n_1531),
.Y(n_1564)
);

OAI22xp33_ASAP7_75t_R g1565 ( 
.A1(n_1523),
.A2(n_1479),
.B1(n_1407),
.B2(n_1442),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1546),
.B(n_1420),
.Y(n_1566)
);

OAI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1558),
.A2(n_1390),
.B1(n_1509),
.B2(n_1439),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1530),
.A2(n_1448),
.B1(n_1491),
.B2(n_1487),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_L g1569 ( 
.A(n_1483),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1396),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1535),
.Y(n_1571)
);

CKINVDCx20_ASAP7_75t_R g1572 ( 
.A(n_1503),
.Y(n_1572)
);

INVx1_ASAP7_75t_SL g1573 ( 
.A(n_1496),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1450),
.A2(n_1423),
.B1(n_1443),
.B2(n_1411),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_SL g1575 ( 
.A1(n_1493),
.A2(n_1456),
.B1(n_1483),
.B2(n_1454),
.Y(n_1575)
);

CKINVDCx6p67_ASAP7_75t_R g1576 ( 
.A(n_1519),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_1516),
.Y(n_1577)
);

OAI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1520),
.A2(n_1522),
.B1(n_1431),
.B2(n_1476),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1432),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1408),
.A2(n_1515),
.B1(n_1397),
.B2(n_1478),
.Y(n_1580)
);

INVx8_ASAP7_75t_L g1581 ( 
.A(n_1492),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_SL g1582 ( 
.A1(n_1466),
.A2(n_1408),
.B1(n_1431),
.B2(n_1397),
.Y(n_1582)
);

CKINVDCx11_ASAP7_75t_R g1583 ( 
.A(n_1519),
.Y(n_1583)
);

CKINVDCx14_ASAP7_75t_R g1584 ( 
.A(n_1539),
.Y(n_1584)
);

AOI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1498),
.A2(n_1507),
.B1(n_1502),
.B2(n_1497),
.Y(n_1585)
);

BUFx2_ASAP7_75t_L g1586 ( 
.A(n_1379),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1445),
.Y(n_1587)
);

OAI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1381),
.A2(n_1410),
.B1(n_1511),
.B2(n_1472),
.Y(n_1588)
);

INVx1_ASAP7_75t_SL g1589 ( 
.A(n_1421),
.Y(n_1589)
);

BUFx3_ASAP7_75t_L g1590 ( 
.A(n_1379),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1505),
.A2(n_1461),
.B1(n_1420),
.B2(n_1438),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_1517),
.Y(n_1592)
);

CKINVDCx11_ASAP7_75t_R g1593 ( 
.A(n_1430),
.Y(n_1593)
);

BUFx3_ASAP7_75t_L g1594 ( 
.A(n_1508),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1444),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1505),
.A2(n_1430),
.B1(n_1398),
.B2(n_1446),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1464),
.Y(n_1597)
);

INVx8_ASAP7_75t_L g1598 ( 
.A(n_1492),
.Y(n_1598)
);

INVx5_ASAP7_75t_SL g1599 ( 
.A(n_1386),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1464),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1467),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1446),
.A2(n_1403),
.B1(n_1395),
.B2(n_1480),
.Y(n_1602)
);

INVx4_ASAP7_75t_L g1603 ( 
.A(n_1386),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_1386),
.Y(n_1604)
);

BUFx4f_ASAP7_75t_L g1605 ( 
.A(n_1402),
.Y(n_1605)
);

BUFx12f_ASAP7_75t_L g1606 ( 
.A(n_1402),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1467),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1452),
.Y(n_1608)
);

BUFx8_ASAP7_75t_L g1609 ( 
.A(n_1402),
.Y(n_1609)
);

AOI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1501),
.A2(n_1435),
.B1(n_1477),
.B2(n_1384),
.Y(n_1610)
);

BUFx12f_ASAP7_75t_L g1611 ( 
.A(n_1521),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1481),
.A2(n_1504),
.B1(n_1449),
.B2(n_1470),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1382),
.Y(n_1613)
);

BUFx3_ASAP7_75t_L g1614 ( 
.A(n_1521),
.Y(n_1614)
);

OAI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1414),
.A2(n_1428),
.B1(n_1457),
.B2(n_1412),
.Y(n_1615)
);

BUFx3_ASAP7_75t_L g1616 ( 
.A(n_1521),
.Y(n_1616)
);

BUFx4f_ASAP7_75t_SL g1617 ( 
.A(n_1552),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1524),
.Y(n_1618)
);

CKINVDCx11_ASAP7_75t_R g1619 ( 
.A(n_1552),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1485),
.B(n_1500),
.Y(n_1620)
);

AOI21xp33_ASAP7_75t_L g1621 ( 
.A1(n_1394),
.A2(n_1441),
.B(n_1453),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1533),
.B(n_1541),
.Y(n_1622)
);

BUFx8_ASAP7_75t_L g1623 ( 
.A(n_1546),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_SL g1624 ( 
.A1(n_1391),
.A2(n_1468),
.B1(n_1463),
.B2(n_1547),
.Y(n_1624)
);

BUFx10_ASAP7_75t_L g1625 ( 
.A(n_1383),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1385),
.Y(n_1626)
);

BUFx12f_ASAP7_75t_L g1627 ( 
.A(n_1383),
.Y(n_1627)
);

BUFx8_ASAP7_75t_SL g1628 ( 
.A(n_1387),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1544),
.Y(n_1629)
);

CKINVDCx11_ASAP7_75t_R g1630 ( 
.A(n_1429),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1425),
.A2(n_1424),
.B(n_1555),
.Y(n_1631)
);

INVx8_ASAP7_75t_L g1632 ( 
.A(n_1514),
.Y(n_1632)
);

OAI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1545),
.A2(n_1556),
.B1(n_1469),
.B2(n_1494),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_SL g1634 ( 
.A1(n_1468),
.A2(n_1549),
.B1(n_1547),
.B2(n_1525),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1556),
.B(n_1553),
.Y(n_1635)
);

INVx6_ASAP7_75t_L g1636 ( 
.A(n_1458),
.Y(n_1636)
);

BUFx4f_ASAP7_75t_SL g1637 ( 
.A(n_1458),
.Y(n_1637)
);

BUFx6f_ASAP7_75t_L g1638 ( 
.A(n_1512),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1429),
.Y(n_1639)
);

BUFx2_ASAP7_75t_SL g1640 ( 
.A(n_1512),
.Y(n_1640)
);

AOI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1455),
.A2(n_1489),
.B1(n_1419),
.B2(n_1495),
.Y(n_1641)
);

OAI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1499),
.A2(n_1495),
.B1(n_1462),
.B2(n_1536),
.Y(n_1642)
);

BUFx10_ASAP7_75t_L g1643 ( 
.A(n_1471),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1482),
.A2(n_1405),
.B1(n_1542),
.B2(n_1543),
.Y(n_1644)
);

CKINVDCx11_ASAP7_75t_R g1645 ( 
.A(n_1440),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1387),
.Y(n_1646)
);

BUFx6f_ASAP7_75t_L g1647 ( 
.A(n_1510),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1433),
.Y(n_1648)
);

CKINVDCx11_ASAP7_75t_R g1649 ( 
.A(n_1440),
.Y(n_1649)
);

BUFx3_ASAP7_75t_L g1650 ( 
.A(n_1506),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1433),
.Y(n_1651)
);

INVx4_ASAP7_75t_L g1652 ( 
.A(n_1518),
.Y(n_1652)
);

CKINVDCx8_ASAP7_75t_R g1653 ( 
.A(n_1518),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1433),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1427),
.Y(n_1655)
);

INVx6_ASAP7_75t_L g1656 ( 
.A(n_1537),
.Y(n_1656)
);

INVx6_ASAP7_75t_L g1657 ( 
.A(n_1413),
.Y(n_1657)
);

OAI22xp5_ASAP7_75t_SL g1658 ( 
.A1(n_1465),
.A2(n_1532),
.B1(n_1549),
.B2(n_1547),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1534),
.B(n_1400),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1473),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_1488),
.Y(n_1661)
);

INVx1_ASAP7_75t_SL g1662 ( 
.A(n_1532),
.Y(n_1662)
);

INVx6_ASAP7_75t_L g1663 ( 
.A(n_1465),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1465),
.B(n_1440),
.Y(n_1664)
);

BUFx6f_ASAP7_75t_L g1665 ( 
.A(n_1451),
.Y(n_1665)
);

CKINVDCx20_ASAP7_75t_R g1666 ( 
.A(n_1406),
.Y(n_1666)
);

BUFx6f_ASAP7_75t_L g1667 ( 
.A(n_1513),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_SL g1668 ( 
.A1(n_1525),
.A2(n_1549),
.B1(n_1484),
.B2(n_1399),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1436),
.Y(n_1669)
);

BUFx8_ASAP7_75t_L g1670 ( 
.A(n_1484),
.Y(n_1670)
);

CKINVDCx20_ASAP7_75t_R g1671 ( 
.A(n_1417),
.Y(n_1671)
);

INVx3_ASAP7_75t_SL g1672 ( 
.A(n_1389),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1422),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_SL g1674 ( 
.A1(n_1525),
.A2(n_1484),
.B1(n_1418),
.B2(n_1426),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1393),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1422),
.Y(n_1676)
);

AOI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1392),
.A2(n_1409),
.B1(n_1401),
.B2(n_1380),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1527),
.A2(n_1540),
.B1(n_1538),
.B2(n_1474),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_SL g1679 ( 
.A1(n_1548),
.A2(n_1551),
.B1(n_1550),
.B2(n_1474),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1393),
.Y(n_1680)
);

CKINVDCx11_ASAP7_75t_R g1681 ( 
.A(n_1548),
.Y(n_1681)
);

CKINVDCx11_ASAP7_75t_R g1682 ( 
.A(n_1548),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1416),
.A2(n_1550),
.B1(n_1551),
.B2(n_1474),
.Y(n_1683)
);

OAI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1550),
.A2(n_1551),
.B1(n_1393),
.B2(n_1475),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1490),
.Y(n_1685)
);

OAI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1475),
.A2(n_1526),
.B1(n_1447),
.B2(n_1057),
.Y(n_1686)
);

BUFx4_ASAP7_75t_SL g1687 ( 
.A(n_1490),
.Y(n_1687)
);

BUFx2_ASAP7_75t_L g1688 ( 
.A(n_1490),
.Y(n_1688)
);

BUFx2_ASAP7_75t_SL g1689 ( 
.A(n_1415),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1415),
.B(n_1529),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1526),
.A2(n_1528),
.B1(n_1447),
.B2(n_1057),
.Y(n_1691)
);

INVx6_ASAP7_75t_L g1692 ( 
.A(n_1379),
.Y(n_1692)
);

INVx5_ASAP7_75t_L g1693 ( 
.A(n_1492),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1526),
.A2(n_1528),
.B1(n_1447),
.B2(n_1057),
.Y(n_1694)
);

INVx6_ASAP7_75t_L g1695 ( 
.A(n_1379),
.Y(n_1695)
);

INVx6_ASAP7_75t_L g1696 ( 
.A(n_1379),
.Y(n_1696)
);

BUFx3_ASAP7_75t_L g1697 ( 
.A(n_1379),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1526),
.A2(n_1528),
.B1(n_1447),
.B2(n_1057),
.Y(n_1698)
);

INVx3_ASAP7_75t_L g1699 ( 
.A(n_1386),
.Y(n_1699)
);

OAI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1528),
.A2(n_1526),
.B1(n_1229),
.B2(n_1147),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1388),
.Y(n_1701)
);

INVxp67_ASAP7_75t_SL g1702 ( 
.A(n_1486),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1526),
.A2(n_1528),
.B1(n_1447),
.B2(n_1057),
.Y(n_1703)
);

CKINVDCx6p67_ASAP7_75t_R g1704 ( 
.A(n_1519),
.Y(n_1704)
);

CKINVDCx6p67_ASAP7_75t_R g1705 ( 
.A(n_1519),
.Y(n_1705)
);

AOI21xp33_ASAP7_75t_L g1706 ( 
.A1(n_1528),
.A2(n_1526),
.B(n_1390),
.Y(n_1706)
);

AOI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1528),
.A2(n_1526),
.B1(n_1057),
.B2(n_1068),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1526),
.A2(n_1528),
.B1(n_1447),
.B2(n_1057),
.Y(n_1708)
);

BUFx3_ASAP7_75t_L g1709 ( 
.A(n_1379),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1528),
.A2(n_1526),
.B1(n_1229),
.B2(n_1147),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_1434),
.Y(n_1711)
);

INVx4_ASAP7_75t_L g1712 ( 
.A(n_1492),
.Y(n_1712)
);

CKINVDCx20_ASAP7_75t_R g1713 ( 
.A(n_1434),
.Y(n_1713)
);

CKINVDCx11_ASAP7_75t_R g1714 ( 
.A(n_1519),
.Y(n_1714)
);

BUFx3_ASAP7_75t_L g1715 ( 
.A(n_1379),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1388),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_SL g1717 ( 
.A1(n_1447),
.A2(n_1057),
.B1(n_1068),
.B2(n_1216),
.Y(n_1717)
);

OAI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1526),
.A2(n_1447),
.B1(n_1057),
.B2(n_1068),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1388),
.Y(n_1719)
);

AOI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1391),
.A2(n_1448),
.B(n_1493),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_SL g1721 ( 
.A1(n_1447),
.A2(n_1057),
.B1(n_1068),
.B2(n_1216),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1526),
.A2(n_1528),
.B1(n_1447),
.B2(n_1057),
.Y(n_1722)
);

INVx6_ASAP7_75t_L g1723 ( 
.A(n_1379),
.Y(n_1723)
);

BUFx2_ASAP7_75t_L g1724 ( 
.A(n_1496),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1388),
.Y(n_1725)
);

BUFx10_ASAP7_75t_L g1726 ( 
.A(n_1434),
.Y(n_1726)
);

INVx6_ASAP7_75t_L g1727 ( 
.A(n_1379),
.Y(n_1727)
);

BUFx2_ASAP7_75t_L g1728 ( 
.A(n_1496),
.Y(n_1728)
);

CKINVDCx20_ASAP7_75t_R g1729 ( 
.A(n_1434),
.Y(n_1729)
);

CKINVDCx5p33_ASAP7_75t_R g1730 ( 
.A(n_1434),
.Y(n_1730)
);

INVx1_ASAP7_75t_SL g1731 ( 
.A(n_1437),
.Y(n_1731)
);

INVx6_ASAP7_75t_L g1732 ( 
.A(n_1379),
.Y(n_1732)
);

INVx1_ASAP7_75t_SL g1733 ( 
.A(n_1437),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1526),
.A2(n_1528),
.B1(n_1447),
.B2(n_1057),
.Y(n_1734)
);

INVx8_ASAP7_75t_L g1735 ( 
.A(n_1492),
.Y(n_1735)
);

BUFx6f_ASAP7_75t_L g1736 ( 
.A(n_1483),
.Y(n_1736)
);

INVx6_ASAP7_75t_L g1737 ( 
.A(n_1379),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1388),
.Y(n_1738)
);

OAI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1526),
.A2(n_1447),
.B1(n_1057),
.B2(n_1068),
.Y(n_1739)
);

INVx6_ASAP7_75t_L g1740 ( 
.A(n_1379),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1664),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1690),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1690),
.Y(n_1743)
);

OAI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1691),
.A2(n_1698),
.B(n_1694),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_SL g1745 ( 
.A(n_1718),
.B(n_1739),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1635),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1613),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1635),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1618),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1648),
.Y(n_1750)
);

AO31x2_ASAP7_75t_L g1751 ( 
.A1(n_1720),
.A2(n_1683),
.A3(n_1652),
.B(n_1688),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1651),
.Y(n_1752)
);

OA21x2_ASAP7_75t_L g1753 ( 
.A1(n_1720),
.A2(n_1631),
.B(n_1659),
.Y(n_1753)
);

INVxp67_ASAP7_75t_SL g1754 ( 
.A(n_1561),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1579),
.Y(n_1755)
);

BUFx3_ASAP7_75t_L g1756 ( 
.A(n_1628),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1654),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1675),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1595),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1661),
.B(n_1597),
.Y(n_1760)
);

BUFx3_ASAP7_75t_L g1761 ( 
.A(n_1609),
.Y(n_1761)
);

BUFx6f_ASAP7_75t_L g1762 ( 
.A(n_1569),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1658),
.Y(n_1763)
);

CKINVDCx10_ASAP7_75t_R g1764 ( 
.A(n_1584),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1600),
.B(n_1601),
.Y(n_1765)
);

BUFx2_ASAP7_75t_L g1766 ( 
.A(n_1685),
.Y(n_1766)
);

BUFx6f_ASAP7_75t_L g1767 ( 
.A(n_1569),
.Y(n_1767)
);

INVx3_ASAP7_75t_L g1768 ( 
.A(n_1667),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1622),
.Y(n_1769)
);

OA21x2_ASAP7_75t_L g1770 ( 
.A1(n_1631),
.A2(n_1659),
.B(n_1644),
.Y(n_1770)
);

OAI21x1_ASAP7_75t_L g1771 ( 
.A1(n_1678),
.A2(n_1660),
.B(n_1655),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1607),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1622),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1683),
.B(n_1680),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1639),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1702),
.B(n_1673),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1676),
.B(n_1684),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1560),
.A2(n_1722),
.B1(n_1703),
.B2(n_1734),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1663),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1668),
.B(n_1620),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1573),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1668),
.B(n_1663),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1571),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1681),
.B(n_1682),
.Y(n_1784)
);

AOI21x1_ASAP7_75t_L g1785 ( 
.A1(n_1669),
.A2(n_1578),
.B(n_1633),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1608),
.Y(n_1786)
);

AOI21xp33_ASAP7_75t_L g1787 ( 
.A1(n_1560),
.A2(n_1686),
.B(n_1708),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1626),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1647),
.Y(n_1789)
);

INVx2_ASAP7_75t_SL g1790 ( 
.A(n_1632),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1578),
.B(n_1563),
.Y(n_1791)
);

INVx3_ASAP7_75t_L g1792 ( 
.A(n_1667),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1647),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1647),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1687),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1629),
.Y(n_1796)
);

BUFx3_ASAP7_75t_L g1797 ( 
.A(n_1609),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1706),
.A2(n_1721),
.B1(n_1717),
.B2(n_1707),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1650),
.Y(n_1799)
);

BUFx2_ASAP7_75t_L g1800 ( 
.A(n_1671),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1689),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1662),
.Y(n_1802)
);

AO21x1_ASAP7_75t_SL g1803 ( 
.A1(n_1621),
.A2(n_1641),
.B(n_1568),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1662),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1679),
.B(n_1634),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1653),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1679),
.Y(n_1807)
);

INVx3_ASAP7_75t_L g1808 ( 
.A(n_1667),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1652),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1670),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1670),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1634),
.Y(n_1812)
);

AND2x6_ASAP7_75t_L g1813 ( 
.A(n_1599),
.B(n_1610),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1656),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_L g1815 ( 
.A(n_1573),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1564),
.B(n_1624),
.Y(n_1816)
);

OAI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1717),
.A2(n_1721),
.B1(n_1574),
.B2(n_1580),
.Y(n_1817)
);

HB1xp67_ASAP7_75t_L g1818 ( 
.A(n_1577),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1559),
.B(n_1731),
.Y(n_1819)
);

INVxp67_ASAP7_75t_L g1820 ( 
.A(n_1724),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1656),
.Y(n_1821)
);

INVx2_ASAP7_75t_SL g1822 ( 
.A(n_1632),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1559),
.B(n_1731),
.Y(n_1823)
);

AOI21x1_ASAP7_75t_L g1824 ( 
.A1(n_1633),
.A2(n_1710),
.B(n_1700),
.Y(n_1824)
);

HB1xp67_ASAP7_75t_L g1825 ( 
.A(n_1577),
.Y(n_1825)
);

OAI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1706),
.A2(n_1710),
.B(n_1700),
.Y(n_1826)
);

OAI21x1_ASAP7_75t_L g1827 ( 
.A1(n_1677),
.A2(n_1612),
.B(n_1596),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1728),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1656),
.Y(n_1829)
);

AO21x1_ASAP7_75t_SL g1830 ( 
.A1(n_1621),
.A2(n_1591),
.B(n_1602),
.Y(n_1830)
);

BUFx6f_ASAP7_75t_L g1831 ( 
.A(n_1569),
.Y(n_1831)
);

AOI22xp33_ASAP7_75t_L g1832 ( 
.A1(n_1567),
.A2(n_1575),
.B1(n_1643),
.B2(n_1565),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1666),
.B(n_1736),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1738),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1674),
.Y(n_1835)
);

INVx3_ASAP7_75t_L g1836 ( 
.A(n_1665),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1570),
.Y(n_1837)
);

BUFx2_ASAP7_75t_L g1838 ( 
.A(n_1672),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1624),
.B(n_1674),
.Y(n_1839)
);

BUFx3_ASAP7_75t_L g1840 ( 
.A(n_1736),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1657),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1575),
.A2(n_1643),
.B1(n_1582),
.B2(n_1649),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1657),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_1583),
.Y(n_1844)
);

AO21x2_ASAP7_75t_L g1845 ( 
.A1(n_1642),
.A2(n_1615),
.B(n_1588),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1657),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1701),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1716),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1719),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1725),
.Y(n_1850)
);

OAI21x1_ASAP7_75t_L g1851 ( 
.A1(n_1646),
.A2(n_1699),
.B(n_1665),
.Y(n_1851)
);

BUFx2_ASAP7_75t_L g1852 ( 
.A(n_1589),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1645),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1582),
.Y(n_1854)
);

BUFx2_ASAP7_75t_L g1855 ( 
.A(n_1733),
.Y(n_1855)
);

BUFx3_ASAP7_75t_L g1856 ( 
.A(n_1627),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1638),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1640),
.Y(n_1858)
);

BUFx2_ASAP7_75t_L g1859 ( 
.A(n_1733),
.Y(n_1859)
);

BUFx2_ASAP7_75t_L g1860 ( 
.A(n_1699),
.Y(n_1860)
);

BUFx2_ASAP7_75t_L g1861 ( 
.A(n_1632),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1585),
.B(n_1566),
.Y(n_1862)
);

AOI22xp33_ASAP7_75t_L g1863 ( 
.A1(n_1593),
.A2(n_1630),
.B1(n_1740),
.B2(n_1723),
.Y(n_1863)
);

HB1xp67_ASAP7_75t_SL g1864 ( 
.A(n_1590),
.Y(n_1864)
);

BUFx2_ASAP7_75t_SL g1865 ( 
.A(n_1693),
.Y(n_1865)
);

OA21x2_ASAP7_75t_L g1866 ( 
.A1(n_1604),
.A2(n_1566),
.B(n_1586),
.Y(n_1866)
);

BUFx6f_ASAP7_75t_L g1867 ( 
.A(n_1619),
.Y(n_1867)
);

INVxp67_ASAP7_75t_L g1868 ( 
.A(n_1594),
.Y(n_1868)
);

OAI22xp33_ASAP7_75t_L g1869 ( 
.A1(n_1723),
.A2(n_1740),
.B1(n_1737),
.B2(n_1732),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1636),
.Y(n_1870)
);

HB1xp67_ASAP7_75t_L g1871 ( 
.A(n_1614),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1636),
.Y(n_1872)
);

INVxp67_ASAP7_75t_L g1873 ( 
.A(n_1592),
.Y(n_1873)
);

AOI21xp5_ASAP7_75t_L g1874 ( 
.A1(n_1605),
.A2(n_1735),
.B(n_1581),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1603),
.Y(n_1875)
);

OA21x2_ASAP7_75t_L g1876 ( 
.A1(n_1599),
.A2(n_1598),
.B(n_1735),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1587),
.B(n_1572),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1625),
.Y(n_1878)
);

AOI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1723),
.A2(n_1740),
.B1(n_1737),
.B2(n_1695),
.Y(n_1879)
);

CKINVDCx5p33_ASAP7_75t_R g1880 ( 
.A(n_1714),
.Y(n_1880)
);

OR2x6_ASAP7_75t_L g1881 ( 
.A(n_1692),
.B(n_1696),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1616),
.Y(n_1882)
);

AO21x1_ASAP7_75t_L g1883 ( 
.A1(n_1712),
.A2(n_1617),
.B(n_1637),
.Y(n_1883)
);

HB1xp67_ASAP7_75t_L g1884 ( 
.A(n_1623),
.Y(n_1884)
);

INVx3_ASAP7_75t_L g1885 ( 
.A(n_1606),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1611),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1623),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1697),
.B(n_1715),
.Y(n_1888)
);

INVx2_ASAP7_75t_SL g1889 ( 
.A(n_1692),
.Y(n_1889)
);

INVxp67_ASAP7_75t_SL g1890 ( 
.A(n_1709),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1695),
.Y(n_1891)
);

AOI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1745),
.A2(n_1732),
.B1(n_1727),
.B2(n_1696),
.Y(n_1892)
);

AOI22xp5_ASAP7_75t_L g1893 ( 
.A1(n_1817),
.A2(n_1727),
.B1(n_1576),
.B2(n_1705),
.Y(n_1893)
);

NAND2x1_ASAP7_75t_L g1894 ( 
.A(n_1866),
.B(n_1704),
.Y(n_1894)
);

NOR2xp33_ASAP7_75t_SL g1895 ( 
.A(n_1787),
.B(n_1711),
.Y(n_1895)
);

OA21x2_ASAP7_75t_L g1896 ( 
.A1(n_1827),
.A2(n_1730),
.B(n_1726),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1760),
.B(n_1562),
.Y(n_1897)
);

NOR2xp33_ASAP7_75t_L g1898 ( 
.A(n_1800),
.B(n_1713),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1766),
.B(n_1726),
.Y(n_1899)
);

AOI22xp5_ASAP7_75t_L g1900 ( 
.A1(n_1778),
.A2(n_1729),
.B1(n_1744),
.B2(n_1798),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1780),
.B(n_1766),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1852),
.B(n_1855),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1852),
.B(n_1859),
.Y(n_1903)
);

A2O1A1Ixp33_ASAP7_75t_L g1904 ( 
.A1(n_1826),
.A2(n_1832),
.B(n_1842),
.C(n_1816),
.Y(n_1904)
);

AND2x4_ASAP7_75t_L g1905 ( 
.A(n_1795),
.B(n_1789),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1819),
.B(n_1823),
.Y(n_1906)
);

AOI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1770),
.A2(n_1753),
.B(n_1748),
.Y(n_1907)
);

OR2x6_ASAP7_75t_L g1908 ( 
.A(n_1881),
.B(n_1865),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1750),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1853),
.B(n_1800),
.Y(n_1910)
);

A2O1A1Ixp33_ASAP7_75t_L g1911 ( 
.A1(n_1816),
.A2(n_1784),
.B(n_1791),
.C(n_1853),
.Y(n_1911)
);

OAI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1824),
.A2(n_1838),
.B(n_1754),
.Y(n_1912)
);

OA21x2_ASAP7_75t_L g1913 ( 
.A1(n_1771),
.A2(n_1785),
.B(n_1801),
.Y(n_1913)
);

AOI22xp5_ASAP7_75t_L g1914 ( 
.A1(n_1845),
.A2(n_1813),
.B1(n_1784),
.B2(n_1791),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1776),
.B(n_1741),
.Y(n_1915)
);

AND2x4_ASAP7_75t_L g1916 ( 
.A(n_1795),
.B(n_1789),
.Y(n_1916)
);

O2A1O1Ixp33_ASAP7_75t_L g1917 ( 
.A1(n_1845),
.A2(n_1781),
.B(n_1825),
.C(n_1815),
.Y(n_1917)
);

BUFx2_ASAP7_75t_L g1918 ( 
.A(n_1866),
.Y(n_1918)
);

AO22x2_ASAP7_75t_L g1919 ( 
.A1(n_1741),
.A2(n_1763),
.B1(n_1807),
.B2(n_1758),
.Y(n_1919)
);

AOI22xp5_ASAP7_75t_L g1920 ( 
.A1(n_1845),
.A2(n_1813),
.B1(n_1869),
.B2(n_1833),
.Y(n_1920)
);

AO32x2_ASAP7_75t_L g1921 ( 
.A1(n_1812),
.A2(n_1805),
.A3(n_1763),
.B1(n_1807),
.B2(n_1835),
.Y(n_1921)
);

INVx5_ASAP7_75t_SL g1922 ( 
.A(n_1867),
.Y(n_1922)
);

AOI21xp5_ASAP7_75t_L g1923 ( 
.A1(n_1770),
.A2(n_1753),
.B(n_1748),
.Y(n_1923)
);

OAI21x1_ASAP7_75t_SL g1924 ( 
.A1(n_1824),
.A2(n_1883),
.B(n_1866),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1810),
.B(n_1811),
.Y(n_1925)
);

OAI211xp5_ASAP7_75t_L g1926 ( 
.A1(n_1854),
.A2(n_1838),
.B(n_1818),
.C(n_1839),
.Y(n_1926)
);

A2O1A1Ixp33_ASAP7_75t_L g1927 ( 
.A1(n_1854),
.A2(n_1839),
.B(n_1833),
.C(n_1843),
.Y(n_1927)
);

OAI21xp5_ASAP7_75t_L g1928 ( 
.A1(n_1813),
.A2(n_1868),
.B(n_1843),
.Y(n_1928)
);

AOI211xp5_ASAP7_75t_L g1929 ( 
.A1(n_1883),
.A2(n_1835),
.B(n_1862),
.C(n_1820),
.Y(n_1929)
);

INVx3_ASAP7_75t_L g1930 ( 
.A(n_1866),
.Y(n_1930)
);

CKINVDCx5p33_ASAP7_75t_R g1931 ( 
.A(n_1764),
.Y(n_1931)
);

OR2x2_ASAP7_75t_L g1932 ( 
.A(n_1746),
.B(n_1783),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1750),
.Y(n_1933)
);

AOI221xp5_ASAP7_75t_L g1934 ( 
.A1(n_1805),
.A2(n_1828),
.B1(n_1746),
.B2(n_1743),
.C(n_1742),
.Y(n_1934)
);

OAI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1862),
.A2(n_1863),
.B1(n_1879),
.B2(n_1829),
.Y(n_1935)
);

A2O1A1Ixp33_ASAP7_75t_L g1936 ( 
.A1(n_1833),
.A2(n_1846),
.B(n_1841),
.C(n_1879),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1752),
.Y(n_1937)
);

OR2x2_ASAP7_75t_L g1938 ( 
.A(n_1783),
.B(n_1786),
.Y(n_1938)
);

OA21x2_ASAP7_75t_L g1939 ( 
.A1(n_1801),
.A2(n_1809),
.B(n_1851),
.Y(n_1939)
);

AOI221xp5_ASAP7_75t_L g1940 ( 
.A1(n_1742),
.A2(n_1743),
.B1(n_1782),
.B2(n_1834),
.C(n_1890),
.Y(n_1940)
);

BUFx12f_ASAP7_75t_L g1941 ( 
.A(n_1844),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1786),
.B(n_1765),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1752),
.Y(n_1943)
);

BUFx2_ASAP7_75t_L g1944 ( 
.A(n_1860),
.Y(n_1944)
);

AOI22xp33_ASAP7_75t_L g1945 ( 
.A1(n_1803),
.A2(n_1830),
.B1(n_1813),
.B2(n_1806),
.Y(n_1945)
);

AO32x2_ASAP7_75t_L g1946 ( 
.A1(n_1790),
.A2(n_1822),
.A3(n_1782),
.B1(n_1751),
.B2(n_1889),
.Y(n_1946)
);

AO32x2_ASAP7_75t_L g1947 ( 
.A1(n_1790),
.A2(n_1822),
.A3(n_1751),
.B1(n_1889),
.B2(n_1774),
.Y(n_1947)
);

OAI21xp5_ASAP7_75t_L g1948 ( 
.A1(n_1813),
.A2(n_1841),
.B(n_1846),
.Y(n_1948)
);

OR2x6_ASAP7_75t_L g1949 ( 
.A(n_1881),
.B(n_1865),
.Y(n_1949)
);

A2O1A1Ixp33_ASAP7_75t_L g1950 ( 
.A1(n_1814),
.A2(n_1821),
.B(n_1829),
.C(n_1803),
.Y(n_1950)
);

OR2x2_ASAP7_75t_L g1951 ( 
.A(n_1747),
.B(n_1749),
.Y(n_1951)
);

AOI22xp33_ASAP7_75t_SL g1952 ( 
.A1(n_1813),
.A2(n_1830),
.B1(n_1770),
.B2(n_1806),
.Y(n_1952)
);

INVxp67_ASAP7_75t_L g1953 ( 
.A(n_1871),
.Y(n_1953)
);

HB1xp67_ASAP7_75t_L g1954 ( 
.A(n_1860),
.Y(n_1954)
);

NAND2xp33_ASAP7_75t_L g1955 ( 
.A(n_1844),
.B(n_1880),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1769),
.B(n_1773),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1757),
.Y(n_1957)
);

INVxp67_ASAP7_75t_L g1958 ( 
.A(n_1882),
.Y(n_1958)
);

BUFx6f_ASAP7_75t_L g1959 ( 
.A(n_1762),
.Y(n_1959)
);

NOR2xp33_ASAP7_75t_L g1960 ( 
.A(n_1873),
.B(n_1877),
.Y(n_1960)
);

BUFx2_ASAP7_75t_L g1961 ( 
.A(n_1881),
.Y(n_1961)
);

OR2x6_ASAP7_75t_L g1962 ( 
.A(n_1881),
.B(n_1867),
.Y(n_1962)
);

OR2x2_ASAP7_75t_L g1963 ( 
.A(n_1747),
.B(n_1749),
.Y(n_1963)
);

AO32x2_ASAP7_75t_L g1964 ( 
.A1(n_1751),
.A2(n_1774),
.A3(n_1802),
.B1(n_1804),
.B2(n_1777),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1769),
.B(n_1773),
.Y(n_1965)
);

OR2x6_ASAP7_75t_L g1966 ( 
.A(n_1881),
.B(n_1867),
.Y(n_1966)
);

AND2x4_ASAP7_75t_L g1967 ( 
.A(n_1793),
.B(n_1794),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1847),
.Y(n_1968)
);

INVxp67_ASAP7_75t_L g1969 ( 
.A(n_1872),
.Y(n_1969)
);

O2A1O1Ixp33_ASAP7_75t_L g1970 ( 
.A1(n_1814),
.A2(n_1821),
.B(n_1891),
.C(n_1858),
.Y(n_1970)
);

OAI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1813),
.A2(n_1858),
.B(n_1770),
.Y(n_1971)
);

AOI22xp5_ASAP7_75t_L g1972 ( 
.A1(n_1891),
.A2(n_1887),
.B1(n_1884),
.B2(n_1880),
.Y(n_1972)
);

AOI221xp5_ASAP7_75t_L g1973 ( 
.A1(n_1847),
.A2(n_1850),
.B1(n_1886),
.B2(n_1870),
.C(n_1788),
.Y(n_1973)
);

AOI221xp5_ASAP7_75t_L g1974 ( 
.A1(n_1850),
.A2(n_1886),
.B1(n_1870),
.B2(n_1796),
.C(n_1837),
.Y(n_1974)
);

NOR2xp33_ASAP7_75t_L g1975 ( 
.A(n_1872),
.B(n_1887),
.Y(n_1975)
);

INVxp67_ASAP7_75t_L g1976 ( 
.A(n_1857),
.Y(n_1976)
);

HB1xp67_ASAP7_75t_L g1977 ( 
.A(n_1755),
.Y(n_1977)
);

AO32x2_ASAP7_75t_L g1978 ( 
.A1(n_1751),
.A2(n_1777),
.A3(n_1772),
.B1(n_1759),
.B2(n_1753),
.Y(n_1978)
);

OA21x2_ASAP7_75t_L g1979 ( 
.A1(n_1851),
.A2(n_1799),
.B(n_1779),
.Y(n_1979)
);

OR2x2_ASAP7_75t_L g1980 ( 
.A(n_1772),
.B(n_1775),
.Y(n_1980)
);

BUFx8_ASAP7_75t_L g1981 ( 
.A(n_1867),
.Y(n_1981)
);

OR2x6_ASAP7_75t_L g1982 ( 
.A(n_1867),
.B(n_1861),
.Y(n_1982)
);

INVx3_ASAP7_75t_L g1983 ( 
.A(n_1875),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1909),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1901),
.B(n_1751),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1894),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1933),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1942),
.B(n_1753),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1937),
.Y(n_1989)
);

NOR2x1p5_ASAP7_75t_L g1990 ( 
.A(n_1899),
.B(n_1797),
.Y(n_1990)
);

AOI22xp33_ASAP7_75t_L g1991 ( 
.A1(n_1900),
.A2(n_1856),
.B1(n_1888),
.B2(n_1797),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1943),
.Y(n_1992)
);

CKINVDCx20_ASAP7_75t_R g1993 ( 
.A(n_1931),
.Y(n_1993)
);

INVxp67_ASAP7_75t_L g1994 ( 
.A(n_1919),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1957),
.Y(n_1995)
);

NOR2xp33_ASAP7_75t_L g1996 ( 
.A(n_1960),
.B(n_1856),
.Y(n_1996)
);

AND2x4_ASAP7_75t_L g1997 ( 
.A(n_1971),
.B(n_1808),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1947),
.B(n_1946),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1946),
.B(n_1792),
.Y(n_1999)
);

OR2x2_ASAP7_75t_L g2000 ( 
.A(n_1918),
.B(n_1792),
.Y(n_2000)
);

HB1xp67_ASAP7_75t_L g2001 ( 
.A(n_1977),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1946),
.B(n_1792),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1921),
.B(n_1792),
.Y(n_2003)
);

INVxp67_ASAP7_75t_SL g2004 ( 
.A(n_1930),
.Y(n_2004)
);

AOI22xp33_ASAP7_75t_L g2005 ( 
.A1(n_1900),
.A2(n_1888),
.B1(n_1797),
.B2(n_1761),
.Y(n_2005)
);

OR2x2_ASAP7_75t_L g2006 ( 
.A(n_1915),
.B(n_1808),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1978),
.B(n_1964),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1964),
.B(n_1768),
.Y(n_2008)
);

INVx1_ASAP7_75t_SL g2009 ( 
.A(n_1944),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1921),
.B(n_1768),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1951),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1963),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1921),
.B(n_1836),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1902),
.B(n_1903),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1934),
.B(n_1849),
.Y(n_2015)
);

BUFx3_ASAP7_75t_L g2016 ( 
.A(n_1981),
.Y(n_2016)
);

INVxp67_ASAP7_75t_L g2017 ( 
.A(n_1919),
.Y(n_2017)
);

BUFx2_ASAP7_75t_L g2018 ( 
.A(n_1954),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1980),
.Y(n_2019)
);

OR2x2_ASAP7_75t_L g2020 ( 
.A(n_1938),
.B(n_1932),
.Y(n_2020)
);

NOR2x1p5_ASAP7_75t_L g2021 ( 
.A(n_1941),
.B(n_1761),
.Y(n_2021)
);

AOI22xp5_ASAP7_75t_L g2022 ( 
.A1(n_1895),
.A2(n_1885),
.B1(n_1878),
.B2(n_1864),
.Y(n_2022)
);

HB1xp67_ASAP7_75t_L g2023 ( 
.A(n_1939),
.Y(n_2023)
);

AND2x4_ASAP7_75t_L g2024 ( 
.A(n_1967),
.B(n_1796),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1925),
.B(n_1848),
.Y(n_2025)
);

OR2x2_ASAP7_75t_L g2026 ( 
.A(n_1907),
.B(n_1837),
.Y(n_2026)
);

BUFx6f_ASAP7_75t_L g2027 ( 
.A(n_1908),
.Y(n_2027)
);

NOR2xp33_ASAP7_75t_L g2028 ( 
.A(n_1897),
.B(n_1885),
.Y(n_2028)
);

HB1xp67_ASAP7_75t_L g2029 ( 
.A(n_2001),
.Y(n_2029)
);

NOR2xp33_ASAP7_75t_L g2030 ( 
.A(n_1996),
.B(n_1898),
.Y(n_2030)
);

INVx2_ASAP7_75t_SL g2031 ( 
.A(n_1990),
.Y(n_2031)
);

INVx1_ASAP7_75t_SL g2032 ( 
.A(n_2009),
.Y(n_2032)
);

NOR2xp33_ASAP7_75t_L g2033 ( 
.A(n_2028),
.B(n_1972),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_2014),
.B(n_1914),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_2014),
.B(n_1914),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1985),
.B(n_1910),
.Y(n_2036)
);

INVxp67_ASAP7_75t_L g2037 ( 
.A(n_2018),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1984),
.Y(n_2038)
);

AND2x4_ASAP7_75t_L g2039 ( 
.A(n_1997),
.B(n_1908),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1987),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1987),
.Y(n_2041)
);

INVxp67_ASAP7_75t_L g2042 ( 
.A(n_2018),
.Y(n_2042)
);

INVxp67_ASAP7_75t_L g2043 ( 
.A(n_2025),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_2011),
.B(n_2012),
.Y(n_2044)
);

INVxp67_ASAP7_75t_SL g2045 ( 
.A(n_2001),
.Y(n_2045)
);

OAI211xp5_ASAP7_75t_SL g2046 ( 
.A1(n_1994),
.A2(n_1911),
.B(n_1929),
.C(n_1904),
.Y(n_2046)
);

HB1xp67_ASAP7_75t_L g2047 ( 
.A(n_2000),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1985),
.B(n_1896),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1989),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1999),
.B(n_1896),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1989),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_2002),
.B(n_1905),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_2002),
.B(n_1916),
.Y(n_2053)
);

BUFx2_ASAP7_75t_L g2054 ( 
.A(n_1986),
.Y(n_2054)
);

NAND2x1_ASAP7_75t_L g2055 ( 
.A(n_1986),
.B(n_1924),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1992),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1992),
.Y(n_2057)
);

OAI21xp5_ASAP7_75t_L g2058 ( 
.A1(n_2022),
.A2(n_1893),
.B(n_1917),
.Y(n_2058)
);

AND4x1_ASAP7_75t_L g2059 ( 
.A(n_2005),
.B(n_1895),
.C(n_1893),
.D(n_1929),
.Y(n_2059)
);

NOR2xp33_ASAP7_75t_L g2060 ( 
.A(n_2016),
.B(n_1972),
.Y(n_2060)
);

NOR3xp33_ASAP7_75t_L g2061 ( 
.A(n_2022),
.B(n_1935),
.C(n_1926),
.Y(n_2061)
);

AND2x4_ASAP7_75t_SL g2062 ( 
.A(n_2027),
.B(n_1949),
.Y(n_2062)
);

OAI22xp33_ASAP7_75t_L g2063 ( 
.A1(n_2027),
.A2(n_1920),
.B1(n_1962),
.B2(n_1966),
.Y(n_2063)
);

INVx3_ASAP7_75t_L g2064 ( 
.A(n_1995),
.Y(n_2064)
);

INVx2_ASAP7_75t_SL g2065 ( 
.A(n_1990),
.Y(n_2065)
);

OAI33xp33_ASAP7_75t_L g2066 ( 
.A1(n_1994),
.A2(n_1906),
.A3(n_1953),
.B1(n_1958),
.B2(n_1969),
.B3(n_1970),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_2011),
.B(n_1912),
.Y(n_2067)
);

OR2x2_ASAP7_75t_L g2068 ( 
.A(n_1988),
.B(n_1923),
.Y(n_2068)
);

BUFx4f_ASAP7_75t_L g2069 ( 
.A(n_1986),
.Y(n_2069)
);

OAI22xp5_ASAP7_75t_L g2070 ( 
.A1(n_1991),
.A2(n_1920),
.B1(n_1945),
.B2(n_1892),
.Y(n_2070)
);

BUFx2_ASAP7_75t_L g2071 ( 
.A(n_1986),
.Y(n_2071)
);

AO21x2_ASAP7_75t_L g2072 ( 
.A1(n_2023),
.A2(n_1928),
.B(n_1948),
.Y(n_2072)
);

OAI211xp5_ASAP7_75t_L g2073 ( 
.A1(n_2017),
.A2(n_1940),
.B(n_1927),
.C(n_1892),
.Y(n_2073)
);

AO221x1_ASAP7_75t_L g2074 ( 
.A1(n_2017),
.A2(n_1961),
.B1(n_1959),
.B2(n_1983),
.C(n_1976),
.Y(n_2074)
);

OR2x2_ASAP7_75t_L g2075 ( 
.A(n_1988),
.B(n_1913),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_2003),
.B(n_1979),
.Y(n_2076)
);

AO21x2_ASAP7_75t_L g2077 ( 
.A1(n_2023),
.A2(n_1950),
.B(n_1956),
.Y(n_2077)
);

BUFx2_ASAP7_75t_L g2078 ( 
.A(n_1986),
.Y(n_2078)
);

OAI31xp33_ASAP7_75t_L g2079 ( 
.A1(n_2005),
.A2(n_1936),
.A3(n_1975),
.B(n_1756),
.Y(n_2079)
);

OAI211xp5_ASAP7_75t_L g2080 ( 
.A1(n_1991),
.A2(n_1952),
.B(n_1973),
.C(n_1974),
.Y(n_2080)
);

BUFx2_ASAP7_75t_L g2081 ( 
.A(n_1986),
.Y(n_2081)
);

AO21x2_ASAP7_75t_L g2082 ( 
.A1(n_2004),
.A2(n_1965),
.B(n_1968),
.Y(n_2082)
);

AOI22xp33_ASAP7_75t_L g2083 ( 
.A1(n_1997),
.A2(n_1962),
.B1(n_1966),
.B2(n_1982),
.Y(n_2083)
);

BUFx6f_ASAP7_75t_L g2084 ( 
.A(n_2016),
.Y(n_2084)
);

HB1xp67_ASAP7_75t_L g2085 ( 
.A(n_2000),
.Y(n_2085)
);

BUFx3_ASAP7_75t_L g2086 ( 
.A(n_2016),
.Y(n_2086)
);

INVx4_ASAP7_75t_L g2087 ( 
.A(n_2084),
.Y(n_2087)
);

NOR2xp33_ASAP7_75t_L g2088 ( 
.A(n_2033),
.B(n_1955),
.Y(n_2088)
);

AND2x2_ASAP7_75t_L g2089 ( 
.A(n_2034),
.B(n_2010),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2038),
.Y(n_2090)
);

OR2x2_ASAP7_75t_L g2091 ( 
.A(n_2068),
.B(n_2020),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2034),
.B(n_2013),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2038),
.Y(n_2093)
);

OR2x2_ASAP7_75t_L g2094 ( 
.A(n_2068),
.B(n_2020),
.Y(n_2094)
);

BUFx2_ASAP7_75t_L g2095 ( 
.A(n_2054),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_2035),
.B(n_2013),
.Y(n_2096)
);

INVxp33_ASAP7_75t_SL g2097 ( 
.A(n_2060),
.Y(n_2097)
);

AND2x4_ASAP7_75t_L g2098 ( 
.A(n_2031),
.B(n_1997),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2040),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_2035),
.B(n_1998),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_2082),
.Y(n_2101)
);

NOR2x1_ASAP7_75t_SL g2102 ( 
.A(n_2077),
.B(n_1998),
.Y(n_2102)
);

HB1xp67_ASAP7_75t_L g2103 ( 
.A(n_2029),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2067),
.B(n_2009),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2040),
.Y(n_2105)
);

INVx2_ASAP7_75t_SL g2106 ( 
.A(n_2086),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2031),
.B(n_2008),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_2032),
.B(n_2025),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_2082),
.Y(n_2109)
);

INVx1_ASAP7_75t_SL g2110 ( 
.A(n_2086),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2041),
.Y(n_2111)
);

OR2x2_ASAP7_75t_L g2112 ( 
.A(n_2047),
.B(n_2026),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2041),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_2082),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_2037),
.B(n_2012),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2042),
.B(n_2019),
.Y(n_2116)
);

AND2x4_ASAP7_75t_L g2117 ( 
.A(n_2065),
.B(n_2027),
.Y(n_2117)
);

INVxp67_ASAP7_75t_L g2118 ( 
.A(n_2044),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_2065),
.B(n_2008),
.Y(n_2119)
);

OAI22xp5_ASAP7_75t_L g2120 ( 
.A1(n_2061),
.A2(n_1982),
.B1(n_1922),
.B2(n_2027),
.Y(n_2120)
);

OR2x2_ASAP7_75t_L g2121 ( 
.A(n_2085),
.B(n_2026),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2049),
.Y(n_2122)
);

INVx4_ASAP7_75t_L g2123 ( 
.A(n_2084),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_2036),
.B(n_2019),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2049),
.Y(n_2125)
);

AND2x4_ASAP7_75t_L g2126 ( 
.A(n_2039),
.B(n_2027),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2051),
.Y(n_2127)
);

HB1xp67_ASAP7_75t_L g2128 ( 
.A(n_2077),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2052),
.B(n_2053),
.Y(n_2129)
);

INVx3_ASAP7_75t_L g2130 ( 
.A(n_2064),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_2036),
.B(n_2024),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_2064),
.Y(n_2132)
);

HB1xp67_ASAP7_75t_L g2133 ( 
.A(n_2077),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2056),
.Y(n_2134)
);

OR2x2_ASAP7_75t_L g2135 ( 
.A(n_2075),
.B(n_2045),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2043),
.B(n_2024),
.Y(n_2136)
);

OAI22xp5_ASAP7_75t_L g2137 ( 
.A1(n_2058),
.A2(n_1922),
.B1(n_2027),
.B2(n_2015),
.Y(n_2137)
);

OR2x2_ASAP7_75t_L g2138 ( 
.A(n_2075),
.B(n_2006),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2056),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2057),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2090),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2115),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_2126),
.B(n_2048),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2090),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2126),
.B(n_2048),
.Y(n_2145)
);

OR2x2_ASAP7_75t_L g2146 ( 
.A(n_2091),
.B(n_2094),
.Y(n_2146)
);

AOI21xp5_ASAP7_75t_L g2147 ( 
.A1(n_2097),
.A2(n_2046),
.B(n_2079),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2093),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_2132),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2132),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_2118),
.B(n_2073),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_2126),
.B(n_2050),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2116),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_2104),
.B(n_2050),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2093),
.Y(n_2155)
);

OR2x6_ASAP7_75t_L g2156 ( 
.A(n_2087),
.B(n_2084),
.Y(n_2156)
);

HB1xp67_ASAP7_75t_L g2157 ( 
.A(n_2103),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2099),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2099),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2089),
.B(n_2054),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_2089),
.B(n_2071),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2105),
.Y(n_2162)
);

NOR2x1_ASAP7_75t_L g2163 ( 
.A(n_2087),
.B(n_2086),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2092),
.B(n_2071),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_2101),
.Y(n_2165)
);

NOR2xp67_ASAP7_75t_R g2166 ( 
.A(n_2087),
.B(n_2123),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2105),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_2092),
.B(n_2078),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_2097),
.B(n_2084),
.Y(n_2169)
);

OR2x2_ASAP7_75t_L g2170 ( 
.A(n_2091),
.B(n_2072),
.Y(n_2170)
);

OR2x2_ASAP7_75t_L g2171 ( 
.A(n_2094),
.B(n_2072),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2101),
.Y(n_2172)
);

OR2x2_ASAP7_75t_L g2173 ( 
.A(n_2135),
.B(n_2138),
.Y(n_2173)
);

NAND2x1_ASAP7_75t_SL g2174 ( 
.A(n_2128),
.B(n_2007),
.Y(n_2174)
);

OR2x2_ASAP7_75t_L g2175 ( 
.A(n_2135),
.B(n_2072),
.Y(n_2175)
);

NAND2x1_ASAP7_75t_L g2176 ( 
.A(n_2095),
.B(n_2074),
.Y(n_2176)
);

HB1xp67_ASAP7_75t_L g2177 ( 
.A(n_2095),
.Y(n_2177)
);

INVx3_ASAP7_75t_L g2178 ( 
.A(n_2123),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_2096),
.B(n_2078),
.Y(n_2179)
);

NOR2xp33_ASAP7_75t_L g2180 ( 
.A(n_2088),
.B(n_1993),
.Y(n_2180)
);

AND2x4_ASAP7_75t_L g2181 ( 
.A(n_2123),
.B(n_2039),
.Y(n_2181)
);

AND2x4_ASAP7_75t_L g2182 ( 
.A(n_2117),
.B(n_2039),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2111),
.Y(n_2183)
);

OR2x2_ASAP7_75t_L g2184 ( 
.A(n_2138),
.B(n_2076),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2110),
.B(n_2084),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2096),
.B(n_2081),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2111),
.Y(n_2187)
);

NOR2xp33_ASAP7_75t_L g2188 ( 
.A(n_2137),
.B(n_1756),
.Y(n_2188)
);

NAND5xp2_ASAP7_75t_L g2189 ( 
.A(n_2107),
.B(n_2079),
.C(n_2080),
.D(n_2083),
.E(n_2030),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_2109),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_2106),
.B(n_2076),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2113),
.Y(n_2192)
);

INVx3_ASAP7_75t_L g2193 ( 
.A(n_2130),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2113),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2122),
.Y(n_2195)
);

AND2x2_ASAP7_75t_L g2196 ( 
.A(n_2100),
.B(n_2081),
.Y(n_2196)
);

AOI22xp5_ASAP7_75t_L g2197 ( 
.A1(n_2147),
.A2(n_2070),
.B1(n_2120),
.B2(n_2066),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_2196),
.B(n_2102),
.Y(n_2198)
);

NAND4xp75_ASAP7_75t_L g2199 ( 
.A(n_2163),
.B(n_2106),
.C(n_2059),
.D(n_2007),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_2196),
.Y(n_2200)
);

OR2x2_ASAP7_75t_L g2201 ( 
.A(n_2146),
.B(n_2112),
.Y(n_2201)
);

INVx1_ASAP7_75t_SL g2202 ( 
.A(n_2169),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_2160),
.B(n_2102),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2141),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2141),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_2160),
.B(n_2100),
.Y(n_2206)
);

OR2x2_ASAP7_75t_L g2207 ( 
.A(n_2146),
.B(n_2112),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_2161),
.B(n_2117),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2144),
.Y(n_2209)
);

INVx2_ASAP7_75t_SL g2210 ( 
.A(n_2156),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2144),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2161),
.Y(n_2212)
);

OR2x2_ASAP7_75t_L g2213 ( 
.A(n_2173),
.B(n_2121),
.Y(n_2213)
);

INVxp67_ASAP7_75t_L g2214 ( 
.A(n_2157),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2164),
.B(n_2117),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_2151),
.B(n_2129),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_L g2217 ( 
.A(n_2188),
.B(n_1764),
.Y(n_2217)
);

AOI21xp5_ASAP7_75t_L g2218 ( 
.A1(n_2189),
.A2(n_2133),
.B(n_2055),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_2142),
.B(n_2129),
.Y(n_2219)
);

INVx1_ASAP7_75t_SL g2220 ( 
.A(n_2182),
.Y(n_2220)
);

INVx2_ASAP7_75t_SL g2221 ( 
.A(n_2156),
.Y(n_2221)
);

INVx2_ASAP7_75t_SL g2222 ( 
.A(n_2156),
.Y(n_2222)
);

OR2x2_ASAP7_75t_L g2223 ( 
.A(n_2173),
.B(n_2121),
.Y(n_2223)
);

INVxp67_ASAP7_75t_L g2224 ( 
.A(n_2177),
.Y(n_2224)
);

OR2x2_ASAP7_75t_L g2225 ( 
.A(n_2153),
.B(n_2124),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2143),
.B(n_2131),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_2164),
.B(n_2098),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_2168),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_2168),
.Y(n_2229)
);

OAI31xp33_ASAP7_75t_L g2230 ( 
.A1(n_2175),
.A2(n_2063),
.A3(n_2059),
.B(n_2021),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_2143),
.B(n_2107),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_2179),
.B(n_2098),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2148),
.Y(n_2233)
);

BUFx2_ASAP7_75t_L g2234 ( 
.A(n_2156),
.Y(n_2234)
);

AND2x2_ASAP7_75t_L g2235 ( 
.A(n_2179),
.B(n_2098),
.Y(n_2235)
);

OR2x2_ASAP7_75t_L g2236 ( 
.A(n_2184),
.B(n_2122),
.Y(n_2236)
);

O2A1O1Ixp33_ASAP7_75t_L g2237 ( 
.A1(n_2176),
.A2(n_2055),
.B(n_2109),
.C(n_2114),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2148),
.Y(n_2238)
);

OR2x2_ASAP7_75t_L g2239 ( 
.A(n_2216),
.B(n_2214),
.Y(n_2239)
);

AOI211xp5_ASAP7_75t_L g2240 ( 
.A1(n_2230),
.A2(n_2175),
.B(n_2171),
.C(n_2170),
.Y(n_2240)
);

AND2x2_ASAP7_75t_SL g2241 ( 
.A(n_2197),
.B(n_2180),
.Y(n_2241)
);

OAI21xp5_ASAP7_75t_L g2242 ( 
.A1(n_2199),
.A2(n_2176),
.B(n_2174),
.Y(n_2242)
);

NAND3xp33_ASAP7_75t_L g2243 ( 
.A(n_2230),
.B(n_2178),
.C(n_2185),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2208),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2204),
.Y(n_2245)
);

NOR4xp25_ASAP7_75t_SL g2246 ( 
.A(n_2234),
.B(n_2166),
.C(n_2194),
.D(n_2162),
.Y(n_2246)
);

NOR2x1_ASAP7_75t_L g2247 ( 
.A(n_2199),
.B(n_2178),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2204),
.Y(n_2248)
);

NOR2xp33_ASAP7_75t_L g2249 ( 
.A(n_2217),
.B(n_2182),
.Y(n_2249)
);

O2A1O1Ixp33_ASAP7_75t_L g2250 ( 
.A1(n_2218),
.A2(n_2178),
.B(n_2171),
.C(n_2170),
.Y(n_2250)
);

AND2x4_ASAP7_75t_L g2251 ( 
.A(n_2208),
.B(n_2182),
.Y(n_2251)
);

AOI21xp33_ASAP7_75t_L g2252 ( 
.A1(n_2197),
.A2(n_2114),
.B(n_2155),
.Y(n_2252)
);

AOI22xp5_ASAP7_75t_L g2253 ( 
.A1(n_2220),
.A2(n_2181),
.B1(n_2152),
.B2(n_2145),
.Y(n_2253)
);

INVxp33_ASAP7_75t_L g2254 ( 
.A(n_2215),
.Y(n_2254)
);

NOR2x1_ASAP7_75t_L g2255 ( 
.A(n_2234),
.B(n_2021),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2205),
.Y(n_2256)
);

NOR2xp33_ASAP7_75t_L g2257 ( 
.A(n_2202),
.B(n_2181),
.Y(n_2257)
);

HB1xp67_ASAP7_75t_L g2258 ( 
.A(n_2200),
.Y(n_2258)
);

OAI22xp33_ASAP7_75t_SL g2259 ( 
.A1(n_2210),
.A2(n_2181),
.B1(n_2191),
.B2(n_2184),
.Y(n_2259)
);

AOI22xp5_ASAP7_75t_L g2260 ( 
.A1(n_2215),
.A2(n_2152),
.B1(n_2145),
.B2(n_2186),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2205),
.Y(n_2261)
);

OAI221xp5_ASAP7_75t_L g2262 ( 
.A1(n_2224),
.A2(n_2174),
.B1(n_2154),
.B2(n_2069),
.C(n_2186),
.Y(n_2262)
);

OAI211xp5_ASAP7_75t_L g2263 ( 
.A1(n_2237),
.A2(n_2195),
.B(n_2194),
.C(n_2155),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2209),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2209),
.Y(n_2265)
);

AOI21xp33_ASAP7_75t_L g2266 ( 
.A1(n_2210),
.A2(n_2159),
.B(n_2158),
.Y(n_2266)
);

OR2x2_ASAP7_75t_L g2267 ( 
.A(n_2213),
.B(n_2136),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2211),
.Y(n_2268)
);

XNOR2xp5_ASAP7_75t_L g2269 ( 
.A(n_2227),
.B(n_2062),
.Y(n_2269)
);

INVx3_ASAP7_75t_L g2270 ( 
.A(n_2251),
.Y(n_2270)
);

AOI21xp33_ASAP7_75t_SL g2271 ( 
.A1(n_2241),
.A2(n_2222),
.B(n_2221),
.Y(n_2271)
);

OAI21xp33_ASAP7_75t_SL g2272 ( 
.A1(n_2242),
.A2(n_2222),
.B(n_2221),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_2244),
.B(n_2200),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2257),
.B(n_2212),
.Y(n_2274)
);

NAND3xp33_ASAP7_75t_SL g2275 ( 
.A(n_2246),
.B(n_2203),
.C(n_2198),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2251),
.Y(n_2276)
);

OAI211xp5_ASAP7_75t_SL g2277 ( 
.A1(n_2252),
.A2(n_2240),
.B(n_2250),
.C(n_2242),
.Y(n_2277)
);

AOI21xp33_ASAP7_75t_L g2278 ( 
.A1(n_2255),
.A2(n_2223),
.B(n_2213),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2258),
.Y(n_2279)
);

OAI21xp5_ASAP7_75t_L g2280 ( 
.A1(n_2247),
.A2(n_2203),
.B(n_2198),
.Y(n_2280)
);

AOI21xp5_ASAP7_75t_L g2281 ( 
.A1(n_2252),
.A2(n_2228),
.B(n_2212),
.Y(n_2281)
);

AOI211x1_ASAP7_75t_L g2282 ( 
.A1(n_2262),
.A2(n_2227),
.B(n_2235),
.C(n_2232),
.Y(n_2282)
);

NOR2x1_ASAP7_75t_L g2283 ( 
.A(n_2243),
.B(n_2211),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2254),
.B(n_2228),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_2249),
.B(n_2232),
.Y(n_2285)
);

NAND3xp33_ASAP7_75t_L g2286 ( 
.A(n_2239),
.B(n_2229),
.C(n_2233),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_2253),
.B(n_2229),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_2267),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2245),
.Y(n_2289)
);

O2A1O1Ixp33_ASAP7_75t_L g2290 ( 
.A1(n_2259),
.A2(n_2238),
.B(n_2233),
.C(n_2219),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2248),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2256),
.Y(n_2292)
);

HB1xp67_ASAP7_75t_L g2293 ( 
.A(n_2270),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2279),
.Y(n_2294)
);

AOI21xp5_ASAP7_75t_L g2295 ( 
.A1(n_2277),
.A2(n_2266),
.B(n_2262),
.Y(n_2295)
);

NAND3xp33_ASAP7_75t_L g2296 ( 
.A(n_2283),
.B(n_2266),
.C(n_2264),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2276),
.B(n_2206),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2276),
.B(n_2206),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2288),
.Y(n_2299)
);

INVxp67_ASAP7_75t_SL g2300 ( 
.A(n_2270),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2292),
.Y(n_2301)
);

AOI22xp33_ASAP7_75t_L g2302 ( 
.A1(n_2278),
.A2(n_2268),
.B1(n_2265),
.B2(n_2261),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2270),
.B(n_2260),
.Y(n_2303)
);

INVxp67_ASAP7_75t_SL g2304 ( 
.A(n_2280),
.Y(n_2304)
);

OAI221xp5_ASAP7_75t_SL g2305 ( 
.A1(n_2272),
.A2(n_2263),
.B1(n_2269),
.B2(n_2223),
.C(n_2201),
.Y(n_2305)
);

OAI321xp33_ASAP7_75t_L g2306 ( 
.A1(n_2275),
.A2(n_2201),
.A3(n_2207),
.B1(n_2231),
.B2(n_2238),
.C(n_2235),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2271),
.B(n_2226),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2300),
.B(n_2285),
.Y(n_2308)
);

AND2x2_ASAP7_75t_L g2309 ( 
.A(n_2293),
.B(n_2285),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2299),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2304),
.B(n_2288),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2299),
.Y(n_2312)
);

NOR3xp33_ASAP7_75t_L g2313 ( 
.A(n_2305),
.B(n_2306),
.C(n_2295),
.Y(n_2313)
);

AOI21xp5_ASAP7_75t_L g2314 ( 
.A1(n_2296),
.A2(n_2290),
.B(n_2281),
.Y(n_2314)
);

OR2x2_ASAP7_75t_L g2315 ( 
.A(n_2297),
.B(n_2298),
.Y(n_2315)
);

AND2x4_ASAP7_75t_L g2316 ( 
.A(n_2294),
.B(n_2286),
.Y(n_2316)
);

NAND2x1_ASAP7_75t_L g2317 ( 
.A(n_2301),
.B(n_2282),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2303),
.Y(n_2318)
);

AOI221xp5_ASAP7_75t_L g2319 ( 
.A1(n_2302),
.A2(n_2287),
.B1(n_2274),
.B2(n_2284),
.C(n_2273),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_2307),
.B(n_2289),
.Y(n_2320)
);

OA22x2_ASAP7_75t_L g2321 ( 
.A1(n_2317),
.A2(n_2291),
.B1(n_2292),
.B2(n_2302),
.Y(n_2321)
);

NAND3xp33_ASAP7_75t_SL g2322 ( 
.A(n_2313),
.B(n_2207),
.C(n_2225),
.Y(n_2322)
);

NAND3xp33_ASAP7_75t_SL g2323 ( 
.A(n_2314),
.B(n_2225),
.C(n_2236),
.Y(n_2323)
);

NOR2x1_ASAP7_75t_L g2324 ( 
.A(n_2311),
.B(n_1885),
.Y(n_2324)
);

AOI211xp5_ASAP7_75t_L g2325 ( 
.A1(n_2319),
.A2(n_2236),
.B(n_2165),
.C(n_2172),
.Y(n_2325)
);

OAI211xp5_ASAP7_75t_L g2326 ( 
.A1(n_2308),
.A2(n_1885),
.B(n_2165),
.C(n_2172),
.Y(n_2326)
);

AOI221xp5_ASAP7_75t_L g2327 ( 
.A1(n_2316),
.A2(n_2190),
.B1(n_2159),
.B2(n_2158),
.C(n_2195),
.Y(n_2327)
);

A2O1A1Ixp33_ASAP7_75t_L g2328 ( 
.A1(n_2316),
.A2(n_2069),
.B(n_2193),
.C(n_2167),
.Y(n_2328)
);

AOI21xp5_ASAP7_75t_L g2329 ( 
.A1(n_2321),
.A2(n_2323),
.B(n_2322),
.Y(n_2329)
);

NAND3xp33_ASAP7_75t_SL g2330 ( 
.A(n_2328),
.B(n_2309),
.C(n_2318),
.Y(n_2330)
);

NAND4xp25_ASAP7_75t_L g2331 ( 
.A(n_2324),
.B(n_2315),
.C(n_2320),
.D(n_2312),
.Y(n_2331)
);

CKINVDCx16_ASAP7_75t_R g2332 ( 
.A(n_2326),
.Y(n_2332)
);

NAND3xp33_ASAP7_75t_SL g2333 ( 
.A(n_2325),
.B(n_2310),
.C(n_1981),
.Y(n_2333)
);

AOI21xp5_ASAP7_75t_L g2334 ( 
.A1(n_2327),
.A2(n_2190),
.B(n_2167),
.Y(n_2334)
);

AOI221xp5_ASAP7_75t_L g2335 ( 
.A1(n_2323),
.A2(n_2183),
.B1(n_2162),
.B2(n_2187),
.C(n_2192),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2321),
.Y(n_2336)
);

AOI221xp5_ASAP7_75t_L g2337 ( 
.A1(n_2323),
.A2(n_2183),
.B1(n_2193),
.B2(n_2150),
.C(n_2149),
.Y(n_2337)
);

AOI22xp33_ASAP7_75t_SL g2338 ( 
.A1(n_2336),
.A2(n_2069),
.B1(n_2193),
.B2(n_2074),
.Y(n_2338)
);

NOR2x1p5_ASAP7_75t_L g2339 ( 
.A(n_2330),
.B(n_1840),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2329),
.B(n_2150),
.Y(n_2340)
);

NAND4xp75_ASAP7_75t_L g2341 ( 
.A(n_2334),
.B(n_1874),
.C(n_2119),
.D(n_2149),
.Y(n_2341)
);

AND2x4_ASAP7_75t_L g2342 ( 
.A(n_2331),
.B(n_2119),
.Y(n_2342)
);

OR2x2_ASAP7_75t_L g2343 ( 
.A(n_2332),
.B(n_2108),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2342),
.Y(n_2344)
);

AO22x2_ASAP7_75t_L g2345 ( 
.A1(n_2340),
.A2(n_2333),
.B1(n_2335),
.B2(n_2337),
.Y(n_2345)
);

NAND3xp33_ASAP7_75t_L g2346 ( 
.A(n_2343),
.B(n_1762),
.C(n_1767),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2339),
.B(n_2125),
.Y(n_2347)
);

OAI22xp5_ASAP7_75t_L g2348 ( 
.A1(n_2344),
.A2(n_2338),
.B1(n_2341),
.B2(n_2130),
.Y(n_2348)
);

AOI22xp5_ASAP7_75t_L g2349 ( 
.A1(n_2348),
.A2(n_2345),
.B1(n_2346),
.B2(n_2347),
.Y(n_2349)
);

AOI22x1_ASAP7_75t_L g2350 ( 
.A1(n_2349),
.A2(n_1762),
.B1(n_1767),
.B2(n_1831),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_2349),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2351),
.Y(n_2352)
);

XNOR2x1_ASAP7_75t_L g2353 ( 
.A(n_2350),
.B(n_1840),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2352),
.B(n_2353),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2352),
.Y(n_2355)
);

OAI21x1_ASAP7_75t_SL g2356 ( 
.A1(n_2354),
.A2(n_1876),
.B(n_2015),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_SL g2357 ( 
.A(n_2356),
.B(n_2355),
.Y(n_2357)
);

AOI22xp5_ASAP7_75t_L g2358 ( 
.A1(n_2357),
.A2(n_2130),
.B1(n_2140),
.B2(n_2139),
.Y(n_2358)
);

AOI221xp5_ASAP7_75t_L g2359 ( 
.A1(n_2358),
.A2(n_2127),
.B1(n_2140),
.B2(n_2139),
.C(n_2134),
.Y(n_2359)
);

AOI211xp5_ASAP7_75t_L g2360 ( 
.A1(n_2359),
.A2(n_1762),
.B(n_1767),
.C(n_1831),
.Y(n_2360)
);


endmodule