module fake_jpeg_17332_n_227 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_37),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_22),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_24),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_45),
.B(n_42),
.Y(n_75)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_53),
.Y(n_62)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx4f_ASAP7_75t_SL g52 ( 
.A(n_35),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_52),
.Y(n_63)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_54),
.Y(n_82)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_19),
.B1(n_33),
.B2(n_18),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_34),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_64),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_34),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_61),
.A2(n_74),
.B(n_36),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_34),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_41),
.B(n_42),
.C(n_38),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_65),
.A2(n_80),
.B1(n_18),
.B2(n_23),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_56),
.A2(n_27),
.B1(n_32),
.B2(n_20),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_34),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_72),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_57),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_37),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_86),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_36),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_75),
.B(n_83),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_81),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_38),
.B1(n_30),
.B2(n_17),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_79),
.A2(n_26),
.B1(n_30),
.B2(n_17),
.Y(n_112)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_25),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_54),
.A2(n_25),
.B(n_20),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_31),
.C(n_23),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_43),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_87),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_36),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_92),
.B(n_1),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_97),
.Y(n_114)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_75),
.B(n_60),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_98),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_49),
.B1(n_46),
.B2(n_53),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_102),
.B1(n_74),
.B2(n_67),
.Y(n_116)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_105),
.Y(n_120)
);

O2A1O1Ixp33_ASAP7_75t_SL g102 ( 
.A1(n_64),
.A2(n_54),
.B(n_52),
.C(n_36),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_71),
.B(n_24),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_104),
.Y(n_123)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_112),
.B1(n_26),
.B2(n_28),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_28),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_107),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_111),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_61),
.A2(n_43),
.B(n_47),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_73),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_119),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_121),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_116),
.A2(n_118),
.B1(n_126),
.B2(n_105),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_74),
.B1(n_61),
.B2(n_80),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_69),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_62),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_89),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_125),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_89),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_90),
.A2(n_86),
.B1(n_76),
.B2(n_59),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_127),
.A2(n_30),
.B1(n_17),
.B2(n_21),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_101),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_134),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_65),
.Y(n_130)
);

AOI221xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_93),
.B1(n_98),
.B2(n_104),
.C(n_112),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_84),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_91),
.C(n_108),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_92),
.B1(n_91),
.B2(n_108),
.Y(n_144)
);

NAND2xp33_ASAP7_75t_SL g133 ( 
.A(n_102),
.B(n_77),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_133),
.A2(n_103),
.B(n_101),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_103),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_63),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_135),
.Y(n_139)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_140),
.Y(n_163)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_136),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_142),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_133),
.A2(n_111),
.B(n_95),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_143),
.A2(n_144),
.B(n_149),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_148),
.C(n_131),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_99),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_151),
.B1(n_123),
.B2(n_132),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_117),
.A2(n_93),
.B1(n_97),
.B2(n_63),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_157),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_114),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_158),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_116),
.A2(n_68),
.B1(n_85),
.B2(n_100),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_142),
.B1(n_134),
.B2(n_122),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_115),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_124),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_160),
.C(n_164),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_161),
.B(n_149),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_156),
.B(n_128),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_162),
.B(n_166),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_113),
.C(n_118),
.Y(n_164)
);

NAND3xp33_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_152),
.C(n_153),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_143),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_125),
.Y(n_170)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_170),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_139),
.B(n_132),
.Y(n_171)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_171),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_130),
.C(n_77),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_174),
.C(n_151),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_87),
.C(n_78),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_13),
.Y(n_176)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_179),
.A2(n_182),
.B1(n_161),
.B2(n_172),
.Y(n_195)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_163),
.Y(n_181)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_187),
.C(n_189),
.Y(n_193)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_175),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_186),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_144),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_188),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_155),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_140),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_138),
.Y(n_191)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

A2O1A1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_167),
.B(n_141),
.C(n_168),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_199),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_31),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_164),
.C(n_167),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_31),
.C(n_4),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_181),
.A2(n_174),
.B(n_2),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_183),
.A2(n_1),
.B(n_2),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_200),
.A2(n_201),
.B1(n_185),
.B2(n_3),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_177),
.A2(n_12),
.B1(n_21),
.B2(n_16),
.Y(n_201)
);

AO22x1_ASAP7_75t_L g202 ( 
.A1(n_192),
.A2(n_184),
.B1(n_189),
.B2(n_180),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_203),
.B(n_205),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_194),
.A2(n_178),
.B1(n_187),
.B2(n_21),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_207),
.C(n_208),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_31),
.C(n_12),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_2),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_210),
.Y(n_211)
);

OAI211xp5_ASAP7_75t_L g215 ( 
.A1(n_209),
.A2(n_196),
.B(n_200),
.C(n_199),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_215),
.A2(n_4),
.B(n_5),
.Y(n_219)
);

NAND4xp25_ASAP7_75t_SL g216 ( 
.A(n_204),
.B(n_191),
.C(n_31),
.D(n_6),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_4),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_213),
.A2(n_206),
.B1(n_202),
.B2(n_207),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_220),
.Y(n_221)
);

OAI321xp33_ASAP7_75t_L g218 ( 
.A1(n_214),
.A2(n_208),
.A3(n_205),
.B1(n_197),
.B2(n_193),
.C(n_10),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_SL g222 ( 
.A1(n_218),
.A2(n_211),
.B(n_7),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_219),
.A2(n_5),
.B(n_9),
.Y(n_223)
);

AOI322xp5_ASAP7_75t_L g225 ( 
.A1(n_222),
.A2(n_223),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_203),
.C2(n_127),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_212),
.C(n_214),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_225),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_9),
.Y(n_227)
);


endmodule