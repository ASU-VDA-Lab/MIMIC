module fake_jpeg_21203_n_273 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_273);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_100;
wire n_258;
wire n_96;

BUFx16f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_19),
.Y(n_28)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_12),
.B(n_10),
.Y(n_29)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_32),
.A2(n_33),
.B1(n_14),
.B2(n_11),
.Y(n_35)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_33),
.A2(n_14),
.B1(n_20),
.B2(n_19),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_28),
.B1(n_26),
.B2(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_49),
.Y(n_63)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_33),
.B1(n_26),
.B2(n_14),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_46),
.A2(n_47),
.B1(n_51),
.B2(n_56),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_28),
.B1(n_31),
.B2(n_16),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_16),
.B1(n_14),
.B2(n_31),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_29),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_55),
.B(n_60),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_31),
.B1(n_16),
.B2(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_29),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_17),
.Y(n_79)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_61),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_11),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_69),
.Y(n_84)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_68),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_59),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_36),
.B(n_1),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_48),
.A2(n_21),
.B1(n_18),
.B2(n_20),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_79),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_11),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_36),
.Y(n_93)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_48),
.B1(n_44),
.B2(n_47),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_83),
.A2(n_92),
.B1(n_40),
.B2(n_36),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_63),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_56),
.B1(n_51),
.B2(n_40),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_90),
.A2(n_69),
.B1(n_78),
.B2(n_75),
.Y(n_104)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_40),
.B1(n_60),
.B2(n_53),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_55),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_95),
.Y(n_120)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_96),
.Y(n_106)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_42),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_98),
.B(n_32),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_116),
.B1(n_90),
.B2(n_96),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_98),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_105),
.B(n_109),
.Y(n_128)
);

OAI32xp33_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_79),
.A3(n_73),
.B1(n_75),
.B2(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_113),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_84),
.B(n_64),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_112),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_80),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_99),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_64),
.B(n_62),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_122),
.B(n_23),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_66),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_93),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_121),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_86),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_118),
.B(n_119),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_91),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_65),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_85),
.A2(n_12),
.B(n_13),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_115),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_131),
.Y(n_152)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_125),
.A2(n_147),
.B1(n_42),
.B2(n_74),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_122),
.B(n_95),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_126),
.B(n_151),
.Y(n_175)
);

INVxp33_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_149),
.Y(n_164)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_92),
.C(n_82),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_150),
.C(n_11),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_111),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_82),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_141),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_121),
.A2(n_92),
.B1(n_97),
.B2(n_40),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_137),
.A2(n_34),
.B1(n_25),
.B2(n_27),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_107),
.A2(n_89),
.B(n_67),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_138),
.A2(n_19),
.B(n_20),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_139),
.A2(n_146),
.B1(n_19),
.B2(n_23),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_116),
.A2(n_65),
.B1(n_16),
.B2(n_81),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_143),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_145),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_102),
.A2(n_16),
.B1(n_89),
.B2(n_18),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_100),
.A2(n_42),
.B1(n_32),
.B2(n_25),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_34),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_108),
.B(n_109),
.C(n_100),
.Y(n_150)
);

NAND3xp33_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_21),
.C(n_20),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_138),
.A2(n_67),
.B(n_1),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_153),
.A2(n_157),
.B(n_172),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_74),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_155),
.B(n_174),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_156),
.A2(n_159),
.B1(n_164),
.B2(n_136),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_163),
.Y(n_185)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_21),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_154),
.Y(n_180)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_167),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_11),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_171),
.C(n_129),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_12),
.Y(n_170)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_30),
.C(n_24),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_134),
.A2(n_0),
.B(n_1),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_135),
.B(n_15),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_34),
.Y(n_176)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_137),
.B1(n_125),
.B2(n_141),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_183),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_152),
.Y(n_199)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_180),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_128),
.C(n_139),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_186),
.C(n_187),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_149),
.Y(n_182)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

FAx1_ASAP7_75t_SL g183 ( 
.A(n_163),
.B(n_128),
.CI(n_147),
.CON(n_183),
.SN(n_183)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_148),
.C(n_30),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_174),
.C(n_168),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_173),
.Y(n_191)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_30),
.C(n_25),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_197),
.C(n_162),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_127),
.Y(n_193)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_194),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_30),
.C(n_27),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_210),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_161),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_200),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_197),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_205),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_172),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_204),
.B(n_209),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_153),
.C(n_157),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_212),
.C(n_184),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_195),
.A2(n_159),
.B(n_167),
.Y(n_209)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_181),
.B(n_169),
.CI(n_15),
.CON(n_210),
.SN(n_210)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_185),
.B(n_136),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_184),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_30),
.C(n_27),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_221),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_220),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_214),
.A2(n_188),
.B1(n_196),
.B2(n_179),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_218),
.A2(n_203),
.B1(n_202),
.B2(n_210),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_211),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_186),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_192),
.C(n_177),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_30),
.C(n_27),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_206),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_212),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_213),
.A2(n_189),
.B1(n_183),
.B2(n_23),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_225),
.A2(n_226),
.B1(n_0),
.B2(n_1),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_207),
.A2(n_17),
.B1(n_13),
.B2(n_24),
.Y(n_226)
);

AOI21xp33_ASAP7_75t_L g228 ( 
.A1(n_198),
.A2(n_17),
.B(n_13),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_228),
.A2(n_2),
.B(n_3),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_235),
.Y(n_250)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_234),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_15),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_237),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_224),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_15),
.C(n_24),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_239),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_217),
.C(n_219),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_227),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_240),
.B(n_3),
.Y(n_247)
);

MAJx2_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_223),
.C(n_3),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_235),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_237),
.A2(n_24),
.B(n_3),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_247),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_2),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_246),
.A2(n_6),
.B(n_7),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_4),
.Y(n_253)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_251),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_243),
.A2(n_229),
.B1(n_5),
.B2(n_6),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_253),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_4),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_254),
.B(n_255),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_5),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_5),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_256),
.A2(n_258),
.B(n_259),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_5),
.C(n_6),
.Y(n_258)
);

OAI21x1_ASAP7_75t_L g261 ( 
.A1(n_259),
.A2(n_6),
.B(n_7),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_260),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_262),
.Y(n_265)
);

AO21x1_ASAP7_75t_L g268 ( 
.A1(n_265),
.A2(n_267),
.B(n_264),
.Y(n_268)
);

A2O1A1O1Ixp25_ASAP7_75t_L g267 ( 
.A1(n_263),
.A2(n_245),
.B(n_246),
.C(n_257),
.D(n_9),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_268),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_8),
.C(n_9),
.Y(n_269)
);

BUFx24_ASAP7_75t_SL g271 ( 
.A(n_270),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_271),
.B(n_269),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_9),
.Y(n_273)
);


endmodule