module real_jpeg_23559_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_1),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_1),
.A2(n_20),
.B1(n_53),
.B2(n_56),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_1),
.A2(n_20),
.B1(n_28),
.B2(n_29),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_2),
.A2(n_19),
.B1(n_21),
.B2(n_57),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_2),
.B(n_24),
.C(n_29),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_2),
.A2(n_39),
.B1(n_90),
.B2(n_97),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_5),
.A2(n_19),
.B1(n_21),
.B2(n_44),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_6),
.A2(n_19),
.B1(n_21),
.B2(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_11),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_74),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_72),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_50),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_15),
.B(n_50),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_33),
.C(n_38),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_16),
.A2(n_17),
.B1(n_33),
.B2(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_22),
.B1(n_30),
.B2(n_31),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_18),
.A2(n_22),
.B1(n_30),
.B2(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_19),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_21),
.B1(n_24),
.B2(n_26),
.Y(n_23)
);

AO22x1_ASAP7_75t_L g35 ( 
.A1(n_19),
.A2(n_21),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

OAI32xp33_ASAP7_75t_L g52 ( 
.A1(n_19),
.A2(n_36),
.A3(n_53),
.B1(n_55),
.B2(n_58),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_19),
.B(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_21),
.B(n_37),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_22),
.A2(n_30),
.B1(n_31),
.B2(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_27),
.Y(n_22)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_27),
.B(n_57),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_28),
.B(n_103),
.Y(n_102)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_35),
.A2(n_55),
.B1(n_69),
.B2(n_71),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_35),
.B(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_36),
.A2(n_37),
.B1(n_53),
.B2(n_56),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_38),
.B(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_43),
.B(n_45),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_60),
.B(n_61),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_39),
.A2(n_87),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_40),
.A2(n_86),
.B1(n_88),
.B2(n_89),
.Y(n_85)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_48),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_65),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_59),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_53),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

HAxp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_57),
.CON(n_55),
.SN(n_55)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_57),
.B(n_98),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_83),
.B(n_106),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_81),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_76),
.B(n_81),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_79),
.Y(n_92)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_93),
.B(n_105),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_92),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_92),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_100),
.B(n_104),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_95),
.B(n_96),
.Y(n_104)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);


endmodule