module fake_aes_4387_n_545 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_545);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_545;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_10), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_68), .Y(n_79) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_74), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_22), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_58), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_59), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_14), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_35), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_30), .Y(n_86) );
HB1xp67_ASAP7_75t_L g87 ( .A(n_34), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_23), .Y(n_88) );
BUFx2_ASAP7_75t_L g89 ( .A(n_53), .Y(n_89) );
INVxp33_ASAP7_75t_SL g90 ( .A(n_3), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_27), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_10), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_0), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_66), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_32), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_0), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_8), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_6), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_70), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_45), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_48), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_9), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_64), .Y(n_103) );
BUFx2_ASAP7_75t_L g104 ( .A(n_21), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_44), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_19), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_9), .Y(n_107) );
INVxp67_ASAP7_75t_SL g108 ( .A(n_61), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_52), .Y(n_109) );
BUFx3_ASAP7_75t_L g110 ( .A(n_41), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_63), .Y(n_111) );
BUFx3_ASAP7_75t_L g112 ( .A(n_8), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_72), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_7), .Y(n_114) );
CKINVDCx6p67_ASAP7_75t_R g115 ( .A(n_110), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_82), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_79), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_84), .Y(n_118) );
AND2x2_ASAP7_75t_L g119 ( .A(n_89), .B(n_1), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_82), .Y(n_120) );
INVx3_ASAP7_75t_L g121 ( .A(n_112), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_89), .B(n_1), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_84), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_112), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_85), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_114), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_104), .B(n_2), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_85), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_105), .Y(n_129) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_90), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_86), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_104), .B(n_4), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_80), .B(n_5), .Y(n_133) );
INVx3_ASAP7_75t_L g134 ( .A(n_114), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_86), .Y(n_135) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_88), .A2(n_40), .B(n_76), .Y(n_136) );
INVx6_ASAP7_75t_L g137 ( .A(n_110), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_121), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_121), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_119), .Y(n_140) );
INVx4_ASAP7_75t_L g141 ( .A(n_115), .Y(n_141) );
NAND2x1p5_ASAP7_75t_L g142 ( .A(n_119), .B(n_78), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_119), .Y(n_143) );
NAND2x1p5_ASAP7_75t_L g144 ( .A(n_132), .B(n_78), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_115), .B(n_87), .Y(n_145) );
XOR2x2_ASAP7_75t_L g146 ( .A(n_130), .B(n_5), .Y(n_146) );
AND2x6_ASAP7_75t_L g147 ( .A(n_132), .B(n_88), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_121), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_121), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_124), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_124), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_132), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_118), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_124), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_124), .Y(n_155) );
NAND2x1p5_ASAP7_75t_L g156 ( .A(n_118), .B(n_94), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_123), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_129), .Y(n_158) );
INVxp67_ASAP7_75t_SL g159 ( .A(n_122), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_126), .Y(n_160) );
BUFx2_ASAP7_75t_L g161 ( .A(n_115), .Y(n_161) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_122), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_126), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_159), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_162), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_158), .Y(n_166) );
AND2x4_ASAP7_75t_SL g167 ( .A(n_141), .B(n_133), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_156), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_139), .Y(n_169) );
INVx5_ASAP7_75t_L g170 ( .A(n_141), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_156), .B(n_133), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_156), .B(n_133), .Y(n_172) );
NOR3xp33_ASAP7_75t_SL g173 ( .A(n_158), .B(n_117), .C(n_130), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_140), .B(n_127), .Y(n_174) );
O2A1O1Ixp5_ASAP7_75t_L g175 ( .A1(n_143), .A2(n_127), .B(n_123), .C(n_135), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_152), .B(n_125), .Y(n_176) );
OAI22xp33_ASAP7_75t_L g177 ( .A1(n_142), .A2(n_97), .B1(n_125), .B2(n_135), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_142), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_144), .Y(n_179) );
HB1xp67_ASAP7_75t_L g180 ( .A(n_144), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_145), .B(n_128), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_161), .B(n_97), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_147), .B(n_128), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_147), .B(n_131), .Y(n_184) );
OR2x6_ASAP7_75t_L g185 ( .A(n_141), .B(n_92), .Y(n_185) );
BUFx3_ASAP7_75t_L g186 ( .A(n_161), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_147), .B(n_131), .Y(n_187) );
OR2x6_ASAP7_75t_SL g188 ( .A(n_146), .B(n_105), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_138), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_153), .B(n_81), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_147), .B(n_126), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_139), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_138), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_139), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_146), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_147), .B(n_92), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_164), .Y(n_197) );
INVx4_ASAP7_75t_L g198 ( .A(n_170), .Y(n_198) );
INVx4_ASAP7_75t_L g199 ( .A(n_170), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_181), .B(n_147), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_176), .Y(n_201) );
BUFx2_ASAP7_75t_L g202 ( .A(n_185), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_189), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_170), .Y(n_204) );
CKINVDCx16_ASAP7_75t_R g205 ( .A(n_188), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_189), .Y(n_206) );
OAI221xp5_ASAP7_75t_L g207 ( .A1(n_165), .A2(n_174), .B1(n_178), .B2(n_179), .C(n_180), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_186), .B(n_163), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_186), .B(n_163), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g210 ( .A1(n_168), .A2(n_157), .B1(n_163), .B2(n_160), .Y(n_210) );
INVxp67_ASAP7_75t_L g211 ( .A(n_185), .Y(n_211) );
BUFx4f_ASAP7_75t_L g212 ( .A(n_185), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g213 ( .A1(n_175), .A2(n_120), .B(n_116), .C(n_154), .Y(n_213) );
AOI22xp33_ASAP7_75t_SL g214 ( .A1(n_166), .A2(n_113), .B1(n_126), .B2(n_134), .Y(n_214) );
NOR2x1_ASAP7_75t_SL g215 ( .A(n_185), .B(n_94), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_171), .A2(n_160), .B(n_155), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_170), .Y(n_217) );
BUFx2_ASAP7_75t_L g218 ( .A(n_166), .Y(n_218) );
O2A1O1Ixp33_ASAP7_75t_L g219 ( .A1(n_177), .A2(n_102), .B(n_96), .C(n_107), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_184), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_167), .B(n_148), .Y(n_221) );
AOI22xp33_ASAP7_75t_SL g222 ( .A1(n_167), .A2(n_113), .B1(n_134), .B2(n_93), .Y(n_222) );
INVx2_ASAP7_75t_SL g223 ( .A(n_170), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_184), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_184), .B(n_148), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_193), .Y(n_226) );
INVx3_ASAP7_75t_L g227 ( .A(n_169), .Y(n_227) );
INVx5_ASAP7_75t_L g228 ( .A(n_196), .Y(n_228) );
BUFx2_ASAP7_75t_L g229 ( .A(n_182), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_203), .Y(n_230) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_213), .A2(n_191), .B(n_171), .Y(n_231) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_212), .A2(n_196), .B1(n_172), .B2(n_183), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_203), .Y(n_233) );
AND2x4_ASAP7_75t_L g234 ( .A(n_201), .B(n_196), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_197), .Y(n_235) );
NAND2x1p5_ASAP7_75t_L g236 ( .A(n_212), .B(n_172), .Y(n_236) );
NAND3xp33_ASAP7_75t_L g237 ( .A(n_213), .B(n_173), .C(n_190), .Y(n_237) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_202), .Y(n_238) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_216), .A2(n_111), .B(n_95), .Y(n_239) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_206), .A2(n_111), .B(n_95), .Y(n_240) );
AOI21x1_ASAP7_75t_L g241 ( .A1(n_200), .A2(n_136), .B(n_116), .Y(n_241) );
AOI21x1_ASAP7_75t_L g242 ( .A1(n_206), .A2(n_136), .B(n_116), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_205), .Y(n_243) );
INVx3_ASAP7_75t_SL g244 ( .A(n_198), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_226), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_211), .B(n_187), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_226), .Y(n_247) );
INVx3_ASAP7_75t_L g248 ( .A(n_204), .Y(n_248) );
OAI21x1_ASAP7_75t_L g249 ( .A1(n_217), .A2(n_136), .B(n_190), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_227), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_211), .B(n_169), .Y(n_251) );
CKINVDCx6p67_ASAP7_75t_R g252 ( .A(n_228), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_207), .B(n_188), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_204), .Y(n_254) );
AO21x2_ASAP7_75t_L g255 ( .A1(n_215), .A2(n_120), .B(n_109), .Y(n_255) );
NOR2xp33_ASAP7_75t_SL g256 ( .A(n_198), .B(n_192), .Y(n_256) );
BUFx12f_ASAP7_75t_L g257 ( .A(n_243), .Y(n_257) );
OAI21x1_ASAP7_75t_L g258 ( .A1(n_241), .A2(n_136), .B(n_217), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_234), .Y(n_259) );
OR2x2_ASAP7_75t_L g260 ( .A(n_245), .B(n_229), .Y(n_260) );
OR2x6_ASAP7_75t_L g261 ( .A(n_236), .B(n_204), .Y(n_261) );
AOI221xp5_ASAP7_75t_L g262 ( .A1(n_253), .A2(n_219), .B1(n_195), .B2(n_218), .C(n_222), .Y(n_262) );
INVxp67_ASAP7_75t_L g263 ( .A(n_238), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_237), .A2(n_195), .B1(n_214), .B2(n_208), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_232), .A2(n_210), .B1(n_228), .B2(n_209), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_237), .A2(n_208), .B1(n_209), .B2(n_220), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_256), .B(n_204), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_235), .B(n_208), .Y(n_268) );
OAI21x1_ASAP7_75t_L g269 ( .A1(n_241), .A2(n_136), .B(n_227), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_230), .A2(n_223), .B(n_227), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_235), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_232), .A2(n_228), .B1(n_209), .B2(n_221), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_230), .Y(n_273) );
AOI21xp33_ASAP7_75t_L g274 ( .A1(n_231), .A2(n_223), .B(n_199), .Y(n_274) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_244), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_245), .Y(n_276) );
OAI21xp5_ASAP7_75t_L g277 ( .A1(n_249), .A2(n_225), .B(n_194), .Y(n_277) );
OAI211xp5_ASAP7_75t_L g278 ( .A1(n_251), .A2(n_93), .B(n_96), .C(n_107), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_275), .B(n_256), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_273), .Y(n_280) );
AO21x2_ASAP7_75t_L g281 ( .A1(n_274), .A2(n_242), .B(n_249), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_276), .Y(n_282) );
NAND2x1p5_ASAP7_75t_SL g283 ( .A(n_267), .B(n_254), .Y(n_283) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_260), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_273), .B(n_247), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g286 ( .A1(n_262), .A2(n_234), .B1(n_236), .B2(n_244), .Y(n_286) );
AOI21xp5_ASAP7_75t_SL g287 ( .A1(n_267), .A2(n_240), .B(n_239), .Y(n_287) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_260), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_271), .B(n_247), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_269), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_269), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_268), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_258), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_277), .Y(n_294) );
OA21x2_ASAP7_75t_L g295 ( .A1(n_258), .A2(n_249), .B(n_242), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_261), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_259), .B(n_230), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_261), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_275), .B(n_233), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_261), .Y(n_300) );
BUFx3_ASAP7_75t_L g301 ( .A(n_299), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_285), .B(n_240), .Y(n_302) );
INVx3_ASAP7_75t_L g303 ( .A(n_293), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_285), .B(n_240), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_280), .B(n_240), .Y(n_305) );
INVx1_ASAP7_75t_SL g306 ( .A(n_299), .Y(n_306) );
INVx5_ASAP7_75t_L g307 ( .A(n_280), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_284), .B(n_263), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_288), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_298), .B(n_261), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_293), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_289), .B(n_233), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_282), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_298), .B(n_275), .Y(n_314) );
AOI211xp5_ASAP7_75t_L g315 ( .A1(n_287), .A2(n_278), .B(n_244), .C(n_275), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_282), .Y(n_316) );
AOI322xp5_ASAP7_75t_L g317 ( .A1(n_286), .A2(n_264), .A3(n_98), .B1(n_257), .B2(n_120), .C1(n_109), .C2(n_266), .Y(n_317) );
INVx1_ASAP7_75t_SL g318 ( .A(n_279), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_294), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_297), .B(n_233), .Y(n_320) );
AOI22xp33_ASAP7_75t_SL g321 ( .A1(n_292), .A2(n_272), .B1(n_265), .B2(n_236), .Y(n_321) );
INVx2_ASAP7_75t_SL g322 ( .A(n_297), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_289), .Y(n_323) );
INVxp67_ASAP7_75t_SL g324 ( .A(n_292), .Y(n_324) );
INVx4_ASAP7_75t_L g325 ( .A(n_296), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_294), .Y(n_326) );
BUFx3_ASAP7_75t_L g327 ( .A(n_296), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_300), .B(n_231), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_300), .B(n_231), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_283), .Y(n_330) );
AOI221xp5_ASAP7_75t_L g331 ( .A1(n_308), .A2(n_98), .B1(n_103), .B2(n_101), .C(n_99), .Y(n_331) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_315), .B(n_257), .Y(n_332) );
AOI33xp33_ASAP7_75t_L g333 ( .A1(n_313), .A2(n_100), .A3(n_106), .B1(n_83), .B2(n_91), .B3(n_234), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_324), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_323), .B(n_283), .Y(n_335) );
NOR3xp33_ASAP7_75t_L g336 ( .A(n_315), .B(n_134), .C(n_108), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_311), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_328), .B(n_281), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_322), .B(n_281), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_322), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_311), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_311), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_313), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_316), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_316), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_328), .B(n_281), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_312), .B(n_287), .Y(n_347) );
AND2x4_ASAP7_75t_L g348 ( .A(n_310), .B(n_290), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_329), .B(n_290), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_306), .B(n_291), .Y(n_350) );
BUFx3_ASAP7_75t_L g351 ( .A(n_307), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_329), .B(n_291), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_301), .B(n_295), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_309), .B(n_248), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_312), .B(n_231), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_302), .B(n_239), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_302), .B(n_239), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_303), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_301), .B(n_295), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_319), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_301), .B(n_6), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_303), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_303), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_319), .B(n_295), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_326), .Y(n_365) );
INVx1_ASAP7_75t_SL g366 ( .A(n_306), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_326), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_304), .B(n_295), .Y(n_368) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_320), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_320), .B(n_239), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_304), .B(n_7), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_327), .B(n_325), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_303), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_305), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_369), .B(n_305), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_343), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_343), .Y(n_377) );
OAI21xp5_ASAP7_75t_L g378 ( .A1(n_333), .A2(n_332), .B(n_334), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_340), .B(n_327), .Y(n_379) );
INVxp67_ASAP7_75t_SL g380 ( .A(n_334), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_344), .B(n_310), .Y(n_381) );
BUFx2_ASAP7_75t_L g382 ( .A(n_351), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_344), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_345), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_345), .B(n_310), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_360), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_368), .B(n_310), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_366), .B(n_327), .Y(n_388) );
INVxp67_ASAP7_75t_L g389 ( .A(n_361), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_360), .Y(n_390) );
AND3x2_ASAP7_75t_L g391 ( .A(n_336), .B(n_314), .C(n_330), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_374), .B(n_366), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_365), .Y(n_393) );
AND2x4_ASAP7_75t_SL g394 ( .A(n_372), .B(n_314), .Y(n_394) );
INVx1_ASAP7_75t_SL g395 ( .A(n_351), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_374), .B(n_325), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_368), .B(n_314), .Y(n_397) );
INVx1_ASAP7_75t_SL g398 ( .A(n_351), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_365), .Y(n_399) );
INVx1_ASAP7_75t_SL g400 ( .A(n_372), .Y(n_400) );
OR2x6_ASAP7_75t_L g401 ( .A(n_335), .B(n_325), .Y(n_401) );
INVx1_ASAP7_75t_SL g402 ( .A(n_353), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_349), .B(n_314), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_349), .B(n_325), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_367), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_367), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_335), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_352), .B(n_330), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_354), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_339), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_371), .B(n_307), .Y(n_411) );
INVx1_ASAP7_75t_SL g412 ( .A(n_353), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_338), .B(n_307), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_339), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_352), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_347), .A2(n_321), .B1(n_318), .B2(n_255), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_338), .B(n_307), .Y(n_417) );
INVx2_ASAP7_75t_SL g418 ( .A(n_350), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_350), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_331), .A2(n_318), .B1(n_307), .B2(n_255), .Y(n_420) );
NAND2xp33_ASAP7_75t_L g421 ( .A(n_370), .B(n_307), .Y(n_421) );
INVx1_ASAP7_75t_SL g422 ( .A(n_359), .Y(n_422) );
NOR2xp67_ASAP7_75t_SL g423 ( .A(n_370), .B(n_228), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_359), .B(n_317), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_346), .B(n_317), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_364), .Y(n_426) );
INVxp67_ASAP7_75t_L g427 ( .A(n_380), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_376), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_377), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_403), .B(n_346), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_424), .A2(n_348), .B1(n_355), .B2(n_356), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_402), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_407), .B(n_364), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_426), .B(n_357), .Y(n_434) );
OAI21xp5_ASAP7_75t_SL g435 ( .A1(n_378), .A2(n_348), .B(n_363), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_402), .Y(n_436) );
OAI22xp33_ASAP7_75t_L g437 ( .A1(n_378), .A2(n_373), .B1(n_363), .B2(n_362), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_425), .A2(n_348), .B1(n_373), .B2(n_358), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_409), .A2(n_348), .B1(n_337), .B2(n_341), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_383), .Y(n_440) );
INVx3_ASAP7_75t_SL g441 ( .A(n_394), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_384), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_386), .Y(n_443) );
AOI32xp33_ASAP7_75t_L g444 ( .A1(n_421), .A2(n_358), .A3(n_362), .B1(n_134), .B2(n_341), .Y(n_444) );
OAI21xp5_ASAP7_75t_SL g445 ( .A1(n_391), .A2(n_342), .B(n_337), .Y(n_445) );
AOI32xp33_ASAP7_75t_L g446 ( .A1(n_400), .A2(n_342), .A3(n_83), .B1(n_91), .B2(n_248), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_389), .A2(n_255), .B1(n_248), .B2(n_254), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_423), .A2(n_255), .B1(n_248), .B2(n_254), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_390), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_393), .Y(n_450) );
OAI221xp5_ASAP7_75t_L g451 ( .A1(n_416), .A2(n_137), .B1(n_251), .B2(n_250), .C(n_246), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_415), .B(n_11), .Y(n_452) );
NAND3xp33_ASAP7_75t_SL g453 ( .A(n_395), .B(n_270), .C(n_199), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_399), .Y(n_454) );
OAI21xp33_ASAP7_75t_L g455 ( .A1(n_387), .A2(n_250), .B(n_234), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_410), .B(n_11), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_382), .Y(n_457) );
XOR2x2_ASAP7_75t_L g458 ( .A(n_400), .B(n_12), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_405), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_411), .A2(n_252), .B1(n_137), .B2(n_246), .Y(n_460) );
INVxp67_ASAP7_75t_SL g461 ( .A(n_413), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_406), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_414), .B(n_12), .Y(n_463) );
OAI22xp5_ASAP7_75t_SL g464 ( .A1(n_401), .A2(n_252), .B1(n_199), .B2(n_198), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_381), .Y(n_465) );
OAI22xp33_ASAP7_75t_L g466 ( .A1(n_401), .A2(n_252), .B1(n_137), .B2(n_224), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_408), .B(n_137), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_417), .A2(n_137), .B1(n_169), .B2(n_155), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_385), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_404), .B(n_13), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_392), .Y(n_471) );
INVx2_ASAP7_75t_SL g472 ( .A(n_441), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_457), .B(n_397), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_431), .B(n_418), .Y(n_474) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_436), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_465), .B(n_422), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_428), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_461), .B(n_422), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_435), .A2(n_398), .B(n_395), .C(n_412), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_429), .Y(n_480) );
OAI211xp5_ASAP7_75t_SL g481 ( .A1(n_435), .A2(n_420), .B(n_398), .C(n_412), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_458), .A2(n_401), .B1(n_379), .B2(n_375), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_440), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_469), .B(n_419), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_471), .B(n_388), .Y(n_485) );
INVxp67_ASAP7_75t_L g486 ( .A(n_427), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_442), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_439), .A2(n_396), .B1(n_154), .B2(n_151), .Y(n_488) );
BUFx3_ASAP7_75t_L g489 ( .A(n_470), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_443), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_434), .B(n_15), .Y(n_491) );
AOI21xp33_ASAP7_75t_SL g492 ( .A1(n_445), .A2(n_16), .B(n_17), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_433), .B(n_18), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_430), .B(n_20), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_449), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_438), .B(n_24), .Y(n_496) );
INVxp67_ASAP7_75t_L g497 ( .A(n_456), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_445), .A2(n_151), .B(n_150), .Y(n_498) );
AOI21xp5_ASAP7_75t_SL g499 ( .A1(n_439), .A2(n_25), .B(n_26), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_455), .A2(n_150), .B1(n_149), .B2(n_193), .Y(n_500) );
NAND2xp33_ASAP7_75t_SL g501 ( .A(n_432), .B(n_28), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_475), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_475), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_477), .Y(n_504) );
NAND3xp33_ASAP7_75t_L g505 ( .A(n_482), .B(n_446), .C(n_437), .Y(n_505) );
AOI211xp5_ASAP7_75t_SL g506 ( .A1(n_499), .A2(n_466), .B(n_451), .C(n_464), .Y(n_506) );
OAI311xp33_ASAP7_75t_L g507 ( .A1(n_482), .A2(n_452), .A3(n_463), .B1(n_444), .C1(n_447), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_492), .A2(n_467), .B(n_453), .C(n_462), .Y(n_508) );
INVxp67_ASAP7_75t_SL g509 ( .A(n_488), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_479), .A2(n_472), .B1(n_489), .B2(n_478), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_480), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_483), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_481), .A2(n_459), .B1(n_454), .B2(n_450), .Y(n_513) );
OAI211xp5_ASAP7_75t_L g514 ( .A1(n_486), .A2(n_460), .B(n_448), .C(n_468), .Y(n_514) );
NAND4xp25_ASAP7_75t_L g515 ( .A(n_494), .B(n_149), .C(n_31), .D(n_33), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_474), .A2(n_29), .B1(n_36), .B2(n_37), .Y(n_516) );
AOI21xp33_ASAP7_75t_SL g517 ( .A1(n_473), .A2(n_497), .B(n_476), .Y(n_517) );
OAI21xp5_ASAP7_75t_SL g518 ( .A1(n_500), .A2(n_38), .B(n_39), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_487), .B(n_42), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_504), .Y(n_520) );
OAI22xp33_ASAP7_75t_L g521 ( .A1(n_510), .A2(n_485), .B1(n_484), .B2(n_490), .Y(n_521) );
AOI321xp33_ASAP7_75t_L g522 ( .A1(n_509), .A2(n_496), .A3(n_500), .B1(n_495), .B2(n_491), .C(n_493), .Y(n_522) );
NAND5xp2_ASAP7_75t_L g523 ( .A(n_506), .B(n_498), .C(n_501), .D(n_47), .E(n_49), .Y(n_523) );
AO21x1_ASAP7_75t_L g524 ( .A1(n_508), .A2(n_43), .B(n_46), .Y(n_524) );
AOI222xp33_ASAP7_75t_L g525 ( .A1(n_509), .A2(n_50), .B1(n_51), .B2(n_54), .C1(n_55), .C2(n_56), .Y(n_525) );
AOI211x1_ASAP7_75t_L g526 ( .A1(n_505), .A2(n_57), .B(n_60), .C(n_62), .Y(n_526) );
AOI221xp5_ASAP7_75t_L g527 ( .A1(n_507), .A2(n_65), .B1(n_67), .B2(n_69), .C(n_71), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_508), .A2(n_73), .B(n_75), .Y(n_528) );
XOR2xp5_ASAP7_75t_L g529 ( .A(n_515), .B(n_77), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_520), .B(n_513), .Y(n_530) );
OAI21x1_ASAP7_75t_SL g531 ( .A1(n_524), .A2(n_517), .B(n_513), .Y(n_531) );
AND2x4_ASAP7_75t_L g532 ( .A(n_528), .B(n_502), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_522), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_521), .B(n_503), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_534), .Y(n_535) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_533), .Y(n_536) );
OR4x2_ASAP7_75t_L g537 ( .A(n_531), .B(n_523), .C(n_526), .D(n_527), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_536), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_535), .B(n_530), .Y(n_539) );
INVxp67_ASAP7_75t_SL g540 ( .A(n_538), .Y(n_540) );
INVx3_ASAP7_75t_L g541 ( .A(n_539), .Y(n_541) );
INVx4_ASAP7_75t_L g542 ( .A(n_541), .Y(n_542) );
AOI222xp33_ASAP7_75t_SL g543 ( .A1(n_542), .A2(n_541), .B1(n_536), .B2(n_540), .C1(n_537), .C2(n_518), .Y(n_543) );
AOI322xp5_ASAP7_75t_L g544 ( .A1(n_543), .A2(n_532), .A3(n_519), .B1(n_512), .B2(n_511), .C1(n_516), .C2(n_525), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_544), .A2(n_529), .B(n_514), .Y(n_545) );
endmodule