module real_jpeg_25563_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_1),
.A2(n_42),
.B1(n_44),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_1),
.A2(n_28),
.B1(n_36),
.B2(n_51),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_1),
.A2(n_51),
.B1(n_63),
.B2(n_68),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_1),
.A2(n_51),
.B1(n_72),
.B2(n_138),
.Y(n_344)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_3),
.A2(n_63),
.B1(n_68),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_3),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_3),
.A2(n_42),
.B1(n_44),
.B2(n_86),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_3),
.A2(n_86),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_3),
.A2(n_28),
.B1(n_36),
.B2(n_86),
.Y(n_192)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_5),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_5),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_5),
.A2(n_60),
.B1(n_63),
.B2(n_68),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_5),
.A2(n_42),
.B1(n_44),
.B2(n_60),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_5),
.A2(n_28),
.B1(n_36),
.B2(n_60),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_7),
.A2(n_113),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_7),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_7),
.A2(n_63),
.B1(n_68),
.B2(n_164),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_7),
.A2(n_42),
.B1(n_44),
.B2(n_164),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_7),
.A2(n_28),
.B1(n_36),
.B2(n_164),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_8),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_8),
.A2(n_41),
.B1(n_63),
.B2(n_68),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_8),
.A2(n_41),
.B1(n_72),
.B2(n_111),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_8),
.A2(n_28),
.B1(n_36),
.B2(n_41),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_9),
.Y(n_82)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_11),
.A2(n_59),
.B1(n_72),
.B2(n_74),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_11),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_11),
.A2(n_63),
.B1(n_68),
.B2(n_74),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_11),
.A2(n_42),
.B1(n_44),
.B2(n_74),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_11),
.A2(n_28),
.B1(n_36),
.B2(n_74),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_12),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_12),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_12),
.A2(n_63),
.B1(n_68),
.B2(n_110),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_12),
.A2(n_42),
.B1(n_44),
.B2(n_110),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_12),
.A2(n_28),
.B1(n_36),
.B2(n_110),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_13),
.B(n_137),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_13),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_13),
.B(n_62),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_13),
.B(n_42),
.C(n_82),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_13),
.A2(n_63),
.B1(n_68),
.B2(n_216),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_13),
.B(n_128),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_13),
.A2(n_42),
.B1(n_44),
.B2(n_216),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_13),
.B(n_28),
.C(n_47),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_13),
.A2(n_27),
.B(n_276),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_15),
.A2(n_28),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_15),
.A2(n_37),
.B1(n_42),
.B2(n_44),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_15),
.A2(n_37),
.B1(n_63),
.B2(n_68),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_15),
.A2(n_37),
.B1(n_59),
.B2(n_137),
.Y(n_351)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_16),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_16),
.B(n_277),
.Y(n_276)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_16),
.Y(n_290)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI21xp33_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_354),
.B(n_357),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_349),
.B(n_353),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_336),
.B(n_348),
.Y(n_20)
);

OAI31xp33_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_140),
.A3(n_154),
.B(n_333),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_117),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_23),
.B(n_117),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_77),
.C(n_93),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_24),
.A2(n_77),
.B1(n_78),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_24),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_53),
.Y(n_24)
);

AOI21xp33_ASAP7_75t_L g118 ( 
.A1(n_25),
.A2(n_26),
.B(n_55),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_38),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_26),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_26),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_26),
.A2(n_38),
.B1(n_39),
.B2(n_54),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_32),
.B(n_35),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_27),
.A2(n_35),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_27),
.A2(n_98),
.B1(n_99),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_27),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_27),
.A2(n_192),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_27),
.B(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_27),
.A2(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_28),
.A2(n_36),
.B1(n_47),
.B2(n_48),
.Y(n_49)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_29),
.Y(n_193)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_34),
.B(n_216),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_36),
.B(n_301),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_45),
.B1(n_50),
.B2(n_52),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_40),
.A2(n_45),
.B1(n_52),
.B2(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_42),
.A2(n_44),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_42),
.B(n_283),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_45),
.A2(n_52),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_45),
.B(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_45),
.A2(n_52),
.B1(n_248),
.B2(n_250),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_49),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_49),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_49),
.A2(n_89),
.B1(n_104),
.B2(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_49),
.A2(n_175),
.B(n_212),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_49),
.A2(n_212),
.B(n_249),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_49),
.B(n_216),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_50),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_52),
.B(n_213),
.Y(n_264)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_61),
.B(n_69),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_57),
.A2(n_61),
.B1(n_114),
.B2(n_136),
.Y(n_135)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_59),
.B1(n_66),
.B2(n_67),
.Y(n_76)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_61),
.B(n_71),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_61),
.A2(n_114),
.B1(n_136),
.B2(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_61),
.A2(n_69),
.B(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_62),
.A2(n_75),
.B1(n_109),
.B2(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_62),
.A2(n_75),
.B1(n_343),
.B2(n_344),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_62),
.A2(n_75),
.B1(n_344),
.B2(n_351),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_62),
.A2(n_75),
.B(n_351),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_62)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_68),
.B1(n_82),
.B2(n_83),
.Y(n_84)
);

NAND2xp33_ASAP7_75t_SL g188 ( 
.A(n_63),
.B(n_67),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_63),
.B(n_242),
.Y(n_241)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI32xp33_ASAP7_75t_L g186 ( 
.A1(n_66),
.A2(n_68),
.A3(n_111),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_75),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_75),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_75),
.A2(n_116),
.B(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_88),
.B(n_92),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_88),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_85),
.B2(n_87),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_80),
.A2(n_81),
.B1(n_85),
.B2(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_80),
.A2(n_81),
.B1(n_130),
.B2(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_80),
.A2(n_182),
.B(n_184),
.Y(n_181)
);

OAI21xp33_ASAP7_75t_L g252 ( 
.A1(n_80),
.A2(n_184),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_81),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_81),
.A2(n_106),
.B(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_81),
.A2(n_168),
.B(n_221),
.Y(n_220)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_87),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_89),
.A2(n_263),
.B(n_264),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_89),
.A2(n_264),
.B(n_281),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_91),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_93),
.A2(n_94),
.B1(n_328),
.B2(n_330),
.Y(n_327)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_105),
.C(n_107),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_95),
.A2(n_96),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_101),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_97),
.A2(n_101),
.B1(n_102),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_97),
.Y(n_177)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_105),
.B(n_107),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_114),
.B(n_115),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_111),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_L g215 ( 
.A1(n_111),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_120),
.C(n_122),
.Y(n_153)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_135),
.B2(n_139),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_131),
.B1(n_132),
.B2(n_134),
.Y(n_124)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_132),
.C(n_135),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_127),
.A2(n_128),
.B1(n_183),
.B2(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_127),
.A2(n_128),
.B(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_128),
.B(n_169),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_132),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_132),
.B(n_147),
.C(n_151),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_135),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_135),
.A2(n_139),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_135),
.B(n_143),
.C(n_146),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_141),
.A2(n_334),
.B(n_335),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_153),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_142),
.B(n_153),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_148),
.Y(n_343)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_152),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_326),
.B(n_332),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_201),
.B(n_325),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_194),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_157),
.B(n_194),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_176),
.C(n_178),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_158),
.A2(n_159),
.B1(n_176),
.B2(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_170),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_166),
.B2(n_167),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_166),
.C(n_170),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_163),
.Y(n_180)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_171),
.B(n_174),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_173),
.A2(n_190),
.B1(n_191),
.B2(n_193),
.Y(n_189)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_176),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_178),
.B(n_322),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.C(n_185),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_179),
.B(n_181),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_185),
.B(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_189),
.Y(n_218)
);

INVxp33_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_190),
.A2(n_287),
.B1(n_289),
.B2(n_291),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_193),
.A2(n_244),
.B(n_245),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_200),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_196),
.B(n_197),
.C(n_200),
.Y(n_331)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

O2A1O1Ixp33_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_234),
.B(n_319),
.C(n_324),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_228),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_228),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_218),
.C(n_219),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_204),
.A2(n_205),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_214),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_210),
.B2(n_211),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_210),
.C(n_214),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_209),
.Y(n_221)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_218),
.B(n_219),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.C(n_224),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_258),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_224),
.Y(n_258)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_229),
.B(n_232),
.C(n_233),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_313),
.B(n_318),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_265),
.B(n_312),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_254),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_239),
.B(n_254),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_247),
.C(n_251),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_240),
.B(n_308),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_243),
.Y(n_261)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_245),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_246),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_247),
.A2(n_251),
.B1(n_252),
.B2(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_247),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_250),
.Y(n_263)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_259),
.B2(n_260),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_255),
.B(n_261),
.C(n_262),
.Y(n_317)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_306),
.B(n_311),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_284),
.B(n_305),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_278),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_268),
.B(n_278),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_274),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_270),
.B(n_273),
.C(n_274),
.Y(n_310)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_275),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_282),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_279),
.A2(n_280),
.B1(n_282),
.B2(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_282),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_294),
.B(n_304),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_292),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_292),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_288),
.A2(n_290),
.B(n_298),
.Y(n_297)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_299),
.B(n_303),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_297),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_310),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_310),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_317),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_317),
.Y(n_318)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_321),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_331),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_331),
.Y(n_332)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_328),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_338),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_347),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_342),
.B1(n_345),
.B2(n_346),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_340),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_342),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_345),
.C(n_347),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_352),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_350),
.B(n_352),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_350),
.B(n_355),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_350),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_356),
.B(n_359),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_358),
.Y(n_357)
);


endmodule