module fake_jpeg_5145_n_180 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_180);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_13),
.B(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_33),
.Y(n_46)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_35),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_39),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_44),
.Y(n_66)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_52),
.Y(n_71)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_54),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_31),
.A2(n_27),
.B1(n_25),
.B2(n_17),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_20),
.Y(n_72)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_57),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_44),
.A2(n_31),
.B1(n_27),
.B2(n_25),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_58),
.A2(n_64),
.B1(n_16),
.B2(n_21),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_50),
.B(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_68),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_25),
.B1(n_32),
.B2(n_19),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_38),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_24),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_76),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_70),
.Y(n_79)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_16),
.Y(n_73)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_45),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_74),
.B(n_26),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_36),
.C(n_32),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_37),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_24),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_87),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_47),
.B1(n_28),
.B2(n_22),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_80),
.A2(n_81),
.B1(n_85),
.B2(n_88),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_75),
.A2(n_56),
.B1(n_52),
.B2(n_28),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_42),
.Y(n_82)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_84),
.A2(n_61),
.B(n_71),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_19),
.B1(n_22),
.B2(n_16),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_26),
.B1(n_15),
.B2(n_64),
.Y(n_111)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_30),
.B1(n_23),
.B2(n_29),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_92),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_42),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_76),
.B1(n_63),
.B2(n_68),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_93),
.B(n_73),
.Y(n_98)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_65),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_72),
.A2(n_29),
.B1(n_21),
.B2(n_23),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_96),
.A2(n_89),
.B1(n_86),
.B2(n_30),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_71),
.C(n_61),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_113),
.C(n_60),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_104),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_79),
.Y(n_100)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_109),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_58),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_103),
.A2(n_106),
.B(n_113),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_66),
.Y(n_104)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_90),
.B(n_59),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_59),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_60),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_111),
.B(n_96),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_37),
.C(n_51),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_106),
.A2(n_77),
.B(n_89),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_101),
.B1(n_103),
.B2(n_112),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_77),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_123),
.C(n_125),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_117),
.B(n_120),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_119),
.A2(n_101),
.B1(n_105),
.B2(n_111),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_L g120 ( 
.A1(n_104),
.A2(n_83),
.B(n_94),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_94),
.B1(n_85),
.B2(n_60),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_79),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_51),
.Y(n_126)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_129),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_0),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_115),
.B(n_112),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_128),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_1),
.Y(n_152)
);

INVxp33_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_134),
.A2(n_135),
.B(n_137),
.Y(n_144)
);

OA21x2_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_37),
.B(n_33),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_108),
.C(n_33),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_140),
.C(n_136),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_33),
.C(n_15),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_132),
.A2(n_114),
.B(n_127),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_143),
.A2(n_145),
.B(n_151),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_139),
.A2(n_127),
.B(n_129),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_147),
.C(n_149),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_121),
.C(n_125),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_141),
.B(n_115),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_150),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_118),
.C(n_117),
.Y(n_149)
);

XOR2x2_ASAP7_75t_SL g151 ( 
.A(n_137),
.B(n_0),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_151),
.B(n_135),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_142),
.Y(n_155)
);

OAI322xp33_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_14),
.A3(n_10),
.B1(n_3),
.B2(n_5),
.C1(n_1),
.C2(n_8),
.Y(n_153)
);

OA21x2_ASAP7_75t_SL g158 ( 
.A1(n_153),
.A2(n_10),
.B(n_3),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_155),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_156),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_144),
.A2(n_139),
.B(n_133),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_157),
.B(n_158),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_147),
.A2(n_140),
.B(n_134),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_146),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_166),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_156),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_2),
.C(n_3),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_167),
.A2(n_7),
.B(n_8),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g169 ( 
.A1(n_166),
.A2(n_155),
.A3(n_161),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_2),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_170),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_5),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_171),
.Y(n_173)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_167),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_172),
.A2(n_164),
.B1(n_165),
.B2(n_163),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_168),
.C(n_169),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_173),
.C(n_9),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_9),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_177),
.Y(n_180)
);


endmodule