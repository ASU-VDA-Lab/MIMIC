module fake_netlist_5_2583_n_426 (n_91, n_82, n_10, n_24, n_86, n_83, n_61, n_90, n_75, n_101, n_65, n_78, n_74, n_57, n_96, n_37, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_0, n_58, n_9, n_69, n_18, n_42, n_22, n_1, n_45, n_46, n_21, n_94, n_38, n_105, n_80, n_4, n_35, n_73, n_17, n_92, n_19, n_30, n_5, n_33, n_14, n_84, n_23, n_29, n_79, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_71, n_85, n_95, n_59, n_26, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_81, n_28, n_89, n_70, n_68, n_93, n_72, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_426);

input n_91;
input n_82;
input n_10;
input n_24;
input n_86;
input n_83;
input n_61;
input n_90;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_57;
input n_96;
input n_37;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_42;
input n_22;
input n_1;
input n_45;
input n_46;
input n_21;
input n_94;
input n_38;
input n_105;
input n_80;
input n_4;
input n_35;
input n_73;
input n_17;
input n_92;
input n_19;
input n_30;
input n_5;
input n_33;
input n_14;
input n_84;
input n_23;
input n_29;
input n_79;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_71;
input n_85;
input n_95;
input n_59;
input n_26;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_81;
input n_28;
input n_89;
input n_70;
input n_68;
input n_93;
input n_72;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;

output n_426;

wire n_137;
wire n_294;
wire n_318;
wire n_380;
wire n_419;
wire n_194;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_124;
wire n_146;
wire n_136;
wire n_315;
wire n_268;
wire n_408;
wire n_376;
wire n_127;
wire n_235;
wire n_226;
wire n_353;
wire n_351;
wire n_367;
wire n_397;
wire n_111;
wire n_155;
wire n_116;
wire n_423;
wire n_284;
wire n_245;
wire n_139;
wire n_280;
wire n_378;
wire n_382;
wire n_254;
wire n_302;
wire n_265;
wire n_293;
wire n_372;
wire n_244;
wire n_173;
wire n_198;
wire n_247;
wire n_314;
wire n_368;
wire n_321;
wire n_292;
wire n_417;
wire n_212;
wire n_385;
wire n_119;
wire n_275;
wire n_252;
wire n_295;
wire n_133;
wire n_330;
wire n_147;
wire n_373;
wire n_307;
wire n_150;
wire n_106;
wire n_209;
wire n_259;
wire n_375;
wire n_301;
wire n_186;
wire n_134;
wire n_191;
wire n_171;
wire n_153;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_260;
wire n_298;
wire n_320;
wire n_286;
wire n_122;
wire n_282;
wire n_331;
wire n_406;
wire n_325;
wire n_132;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_371;
wire n_152;
wire n_317;
wire n_323;
wire n_195;
wire n_356;
wire n_227;
wire n_271;
wire n_335;
wire n_123;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_267;
wire n_297;
wire n_156;
wire n_225;
wire n_377;
wire n_219;
wire n_157;
wire n_131;
wire n_192;
wire n_223;
wire n_392;
wire n_158;
wire n_138;
wire n_264;
wire n_109;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_185;
wire n_183;
wire n_243;
wire n_398;
wire n_396;
wire n_347;
wire n_169;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_290;
wire n_221;
wire n_178;
wire n_386;
wire n_287;
wire n_344;
wire n_422;
wire n_415;
wire n_141;
wire n_355;
wire n_336;
wire n_145;
wire n_337;
wire n_313;
wire n_216;
wire n_168;
wire n_395;
wire n_164;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_328;
wire n_140;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_241;
wire n_357;
wire n_184;
wire n_144;
wire n_114;
wire n_165;
wire n_213;
wire n_129;
wire n_342;
wire n_361;
wire n_363;
wire n_402;
wire n_413;
wire n_197;
wire n_107;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_384;
wire n_277;
wire n_338;
wire n_149;
wire n_333;
wire n_309;
wire n_130;
wire n_322;
wire n_258;
wire n_151;
wire n_306;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_112;
wire n_239;
wire n_420;
wire n_310;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_270;
wire n_230;
wire n_118;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_206;
wire n_172;
wire n_217;
wire n_312;
wire n_345;
wire n_210;
wire n_365;
wire n_176;
wire n_182;
wire n_143;
wire n_354;
wire n_237;
wire n_425;
wire n_407;
wire n_180;
wire n_340;
wire n_207;
wire n_346;
wire n_393;
wire n_229;
wire n_108;
wire n_177;
wire n_403;
wire n_421;
wire n_405;
wire n_359;
wire n_117;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_113;
wire n_246;
wire n_179;
wire n_125;
wire n_410;
wire n_269;
wire n_128;
wire n_285;
wire n_412;
wire n_120;
wire n_232;
wire n_327;
wire n_135;
wire n_126;
wire n_202;
wire n_266;
wire n_272;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_409;
wire n_154;
wire n_148;
wire n_300;
wire n_159;
wire n_334;
wire n_391;
wire n_175;
wire n_262;
wire n_238;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_121;
wire n_242;
wire n_360;
wire n_200;
wire n_162;
wire n_222;
wire n_115;
wire n_324;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_424;
wire n_256;
wire n_305;
wire n_278;
wire n_110;

INVx1_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

CKINVDCx5p33_ASAP7_75t_R g108 ( 
.A(n_2),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_28),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

NOR2xp67_ASAP7_75t_L g111 ( 
.A(n_44),
.B(n_54),
.Y(n_111)
);

CKINVDCx5p33_ASAP7_75t_R g112 ( 
.A(n_84),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_42),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_21),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_22),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_19),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_64),
.Y(n_122)
);

INVxp33_ASAP7_75t_SL g123 ( 
.A(n_27),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_40),
.Y(n_124)
);

INVxp33_ASAP7_75t_SL g125 ( 
.A(n_45),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_33),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_23),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_89),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_3),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_24),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_26),
.Y(n_134)
);

INVxp33_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_16),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_11),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_56),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_5),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_52),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_15),
.Y(n_143)
);

INVxp33_ASAP7_75t_SL g144 ( 
.A(n_32),
.Y(n_144)
);

INVxp33_ASAP7_75t_SL g145 ( 
.A(n_51),
.Y(n_145)
);

INVxp33_ASAP7_75t_SL g146 ( 
.A(n_35),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_46),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_53),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_68),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_3),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_1),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_37),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_81),
.Y(n_154)
);

INVxp67_ASAP7_75t_SL g155 ( 
.A(n_29),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_10),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_41),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_93),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_73),
.Y(n_159)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_94),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_1),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_95),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

INVxp67_ASAP7_75t_SL g164 ( 
.A(n_66),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_12),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_39),
.Y(n_166)
);

INVxp67_ASAP7_75t_SL g167 ( 
.A(n_100),
.Y(n_167)
);

INVxp67_ASAP7_75t_SL g168 ( 
.A(n_36),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_75),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_7),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_77),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_30),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_79),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_7),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_20),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_124),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_0),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

OAI21x1_ASAP7_75t_L g182 ( 
.A1(n_128),
.A2(n_139),
.B(n_176),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_124),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_141),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_128),
.B(n_0),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_129),
.B(n_4),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_165),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_106),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_129),
.B(n_4),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_107),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_110),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_108),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_113),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_114),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_115),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_116),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_117),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_118),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_120),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_161),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_121),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_135),
.B(n_5),
.Y(n_211)
);

AND2x4_ASAP7_75t_L g212 ( 
.A(n_140),
.B(n_6),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

AND2x4_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_174),
.Y(n_214)
);

AND2x4_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_155),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_142),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_199),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_135),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

AND2x4_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_155),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

AND2x4_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_164),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_177),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_177),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_211),
.A2(n_109),
.B1(n_122),
.B2(n_160),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_177),
.Y(n_228)
);

INVx8_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_183),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_211),
.A2(n_146),
.B1(n_123),
.B2(n_125),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_183),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_203),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_187),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_188),
.B(n_190),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_187),
.Y(n_238)
);

BUFx10_ASAP7_75t_L g239 ( 
.A(n_191),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_191),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_191),
.Y(n_241)
);

AND2x6_ASAP7_75t_L g242 ( 
.A(n_188),
.B(n_126),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_195),
.B(n_160),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_195),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_185),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_184),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_181),
.A2(n_145),
.B1(n_144),
.B2(n_119),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_195),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_194),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_197),
.Y(n_250)
);

A2O1A1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_218),
.A2(n_182),
.B(n_208),
.C(n_207),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_215),
.B(n_202),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_216),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_190),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_247),
.A2(n_222),
.B1(n_215),
.B2(n_242),
.Y(n_256)
);

NOR2x1_ASAP7_75t_R g257 ( 
.A(n_221),
.B(n_164),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_204),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_205),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_226),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_242),
.A2(n_198),
.B1(n_206),
.B2(n_210),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_225),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_193),
.Y(n_263)
);

BUFx5_ASAP7_75t_L g264 ( 
.A(n_217),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_224),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_233),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_229),
.B(n_196),
.Y(n_267)
);

OR2x2_ASAP7_75t_SL g268 ( 
.A(n_238),
.B(n_198),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_229),
.B(n_196),
.Y(n_269)
);

OR2x6_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_181),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_214),
.B(n_167),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_226),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_231),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_231),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_226),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_228),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_214),
.B(n_167),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_239),
.Y(n_278)
);

AND2x6_ASAP7_75t_L g279 ( 
.A(n_219),
.B(n_127),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_235),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_220),
.B(n_168),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_235),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_235),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_239),
.B(n_112),
.Y(n_284)
);

AND2x4_ASAP7_75t_L g285 ( 
.A(n_240),
.B(n_178),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_223),
.A2(n_230),
.B1(n_234),
.B2(n_237),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_240),
.B(n_244),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_240),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_244),
.B(n_168),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_260),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_265),
.A2(n_213),
.B(n_245),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_262),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_285),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_285),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_254),
.A2(n_157),
.B1(n_131),
.B2(n_133),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_266),
.Y(n_296)
);

AND2x4_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_244),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_253),
.A2(n_256),
.B1(n_261),
.B2(n_277),
.Y(n_298)
);

AND2x4_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_248),
.Y(n_299)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_288),
.Y(n_300)
);

NOR2x1_ASAP7_75t_SL g301 ( 
.A(n_259),
.B(n_134),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_257),
.Y(n_302)
);

A2O1A1Ixp33_ASAP7_75t_L g303 ( 
.A1(n_251),
.A2(n_111),
.B(n_159),
.C(n_163),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_289),
.Y(n_304)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_287),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_271),
.A2(n_162),
.B1(n_136),
.B2(n_138),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_252),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_270),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_263),
.B(n_246),
.Y(n_309)
);

BUFx4_ASAP7_75t_SL g310 ( 
.A(n_278),
.Y(n_310)
);

CKINVDCx8_ASAP7_75t_R g311 ( 
.A(n_270),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_264),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_264),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_250),
.B(n_246),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_258),
.A2(n_213),
.B(n_245),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_255),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_268),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_276),
.Y(n_318)
);

OR2x6_ASAP7_75t_L g319 ( 
.A(n_281),
.B(n_186),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_260),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_279),
.A2(n_153),
.B1(n_143),
.B2(n_147),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_279),
.A2(n_166),
.B1(n_148),
.B2(n_149),
.Y(n_322)
);

AND2x4_ASAP7_75t_L g323 ( 
.A(n_280),
.B(n_248),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_264),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_267),
.A2(n_169),
.B(n_150),
.Y(n_325)
);

CKINVDCx11_ASAP7_75t_R g326 ( 
.A(n_311),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_307),
.A2(n_269),
.B1(n_279),
.B2(n_274),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_292),
.Y(n_328)
);

O2A1O1Ixp33_ASAP7_75t_SL g329 ( 
.A1(n_303),
.A2(n_170),
.B(n_172),
.C(n_173),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_292),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_290),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_294),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_293),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_298),
.B(n_264),
.Y(n_334)
);

OAI21x1_ASAP7_75t_L g335 ( 
.A1(n_291),
.A2(n_286),
.B(n_284),
.Y(n_335)
);

OA21x2_ASAP7_75t_L g336 ( 
.A1(n_325),
.A2(n_189),
.B(n_192),
.Y(n_336)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_290),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_304),
.B(n_273),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_317),
.Y(n_339)
);

OAI221xp5_ASAP7_75t_L g340 ( 
.A1(n_295),
.A2(n_130),
.B1(n_248),
.B2(n_282),
.C(n_283),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_309),
.B(n_282),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_290),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_308),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g344 ( 
.A(n_317),
.B(n_283),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_300),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_314),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_305),
.A2(n_55),
.B1(n_104),
.B2(n_102),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_296),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_315),
.B(n_319),
.Y(n_349)
);

NOR2x1_ASAP7_75t_SL g350 ( 
.A(n_312),
.B(n_13),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_316),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_300),
.A2(n_14),
.B1(n_17),
.B2(n_18),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_318),
.Y(n_353)
);

AO21x2_ASAP7_75t_L g354 ( 
.A1(n_334),
.A2(n_301),
.B(n_324),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_L g355 ( 
.A1(n_348),
.A2(n_306),
.B1(n_319),
.B2(n_321),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_346),
.A2(n_306),
.B1(n_322),
.B2(n_321),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_341),
.B(n_302),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_339),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_334),
.A2(n_313),
.B1(n_322),
.B2(n_320),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_349),
.A2(n_338),
.B(n_335),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_346),
.A2(n_297),
.B1(n_299),
.B2(n_323),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_348),
.A2(n_320),
.B(n_297),
.Y(n_362)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_344),
.Y(n_363)
);

AOI222xp33_ASAP7_75t_L g364 ( 
.A1(n_339),
.A2(n_323),
.B1(n_299),
.B2(n_320),
.C1(n_310),
.C2(n_25),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_333),
.Y(n_365)
);

AND2x4_ASAP7_75t_L g366 ( 
.A(n_351),
.B(n_31),
.Y(n_366)
);

OAI21x1_ASAP7_75t_SL g367 ( 
.A1(n_350),
.A2(n_34),
.B(n_43),
.Y(n_367)
);

OAI221xp5_ASAP7_75t_L g368 ( 
.A1(n_327),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.C(n_50),
.Y(n_368)
);

OAI21xp33_ASAP7_75t_L g369 ( 
.A1(n_356),
.A2(n_353),
.B(n_332),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_328),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_358),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_363),
.Y(n_372)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_366),
.Y(n_373)
);

AOI221xp5_ASAP7_75t_L g374 ( 
.A1(n_356),
.A2(n_343),
.B1(n_329),
.B2(n_347),
.C(n_340),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_365),
.B(n_330),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_361),
.B(n_352),
.Y(n_376)
);

O2A1O1Ixp5_ASAP7_75t_L g377 ( 
.A1(n_360),
.A2(n_337),
.B(n_329),
.C(n_336),
.Y(n_377)
);

OAI211xp5_ASAP7_75t_L g378 ( 
.A1(n_364),
.A2(n_326),
.B(n_345),
.C(n_337),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_362),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_359),
.Y(n_380)
);

OAI22xp33_ASAP7_75t_L g381 ( 
.A1(n_368),
.A2(n_331),
.B1(n_342),
.B2(n_336),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_355),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_375),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_382),
.B(n_354),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_369),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_380),
.Y(n_386)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_373),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_376),
.B(n_361),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g389 ( 
.A(n_372),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_378),
.A2(n_367),
.B1(n_342),
.B2(n_331),
.Y(n_390)
);

OAI33xp33_ASAP7_75t_L g391 ( 
.A1(n_381),
.A2(n_342),
.A3(n_331),
.B1(n_61),
.B2(n_62),
.B3(n_63),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_373),
.B(n_59),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_370),
.B(n_105),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_379),
.A2(n_60),
.B(n_65),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_374),
.B(n_67),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_386),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_386),
.B(n_371),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_384),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_393),
.B(n_69),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_384),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_388),
.B(n_395),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_385),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_388),
.B(n_377),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_389),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_383),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_395),
.B(n_71),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_392),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_402),
.B(n_390),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_397),
.B(n_401),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_396),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_409),
.B(n_405),
.Y(n_411)
);

AO211x2_ASAP7_75t_L g412 ( 
.A1(n_408),
.A2(n_406),
.B(n_407),
.C(n_397),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_411),
.Y(n_413)
);

XNOR2x2_ASAP7_75t_L g414 ( 
.A(n_412),
.B(n_408),
.Y(n_414)
);

OAI322xp33_ASAP7_75t_L g415 ( 
.A1(n_414),
.A2(n_398),
.A3(n_410),
.B1(n_400),
.B2(n_404),
.C1(n_403),
.C2(n_396),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_413),
.Y(n_416)
);

NOR3xp33_ASAP7_75t_L g417 ( 
.A(n_415),
.B(n_399),
.C(n_391),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_416),
.A2(n_394),
.B(n_400),
.Y(n_418)
);

NOR3xp33_ASAP7_75t_L g419 ( 
.A(n_418),
.B(n_387),
.C(n_72),
.Y(n_419)
);

NOR3xp33_ASAP7_75t_L g420 ( 
.A(n_417),
.B(n_387),
.C(n_74),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_420),
.Y(n_421)
);

NOR3x1_ASAP7_75t_L g422 ( 
.A(n_421),
.B(n_419),
.C(n_78),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_422),
.B(n_88),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_423),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_424),
.B(n_90),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_425),
.A2(n_99),
.B(n_96),
.Y(n_426)
);


endmodule