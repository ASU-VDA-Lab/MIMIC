module fake_jpeg_15324_n_137 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

INVx11_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_9),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_25),
.B(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_27),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx2_ASAP7_75t_SL g28 ( 
.A(n_11),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_13),
.B(n_0),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_19),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_15),
.B1(n_21),
.B2(n_20),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_30),
.B1(n_11),
.B2(n_23),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_20),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_SL g52 ( 
.A(n_33),
.B(n_18),
.C(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_14),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_20),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_18),
.B(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_42),
.A2(n_39),
.B1(n_23),
.B2(n_35),
.Y(n_72)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_46),
.B(n_52),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_48),
.B(n_50),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_14),
.Y(n_50)
);

AND2x6_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_0),
.Y(n_51)
);

AND2x6_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_1),
.Y(n_66)
);

CKINVDCx10_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_55),
.Y(n_64)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_56),
.B(n_16),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_58),
.Y(n_65)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_68),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_33),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_63),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_32),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_72),
.B1(n_15),
.B2(n_32),
.Y(n_79)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_38),
.C(n_36),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_36),
.C(n_19),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_58),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_38),
.Y(n_74)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_10),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_78),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_59),
.B1(n_24),
.B2(n_72),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_73),
.A2(n_51),
.B1(n_66),
.B2(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_85),
.Y(n_103)
);

A2O1A1O1Ixp25_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_52),
.B(n_40),
.C(n_48),
.D(n_54),
.Y(n_82)
);

NAND3xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_71),
.C(n_69),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_83),
.B(n_84),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_70),
.B(n_55),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_67),
.C(n_27),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_44),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_88),
.B(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_24),
.Y(n_90)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

XNOR2x1_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_90),
.Y(n_111)
);

NAND3xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_69),
.C(n_61),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_95),
.Y(n_109)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_81),
.C(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_98),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_87),
.C(n_80),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_59),
.B1(n_68),
.B2(n_21),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_27),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_108),
.C(n_110),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_106),
.B(n_101),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_86),
.C(n_78),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_104),
.C(n_102),
.Y(n_110)
);

AOI321xp33_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_77),
.A3(n_97),
.B1(n_83),
.B2(n_19),
.C(n_26),
.Y(n_118)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_112),
.Y(n_115)
);

FAx1_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_96),
.CI(n_99),
.CON(n_114),
.SN(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_110),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_93),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_105),
.C(n_108),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_118),
.A2(n_107),
.B(n_106),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_1),
.B(n_2),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_SL g129 ( 
.A1(n_122),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_119),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_112),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_124),
.B(n_21),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_128),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_120),
.A2(n_21),
.B1(n_109),
.B2(n_19),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_L g130 ( 
.A1(n_126),
.A2(n_123),
.A3(n_26),
.B1(n_6),
.B2(n_8),
.C1(n_9),
.C2(n_5),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_129),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_130),
.A2(n_5),
.B1(n_6),
.B2(n_131),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_4),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_5),
.Y(n_134)
);

AO21x1_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_135),
.B(n_133),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_133),
.Y(n_137)
);


endmodule