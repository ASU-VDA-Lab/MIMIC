module fake_netlist_6_535_n_16688 (n_992, n_2542, n_1671, n_1, n_2817, n_3660, n_3813, n_801, n_3766, n_1613, n_1234, n_1458, n_2576, n_3254, n_3684, n_1199, n_1674, n_3392, n_741, n_1027, n_1351, n_3266, n_3574, n_625, n_1189, n_3152, n_223, n_4154, n_3579, n_1212, n_226, n_208, n_68, n_4251, n_726, n_2157, n_3335, n_2332, n_212, n_3773, n_700, n_3783, n_4177, n_50, n_1307, n_3178, n_2003, n_3849, n_4127, n_1038, n_578, n_1581, n_1003, n_365, n_3844, n_168, n_1237, n_1061, n_2353, n_2534, n_3089, n_3301, n_4099, n_1357, n_4241, n_1853, n_3741, n_77, n_4168, n_783, n_2451, n_1738, n_2243, n_798, n_188, n_1575, n_1854, n_2324, n_3088, n_3443, n_1923, n_3257, n_509, n_1342, n_245, n_1209, n_1348, n_1387, n_2260, n_3222, n_677, n_1708, n_805, n_1151, n_396, n_2977, n_3952, n_1739, n_350, n_78, n_2051, n_2317, n_1380, n_3911, n_2359, n_442, n_480, n_142, n_2847, n_1402, n_2557, n_1688, n_1691, n_3332, n_4134, n_4285, n_3465, n_1975, n_1009, n_1743, n_62, n_1930, n_2405, n_3706, n_4050, n_1160, n_883, n_2647, n_1238, n_1991, n_2570, n_2179, n_2386, n_2997, n_4092, n_1724, n_1032, n_3708, n_2336, n_1247, n_3668, n_4078, n_1547, n_2521, n_3376, n_3046, n_2956, n_1553, n_893, n_1099, n_2491, n_3801, n_4249, n_1264, n_1192, n_471, n_3564, n_1844, n_424, n_3619, n_4087, n_1700, n_1555, n_1415, n_2211, n_1370, n_1786, n_3487, n_369, n_4198, n_287, n_2382, n_3754, n_2672, n_3030, n_4302, n_2291, n_415, n_830, n_2299, n_65, n_230, n_3340, n_4179, n_461, n_873, n_141, n_383, n_1285, n_1371, n_2886, n_2974, n_3946, n_200, n_1985, n_4213, n_2989, n_447, n_2838, n_2184, n_3395, n_2982, n_1803, n_3427, n_1172, n_852, n_2509, n_4065, n_4026, n_71, n_229, n_2513, n_3282, n_1590, n_2645, n_1532, n_2313, n_2628, n_3071, n_3626, n_3757, n_3904, n_4178, n_1393, n_1517, n_1867, n_2926, n_1704, n_1078, n_250, n_544, n_1711, n_2247, n_3106, n_1140, n_2630, n_4273, n_1444, n_1670, n_1603, n_2344, n_1579, n_3275, n_35, n_2365, n_2470, n_2321, n_1263, n_2019, n_3031, n_4029, n_836, n_3345, n_375, n_2074, n_2447, n_522, n_2919, n_3678, n_3440, n_2129, n_2340, n_1261, n_945, n_3879, n_4010, n_2286, n_1649, n_2018, n_2094, n_3080, n_1903, n_1511, n_1143, n_2356, n_2399, n_1422, n_1232, n_1772, n_1572, n_3979, n_616, n_658, n_4308, n_1874, n_3165, n_1119, n_2865, n_2825, n_3463, n_2013, n_428, n_1433, n_1902, n_1842, n_1620, n_2044, n_1954, n_1735, n_2510, n_1541, n_1300, n_641, n_2480, n_2739, n_3023, n_822, n_3232, n_693, n_1313, n_2791, n_3607, n_3750, n_3251, n_1056, n_3877, n_3316, n_2212, n_3929, n_758, n_516, n_3494, n_3048, n_1455, n_2418, n_2864, n_1163, n_2729, n_3063, n_4311, n_1180, n_2256, n_2582, n_943, n_1798, n_4060, n_1550, n_2703, n_491, n_3998, n_2786, n_3371, n_1591, n_42, n_772, n_3632, n_3122, n_2806, n_1344, n_3261, n_2730, n_2495, n_666, n_371, n_4187, n_940, n_770, n_567, n_1781, n_1971, n_2058, n_2090, n_2603, n_405, n_213, n_2660, n_538, n_3028, n_3829, n_3662, n_2981, n_3076, n_2173, n_4164, n_2004, n_1106, n_886, n_1471, n_343, n_953, n_1094, n_3624, n_3077, n_3737, n_1345, n_1820, n_2873, n_3452, n_3655, n_494, n_539, n_493, n_3107, n_155, n_3825, n_2880, n_3225, n_2394, n_2108, n_3532, n_45, n_4117, n_454, n_3948, n_1421, n_2836, n_3664, n_1936, n_638, n_1404, n_1211, n_2124, n_381, n_2378, n_887, n_1660, n_1961, n_3047, n_112, n_1280, n_3765, n_713, n_2655, n_4125, n_1400, n_2625, n_3296, n_2843, n_126, n_4221, n_1467, n_3297, n_4250, n_58, n_976, n_3760, n_3067, n_2155, n_3906, n_224, n_2686, n_48, n_1445, n_2364, n_2551, n_1526, n_1560, n_734, n_1088, n_4262, n_1894, n_196, n_1231, n_2996, n_2599, n_2985, n_1978, n_3803, n_2085, n_3963, n_3368, n_917, n_574, n_3639, n_9, n_3347, n_2370, n_2612, n_3792, n_907, n_4202, n_6, n_1446, n_14, n_3938, n_2591, n_3507, n_659, n_1815, n_2214, n_3351, n_4253, n_407, n_913, n_4110, n_1658, n_2593, n_808, n_867, n_4071, n_4255, n_3506, n_4268, n_3568, n_3269, n_4047, n_3531, n_1230, n_3413, n_3850, n_473, n_1193, n_1967, n_3999, n_1054, n_3928, n_559, n_3412, n_2613, n_3535, n_1333, n_2496, n_44, n_2708, n_3313, n_1648, n_3189, n_1911, n_1956, n_163, n_1644, n_3791, n_4139, n_2011, n_2725, n_2277, n_3164, n_1558, n_1732, n_281, n_551, n_699, n_1986, n_2300, n_3943, n_4320, n_4305, n_564, n_2397, n_3884, n_3931, n_451, n_824, n_279, n_686, n_4102, n_4297, n_757, n_594, n_1641, n_2113, n_1918, n_2190, n_3603, n_3871, n_2907, n_577, n_3438, n_166, n_2735, n_4141, n_1843, n_619, n_3959, n_2268, n_1367, n_1336, n_521, n_2778, n_4227, n_2850, n_572, n_4314, n_395, n_813, n_1909, n_2080, n_1481, n_3822, n_323, n_4163, n_606, n_1441, n_818, n_3373, n_1123, n_1309, n_92, n_2104, n_513, n_645, n_1381, n_2961, n_3812, n_331, n_1699, n_3910, n_916, n_3934, n_2093, n_4033, n_4296, n_4009, n_2633, n_483, n_102, n_3883, n_2207, n_1970, n_2770, n_608, n_261, n_2101, n_2696, n_3482, n_4080, n_630, n_2059, n_32, n_2198, n_3319, n_541, n_512, n_2669, n_2925, n_3728, n_4094, n_2073, n_2273, n_121, n_3484, n_433, n_3748, n_2546, n_3272, n_3193, n_792, n_2522, n_476, n_3949, n_2792, n_2, n_1328, n_3396, n_1957, n_2917, n_219, n_2616, n_3912, n_3118, n_3315, n_3720, n_1907, n_3923, n_2529, n_264, n_263, n_3900, n_1162, n_860, n_1530, n_3798, n_788, n_939, n_3488, n_1543, n_821, n_2811, n_938, n_1302, n_1068, n_1599, n_3732, n_329, n_982, n_4257, n_2674, n_2832, n_4226, n_549, n_1762, n_1910, n_1075, n_3980, n_408, n_932, n_2831, n_2998, n_4318, n_3446, n_4158, n_61, n_3317, n_237, n_3857, n_3978, n_1876, n_4107, n_1895, n_2123, n_1697, n_2143, n_243, n_979, n_4074, n_3716, n_1873, n_4294, n_905, n_3630, n_3518, n_3824, n_3859, n_1866, n_4013, n_1680, n_117, n_175, n_322, n_993, n_2692, n_3842, n_689, n_3248, n_2031, n_354, n_2130, n_1330, n_1413, n_1605, n_3714, n_3514, n_2228, n_3914, n_3397, n_134, n_1988, n_2941, n_1278, n_547, n_3575, n_2455, n_2876, n_558, n_2654, n_3036, n_2469, n_4032, n_1064, n_3099, n_1396, n_634, n_2355, n_3927, n_4147, n_136, n_966, n_3888, n_2908, n_3168, n_764, n_2751, n_2764, n_3357, n_1663, n_4130, n_4161, n_2895, n_2009, n_4172, n_692, n_3403, n_733, n_1793, n_2922, n_3601, n_3882, n_1233, n_1289, n_2714, n_2245, n_487, n_3055, n_3092, n_3492, n_3895, n_241, n_3966, n_30, n_2068, n_1107, n_2866, n_2457, n_3294, n_4119, n_1014, n_3734, n_3686, n_1290, n_1703, n_2580, n_3455, n_4118, n_882, n_2176, n_2072, n_3649, n_1354, n_2821, n_586, n_423, n_1865, n_1875, n_1701, n_2459, n_318, n_3746, n_1111, n_1713, n_2971, n_715, n_3599, n_2678, n_1251, n_3384, n_3935, n_1265, n_4277, n_2711, n_3490, n_4291, n_88, n_4199, n_1726, n_1950, n_530, n_1563, n_1912, n_277, n_2434, n_4319, n_3369, n_3419, n_1982, n_3872, n_2878, n_618, n_3012, n_1297, n_1662, n_1312, n_3772, n_3875, n_199, n_1167, n_1359, n_2818, n_2428, n_3581, n_3794, n_674, n_3247, n_871, n_3069, n_3921, n_922, n_268, n_1335, n_1760, n_1927, n_210, n_2028, n_3715, n_1069, n_2664, n_5, n_1664, n_1722, n_612, n_2641, n_3022, n_3052, n_3725, n_178, n_247, n_1165, n_355, n_3933, n_702, n_347, n_2008, n_2749, n_3298, n_2192, n_3281, n_2254, n_2345, n_3346, n_1926, n_1175, n_3273, n_328, n_1386, n_2311, n_1896, n_429, n_2965, n_1747, n_3058, n_1012, n_195, n_3691, n_780, n_3861, n_675, n_2624, n_4066, n_903, n_4146, n_1540, n_1977, n_1802, n_1504, n_3549, n_2350, n_2804, n_2453, n_286, n_254, n_3891, n_2193, n_3961, n_2676, n_1655, n_3940, n_4072, n_4220, n_242, n_835, n_1214, n_928, n_47, n_690, n_850, n_1801, n_1886, n_2092, n_2347, n_1654, n_816, n_1157, n_3453, n_1750, n_2994, n_1462, n_3410, n_3153, n_3428, n_1188, n_3689, n_1752, n_877, n_1813, n_2514, n_3768, n_2206, n_604, n_4004, n_2810, n_2967, n_2319, n_2519, n_4043, n_825, n_4313, n_728, n_2916, n_3415, n_1063, n_4292, n_1588, n_3785, n_3942, n_3997, n_2963, n_4041, n_2947, n_3918, n_2467, n_26, n_2602, n_2468, n_55, n_267, n_3145, n_1124, n_1624, n_3873, n_3983, n_515, n_2096, n_2980, n_3968, n_1965, n_3538, n_2476, n_3280, n_598, n_3434, n_696, n_1515, n_961, n_3510, n_437, n_1082, n_1317, n_3227, n_2733, n_2824, n_3289, n_593, n_4169, n_514, n_4055, n_687, n_697, n_890, n_637, n_2377, n_295, n_701, n_2178, n_3271, n_950, n_4248, n_388, n_190, n_2812, n_484, n_2644, n_2036, n_3326, n_2976, n_2152, n_1709, n_3009, n_2652, n_4200, n_3460, n_2411, n_3719, n_2525, n_1825, n_2393, n_1757, n_1796, n_170, n_2657, n_1792, n_3827, n_891, n_2067, n_2136, n_2921, n_2409, n_2082, n_3519, n_2252, n_1412, n_2497, n_3889, n_2687, n_3237, n_949, n_1630, n_678, n_2887, n_3809, n_3500, n_3834, n_4245, n_4136, n_3526, n_3707, n_283, n_2075, n_4045, n_2194, n_2972, n_2619, n_3139, n_3542, n_91, n_2763, n_2762, n_4070, n_1987, n_3545, n_507, n_968, n_909, n_1369, n_3578, n_3885, n_881, n_2271, n_1008, n_3192, n_760, n_3993, n_1546, n_2583, n_590, n_4116, n_63, n_2606, n_4031, n_362, n_148, n_2279, n_161, n_22, n_462, n_1033, n_1052, n_2794, n_1296, n_2663, n_1990, n_3352, n_2391, n_3805, n_304, n_2431, n_3073, n_4018, n_2987, n_694, n_2938, n_2150, n_1294, n_2943, n_1420, n_3696, n_3780, n_4082, n_125, n_1634, n_2078, n_3252, n_2932, n_297, n_595, n_627, n_1767, n_1779, n_524, n_1465, n_3253, n_3337, n_3431, n_342, n_3209, n_3450, n_2622, n_1858, n_1044, n_4002, n_2658, n_2665, n_2165, n_2133, n_1712, n_3021, n_1391, n_449, n_131, n_1523, n_2558, n_2750, n_2775, n_1208, n_2893, n_1164, n_1295, n_1627, n_2954, n_3477, n_4288, n_2728, n_2349, n_3128, n_3763, n_4289, n_2684, n_2712, n_1072, n_3146, n_1527, n_1495, n_3733, n_1438, n_495, n_815, n_3953, n_1100, n_585, n_1487, n_2691, n_3421, n_840, n_2913, n_3614, n_874, n_1756, n_3183, n_1128, n_2493, n_382, n_673, n_2230, n_2705, n_1969, n_4019, n_2690, n_1071, n_1067, n_1565, n_1493, n_2145, n_3405, n_1968, n_898, n_255, n_284, n_1952, n_865, n_3616, n_4228, n_2573, n_3423, n_2646, n_4044, n_3436, n_925, n_1932, n_1101, n_15, n_1026, n_1880, n_2535, n_3366, n_3442, n_2631, n_4191, n_38, n_289, n_1364, n_3078, n_3644, n_2436, n_3937, n_615, n_2870, n_1249, n_2706, n_3838, n_59, n_4287, n_1293, n_2693, n_4137, n_1127, n_1512, n_2151, n_3159, n_1451, n_3941, n_320, n_108, n_639, n_963, n_794, n_2767, n_3793, n_727, n_894, n_1839, n_2341, n_685, n_1765, n_3727, n_353, n_2707, n_3240, n_3576, n_3789, n_605, n_1514, n_1863, n_826, n_3385, n_3747, n_3037, n_1646, n_3293, n_872, n_1139, n_1714, n_3922, n_86, n_3179, n_104, n_718, n_1018, n_3400, n_3729, n_1521, n_1366, n_4000, n_542, n_847, n_644, n_682, n_851, n_2537, n_2897, n_3970, n_305, n_72, n_2554, n_996, n_532, n_173, n_1308, n_2089, n_1376, n_3522, n_1513, n_2747, n_3924, n_413, n_3171, n_791, n_1913, n_4216, n_3608, n_510, n_837, n_4315, n_2097, n_79, n_2170, n_3459, n_4156, n_3491, n_4240, n_1488, n_2853, n_1808, n_3053, n_948, n_3358, n_2517, n_2713, n_3499, n_704, n_2148, n_4284, n_4162, n_977, n_2339, n_1005, n_1947, n_2765, n_2861, n_536, n_3158, n_1788, n_3426, n_1999, n_2731, n_622, n_147, n_2590, n_2643, n_3150, n_3018, n_3353, n_3782, n_3975, n_1469, n_2060, n_2608, n_1838, n_2638, n_4011, n_1835, n_3470, n_1766, n_1776, n_1959, n_3133, n_2002, n_581, n_2650, n_2138, n_4098, n_4021, n_765, n_432, n_987, n_1492, n_3700, n_2414, n_1340, n_3014, n_3166, n_1771, n_2316, n_4058, n_4103, n_3104, n_631, n_720, n_3435, n_153, n_842, n_3148, n_2262, n_3229, n_3348, n_4022, n_1707, n_2239, n_3082, n_3611, n_4310, n_1432, n_156, n_145, n_2208, n_843, n_656, n_989, n_2604, n_2407, n_1277, n_2816, n_797, n_2689, n_2933, n_1473, n_2191, n_1723, n_2717, n_1246, n_3799, n_1878, n_2574, n_899, n_189, n_738, n_2012, n_3497, n_1304, n_1035, n_294, n_2842, n_499, n_2675, n_1426, n_3418, n_705, n_3580, n_3775, n_11, n_3537, n_1004, n_1176, n_2134, n_1529, n_2335, n_2473, n_3887, n_1022, n_614, n_529, n_2069, n_2307, n_3704, n_2362, n_425, n_684, n_2539, n_2667, n_2698, n_4096, n_1431, n_4123, n_1615, n_4114, n_1474, n_3312, n_1571, n_3835, n_4286, n_1809, n_3119, n_4280, n_2948, n_1577, n_2958, n_3735, n_2297, n_1181, n_2119, n_3731, n_1822, n_37, n_486, n_947, n_2936, n_3224, n_1117, n_2489, n_1087, n_1448, n_3173, n_1992, n_3677, n_3631, n_648, n_657, n_1049, n_3223, n_3996, n_2771, n_2445, n_3020, n_2057, n_2103, n_3140, n_3185, n_3770, n_2605, n_4097, n_1666, n_2772, n_1505, n_803, n_290, n_4218, n_118, n_1717, n_926, n_1817, n_2449, n_927, n_3557, n_2610, n_3654, n_3129, n_3880, n_1849, n_2848, n_919, n_3685, n_2868, n_3620, n_1698, n_478, n_4100, n_2231, n_3609, n_929, n_107, n_3832, n_2520, n_1228, n_417, n_4264, n_2857, n_446, n_3693, n_3788, n_89, n_1568, n_1490, n_2372, n_777, n_1299, n_272, n_2896, n_526, n_3837, n_2718, n_3019, n_2639, n_3471, n_1183, n_1436, n_2898, n_2251, n_1384, n_69, n_3674, n_2494, n_2959, n_4079, n_2501, n_3203, n_3325, n_2238, n_293, n_4085, n_2368, n_53, n_458, n_1070, n_2403, n_3342, n_2837, n_4175, n_998, n_16, n_717, n_3200, n_1665, n_4306, n_3600, n_18, n_3259, n_2524, n_154, n_3167, n_1383, n_2460, n_4224, n_3390, n_3656, n_1178, n_98, n_2127, n_1424, n_2338, n_3324, n_3593, n_3341, n_3867, n_1073, n_1000, n_796, n_252, n_1195, n_3559, n_3025, n_2137, n_1626, n_3191, n_4005, n_1507, n_2482, n_184, n_552, n_3810, n_3546, n_2532, n_1358, n_1811, n_1388, n_3661, n_3006, n_216, n_4140, n_2481, n_3561, n_912, n_1857, n_3987, n_1519, n_2144, n_3056, n_745, n_1284, n_1604, n_2296, n_2424, n_3201, n_3633, n_3447, n_3971, n_1142, n_2849, n_716, n_1475, n_623, n_1048, n_1201, n_1398, n_884, n_1774, n_2354, n_2682, n_3032, n_3103, n_3638, n_2589, n_1395, n_2110, n_2199, n_2661, n_731, n_2877, n_1502, n_1659, n_1955, n_755, n_931, n_1021, n_3393, n_474, n_527, n_683, n_811, n_1207, n_2442, n_3627, n_312, n_1791, n_1368, n_66, n_3451, n_3480, n_1418, n_958, n_292, n_1250, n_100, n_3331, n_1137, n_3615, n_1897, n_2064, n_880, n_3072, n_3087, n_2053, n_3612, n_3505, n_2259, n_2121, n_2773, n_4222, n_2545, n_3540, n_3577, n_889, n_3509, n_2432, n_2710, n_150, n_1478, n_589, n_3606, n_1310, n_3142, n_3598, n_819, n_2966, n_2294, n_1363, n_2581, n_1334, n_1942, n_1966, n_3591, n_767, n_3641, n_1314, n_600, n_964, n_831, n_1837, n_2218, n_2788, n_477, n_3196, n_3590, n_2435, n_954, n_864, n_2504, n_2797, n_2623, n_1110, n_2213, n_1410, n_399, n_2389, n_1440, n_124, n_2132, n_2892, n_2063, n_4120, n_1382, n_1534, n_3892, n_1564, n_1736, n_4069, n_211, n_2748, n_4053, n_1483, n_3848, n_1834, n_2331, n_1372, n_231, n_2292, n_2860, n_3327, n_2330, n_40, n_3441, n_1457, n_505, n_1719, n_3534, n_3718, n_319, n_1339, n_1787, n_2701, n_2475, n_537, n_2511, n_3964, n_1993, n_2281, n_4167, n_1427, n_311, n_2416, n_2745, n_2617, n_2776, n_1466, n_10, n_403, n_1919, n_1080, n_723, n_1877, n_3144, n_3705, n_3211, n_3244, n_596, n_123, n_3909, n_3944, n_546, n_562, n_1141, n_1268, n_386, n_1939, n_2030, n_1769, n_1220, n_2323, n_1893, n_556, n_2784, n_2209, n_2301, n_3582, n_3605, n_162, n_3287, n_4223, n_2387, n_3322, n_1755, n_1602, n_2421, n_1136, n_3270, n_2618, n_2025, n_2357, n_2846, n_2464, n_3265, n_128, n_1125, n_3755, n_4042, n_970, n_3306, n_2488, n_3640, n_2224, n_1980, n_642, n_995, n_276, n_1159, n_2329, n_1092, n_3481, n_2237, n_3026, n_441, n_221, n_1060, n_1951, n_2250, n_3090, n_4299, n_444, n_3033, n_3724, n_146, n_1252, n_1784, n_3311, n_3571, n_1223, n_3913, n_303, n_4276, n_511, n_2990, n_3847, n_193, n_1286, n_1773, n_1775, n_2115, n_2410, n_2552, n_1053, n_3302, n_2374, n_416, n_1681, n_520, n_418, n_1093, n_113, n_1783, n_1533, n_1597, n_2929, n_2780, n_3226, n_3323, n_3364, n_4, n_4020, n_4176, n_266, n_296, n_2596, n_2274, n_3163, n_775, n_651, n_1153, n_439, n_1618, n_3407, n_217, n_518, n_1531, n_2828, n_1185, n_3856, n_453, n_4236, n_3425, n_215, n_2384, n_3894, n_4204, n_4261, n_1745, n_914, n_759, n_3479, n_3127, n_2724, n_1831, n_426, n_317, n_2585, n_2621, n_3623, n_1653, n_2352, n_1679, n_4063, n_1625, n_90, n_3986, n_4237, n_2601, n_2160, n_3454, n_54, n_1453, n_2146, n_4006, n_2226, n_2131, n_488, n_2502, n_2801, n_3646, n_497, n_2920, n_4015, n_773, n_3547, n_1901, n_3869, n_920, n_99, n_1374, n_2556, n_2648, n_3212, n_1315, n_1647, n_13, n_2575, n_2754, n_1224, n_2783, n_3753, n_2306, n_1614, n_1459, n_1892, n_3188, n_3742, n_1933, n_2462, n_1135, n_1169, n_1179, n_2889, n_3243, n_3683, n_401, n_4034, n_324, n_1617, n_4056, n_3260, n_3370, n_3386, n_3816, n_335, n_3960, n_1470, n_2550, n_463, n_3093, n_3175, n_3214, n_1243, n_3736, n_848, n_120, n_2732, n_301, n_2928, n_274, n_4206, n_1096, n_2249, n_1091, n_1917, n_2000, n_3862, n_4267, n_1580, n_2227, n_4247, n_2270, n_2822, n_1425, n_3169, n_36, n_4180, n_3205, n_1881, n_1267, n_1281, n_1806, n_3284, n_983, n_3109, n_2023, n_3354, n_427, n_2572, n_2204, n_1520, n_496, n_2720, n_3126, n_2159, n_906, n_1390, n_688, n_2289, n_1077, n_1733, n_2315, n_1419, n_2863, n_3299, n_3663, n_4132, n_351, n_2955, n_2995, n_259, n_1731, n_177, n_2158, n_2087, n_1855, n_1636, n_3051, n_1437, n_3360, n_2135, n_3956, n_3367, n_1645, n_1832, n_4001, n_385, n_1687, n_1439, n_2328, n_1323, n_2859, n_2202, n_858, n_2049, n_4149, n_1331, n_613, n_736, n_2627, n_501, n_956, n_960, n_2276, n_3234, n_3917, n_663, n_856, n_2803, n_2100, n_3314, n_3525, n_379, n_2993, n_778, n_1668, n_2777, n_1134, n_3016, n_3566, n_3688, n_3004, n_3202, n_2830, n_2781, n_3220, n_4003, n_410, n_1129, n_3870, n_4126, n_554, n_602, n_1696, n_2829, n_1995, n_1594, n_2181, n_3751, n_664, n_1869, n_171, n_2911, n_3625, n_3804, n_1764, n_169, n_4207, n_1429, n_2826, n_1610, n_3084, n_3429, n_4113, n_1889, n_2379, n_435, n_1905, n_2016, n_2343, n_793, n_326, n_587, n_3466, n_3554, n_1593, n_580, n_762, n_1030, n_1202, n_3901, n_1937, n_465, n_1790, n_1778, n_3749, n_1635, n_2942, n_4014, n_1079, n_341, n_2515, n_1744, n_828, n_2139, n_2142, n_4067, n_4252, n_607, n_316, n_419, n_28, n_1551, n_4028, n_4054, n_2448, n_1103, n_2875, n_3907, n_2555, n_4048, n_3338, n_144, n_4217, n_3586, n_3462, n_3756, n_2219, n_1203, n_3653, n_3636, n_2851, n_3406, n_820, n_2327, n_951, n_106, n_2201, n_725, n_952, n_3919, n_999, n_358, n_1254, n_160, n_2841, n_3349, n_2420, n_3722, n_186, n_2984, n_0, n_368, n_575, n_994, n_2263, n_3539, n_3291, n_2304, n_4024, n_1508, n_2487, n_732, n_974, n_2983, n_2240, n_392, n_2278, n_2656, n_2538, n_724, n_2597, n_2375, n_3113, n_3194, n_3250, n_1934, n_3276, n_1020, n_1042, n_628, n_1273, n_1434, n_1573, n_3981, n_4214, n_1728, n_3973, n_557, n_2756, n_3572, n_1871, n_349, n_3448, n_617, n_3886, n_845, n_807, n_2924, n_1036, n_3595, n_140, n_1138, n_3414, n_1661, n_1275, n_2884, n_485, n_1549, n_67, n_443, n_1510, n_892, n_768, n_3637, n_421, n_3120, n_1468, n_3991, n_2855, n_3651, n_1859, n_2102, n_3516, n_2563, n_3797, n_3926, n_238, n_1095, n_2024, n_1595, n_202, n_2156, n_3449, n_1718, n_1749, n_3474, n_1683, n_1916, n_2598, n_597, n_280, n_1270, n_2549, n_1187, n_610, n_4234, n_4304, n_1403, n_1669, n_1852, n_4101, n_3548, n_3767, n_1024, n_3864, n_4036, n_1768, n_2153, n_2544, n_2381, n_3670, n_3550, n_3974, n_198, n_1847, n_2052, n_3634, n_179, n_248, n_2302, n_517, n_4211, n_4182, n_1667, n_667, n_1206, n_3230, n_4016, n_621, n_1037, n_1397, n_3268, n_3236, n_1279, n_1115, n_750, n_901, n_1499, n_3592, n_468, n_2755, n_3141, n_923, n_504, n_1409, n_4230, n_1841, n_3839, n_2637, n_2823, n_1639, n_1623, n_183, n_1015, n_3967, n_1503, n_3112, n_2819, n_3195, n_466, n_2526, n_3041, n_4274, n_2423, n_1057, n_3277, n_3108, n_2548, n_603, n_991, n_2785, n_1657, n_4189, n_4270, n_235, n_4151, n_1126, n_2412, n_1997, n_3817, n_3417, n_2636, n_3131, n_340, n_710, n_1108, n_1818, n_2439, n_2404, n_1182, n_3730, n_1298, n_4124, n_3659, n_2559, n_2177, n_39, n_2595, n_3399, n_2088, n_3635, n_73, n_1611, n_785, n_4155, n_2740, n_746, n_4238, n_609, n_1601, n_3011, n_1960, n_2694, n_2061, n_3416, n_3648, n_1686, n_3498, n_2757, n_2337, n_2401, n_101, n_167, n_1356, n_1589, n_3042, n_3213, n_127, n_3820, n_2309, n_2900, n_2957, n_2607, n_1740, n_2737, n_3994, n_1497, n_2890, n_1168, n_1216, n_1943, n_3228, n_133, n_1320, n_2716, n_96, n_3249, n_3081, n_3657, n_2452, n_1430, n_3650, n_1316, n_1287, n_2722, n_1452, n_2854, n_3672, n_3010, n_2499, n_4152, n_3533, n_3043, n_1622, n_1586, n_2543, n_2264, n_3464, n_302, n_1694, n_380, n_1535, n_3137, n_3382, n_2486, n_3132, n_3560, n_137, n_3723, n_2571, n_3138, n_1596, n_3177, n_20, n_1190, n_1734, n_3172, n_397, n_2902, n_3217, n_1983, n_1938, n_2498, n_4219, n_122, n_2220, n_2577, n_34, n_1262, n_2472, n_218, n_1891, n_2171, n_1213, n_3238, n_70, n_2235, n_3529, n_4193, n_3570, n_3394, n_2988, n_3136, n_1350, n_1673, n_3828, n_2232, n_1715, n_172, n_3536, n_4109, n_4192, n_1443, n_1272, n_2392, n_2894, n_3424, n_3957, n_4038, n_2790, n_4131, n_239, n_2037, n_97, n_2808, n_3710, n_4159, n_4195, n_3784, n_2298, n_782, n_2326, n_1539, n_490, n_3594, n_220, n_809, n_1043, n_3819, n_4090, n_3040, n_1797, n_3279, n_1608, n_4165, n_986, n_2305, n_2120, n_80, n_1472, n_2050, n_2373, n_2164, n_2402, n_2225, n_1081, n_3628, n_4144, n_402, n_1870, n_352, n_2964, n_4174, n_1692, n_800, n_1084, n_1171, n_460, n_2169, n_3485, n_4077, n_2371, n_1827, n_1361, n_1864, n_2006, n_3402, n_1491, n_2187, n_3475, n_662, n_3501, n_374, n_1152, n_1840, n_1705, n_3905, n_450, n_3262, n_3544, n_4150, n_2904, n_4008, n_2244, n_4290, n_3013, n_3356, n_2586, n_1684, n_921, n_2446, n_1346, n_711, n_1642, n_579, n_1352, n_2789, n_3105, n_3210, n_2872, n_937, n_2257, n_3692, n_3845, n_1682, n_2017, n_370, n_1695, n_1828, n_2046, n_2272, n_2699, n_2200, n_3029, n_4258, n_650, n_3597, n_1046, n_2560, n_1940, n_1979, n_2760, n_2704, n_3329, n_1145, n_330, n_1121, n_1102, n_1963, n_2738, n_972, n_1405, n_2376, n_258, n_3826, n_1406, n_456, n_3790, n_3878, n_2766, n_1332, n_260, n_2670, n_313, n_2700, n_624, n_962, n_1041, n_2346, n_565, n_3134, n_3647, n_356, n_1569, n_3681, n_936, n_3045, n_3115, n_1883, n_3821, n_1288, n_4300, n_3318, n_1186, n_1062, n_885, n_896, n_83, n_3278, n_2342, n_2167, n_2084, n_2970, n_3676, n_2882, n_3666, n_3675, n_4017, n_4260, n_3320, n_2541, n_654, n_2940, n_411, n_2518, n_2458, n_152, n_1222, n_599, n_776, n_321, n_1823, n_2479, n_3050, n_3350, n_105, n_2782, n_3977, n_227, n_1974, n_3988, n_4122, n_2673, n_2456, n_1720, n_3476, n_2527, n_204, n_482, n_934, n_1637, n_2635, n_3307, n_3439, n_1407, n_1795, n_2768, n_3588, n_4135, n_2871, n_4209, n_4279, n_420, n_2688, n_1341, n_394, n_1456, n_1845, n_3858, n_4183, n_1489, n_4321, n_4298, n_164, n_2314, n_3502, n_23, n_942, n_3003, n_2798, n_2852, n_1524, n_4128, n_543, n_2229, n_1964, n_4133, n_2288, n_1920, n_2753, n_2099, n_1496, n_1271, n_3292, n_1545, n_4145, n_2007, n_3121, n_2039, n_3388, n_4271, n_1946, n_1355, n_4181, n_1225, n_3184, n_1544, n_1485, n_2258, n_325, n_1640, n_4040, n_804, n_464, n_1846, n_3437, n_3245, n_3075, n_2406, n_4111, n_533, n_2390, n_4007, n_806, n_3712, n_879, n_959, n_2310, n_2506, n_584, n_2141, n_2562, n_244, n_2642, n_4312, n_1343, n_1522, n_76, n_4239, n_2734, n_548, n_1782, n_94, n_282, n_2383, n_4184, n_2626, n_1676, n_833, n_1830, n_2351, n_1567, n_4037, n_523, n_1319, n_707, n_2986, n_345, n_1900, n_3930, n_3246, n_799, n_1548, n_3381, n_3044, n_3562, n_2973, n_1155, n_2536, n_3915, n_139, n_2196, n_41, n_2629, n_3665, n_273, n_1633, n_2195, n_3208, n_2809, n_3007, n_787, n_2172, n_3528, n_3489, n_2835, n_1416, n_1528, n_2820, n_2293, n_1146, n_3698, n_2021, n_3355, n_2454, n_2114, n_3074, n_3174, n_159, n_1086, n_1066, n_3102, n_1948, n_157, n_2125, n_2026, n_4215, n_1282, n_2561, n_550, n_3321, n_2567, n_2322, n_275, n_652, n_2154, n_2727, n_2962, n_3377, n_2939, n_560, n_1906, n_1484, n_2992, n_3305, n_1241, n_1321, n_1672, n_569, n_2533, n_3157, n_3530, n_4185, n_1758, n_3221, n_3267, n_3752, n_2283, n_2869, n_2422, n_1925, n_737, n_1318, n_1914, n_1235, n_3457, n_1229, n_2759, n_3517, n_2945, n_3061, n_3893, n_2361, n_306, n_1292, n_1373, n_21, n_3762, n_3469, n_3932, n_2266, n_2960, n_3958, n_3005, n_346, n_3, n_3985, n_2427, n_3151, n_3411, n_1029, n_4196, n_3779, n_1447, n_2388, n_3984, n_2056, n_790, n_2611, n_2901, n_138, n_3258, n_1706, n_4242, n_3389, n_1498, n_3143, n_2653, n_2417, n_4232, n_4190, n_3000, n_1210, n_49, n_299, n_1248, n_1556, n_902, n_333, n_2189, n_2680, n_4052, n_2246, n_1047, n_3149, n_3375, n_3899, n_4084, n_3558, n_1984, n_3365, n_2236, n_1385, n_3713, n_431, n_3379, n_3156, n_24, n_459, n_1269, n_1931, n_2083, n_2834, n_3207, n_502, n_2668, n_672, n_2441, n_1257, n_3008, n_1751, n_3401, n_2840, n_3197, n_3242, n_285, n_3939, n_1375, n_1941, n_3483, n_3613, n_3972, n_4153, n_85, n_2128, n_655, n_706, n_1045, n_1650, n_786, n_1794, n_1236, n_1962, n_1559, n_1725, n_1928, n_2398, n_3743, n_3855, n_1872, n_3091, n_4317, n_834, n_19, n_29, n_2695, n_4035, n_3818, n_75, n_4269, n_743, n_766, n_3124, n_430, n_1741, n_1325, n_1002, n_1746, n_4088, n_1949, n_3398, n_3761, n_3759, n_545, n_3524, n_2671, n_489, n_2761, n_2885, n_2793, n_2715, n_2888, n_1804, n_2923, n_3711, n_3776, n_4235, n_1727, n_251, n_2508, n_1019, n_636, n_4301, n_3511, n_2054, n_4143, n_4170, n_729, n_110, n_151, n_876, n_774, n_3744, n_3642, n_2845, n_1337, n_3097, n_660, n_2062, n_2041, n_2975, n_438, n_1477, n_1360, n_2839, n_1860, n_2856, n_1904, n_2874, n_1200, n_2070, n_2588, n_479, n_3814, n_1607, n_3781, n_1353, n_1777, n_1908, n_1454, n_2484, n_2348, n_2944, n_2614, n_2126, n_3831, n_869, n_1154, n_3308, n_1113, n_1600, n_2833, n_2253, n_2758, n_3843, n_2366, n_646, n_528, n_391, n_1098, n_3694, n_2937, n_1329, n_2045, n_817, n_2261, n_3687, n_2216, n_3589, n_2210, n_262, n_3602, n_187, n_897, n_846, n_3300, n_2978, n_2066, n_3543, n_841, n_1476, n_3621, n_2516, n_3391, n_1001, n_508, n_1800, n_2241, n_1050, n_1411, n_1463, n_2903, n_3777, n_2827, n_1177, n_3216, n_3458, n_332, n_3515, n_1150, n_4203, n_3808, n_1742, n_3190, n_1562, n_1690, n_398, n_1191, n_1826, n_566, n_1023, n_1882, n_2951, n_1076, n_1118, n_194, n_2949, n_3726, n_57, n_1007, n_1807, n_1929, n_1378, n_2369, n_855, n_1592, n_1759, n_2719, n_1814, n_1631, n_52, n_591, n_1377, n_3758, n_1879, n_256, n_853, n_440, n_695, n_3806, n_4081, n_1542, n_2587, n_3199, n_2931, n_875, n_209, n_367, n_680, n_3339, n_1678, n_2569, n_661, n_2400, n_1716, n_3866, n_278, n_3787, n_1256, n_3585, n_671, n_3565, n_1953, n_7, n_933, n_740, n_703, n_3343, n_3303, n_978, n_4157, n_2752, n_4173, n_384, n_3135, n_1976, n_4229, n_2905, n_1291, n_1217, n_3990, n_751, n_749, n_3865, n_1824, n_310, n_3954, n_1628, n_4073, n_1324, n_3890, n_1399, n_2122, n_2109, n_3629, n_1435, n_3920, n_969, n_988, n_2140, n_3503, n_3160, n_1065, n_2796, n_3255, n_2507, n_84, n_1401, n_2358, n_1255, n_568, n_3658, n_1516, n_143, n_1536, n_3846, n_180, n_2163, n_2186, n_3512, n_2029, n_2815, n_1204, n_3951, n_3034, n_823, n_1132, n_643, n_233, n_698, n_1074, n_1394, n_3569, n_1327, n_1326, n_739, n_400, n_955, n_337, n_3874, n_1379, n_2528, n_2814, n_214, n_246, n_2787, n_1338, n_1097, n_2969, n_2395, n_935, n_3027, n_781, n_789, n_1554, n_3231, n_4083, n_1130, n_3083, n_4212, n_2979, n_181, n_1810, n_182, n_2953, n_573, n_769, n_2380, n_676, n_327, n_4295, n_1120, n_832, n_1583, n_3049, n_1730, n_2295, n_555, n_389, n_814, n_2746, n_2946, n_1643, n_2020, n_2500, n_3430, n_2269, n_1729, n_669, n_2290, n_4225, n_4171, n_2048, n_3652, n_176, n_114, n_300, n_222, n_3830, n_3679, n_2005, n_747, n_3541, n_74, n_2565, n_4023, n_1389, n_1105, n_3117, n_721, n_1461, n_742, n_3432, n_535, n_691, n_3617, n_372, n_2076, n_2736, n_111, n_2883, n_3583, n_314, n_3860, n_1408, n_378, n_3851, n_3567, n_1196, n_4282, n_377, n_1598, n_3493, n_2935, n_4046, n_3807, n_863, n_3015, n_2175, n_601, n_2182, n_3774, n_338, n_2910, n_1283, n_2385, n_4112, n_918, n_748, n_506, n_1114, n_1785, n_56, n_763, n_1147, n_1848, n_360, n_1754, n_2149, n_3057, n_3154, n_3701, n_2396, n_1506, n_119, n_2584, n_1652, n_1812, n_957, n_1994, n_3473, n_895, n_866, n_1227, n_2450, n_2485, n_3739, n_2284, n_3898, n_3520, n_191, n_2566, n_387, n_2287, n_452, n_744, n_971, n_2702, n_3241, n_946, n_344, n_2906, n_761, n_1303, n_2769, n_3622, n_1205, n_2492, n_1258, n_3778, n_4095, n_2438, n_2914, n_1392, n_174, n_1173, n_1924, n_525, n_2463, n_3363, n_2881, n_1677, n_1116, n_611, n_1570, n_1702, n_1219, n_3551, n_3064, n_1780, n_3100, n_3897, n_3721, n_1689, n_8, n_2180, n_3372, n_2858, n_3062, n_2679, n_1174, n_3573, n_1944, n_1016, n_1347, n_4106, n_795, n_1501, n_3604, n_1221, n_3334, n_4027, n_1245, n_838, n_3215, n_3969, n_129, n_3336, n_647, n_4160, n_197, n_4231, n_844, n_17, n_448, n_2952, n_1017, n_3068, n_3853, n_2117, n_2234, n_4256, n_2779, n_2685, n_3823, n_1083, n_109, n_445, n_3553, n_1561, n_2741, n_3114, n_930, n_888, n_2275, n_1112, n_2465, n_2620, n_2081, n_2168, n_2568, n_234, n_2022, n_1945, n_2203, n_910, n_3811, n_1656, n_1721, n_1460, n_911, n_2112, n_2255, n_82, n_1464, n_27, n_236, n_653, n_1737, n_2430, n_1414, n_3486, n_4086, n_752, n_908, n_2649, n_2721, n_944, n_3556, n_2034, n_576, n_1028, n_3836, n_2106, n_472, n_2862, n_270, n_2265, n_2615, n_414, n_2683, n_1922, n_563, n_4068, n_2032, n_2744, n_4309, n_1011, n_2474, n_3703, n_1566, n_1215, n_2437, n_25, n_93, n_839, n_2444, n_2743, n_3962, n_708, n_1973, n_3181, n_2267, n_3456, n_3035, n_668, n_4166, n_626, n_990, n_1500, n_779, n_1537, n_1821, n_2205, n_3699, n_4243, n_3204, n_1104, n_854, n_1058, n_3378, n_4025, n_2312, n_498, n_3404, n_1122, n_870, n_904, n_1253, n_709, n_1266, n_366, n_2242, n_3362, n_3745, n_4059, n_1509, n_103, n_4188, n_3328, n_1693, n_2934, n_3667, n_3290, n_4121, n_1109, n_3523, n_185, n_2222, n_712, n_3256, n_348, n_1276, n_3802, n_3868, n_3176, n_376, n_3309, n_3671, n_2015, n_2118, n_4142, n_2111, n_2466, n_390, n_3982, n_4266, n_2915, n_2530, n_1148, n_31, n_2188, n_2505, n_334, n_1989, n_1161, n_2609, n_1085, n_232, n_2802, n_3796, n_2999, n_4115, n_3840, n_2014, n_2042, n_46, n_1239, n_3643, n_3697, n_771, n_1584, n_2425, n_470, n_475, n_924, n_3408, n_3461, n_298, n_1582, n_492, n_3680, n_4265, n_2318, n_3286, n_4012, n_2408, n_4246, n_1149, n_3170, n_3513, n_265, n_3468, n_3690, n_1184, n_3645, n_2483, n_2950, n_228, n_719, n_1972, n_3060, n_3304, n_3682, n_2592, n_3771, n_1525, n_3098, n_3995, n_4076, n_2594, n_455, n_2666, n_4105, n_1585, n_1851, n_363, n_1799, n_1090, n_2147, n_2564, n_592, n_4244, n_1816, n_4064, n_2503, n_2433, n_1518, n_4049, n_829, n_1156, n_1362, n_4259, n_3123, n_393, n_984, n_2600, n_3380, n_1829, n_503, n_2035, n_3508, n_3024, n_1450, n_1638, n_3422, n_132, n_868, n_3038, n_570, n_859, n_2033, n_406, n_3086, n_735, n_4104, n_1789, n_2531, n_1770, n_878, n_620, n_130, n_3285, n_519, n_4208, n_2523, n_307, n_469, n_1218, n_2413, n_500, n_3769, n_1482, n_3361, n_981, n_3596, n_714, n_3478, n_3936, n_1349, n_291, n_4089, n_1144, n_2071, n_3669, n_3863, n_357, n_3219, n_2429, n_3130, n_3702, n_985, n_4316, n_2233, n_2440, n_2723, n_481, n_3521, n_3233, n_997, n_1710, n_2800, n_2161, n_3496, n_1301, n_2805, n_802, n_561, n_33, n_3310, n_980, n_2681, n_1306, n_3264, n_2010, n_2282, n_1651, n_1198, n_3096, n_2360, n_3764, n_2047, n_4061, n_2651, n_2095, n_3239, n_1609, n_2174, n_3161, n_2799, n_436, n_4075, n_116, n_3344, n_2334, n_3902, n_4062, n_3881, n_3295, n_3947, n_409, n_1244, n_1685, n_1763, n_1998, n_3066, n_1574, n_2426, n_2490, n_2844, n_3101, n_240, n_3989, n_756, n_2303, n_1619, n_2478, n_1981, n_2285, n_4233, n_1606, n_810, n_4108, n_1133, n_635, n_95, n_1194, n_3374, n_3786, n_3841, n_2742, n_2640, n_3695, n_4051, n_1051, n_253, n_3976, n_4254, n_1552, n_2918, n_583, n_3288, n_1996, n_3563, n_3992, n_2367, n_4307, n_3876, n_249, n_201, n_2867, n_3198, n_1039, n_1442, n_3495, n_2726, n_1034, n_2043, n_4303, n_1480, n_3125, n_1158, n_2909, n_2248, n_754, n_4293, n_941, n_3552, n_975, n_3206, n_1031, n_115, n_1305, n_2363, n_2578, n_553, n_43, n_849, n_2662, n_3116, n_3147, n_3383, n_3709, n_753, n_3925, n_4091, n_1753, n_3095, n_3180, n_3738, n_3359, n_2795, n_3472, n_2471, n_4186, n_467, n_3187, n_2540, n_269, n_359, n_973, n_2807, n_1921, n_3218, n_3610, n_3618, n_3330, n_1479, n_1055, n_1675, n_2197, n_2217, n_582, n_2065, n_2879, n_861, n_3717, n_857, n_967, n_4148, n_571, n_2215, n_2461, n_271, n_404, n_2001, n_158, n_2107, n_1884, n_206, n_2040, n_679, n_4057, n_2968, n_4201, n_633, n_1170, n_665, n_1629, n_2221, n_588, n_4263, n_225, n_1260, n_308, n_309, n_1819, n_2055, n_3555, n_1010, n_3444, n_4210, n_2553, n_149, n_1040, n_915, n_632, n_3059, n_1166, n_2038, n_812, n_2891, n_1131, n_2634, n_1761, n_2709, n_3155, n_3445, n_534, n_1578, n_1006, n_1861, n_373, n_3110, n_87, n_1632, n_1890, n_3017, n_3955, n_1805, n_2477, n_257, n_1557, n_1888, n_2280, n_1833, n_3903, n_730, n_1311, n_3945, n_1494, n_2325, n_670, n_203, n_1850, n_1898, n_2443, n_2697, n_3235, n_3854, n_2308, n_4205, n_2162, n_3908, n_1868, n_207, n_2333, n_2079, n_3467, n_3001, n_3587, n_1089, n_4278, n_1887, n_1587, n_3916, n_3527, n_3795, n_2512, n_3950, n_3433, n_3852, n_1365, n_4138, n_1417, n_205, n_1242, n_2086, n_2185, n_2927, n_3673, n_1836, n_3833, n_4281, n_3815, n_2774, n_3896, n_3039, n_681, n_1226, n_3740, n_3162, n_1274, n_1486, n_2166, n_3094, n_412, n_2899, n_3274, n_3333, n_3186, n_640, n_1322, n_81, n_4129, n_965, n_1899, n_1428, n_4093, n_1616, n_1576, n_1856, n_1862, n_1958, n_2077, n_339, n_784, n_315, n_434, n_64, n_288, n_1059, n_1197, n_3065, n_3965, n_2632, n_422, n_2579, n_722, n_862, n_2105, n_135, n_3079, n_165, n_2098, n_3085, n_540, n_1423, n_2813, n_1935, n_3584, n_4039, n_3387, n_2027, n_457, n_3070, n_3800, n_2223, n_2091, n_364, n_3263, n_4197, n_3420, n_2991, n_1915, n_629, n_1621, n_4275, n_1748, n_2547, n_2415, n_4283, n_900, n_3504, n_4194, n_1449, n_531, n_827, n_2912, n_60, n_361, n_4272, n_2659, n_2930, n_1025, n_3409, n_2419, n_3111, n_2116, n_336, n_2320, n_12, n_1885, n_2677, n_1013, n_3182, n_1259, n_3054, n_3283, n_192, n_2183, n_3002, n_1538, n_51, n_649, n_4030, n_1612, n_1240, n_16688);

input n_992;
input n_2542;
input n_1671;
input n_1;
input n_2817;
input n_3660;
input n_3813;
input n_801;
input n_3766;
input n_1613;
input n_1234;
input n_1458;
input n_2576;
input n_3254;
input n_3684;
input n_1199;
input n_1674;
input n_3392;
input n_741;
input n_1027;
input n_1351;
input n_3266;
input n_3574;
input n_625;
input n_1189;
input n_3152;
input n_223;
input n_4154;
input n_3579;
input n_1212;
input n_226;
input n_208;
input n_68;
input n_4251;
input n_726;
input n_2157;
input n_3335;
input n_2332;
input n_212;
input n_3773;
input n_700;
input n_3783;
input n_4177;
input n_50;
input n_1307;
input n_3178;
input n_2003;
input n_3849;
input n_4127;
input n_1038;
input n_578;
input n_1581;
input n_1003;
input n_365;
input n_3844;
input n_168;
input n_1237;
input n_1061;
input n_2353;
input n_2534;
input n_3089;
input n_3301;
input n_4099;
input n_1357;
input n_4241;
input n_1853;
input n_3741;
input n_77;
input n_4168;
input n_783;
input n_2451;
input n_1738;
input n_2243;
input n_798;
input n_188;
input n_1575;
input n_1854;
input n_2324;
input n_3088;
input n_3443;
input n_1923;
input n_3257;
input n_509;
input n_1342;
input n_245;
input n_1209;
input n_1348;
input n_1387;
input n_2260;
input n_3222;
input n_677;
input n_1708;
input n_805;
input n_1151;
input n_396;
input n_2977;
input n_3952;
input n_1739;
input n_350;
input n_78;
input n_2051;
input n_2317;
input n_1380;
input n_3911;
input n_2359;
input n_442;
input n_480;
input n_142;
input n_2847;
input n_1402;
input n_2557;
input n_1688;
input n_1691;
input n_3332;
input n_4134;
input n_4285;
input n_3465;
input n_1975;
input n_1009;
input n_1743;
input n_62;
input n_1930;
input n_2405;
input n_3706;
input n_4050;
input n_1160;
input n_883;
input n_2647;
input n_1238;
input n_1991;
input n_2570;
input n_2179;
input n_2386;
input n_2997;
input n_4092;
input n_1724;
input n_1032;
input n_3708;
input n_2336;
input n_1247;
input n_3668;
input n_4078;
input n_1547;
input n_2521;
input n_3376;
input n_3046;
input n_2956;
input n_1553;
input n_893;
input n_1099;
input n_2491;
input n_3801;
input n_4249;
input n_1264;
input n_1192;
input n_471;
input n_3564;
input n_1844;
input n_424;
input n_3619;
input n_4087;
input n_1700;
input n_1555;
input n_1415;
input n_2211;
input n_1370;
input n_1786;
input n_3487;
input n_369;
input n_4198;
input n_287;
input n_2382;
input n_3754;
input n_2672;
input n_3030;
input n_4302;
input n_2291;
input n_415;
input n_830;
input n_2299;
input n_65;
input n_230;
input n_3340;
input n_4179;
input n_461;
input n_873;
input n_141;
input n_383;
input n_1285;
input n_1371;
input n_2886;
input n_2974;
input n_3946;
input n_200;
input n_1985;
input n_4213;
input n_2989;
input n_447;
input n_2838;
input n_2184;
input n_3395;
input n_2982;
input n_1803;
input n_3427;
input n_1172;
input n_852;
input n_2509;
input n_4065;
input n_4026;
input n_71;
input n_229;
input n_2513;
input n_3282;
input n_1590;
input n_2645;
input n_1532;
input n_2313;
input n_2628;
input n_3071;
input n_3626;
input n_3757;
input n_3904;
input n_4178;
input n_1393;
input n_1517;
input n_1867;
input n_2926;
input n_1704;
input n_1078;
input n_250;
input n_544;
input n_1711;
input n_2247;
input n_3106;
input n_1140;
input n_2630;
input n_4273;
input n_1444;
input n_1670;
input n_1603;
input n_2344;
input n_1579;
input n_3275;
input n_35;
input n_2365;
input n_2470;
input n_2321;
input n_1263;
input n_2019;
input n_3031;
input n_4029;
input n_836;
input n_3345;
input n_375;
input n_2074;
input n_2447;
input n_522;
input n_2919;
input n_3678;
input n_3440;
input n_2129;
input n_2340;
input n_1261;
input n_945;
input n_3879;
input n_4010;
input n_2286;
input n_1649;
input n_2018;
input n_2094;
input n_3080;
input n_1903;
input n_1511;
input n_1143;
input n_2356;
input n_2399;
input n_1422;
input n_1232;
input n_1772;
input n_1572;
input n_3979;
input n_616;
input n_658;
input n_4308;
input n_1874;
input n_3165;
input n_1119;
input n_2865;
input n_2825;
input n_3463;
input n_2013;
input n_428;
input n_1433;
input n_1902;
input n_1842;
input n_1620;
input n_2044;
input n_1954;
input n_1735;
input n_2510;
input n_1541;
input n_1300;
input n_641;
input n_2480;
input n_2739;
input n_3023;
input n_822;
input n_3232;
input n_693;
input n_1313;
input n_2791;
input n_3607;
input n_3750;
input n_3251;
input n_1056;
input n_3877;
input n_3316;
input n_2212;
input n_3929;
input n_758;
input n_516;
input n_3494;
input n_3048;
input n_1455;
input n_2418;
input n_2864;
input n_1163;
input n_2729;
input n_3063;
input n_4311;
input n_1180;
input n_2256;
input n_2582;
input n_943;
input n_1798;
input n_4060;
input n_1550;
input n_2703;
input n_491;
input n_3998;
input n_2786;
input n_3371;
input n_1591;
input n_42;
input n_772;
input n_3632;
input n_3122;
input n_2806;
input n_1344;
input n_3261;
input n_2730;
input n_2495;
input n_666;
input n_371;
input n_4187;
input n_940;
input n_770;
input n_567;
input n_1781;
input n_1971;
input n_2058;
input n_2090;
input n_2603;
input n_405;
input n_213;
input n_2660;
input n_538;
input n_3028;
input n_3829;
input n_3662;
input n_2981;
input n_3076;
input n_2173;
input n_4164;
input n_2004;
input n_1106;
input n_886;
input n_1471;
input n_343;
input n_953;
input n_1094;
input n_3624;
input n_3077;
input n_3737;
input n_1345;
input n_1820;
input n_2873;
input n_3452;
input n_3655;
input n_494;
input n_539;
input n_493;
input n_3107;
input n_155;
input n_3825;
input n_2880;
input n_3225;
input n_2394;
input n_2108;
input n_3532;
input n_45;
input n_4117;
input n_454;
input n_3948;
input n_1421;
input n_2836;
input n_3664;
input n_1936;
input n_638;
input n_1404;
input n_1211;
input n_2124;
input n_381;
input n_2378;
input n_887;
input n_1660;
input n_1961;
input n_3047;
input n_112;
input n_1280;
input n_3765;
input n_713;
input n_2655;
input n_4125;
input n_1400;
input n_2625;
input n_3296;
input n_2843;
input n_126;
input n_4221;
input n_1467;
input n_3297;
input n_4250;
input n_58;
input n_976;
input n_3760;
input n_3067;
input n_2155;
input n_3906;
input n_224;
input n_2686;
input n_48;
input n_1445;
input n_2364;
input n_2551;
input n_1526;
input n_1560;
input n_734;
input n_1088;
input n_4262;
input n_1894;
input n_196;
input n_1231;
input n_2996;
input n_2599;
input n_2985;
input n_1978;
input n_3803;
input n_2085;
input n_3963;
input n_3368;
input n_917;
input n_574;
input n_3639;
input n_9;
input n_3347;
input n_2370;
input n_2612;
input n_3792;
input n_907;
input n_4202;
input n_6;
input n_1446;
input n_14;
input n_3938;
input n_2591;
input n_3507;
input n_659;
input n_1815;
input n_2214;
input n_3351;
input n_4253;
input n_407;
input n_913;
input n_4110;
input n_1658;
input n_2593;
input n_808;
input n_867;
input n_4071;
input n_4255;
input n_3506;
input n_4268;
input n_3568;
input n_3269;
input n_4047;
input n_3531;
input n_1230;
input n_3413;
input n_3850;
input n_473;
input n_1193;
input n_1967;
input n_3999;
input n_1054;
input n_3928;
input n_559;
input n_3412;
input n_2613;
input n_3535;
input n_1333;
input n_2496;
input n_44;
input n_2708;
input n_3313;
input n_1648;
input n_3189;
input n_1911;
input n_1956;
input n_163;
input n_1644;
input n_3791;
input n_4139;
input n_2011;
input n_2725;
input n_2277;
input n_3164;
input n_1558;
input n_1732;
input n_281;
input n_551;
input n_699;
input n_1986;
input n_2300;
input n_3943;
input n_4320;
input n_4305;
input n_564;
input n_2397;
input n_3884;
input n_3931;
input n_451;
input n_824;
input n_279;
input n_686;
input n_4102;
input n_4297;
input n_757;
input n_594;
input n_1641;
input n_2113;
input n_1918;
input n_2190;
input n_3603;
input n_3871;
input n_2907;
input n_577;
input n_3438;
input n_166;
input n_2735;
input n_4141;
input n_1843;
input n_619;
input n_3959;
input n_2268;
input n_1367;
input n_1336;
input n_521;
input n_2778;
input n_4227;
input n_2850;
input n_572;
input n_4314;
input n_395;
input n_813;
input n_1909;
input n_2080;
input n_1481;
input n_3822;
input n_323;
input n_4163;
input n_606;
input n_1441;
input n_818;
input n_3373;
input n_1123;
input n_1309;
input n_92;
input n_2104;
input n_513;
input n_645;
input n_1381;
input n_2961;
input n_3812;
input n_331;
input n_1699;
input n_3910;
input n_916;
input n_3934;
input n_2093;
input n_4033;
input n_4296;
input n_4009;
input n_2633;
input n_483;
input n_102;
input n_3883;
input n_2207;
input n_1970;
input n_2770;
input n_608;
input n_261;
input n_2101;
input n_2696;
input n_3482;
input n_4080;
input n_630;
input n_2059;
input n_32;
input n_2198;
input n_3319;
input n_541;
input n_512;
input n_2669;
input n_2925;
input n_3728;
input n_4094;
input n_2073;
input n_2273;
input n_121;
input n_3484;
input n_433;
input n_3748;
input n_2546;
input n_3272;
input n_3193;
input n_792;
input n_2522;
input n_476;
input n_3949;
input n_2792;
input n_2;
input n_1328;
input n_3396;
input n_1957;
input n_2917;
input n_219;
input n_2616;
input n_3912;
input n_3118;
input n_3315;
input n_3720;
input n_1907;
input n_3923;
input n_2529;
input n_264;
input n_263;
input n_3900;
input n_1162;
input n_860;
input n_1530;
input n_3798;
input n_788;
input n_939;
input n_3488;
input n_1543;
input n_821;
input n_2811;
input n_938;
input n_1302;
input n_1068;
input n_1599;
input n_3732;
input n_329;
input n_982;
input n_4257;
input n_2674;
input n_2832;
input n_4226;
input n_549;
input n_1762;
input n_1910;
input n_1075;
input n_3980;
input n_408;
input n_932;
input n_2831;
input n_2998;
input n_4318;
input n_3446;
input n_4158;
input n_61;
input n_3317;
input n_237;
input n_3857;
input n_3978;
input n_1876;
input n_4107;
input n_1895;
input n_2123;
input n_1697;
input n_2143;
input n_243;
input n_979;
input n_4074;
input n_3716;
input n_1873;
input n_4294;
input n_905;
input n_3630;
input n_3518;
input n_3824;
input n_3859;
input n_1866;
input n_4013;
input n_1680;
input n_117;
input n_175;
input n_322;
input n_993;
input n_2692;
input n_3842;
input n_689;
input n_3248;
input n_2031;
input n_354;
input n_2130;
input n_1330;
input n_1413;
input n_1605;
input n_3714;
input n_3514;
input n_2228;
input n_3914;
input n_3397;
input n_134;
input n_1988;
input n_2941;
input n_1278;
input n_547;
input n_3575;
input n_2455;
input n_2876;
input n_558;
input n_2654;
input n_3036;
input n_2469;
input n_4032;
input n_1064;
input n_3099;
input n_1396;
input n_634;
input n_2355;
input n_3927;
input n_4147;
input n_136;
input n_966;
input n_3888;
input n_2908;
input n_3168;
input n_764;
input n_2751;
input n_2764;
input n_3357;
input n_1663;
input n_4130;
input n_4161;
input n_2895;
input n_2009;
input n_4172;
input n_692;
input n_3403;
input n_733;
input n_1793;
input n_2922;
input n_3601;
input n_3882;
input n_1233;
input n_1289;
input n_2714;
input n_2245;
input n_487;
input n_3055;
input n_3092;
input n_3492;
input n_3895;
input n_241;
input n_3966;
input n_30;
input n_2068;
input n_1107;
input n_2866;
input n_2457;
input n_3294;
input n_4119;
input n_1014;
input n_3734;
input n_3686;
input n_1290;
input n_1703;
input n_2580;
input n_3455;
input n_4118;
input n_882;
input n_2176;
input n_2072;
input n_3649;
input n_1354;
input n_2821;
input n_586;
input n_423;
input n_1865;
input n_1875;
input n_1701;
input n_2459;
input n_318;
input n_3746;
input n_1111;
input n_1713;
input n_2971;
input n_715;
input n_3599;
input n_2678;
input n_1251;
input n_3384;
input n_3935;
input n_1265;
input n_4277;
input n_2711;
input n_3490;
input n_4291;
input n_88;
input n_4199;
input n_1726;
input n_1950;
input n_530;
input n_1563;
input n_1912;
input n_277;
input n_2434;
input n_4319;
input n_3369;
input n_3419;
input n_1982;
input n_3872;
input n_2878;
input n_618;
input n_3012;
input n_1297;
input n_1662;
input n_1312;
input n_3772;
input n_3875;
input n_199;
input n_1167;
input n_1359;
input n_2818;
input n_2428;
input n_3581;
input n_3794;
input n_674;
input n_3247;
input n_871;
input n_3069;
input n_3921;
input n_922;
input n_268;
input n_1335;
input n_1760;
input n_1927;
input n_210;
input n_2028;
input n_3715;
input n_1069;
input n_2664;
input n_5;
input n_1664;
input n_1722;
input n_612;
input n_2641;
input n_3022;
input n_3052;
input n_3725;
input n_178;
input n_247;
input n_1165;
input n_355;
input n_3933;
input n_702;
input n_347;
input n_2008;
input n_2749;
input n_3298;
input n_2192;
input n_3281;
input n_2254;
input n_2345;
input n_3346;
input n_1926;
input n_1175;
input n_3273;
input n_328;
input n_1386;
input n_2311;
input n_1896;
input n_429;
input n_2965;
input n_1747;
input n_3058;
input n_1012;
input n_195;
input n_3691;
input n_780;
input n_3861;
input n_675;
input n_2624;
input n_4066;
input n_903;
input n_4146;
input n_1540;
input n_1977;
input n_1802;
input n_1504;
input n_3549;
input n_2350;
input n_2804;
input n_2453;
input n_286;
input n_254;
input n_3891;
input n_2193;
input n_3961;
input n_2676;
input n_1655;
input n_3940;
input n_4072;
input n_4220;
input n_242;
input n_835;
input n_1214;
input n_928;
input n_47;
input n_690;
input n_850;
input n_1801;
input n_1886;
input n_2092;
input n_2347;
input n_1654;
input n_816;
input n_1157;
input n_3453;
input n_1750;
input n_2994;
input n_1462;
input n_3410;
input n_3153;
input n_3428;
input n_1188;
input n_3689;
input n_1752;
input n_877;
input n_1813;
input n_2514;
input n_3768;
input n_2206;
input n_604;
input n_4004;
input n_2810;
input n_2967;
input n_2319;
input n_2519;
input n_4043;
input n_825;
input n_4313;
input n_728;
input n_2916;
input n_3415;
input n_1063;
input n_4292;
input n_1588;
input n_3785;
input n_3942;
input n_3997;
input n_2963;
input n_4041;
input n_2947;
input n_3918;
input n_2467;
input n_26;
input n_2602;
input n_2468;
input n_55;
input n_267;
input n_3145;
input n_1124;
input n_1624;
input n_3873;
input n_3983;
input n_515;
input n_2096;
input n_2980;
input n_3968;
input n_1965;
input n_3538;
input n_2476;
input n_3280;
input n_598;
input n_3434;
input n_696;
input n_1515;
input n_961;
input n_3510;
input n_437;
input n_1082;
input n_1317;
input n_3227;
input n_2733;
input n_2824;
input n_3289;
input n_593;
input n_4169;
input n_514;
input n_4055;
input n_687;
input n_697;
input n_890;
input n_637;
input n_2377;
input n_295;
input n_701;
input n_2178;
input n_3271;
input n_950;
input n_4248;
input n_388;
input n_190;
input n_2812;
input n_484;
input n_2644;
input n_2036;
input n_3326;
input n_2976;
input n_2152;
input n_1709;
input n_3009;
input n_2652;
input n_4200;
input n_3460;
input n_2411;
input n_3719;
input n_2525;
input n_1825;
input n_2393;
input n_1757;
input n_1796;
input n_170;
input n_2657;
input n_1792;
input n_3827;
input n_891;
input n_2067;
input n_2136;
input n_2921;
input n_2409;
input n_2082;
input n_3519;
input n_2252;
input n_1412;
input n_2497;
input n_3889;
input n_2687;
input n_3237;
input n_949;
input n_1630;
input n_678;
input n_2887;
input n_3809;
input n_3500;
input n_3834;
input n_4245;
input n_4136;
input n_3526;
input n_3707;
input n_283;
input n_2075;
input n_4045;
input n_2194;
input n_2972;
input n_2619;
input n_3139;
input n_3542;
input n_91;
input n_2763;
input n_2762;
input n_4070;
input n_1987;
input n_3545;
input n_507;
input n_968;
input n_909;
input n_1369;
input n_3578;
input n_3885;
input n_881;
input n_2271;
input n_1008;
input n_3192;
input n_760;
input n_3993;
input n_1546;
input n_2583;
input n_590;
input n_4116;
input n_63;
input n_2606;
input n_4031;
input n_362;
input n_148;
input n_2279;
input n_161;
input n_22;
input n_462;
input n_1033;
input n_1052;
input n_2794;
input n_1296;
input n_2663;
input n_1990;
input n_3352;
input n_2391;
input n_3805;
input n_304;
input n_2431;
input n_3073;
input n_4018;
input n_2987;
input n_694;
input n_2938;
input n_2150;
input n_1294;
input n_2943;
input n_1420;
input n_3696;
input n_3780;
input n_4082;
input n_125;
input n_1634;
input n_2078;
input n_3252;
input n_2932;
input n_297;
input n_595;
input n_627;
input n_1767;
input n_1779;
input n_524;
input n_1465;
input n_3253;
input n_3337;
input n_3431;
input n_342;
input n_3209;
input n_3450;
input n_2622;
input n_1858;
input n_1044;
input n_4002;
input n_2658;
input n_2665;
input n_2165;
input n_2133;
input n_1712;
input n_3021;
input n_1391;
input n_449;
input n_131;
input n_1523;
input n_2558;
input n_2750;
input n_2775;
input n_1208;
input n_2893;
input n_1164;
input n_1295;
input n_1627;
input n_2954;
input n_3477;
input n_4288;
input n_2728;
input n_2349;
input n_3128;
input n_3763;
input n_4289;
input n_2684;
input n_2712;
input n_1072;
input n_3146;
input n_1527;
input n_1495;
input n_3733;
input n_1438;
input n_495;
input n_815;
input n_3953;
input n_1100;
input n_585;
input n_1487;
input n_2691;
input n_3421;
input n_840;
input n_2913;
input n_3614;
input n_874;
input n_1756;
input n_3183;
input n_1128;
input n_2493;
input n_382;
input n_673;
input n_2230;
input n_2705;
input n_1969;
input n_4019;
input n_2690;
input n_1071;
input n_1067;
input n_1565;
input n_1493;
input n_2145;
input n_3405;
input n_1968;
input n_898;
input n_255;
input n_284;
input n_1952;
input n_865;
input n_3616;
input n_4228;
input n_2573;
input n_3423;
input n_2646;
input n_4044;
input n_3436;
input n_925;
input n_1932;
input n_1101;
input n_15;
input n_1026;
input n_1880;
input n_2535;
input n_3366;
input n_3442;
input n_2631;
input n_4191;
input n_38;
input n_289;
input n_1364;
input n_3078;
input n_3644;
input n_2436;
input n_3937;
input n_615;
input n_2870;
input n_1249;
input n_2706;
input n_3838;
input n_59;
input n_4287;
input n_1293;
input n_2693;
input n_4137;
input n_1127;
input n_1512;
input n_2151;
input n_3159;
input n_1451;
input n_3941;
input n_320;
input n_108;
input n_639;
input n_963;
input n_794;
input n_2767;
input n_3793;
input n_727;
input n_894;
input n_1839;
input n_2341;
input n_685;
input n_1765;
input n_3727;
input n_353;
input n_2707;
input n_3240;
input n_3576;
input n_3789;
input n_605;
input n_1514;
input n_1863;
input n_826;
input n_3385;
input n_3747;
input n_3037;
input n_1646;
input n_3293;
input n_872;
input n_1139;
input n_1714;
input n_3922;
input n_86;
input n_3179;
input n_104;
input n_718;
input n_1018;
input n_3400;
input n_3729;
input n_1521;
input n_1366;
input n_4000;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_2537;
input n_2897;
input n_3970;
input n_305;
input n_72;
input n_2554;
input n_996;
input n_532;
input n_173;
input n_1308;
input n_2089;
input n_1376;
input n_3522;
input n_1513;
input n_2747;
input n_3924;
input n_413;
input n_3171;
input n_791;
input n_1913;
input n_4216;
input n_3608;
input n_510;
input n_837;
input n_4315;
input n_2097;
input n_79;
input n_2170;
input n_3459;
input n_4156;
input n_3491;
input n_4240;
input n_1488;
input n_2853;
input n_1808;
input n_3053;
input n_948;
input n_3358;
input n_2517;
input n_2713;
input n_3499;
input n_704;
input n_2148;
input n_4284;
input n_4162;
input n_977;
input n_2339;
input n_1005;
input n_1947;
input n_2765;
input n_2861;
input n_536;
input n_3158;
input n_1788;
input n_3426;
input n_1999;
input n_2731;
input n_622;
input n_147;
input n_2590;
input n_2643;
input n_3150;
input n_3018;
input n_3353;
input n_3782;
input n_3975;
input n_1469;
input n_2060;
input n_2608;
input n_1838;
input n_2638;
input n_4011;
input n_1835;
input n_3470;
input n_1766;
input n_1776;
input n_1959;
input n_3133;
input n_2002;
input n_581;
input n_2650;
input n_2138;
input n_4098;
input n_4021;
input n_765;
input n_432;
input n_987;
input n_1492;
input n_3700;
input n_2414;
input n_1340;
input n_3014;
input n_3166;
input n_1771;
input n_2316;
input n_4058;
input n_4103;
input n_3104;
input n_631;
input n_720;
input n_3435;
input n_153;
input n_842;
input n_3148;
input n_2262;
input n_3229;
input n_3348;
input n_4022;
input n_1707;
input n_2239;
input n_3082;
input n_3611;
input n_4310;
input n_1432;
input n_156;
input n_145;
input n_2208;
input n_843;
input n_656;
input n_989;
input n_2604;
input n_2407;
input n_1277;
input n_2816;
input n_797;
input n_2689;
input n_2933;
input n_1473;
input n_2191;
input n_1723;
input n_2717;
input n_1246;
input n_3799;
input n_1878;
input n_2574;
input n_899;
input n_189;
input n_738;
input n_2012;
input n_3497;
input n_1304;
input n_1035;
input n_294;
input n_2842;
input n_499;
input n_2675;
input n_1426;
input n_3418;
input n_705;
input n_3580;
input n_3775;
input n_11;
input n_3537;
input n_1004;
input n_1176;
input n_2134;
input n_1529;
input n_2335;
input n_2473;
input n_3887;
input n_1022;
input n_614;
input n_529;
input n_2069;
input n_2307;
input n_3704;
input n_2362;
input n_425;
input n_684;
input n_2539;
input n_2667;
input n_2698;
input n_4096;
input n_1431;
input n_4123;
input n_1615;
input n_4114;
input n_1474;
input n_3312;
input n_1571;
input n_3835;
input n_4286;
input n_1809;
input n_3119;
input n_4280;
input n_2948;
input n_1577;
input n_2958;
input n_3735;
input n_2297;
input n_1181;
input n_2119;
input n_3731;
input n_1822;
input n_37;
input n_486;
input n_947;
input n_2936;
input n_3224;
input n_1117;
input n_2489;
input n_1087;
input n_1448;
input n_3173;
input n_1992;
input n_3677;
input n_3631;
input n_648;
input n_657;
input n_1049;
input n_3223;
input n_3996;
input n_2771;
input n_2445;
input n_3020;
input n_2057;
input n_2103;
input n_3140;
input n_3185;
input n_3770;
input n_2605;
input n_4097;
input n_1666;
input n_2772;
input n_1505;
input n_803;
input n_290;
input n_4218;
input n_118;
input n_1717;
input n_926;
input n_1817;
input n_2449;
input n_927;
input n_3557;
input n_2610;
input n_3654;
input n_3129;
input n_3880;
input n_1849;
input n_2848;
input n_919;
input n_3685;
input n_2868;
input n_3620;
input n_1698;
input n_478;
input n_4100;
input n_2231;
input n_3609;
input n_929;
input n_107;
input n_3832;
input n_2520;
input n_1228;
input n_417;
input n_4264;
input n_2857;
input n_446;
input n_3693;
input n_3788;
input n_89;
input n_1568;
input n_1490;
input n_2372;
input n_777;
input n_1299;
input n_272;
input n_2896;
input n_526;
input n_3837;
input n_2718;
input n_3019;
input n_2639;
input n_3471;
input n_1183;
input n_1436;
input n_2898;
input n_2251;
input n_1384;
input n_69;
input n_3674;
input n_2494;
input n_2959;
input n_4079;
input n_2501;
input n_3203;
input n_3325;
input n_2238;
input n_293;
input n_4085;
input n_2368;
input n_53;
input n_458;
input n_1070;
input n_2403;
input n_3342;
input n_2837;
input n_4175;
input n_998;
input n_16;
input n_717;
input n_3200;
input n_1665;
input n_4306;
input n_3600;
input n_18;
input n_3259;
input n_2524;
input n_154;
input n_3167;
input n_1383;
input n_2460;
input n_4224;
input n_3390;
input n_3656;
input n_1178;
input n_98;
input n_2127;
input n_1424;
input n_2338;
input n_3324;
input n_3593;
input n_3341;
input n_3867;
input n_1073;
input n_1000;
input n_796;
input n_252;
input n_1195;
input n_3559;
input n_3025;
input n_2137;
input n_1626;
input n_3191;
input n_4005;
input n_1507;
input n_2482;
input n_184;
input n_552;
input n_3810;
input n_3546;
input n_2532;
input n_1358;
input n_1811;
input n_1388;
input n_3661;
input n_3006;
input n_216;
input n_4140;
input n_2481;
input n_3561;
input n_912;
input n_1857;
input n_3987;
input n_1519;
input n_2144;
input n_3056;
input n_745;
input n_1284;
input n_1604;
input n_2296;
input n_2424;
input n_3201;
input n_3633;
input n_3447;
input n_3971;
input n_1142;
input n_2849;
input n_716;
input n_1475;
input n_623;
input n_1048;
input n_1201;
input n_1398;
input n_884;
input n_1774;
input n_2354;
input n_2682;
input n_3032;
input n_3103;
input n_3638;
input n_2589;
input n_1395;
input n_2110;
input n_2199;
input n_2661;
input n_731;
input n_2877;
input n_1502;
input n_1659;
input n_1955;
input n_755;
input n_931;
input n_1021;
input n_3393;
input n_474;
input n_527;
input n_683;
input n_811;
input n_1207;
input n_2442;
input n_3627;
input n_312;
input n_1791;
input n_1368;
input n_66;
input n_3451;
input n_3480;
input n_1418;
input n_958;
input n_292;
input n_1250;
input n_100;
input n_3331;
input n_1137;
input n_3615;
input n_1897;
input n_2064;
input n_880;
input n_3072;
input n_3087;
input n_2053;
input n_3612;
input n_3505;
input n_2259;
input n_2121;
input n_2773;
input n_4222;
input n_2545;
input n_3540;
input n_3577;
input n_889;
input n_3509;
input n_2432;
input n_2710;
input n_150;
input n_1478;
input n_589;
input n_3606;
input n_1310;
input n_3142;
input n_3598;
input n_819;
input n_2966;
input n_2294;
input n_1363;
input n_2581;
input n_1334;
input n_1942;
input n_1966;
input n_3591;
input n_767;
input n_3641;
input n_1314;
input n_600;
input n_964;
input n_831;
input n_1837;
input n_2218;
input n_2788;
input n_477;
input n_3196;
input n_3590;
input n_2435;
input n_954;
input n_864;
input n_2504;
input n_2797;
input n_2623;
input n_1110;
input n_2213;
input n_1410;
input n_399;
input n_2389;
input n_1440;
input n_124;
input n_2132;
input n_2892;
input n_2063;
input n_4120;
input n_1382;
input n_1534;
input n_3892;
input n_1564;
input n_1736;
input n_4069;
input n_211;
input n_2748;
input n_4053;
input n_1483;
input n_3848;
input n_1834;
input n_2331;
input n_1372;
input n_231;
input n_2292;
input n_2860;
input n_3327;
input n_2330;
input n_40;
input n_3441;
input n_1457;
input n_505;
input n_1719;
input n_3534;
input n_3718;
input n_319;
input n_1339;
input n_1787;
input n_2701;
input n_2475;
input n_537;
input n_2511;
input n_3964;
input n_1993;
input n_2281;
input n_4167;
input n_1427;
input n_311;
input n_2416;
input n_2745;
input n_2617;
input n_2776;
input n_1466;
input n_10;
input n_403;
input n_1919;
input n_1080;
input n_723;
input n_1877;
input n_3144;
input n_3705;
input n_3211;
input n_3244;
input n_596;
input n_123;
input n_3909;
input n_3944;
input n_546;
input n_562;
input n_1141;
input n_1268;
input n_386;
input n_1939;
input n_2030;
input n_1769;
input n_1220;
input n_2323;
input n_1893;
input n_556;
input n_2784;
input n_2209;
input n_2301;
input n_3582;
input n_3605;
input n_162;
input n_3287;
input n_4223;
input n_2387;
input n_3322;
input n_1755;
input n_1602;
input n_2421;
input n_1136;
input n_3270;
input n_2618;
input n_2025;
input n_2357;
input n_2846;
input n_2464;
input n_3265;
input n_128;
input n_1125;
input n_3755;
input n_4042;
input n_970;
input n_3306;
input n_2488;
input n_3640;
input n_2224;
input n_1980;
input n_642;
input n_995;
input n_276;
input n_1159;
input n_2329;
input n_1092;
input n_3481;
input n_2237;
input n_3026;
input n_441;
input n_221;
input n_1060;
input n_1951;
input n_2250;
input n_3090;
input n_4299;
input n_444;
input n_3033;
input n_3724;
input n_146;
input n_1252;
input n_1784;
input n_3311;
input n_3571;
input n_1223;
input n_3913;
input n_303;
input n_4276;
input n_511;
input n_2990;
input n_3847;
input n_193;
input n_1286;
input n_1773;
input n_1775;
input n_2115;
input n_2410;
input n_2552;
input n_1053;
input n_3302;
input n_2374;
input n_416;
input n_1681;
input n_520;
input n_418;
input n_1093;
input n_113;
input n_1783;
input n_1533;
input n_1597;
input n_2929;
input n_2780;
input n_3226;
input n_3323;
input n_3364;
input n_4;
input n_4020;
input n_4176;
input n_266;
input n_296;
input n_2596;
input n_2274;
input n_3163;
input n_775;
input n_651;
input n_1153;
input n_439;
input n_1618;
input n_3407;
input n_217;
input n_518;
input n_1531;
input n_2828;
input n_1185;
input n_3856;
input n_453;
input n_4236;
input n_3425;
input n_215;
input n_2384;
input n_3894;
input n_4204;
input n_4261;
input n_1745;
input n_914;
input n_759;
input n_3479;
input n_3127;
input n_2724;
input n_1831;
input n_426;
input n_317;
input n_2585;
input n_2621;
input n_3623;
input n_1653;
input n_2352;
input n_1679;
input n_4063;
input n_1625;
input n_90;
input n_3986;
input n_4237;
input n_2601;
input n_2160;
input n_3454;
input n_54;
input n_1453;
input n_2146;
input n_4006;
input n_2226;
input n_2131;
input n_488;
input n_2502;
input n_2801;
input n_3646;
input n_497;
input n_2920;
input n_4015;
input n_773;
input n_3547;
input n_1901;
input n_3869;
input n_920;
input n_99;
input n_1374;
input n_2556;
input n_2648;
input n_3212;
input n_1315;
input n_1647;
input n_13;
input n_2575;
input n_2754;
input n_1224;
input n_2783;
input n_3753;
input n_2306;
input n_1614;
input n_1459;
input n_1892;
input n_3188;
input n_3742;
input n_1933;
input n_2462;
input n_1135;
input n_1169;
input n_1179;
input n_2889;
input n_3243;
input n_3683;
input n_401;
input n_4034;
input n_324;
input n_1617;
input n_4056;
input n_3260;
input n_3370;
input n_3386;
input n_3816;
input n_335;
input n_3960;
input n_1470;
input n_2550;
input n_463;
input n_3093;
input n_3175;
input n_3214;
input n_1243;
input n_3736;
input n_848;
input n_120;
input n_2732;
input n_301;
input n_2928;
input n_274;
input n_4206;
input n_1096;
input n_2249;
input n_1091;
input n_1917;
input n_2000;
input n_3862;
input n_4267;
input n_1580;
input n_2227;
input n_4247;
input n_2270;
input n_2822;
input n_1425;
input n_3169;
input n_36;
input n_4180;
input n_3205;
input n_1881;
input n_1267;
input n_1281;
input n_1806;
input n_3284;
input n_983;
input n_3109;
input n_2023;
input n_3354;
input n_427;
input n_2572;
input n_2204;
input n_1520;
input n_496;
input n_2720;
input n_3126;
input n_2159;
input n_906;
input n_1390;
input n_688;
input n_2289;
input n_1077;
input n_1733;
input n_2315;
input n_1419;
input n_2863;
input n_3299;
input n_3663;
input n_4132;
input n_351;
input n_2955;
input n_2995;
input n_259;
input n_1731;
input n_177;
input n_2158;
input n_2087;
input n_1855;
input n_1636;
input n_3051;
input n_1437;
input n_3360;
input n_2135;
input n_3956;
input n_3367;
input n_1645;
input n_1832;
input n_4001;
input n_385;
input n_1687;
input n_1439;
input n_2328;
input n_1323;
input n_2859;
input n_2202;
input n_858;
input n_2049;
input n_4149;
input n_1331;
input n_613;
input n_736;
input n_2627;
input n_501;
input n_956;
input n_960;
input n_2276;
input n_3234;
input n_3917;
input n_663;
input n_856;
input n_2803;
input n_2100;
input n_3314;
input n_3525;
input n_379;
input n_2993;
input n_778;
input n_1668;
input n_2777;
input n_1134;
input n_3016;
input n_3566;
input n_3688;
input n_3004;
input n_3202;
input n_2830;
input n_2781;
input n_3220;
input n_4003;
input n_410;
input n_1129;
input n_3870;
input n_4126;
input n_554;
input n_602;
input n_1696;
input n_2829;
input n_1995;
input n_1594;
input n_2181;
input n_3751;
input n_664;
input n_1869;
input n_171;
input n_2911;
input n_3625;
input n_3804;
input n_1764;
input n_169;
input n_4207;
input n_1429;
input n_2826;
input n_1610;
input n_3084;
input n_3429;
input n_4113;
input n_1889;
input n_2379;
input n_435;
input n_1905;
input n_2016;
input n_2343;
input n_793;
input n_326;
input n_587;
input n_3466;
input n_3554;
input n_1593;
input n_580;
input n_762;
input n_1030;
input n_1202;
input n_3901;
input n_1937;
input n_465;
input n_1790;
input n_1778;
input n_3749;
input n_1635;
input n_2942;
input n_4014;
input n_1079;
input n_341;
input n_2515;
input n_1744;
input n_828;
input n_2139;
input n_2142;
input n_4067;
input n_4252;
input n_607;
input n_316;
input n_419;
input n_28;
input n_1551;
input n_4028;
input n_4054;
input n_2448;
input n_1103;
input n_2875;
input n_3907;
input n_2555;
input n_4048;
input n_3338;
input n_144;
input n_4217;
input n_3586;
input n_3462;
input n_3756;
input n_2219;
input n_1203;
input n_3653;
input n_3636;
input n_2851;
input n_3406;
input n_820;
input n_2327;
input n_951;
input n_106;
input n_2201;
input n_725;
input n_952;
input n_3919;
input n_999;
input n_358;
input n_1254;
input n_160;
input n_2841;
input n_3349;
input n_2420;
input n_3722;
input n_186;
input n_2984;
input n_0;
input n_368;
input n_575;
input n_994;
input n_2263;
input n_3539;
input n_3291;
input n_2304;
input n_4024;
input n_1508;
input n_2487;
input n_732;
input n_974;
input n_2983;
input n_2240;
input n_392;
input n_2278;
input n_2656;
input n_2538;
input n_724;
input n_2597;
input n_2375;
input n_3113;
input n_3194;
input n_3250;
input n_1934;
input n_3276;
input n_1020;
input n_1042;
input n_628;
input n_1273;
input n_1434;
input n_1573;
input n_3981;
input n_4214;
input n_1728;
input n_3973;
input n_557;
input n_2756;
input n_3572;
input n_1871;
input n_349;
input n_3448;
input n_617;
input n_3886;
input n_845;
input n_807;
input n_2924;
input n_1036;
input n_3595;
input n_140;
input n_1138;
input n_3414;
input n_1661;
input n_1275;
input n_2884;
input n_485;
input n_1549;
input n_67;
input n_443;
input n_1510;
input n_892;
input n_768;
input n_3637;
input n_421;
input n_3120;
input n_1468;
input n_3991;
input n_2855;
input n_3651;
input n_1859;
input n_2102;
input n_3516;
input n_2563;
input n_3797;
input n_3926;
input n_238;
input n_1095;
input n_2024;
input n_1595;
input n_202;
input n_2156;
input n_3449;
input n_1718;
input n_1749;
input n_3474;
input n_1683;
input n_1916;
input n_2598;
input n_597;
input n_280;
input n_1270;
input n_2549;
input n_1187;
input n_610;
input n_4234;
input n_4304;
input n_1403;
input n_1669;
input n_1852;
input n_4101;
input n_3548;
input n_3767;
input n_1024;
input n_3864;
input n_4036;
input n_1768;
input n_2153;
input n_2544;
input n_2381;
input n_3670;
input n_3550;
input n_3974;
input n_198;
input n_1847;
input n_2052;
input n_3634;
input n_179;
input n_248;
input n_2302;
input n_517;
input n_4211;
input n_4182;
input n_1667;
input n_667;
input n_1206;
input n_3230;
input n_4016;
input n_621;
input n_1037;
input n_1397;
input n_3268;
input n_3236;
input n_1279;
input n_1115;
input n_750;
input n_901;
input n_1499;
input n_3592;
input n_468;
input n_2755;
input n_3141;
input n_923;
input n_504;
input n_1409;
input n_4230;
input n_1841;
input n_3839;
input n_2637;
input n_2823;
input n_1639;
input n_1623;
input n_183;
input n_1015;
input n_3967;
input n_1503;
input n_3112;
input n_2819;
input n_3195;
input n_466;
input n_2526;
input n_3041;
input n_4274;
input n_2423;
input n_1057;
input n_3277;
input n_3108;
input n_2548;
input n_603;
input n_991;
input n_2785;
input n_1657;
input n_4189;
input n_4270;
input n_235;
input n_4151;
input n_1126;
input n_2412;
input n_1997;
input n_3817;
input n_3417;
input n_2636;
input n_3131;
input n_340;
input n_710;
input n_1108;
input n_1818;
input n_2439;
input n_2404;
input n_1182;
input n_3730;
input n_1298;
input n_4124;
input n_3659;
input n_2559;
input n_2177;
input n_39;
input n_2595;
input n_3399;
input n_2088;
input n_3635;
input n_73;
input n_1611;
input n_785;
input n_4155;
input n_2740;
input n_746;
input n_4238;
input n_609;
input n_1601;
input n_3011;
input n_1960;
input n_2694;
input n_2061;
input n_3416;
input n_3648;
input n_1686;
input n_3498;
input n_2757;
input n_2337;
input n_2401;
input n_101;
input n_167;
input n_1356;
input n_1589;
input n_3042;
input n_3213;
input n_127;
input n_3820;
input n_2309;
input n_2900;
input n_2957;
input n_2607;
input n_1740;
input n_2737;
input n_3994;
input n_1497;
input n_2890;
input n_1168;
input n_1216;
input n_1943;
input n_3228;
input n_133;
input n_1320;
input n_2716;
input n_96;
input n_3249;
input n_3081;
input n_3657;
input n_2452;
input n_1430;
input n_3650;
input n_1316;
input n_1287;
input n_2722;
input n_1452;
input n_2854;
input n_3672;
input n_3010;
input n_2499;
input n_4152;
input n_3533;
input n_3043;
input n_1622;
input n_1586;
input n_2543;
input n_2264;
input n_3464;
input n_302;
input n_1694;
input n_380;
input n_1535;
input n_3137;
input n_3382;
input n_2486;
input n_3132;
input n_3560;
input n_137;
input n_3723;
input n_2571;
input n_3138;
input n_1596;
input n_3177;
input n_20;
input n_1190;
input n_1734;
input n_3172;
input n_397;
input n_2902;
input n_3217;
input n_1983;
input n_1938;
input n_2498;
input n_4219;
input n_122;
input n_2220;
input n_2577;
input n_34;
input n_1262;
input n_2472;
input n_218;
input n_1891;
input n_2171;
input n_1213;
input n_3238;
input n_70;
input n_2235;
input n_3529;
input n_4193;
input n_3570;
input n_3394;
input n_2988;
input n_3136;
input n_1350;
input n_1673;
input n_3828;
input n_2232;
input n_1715;
input n_172;
input n_3536;
input n_4109;
input n_4192;
input n_1443;
input n_1272;
input n_2392;
input n_2894;
input n_3424;
input n_3957;
input n_4038;
input n_2790;
input n_4131;
input n_239;
input n_2037;
input n_97;
input n_2808;
input n_3710;
input n_4159;
input n_4195;
input n_3784;
input n_2298;
input n_782;
input n_2326;
input n_1539;
input n_490;
input n_3594;
input n_220;
input n_809;
input n_1043;
input n_3819;
input n_4090;
input n_3040;
input n_1797;
input n_3279;
input n_1608;
input n_4165;
input n_986;
input n_2305;
input n_2120;
input n_80;
input n_1472;
input n_2050;
input n_2373;
input n_2164;
input n_2402;
input n_2225;
input n_1081;
input n_3628;
input n_4144;
input n_402;
input n_1870;
input n_352;
input n_2964;
input n_4174;
input n_1692;
input n_800;
input n_1084;
input n_1171;
input n_460;
input n_2169;
input n_3485;
input n_4077;
input n_2371;
input n_1827;
input n_1361;
input n_1864;
input n_2006;
input n_3402;
input n_1491;
input n_2187;
input n_3475;
input n_662;
input n_3501;
input n_374;
input n_1152;
input n_1840;
input n_1705;
input n_3905;
input n_450;
input n_3262;
input n_3544;
input n_4150;
input n_2904;
input n_4008;
input n_2244;
input n_4290;
input n_3013;
input n_3356;
input n_2586;
input n_1684;
input n_921;
input n_2446;
input n_1346;
input n_711;
input n_1642;
input n_579;
input n_1352;
input n_2789;
input n_3105;
input n_3210;
input n_2872;
input n_937;
input n_2257;
input n_3692;
input n_3845;
input n_1682;
input n_2017;
input n_370;
input n_1695;
input n_1828;
input n_2046;
input n_2272;
input n_2699;
input n_2200;
input n_3029;
input n_4258;
input n_650;
input n_3597;
input n_1046;
input n_2560;
input n_1940;
input n_1979;
input n_2760;
input n_2704;
input n_3329;
input n_1145;
input n_330;
input n_1121;
input n_1102;
input n_1963;
input n_2738;
input n_972;
input n_1405;
input n_2376;
input n_258;
input n_3826;
input n_1406;
input n_456;
input n_3790;
input n_3878;
input n_2766;
input n_1332;
input n_260;
input n_2670;
input n_313;
input n_2700;
input n_624;
input n_962;
input n_1041;
input n_2346;
input n_565;
input n_3134;
input n_3647;
input n_356;
input n_1569;
input n_3681;
input n_936;
input n_3045;
input n_3115;
input n_1883;
input n_3821;
input n_1288;
input n_4300;
input n_3318;
input n_1186;
input n_1062;
input n_885;
input n_896;
input n_83;
input n_3278;
input n_2342;
input n_2167;
input n_2084;
input n_2970;
input n_3676;
input n_2882;
input n_3666;
input n_3675;
input n_4017;
input n_4260;
input n_3320;
input n_2541;
input n_654;
input n_2940;
input n_411;
input n_2518;
input n_2458;
input n_152;
input n_1222;
input n_599;
input n_776;
input n_321;
input n_1823;
input n_2479;
input n_3050;
input n_3350;
input n_105;
input n_2782;
input n_3977;
input n_227;
input n_1974;
input n_3988;
input n_4122;
input n_2673;
input n_2456;
input n_1720;
input n_3476;
input n_2527;
input n_204;
input n_482;
input n_934;
input n_1637;
input n_2635;
input n_3307;
input n_3439;
input n_1407;
input n_1795;
input n_2768;
input n_3588;
input n_4135;
input n_2871;
input n_4209;
input n_4279;
input n_420;
input n_2688;
input n_1341;
input n_394;
input n_1456;
input n_1845;
input n_3858;
input n_4183;
input n_1489;
input n_4321;
input n_4298;
input n_164;
input n_2314;
input n_3502;
input n_23;
input n_942;
input n_3003;
input n_2798;
input n_2852;
input n_1524;
input n_4128;
input n_543;
input n_2229;
input n_1964;
input n_4133;
input n_2288;
input n_1920;
input n_2753;
input n_2099;
input n_1496;
input n_1271;
input n_3292;
input n_1545;
input n_4145;
input n_2007;
input n_3121;
input n_2039;
input n_3388;
input n_4271;
input n_1946;
input n_1355;
input n_4181;
input n_1225;
input n_3184;
input n_1544;
input n_1485;
input n_2258;
input n_325;
input n_1640;
input n_4040;
input n_804;
input n_464;
input n_1846;
input n_3437;
input n_3245;
input n_3075;
input n_2406;
input n_4111;
input n_533;
input n_2390;
input n_4007;
input n_806;
input n_3712;
input n_879;
input n_959;
input n_2310;
input n_2506;
input n_584;
input n_2141;
input n_2562;
input n_244;
input n_2642;
input n_4312;
input n_1343;
input n_1522;
input n_76;
input n_4239;
input n_2734;
input n_548;
input n_1782;
input n_94;
input n_282;
input n_2383;
input n_4184;
input n_2626;
input n_1676;
input n_833;
input n_1830;
input n_2351;
input n_1567;
input n_4037;
input n_523;
input n_1319;
input n_707;
input n_2986;
input n_345;
input n_1900;
input n_3930;
input n_3246;
input n_799;
input n_1548;
input n_3381;
input n_3044;
input n_3562;
input n_2973;
input n_1155;
input n_2536;
input n_3915;
input n_139;
input n_2196;
input n_41;
input n_2629;
input n_3665;
input n_273;
input n_1633;
input n_2195;
input n_3208;
input n_2809;
input n_3007;
input n_787;
input n_2172;
input n_3528;
input n_3489;
input n_2835;
input n_1416;
input n_1528;
input n_2820;
input n_2293;
input n_1146;
input n_3698;
input n_2021;
input n_3355;
input n_2454;
input n_2114;
input n_3074;
input n_3174;
input n_159;
input n_1086;
input n_1066;
input n_3102;
input n_1948;
input n_157;
input n_2125;
input n_2026;
input n_4215;
input n_1282;
input n_2561;
input n_550;
input n_3321;
input n_2567;
input n_2322;
input n_275;
input n_652;
input n_2154;
input n_2727;
input n_2962;
input n_3377;
input n_2939;
input n_560;
input n_1906;
input n_1484;
input n_2992;
input n_3305;
input n_1241;
input n_1321;
input n_1672;
input n_569;
input n_2533;
input n_3157;
input n_3530;
input n_4185;
input n_1758;
input n_3221;
input n_3267;
input n_3752;
input n_2283;
input n_2869;
input n_2422;
input n_1925;
input n_737;
input n_1318;
input n_1914;
input n_1235;
input n_3457;
input n_1229;
input n_2759;
input n_3517;
input n_2945;
input n_3061;
input n_3893;
input n_2361;
input n_306;
input n_1292;
input n_1373;
input n_21;
input n_3762;
input n_3469;
input n_3932;
input n_2266;
input n_2960;
input n_3958;
input n_3005;
input n_346;
input n_3;
input n_3985;
input n_2427;
input n_3151;
input n_3411;
input n_1029;
input n_4196;
input n_3779;
input n_1447;
input n_2388;
input n_3984;
input n_2056;
input n_790;
input n_2611;
input n_2901;
input n_138;
input n_3258;
input n_1706;
input n_4242;
input n_3389;
input n_1498;
input n_3143;
input n_2653;
input n_2417;
input n_4232;
input n_4190;
input n_3000;
input n_1210;
input n_49;
input n_299;
input n_1248;
input n_1556;
input n_902;
input n_333;
input n_2189;
input n_2680;
input n_4052;
input n_2246;
input n_1047;
input n_3149;
input n_3375;
input n_3899;
input n_4084;
input n_3558;
input n_1984;
input n_3365;
input n_2236;
input n_1385;
input n_3713;
input n_431;
input n_3379;
input n_3156;
input n_24;
input n_459;
input n_1269;
input n_1931;
input n_2083;
input n_2834;
input n_3207;
input n_502;
input n_2668;
input n_672;
input n_2441;
input n_1257;
input n_3008;
input n_1751;
input n_3401;
input n_2840;
input n_3197;
input n_3242;
input n_285;
input n_3939;
input n_1375;
input n_1941;
input n_3483;
input n_3613;
input n_3972;
input n_4153;
input n_85;
input n_2128;
input n_655;
input n_706;
input n_1045;
input n_1650;
input n_786;
input n_1794;
input n_1236;
input n_1962;
input n_1559;
input n_1725;
input n_1928;
input n_2398;
input n_3743;
input n_3855;
input n_1872;
input n_3091;
input n_4317;
input n_834;
input n_19;
input n_29;
input n_2695;
input n_4035;
input n_3818;
input n_75;
input n_4269;
input n_743;
input n_766;
input n_3124;
input n_430;
input n_1741;
input n_1325;
input n_1002;
input n_1746;
input n_4088;
input n_1949;
input n_3398;
input n_3761;
input n_3759;
input n_545;
input n_3524;
input n_2671;
input n_489;
input n_2761;
input n_2885;
input n_2793;
input n_2715;
input n_2888;
input n_1804;
input n_2923;
input n_3711;
input n_3776;
input n_4235;
input n_1727;
input n_251;
input n_2508;
input n_1019;
input n_636;
input n_4301;
input n_3511;
input n_2054;
input n_4143;
input n_4170;
input n_729;
input n_110;
input n_151;
input n_876;
input n_774;
input n_3744;
input n_3642;
input n_2845;
input n_1337;
input n_3097;
input n_660;
input n_2062;
input n_2041;
input n_2975;
input n_438;
input n_1477;
input n_1360;
input n_2839;
input n_1860;
input n_2856;
input n_1904;
input n_2874;
input n_1200;
input n_2070;
input n_2588;
input n_479;
input n_3814;
input n_1607;
input n_3781;
input n_1353;
input n_1777;
input n_1908;
input n_1454;
input n_2484;
input n_2348;
input n_2944;
input n_2614;
input n_2126;
input n_3831;
input n_869;
input n_1154;
input n_3308;
input n_1113;
input n_1600;
input n_2833;
input n_2253;
input n_2758;
input n_3843;
input n_2366;
input n_646;
input n_528;
input n_391;
input n_1098;
input n_3694;
input n_2937;
input n_1329;
input n_2045;
input n_817;
input n_2261;
input n_3687;
input n_2216;
input n_3589;
input n_2210;
input n_262;
input n_3602;
input n_187;
input n_897;
input n_846;
input n_3300;
input n_2978;
input n_2066;
input n_3543;
input n_841;
input n_1476;
input n_3621;
input n_2516;
input n_3391;
input n_1001;
input n_508;
input n_1800;
input n_2241;
input n_1050;
input n_1411;
input n_1463;
input n_2903;
input n_3777;
input n_2827;
input n_1177;
input n_3216;
input n_3458;
input n_332;
input n_3515;
input n_1150;
input n_4203;
input n_3808;
input n_1742;
input n_3190;
input n_1562;
input n_1690;
input n_398;
input n_1191;
input n_1826;
input n_566;
input n_1023;
input n_1882;
input n_2951;
input n_1076;
input n_1118;
input n_194;
input n_2949;
input n_3726;
input n_57;
input n_1007;
input n_1807;
input n_1929;
input n_1378;
input n_2369;
input n_855;
input n_1592;
input n_1759;
input n_2719;
input n_1814;
input n_1631;
input n_52;
input n_591;
input n_1377;
input n_3758;
input n_1879;
input n_256;
input n_853;
input n_440;
input n_695;
input n_3806;
input n_4081;
input n_1542;
input n_2587;
input n_3199;
input n_2931;
input n_875;
input n_209;
input n_367;
input n_680;
input n_3339;
input n_1678;
input n_2569;
input n_661;
input n_2400;
input n_1716;
input n_3866;
input n_278;
input n_3787;
input n_1256;
input n_3585;
input n_671;
input n_3565;
input n_1953;
input n_7;
input n_933;
input n_740;
input n_703;
input n_3343;
input n_3303;
input n_978;
input n_4157;
input n_2752;
input n_4173;
input n_384;
input n_3135;
input n_1976;
input n_4229;
input n_2905;
input n_1291;
input n_1217;
input n_3990;
input n_751;
input n_749;
input n_3865;
input n_1824;
input n_310;
input n_3954;
input n_1628;
input n_4073;
input n_1324;
input n_3890;
input n_1399;
input n_2122;
input n_2109;
input n_3629;
input n_1435;
input n_3920;
input n_969;
input n_988;
input n_2140;
input n_3503;
input n_3160;
input n_1065;
input n_2796;
input n_3255;
input n_2507;
input n_84;
input n_1401;
input n_2358;
input n_1255;
input n_568;
input n_3658;
input n_1516;
input n_143;
input n_1536;
input n_3846;
input n_180;
input n_2163;
input n_2186;
input n_3512;
input n_2029;
input n_2815;
input n_1204;
input n_3951;
input n_3034;
input n_823;
input n_1132;
input n_643;
input n_233;
input n_698;
input n_1074;
input n_1394;
input n_3569;
input n_1327;
input n_1326;
input n_739;
input n_400;
input n_955;
input n_337;
input n_3874;
input n_1379;
input n_2528;
input n_2814;
input n_214;
input n_246;
input n_2787;
input n_1338;
input n_1097;
input n_2969;
input n_2395;
input n_935;
input n_3027;
input n_781;
input n_789;
input n_1554;
input n_3231;
input n_4083;
input n_1130;
input n_3083;
input n_4212;
input n_2979;
input n_181;
input n_1810;
input n_182;
input n_2953;
input n_573;
input n_769;
input n_2380;
input n_676;
input n_327;
input n_4295;
input n_1120;
input n_832;
input n_1583;
input n_3049;
input n_1730;
input n_2295;
input n_555;
input n_389;
input n_814;
input n_2746;
input n_2946;
input n_1643;
input n_2020;
input n_2500;
input n_3430;
input n_2269;
input n_1729;
input n_669;
input n_2290;
input n_4225;
input n_4171;
input n_2048;
input n_3652;
input n_176;
input n_114;
input n_300;
input n_222;
input n_3830;
input n_3679;
input n_2005;
input n_747;
input n_3541;
input n_74;
input n_2565;
input n_4023;
input n_1389;
input n_1105;
input n_3117;
input n_721;
input n_1461;
input n_742;
input n_3432;
input n_535;
input n_691;
input n_3617;
input n_372;
input n_2076;
input n_2736;
input n_111;
input n_2883;
input n_3583;
input n_314;
input n_3860;
input n_1408;
input n_378;
input n_3851;
input n_3567;
input n_1196;
input n_4282;
input n_377;
input n_1598;
input n_3493;
input n_2935;
input n_4046;
input n_3807;
input n_863;
input n_3015;
input n_2175;
input n_601;
input n_2182;
input n_3774;
input n_338;
input n_2910;
input n_1283;
input n_2385;
input n_4112;
input n_918;
input n_748;
input n_506;
input n_1114;
input n_1785;
input n_56;
input n_763;
input n_1147;
input n_1848;
input n_360;
input n_1754;
input n_2149;
input n_3057;
input n_3154;
input n_3701;
input n_2396;
input n_1506;
input n_119;
input n_2584;
input n_1652;
input n_1812;
input n_957;
input n_1994;
input n_3473;
input n_895;
input n_866;
input n_1227;
input n_2450;
input n_2485;
input n_3739;
input n_2284;
input n_3898;
input n_3520;
input n_191;
input n_2566;
input n_387;
input n_2287;
input n_452;
input n_744;
input n_971;
input n_2702;
input n_3241;
input n_946;
input n_344;
input n_2906;
input n_761;
input n_1303;
input n_2769;
input n_3622;
input n_1205;
input n_2492;
input n_1258;
input n_3778;
input n_4095;
input n_2438;
input n_2914;
input n_1392;
input n_174;
input n_1173;
input n_1924;
input n_525;
input n_2463;
input n_3363;
input n_2881;
input n_1677;
input n_1116;
input n_611;
input n_1570;
input n_1702;
input n_1219;
input n_3551;
input n_3064;
input n_1780;
input n_3100;
input n_3897;
input n_3721;
input n_1689;
input n_8;
input n_2180;
input n_3372;
input n_2858;
input n_3062;
input n_2679;
input n_1174;
input n_3573;
input n_1944;
input n_1016;
input n_1347;
input n_4106;
input n_795;
input n_1501;
input n_3604;
input n_1221;
input n_3334;
input n_4027;
input n_1245;
input n_838;
input n_3215;
input n_3969;
input n_129;
input n_3336;
input n_647;
input n_4160;
input n_197;
input n_4231;
input n_844;
input n_17;
input n_448;
input n_2952;
input n_1017;
input n_3068;
input n_3853;
input n_2117;
input n_2234;
input n_4256;
input n_2779;
input n_2685;
input n_3823;
input n_1083;
input n_109;
input n_445;
input n_3553;
input n_1561;
input n_2741;
input n_3114;
input n_930;
input n_888;
input n_2275;
input n_1112;
input n_2465;
input n_2620;
input n_2081;
input n_2168;
input n_2568;
input n_234;
input n_2022;
input n_1945;
input n_2203;
input n_910;
input n_3811;
input n_1656;
input n_1721;
input n_1460;
input n_911;
input n_2112;
input n_2255;
input n_82;
input n_1464;
input n_27;
input n_236;
input n_653;
input n_1737;
input n_2430;
input n_1414;
input n_3486;
input n_4086;
input n_752;
input n_908;
input n_2649;
input n_2721;
input n_944;
input n_3556;
input n_2034;
input n_576;
input n_1028;
input n_3836;
input n_2106;
input n_472;
input n_2862;
input n_270;
input n_2265;
input n_2615;
input n_414;
input n_2683;
input n_1922;
input n_563;
input n_4068;
input n_2032;
input n_2744;
input n_4309;
input n_1011;
input n_2474;
input n_3703;
input n_1566;
input n_1215;
input n_2437;
input n_25;
input n_93;
input n_839;
input n_2444;
input n_2743;
input n_3962;
input n_708;
input n_1973;
input n_3181;
input n_2267;
input n_3456;
input n_3035;
input n_668;
input n_4166;
input n_626;
input n_990;
input n_1500;
input n_779;
input n_1537;
input n_1821;
input n_2205;
input n_3699;
input n_4243;
input n_3204;
input n_1104;
input n_854;
input n_1058;
input n_3378;
input n_4025;
input n_2312;
input n_498;
input n_3404;
input n_1122;
input n_870;
input n_904;
input n_1253;
input n_709;
input n_1266;
input n_366;
input n_2242;
input n_3362;
input n_3745;
input n_4059;
input n_1509;
input n_103;
input n_4188;
input n_3328;
input n_1693;
input n_2934;
input n_3667;
input n_3290;
input n_4121;
input n_1109;
input n_3523;
input n_185;
input n_2222;
input n_712;
input n_3256;
input n_348;
input n_1276;
input n_3802;
input n_3868;
input n_3176;
input n_376;
input n_3309;
input n_3671;
input n_2015;
input n_2118;
input n_4142;
input n_2111;
input n_2466;
input n_390;
input n_3982;
input n_4266;
input n_2915;
input n_2530;
input n_1148;
input n_31;
input n_2188;
input n_2505;
input n_334;
input n_1989;
input n_1161;
input n_2609;
input n_1085;
input n_232;
input n_2802;
input n_3796;
input n_2999;
input n_4115;
input n_3840;
input n_2014;
input n_2042;
input n_46;
input n_1239;
input n_3643;
input n_3697;
input n_771;
input n_1584;
input n_2425;
input n_470;
input n_475;
input n_924;
input n_3408;
input n_3461;
input n_298;
input n_1582;
input n_492;
input n_3680;
input n_4265;
input n_2318;
input n_3286;
input n_4012;
input n_2408;
input n_4246;
input n_1149;
input n_3170;
input n_3513;
input n_265;
input n_3468;
input n_3690;
input n_1184;
input n_3645;
input n_2483;
input n_2950;
input n_228;
input n_719;
input n_1972;
input n_3060;
input n_3304;
input n_3682;
input n_2592;
input n_3771;
input n_1525;
input n_3098;
input n_3995;
input n_4076;
input n_2594;
input n_455;
input n_2666;
input n_4105;
input n_1585;
input n_1851;
input n_363;
input n_1799;
input n_1090;
input n_2147;
input n_2564;
input n_592;
input n_4244;
input n_1816;
input n_4064;
input n_2503;
input n_2433;
input n_1518;
input n_4049;
input n_829;
input n_1156;
input n_1362;
input n_4259;
input n_3123;
input n_393;
input n_984;
input n_2600;
input n_3380;
input n_1829;
input n_503;
input n_2035;
input n_3508;
input n_3024;
input n_1450;
input n_1638;
input n_3422;
input n_132;
input n_868;
input n_3038;
input n_570;
input n_859;
input n_2033;
input n_406;
input n_3086;
input n_735;
input n_4104;
input n_1789;
input n_2531;
input n_1770;
input n_878;
input n_620;
input n_130;
input n_3285;
input n_519;
input n_4208;
input n_2523;
input n_307;
input n_469;
input n_1218;
input n_2413;
input n_500;
input n_3769;
input n_1482;
input n_3361;
input n_981;
input n_3596;
input n_714;
input n_3478;
input n_3936;
input n_1349;
input n_291;
input n_4089;
input n_1144;
input n_2071;
input n_3669;
input n_3863;
input n_357;
input n_3219;
input n_2429;
input n_3130;
input n_3702;
input n_985;
input n_4316;
input n_2233;
input n_2440;
input n_2723;
input n_481;
input n_3521;
input n_3233;
input n_997;
input n_1710;
input n_2800;
input n_2161;
input n_3496;
input n_1301;
input n_2805;
input n_802;
input n_561;
input n_33;
input n_3310;
input n_980;
input n_2681;
input n_1306;
input n_3264;
input n_2010;
input n_2282;
input n_1651;
input n_1198;
input n_3096;
input n_2360;
input n_3764;
input n_2047;
input n_4061;
input n_2651;
input n_2095;
input n_3239;
input n_1609;
input n_2174;
input n_3161;
input n_2799;
input n_436;
input n_4075;
input n_116;
input n_3344;
input n_2334;
input n_3902;
input n_4062;
input n_3881;
input n_3295;
input n_3947;
input n_409;
input n_1244;
input n_1685;
input n_1763;
input n_1998;
input n_3066;
input n_1574;
input n_2426;
input n_2490;
input n_2844;
input n_3101;
input n_240;
input n_3989;
input n_756;
input n_2303;
input n_1619;
input n_2478;
input n_1981;
input n_2285;
input n_4233;
input n_1606;
input n_810;
input n_4108;
input n_1133;
input n_635;
input n_95;
input n_1194;
input n_3374;
input n_3786;
input n_3841;
input n_2742;
input n_2640;
input n_3695;
input n_4051;
input n_1051;
input n_253;
input n_3976;
input n_4254;
input n_1552;
input n_2918;
input n_583;
input n_3288;
input n_1996;
input n_3563;
input n_3992;
input n_2367;
input n_4307;
input n_3876;
input n_249;
input n_201;
input n_2867;
input n_3198;
input n_1039;
input n_1442;
input n_3495;
input n_2726;
input n_1034;
input n_2043;
input n_4303;
input n_1480;
input n_3125;
input n_1158;
input n_2909;
input n_2248;
input n_754;
input n_4293;
input n_941;
input n_3552;
input n_975;
input n_3206;
input n_1031;
input n_115;
input n_1305;
input n_2363;
input n_2578;
input n_553;
input n_43;
input n_849;
input n_2662;
input n_3116;
input n_3147;
input n_3383;
input n_3709;
input n_753;
input n_3925;
input n_4091;
input n_1753;
input n_3095;
input n_3180;
input n_3738;
input n_3359;
input n_2795;
input n_3472;
input n_2471;
input n_4186;
input n_467;
input n_3187;
input n_2540;
input n_269;
input n_359;
input n_973;
input n_2807;
input n_1921;
input n_3218;
input n_3610;
input n_3618;
input n_3330;
input n_1479;
input n_1055;
input n_1675;
input n_2197;
input n_2217;
input n_582;
input n_2065;
input n_2879;
input n_861;
input n_3717;
input n_857;
input n_967;
input n_4148;
input n_571;
input n_2215;
input n_2461;
input n_271;
input n_404;
input n_2001;
input n_158;
input n_2107;
input n_1884;
input n_206;
input n_2040;
input n_679;
input n_4057;
input n_2968;
input n_4201;
input n_633;
input n_1170;
input n_665;
input n_1629;
input n_2221;
input n_588;
input n_4263;
input n_225;
input n_1260;
input n_308;
input n_309;
input n_1819;
input n_2055;
input n_3555;
input n_1010;
input n_3444;
input n_4210;
input n_2553;
input n_149;
input n_1040;
input n_915;
input n_632;
input n_3059;
input n_1166;
input n_2038;
input n_812;
input n_2891;
input n_1131;
input n_2634;
input n_1761;
input n_2709;
input n_3155;
input n_3445;
input n_534;
input n_1578;
input n_1006;
input n_1861;
input n_373;
input n_3110;
input n_87;
input n_1632;
input n_1890;
input n_3017;
input n_3955;
input n_1805;
input n_2477;
input n_257;
input n_1557;
input n_1888;
input n_2280;
input n_1833;
input n_3903;
input n_730;
input n_1311;
input n_3945;
input n_1494;
input n_2325;
input n_670;
input n_203;
input n_1850;
input n_1898;
input n_2443;
input n_2697;
input n_3235;
input n_3854;
input n_2308;
input n_4205;
input n_2162;
input n_3908;
input n_1868;
input n_207;
input n_2333;
input n_2079;
input n_3467;
input n_3001;
input n_3587;
input n_1089;
input n_4278;
input n_1887;
input n_1587;
input n_3916;
input n_3527;
input n_3795;
input n_2512;
input n_3950;
input n_3433;
input n_3852;
input n_1365;
input n_4138;
input n_1417;
input n_205;
input n_1242;
input n_2086;
input n_2185;
input n_2927;
input n_3673;
input n_1836;
input n_3833;
input n_4281;
input n_3815;
input n_2774;
input n_3896;
input n_3039;
input n_681;
input n_1226;
input n_3740;
input n_3162;
input n_1274;
input n_1486;
input n_2166;
input n_3094;
input n_412;
input n_2899;
input n_3274;
input n_3333;
input n_3186;
input n_640;
input n_1322;
input n_81;
input n_4129;
input n_965;
input n_1899;
input n_1428;
input n_4093;
input n_1616;
input n_1576;
input n_1856;
input n_1862;
input n_1958;
input n_2077;
input n_339;
input n_784;
input n_315;
input n_434;
input n_64;
input n_288;
input n_1059;
input n_1197;
input n_3065;
input n_3965;
input n_2632;
input n_422;
input n_2579;
input n_722;
input n_862;
input n_2105;
input n_135;
input n_3079;
input n_165;
input n_2098;
input n_3085;
input n_540;
input n_1423;
input n_2813;
input n_1935;
input n_3584;
input n_4039;
input n_3387;
input n_2027;
input n_457;
input n_3070;
input n_3800;
input n_2223;
input n_2091;
input n_364;
input n_3263;
input n_4197;
input n_3420;
input n_2991;
input n_1915;
input n_629;
input n_1621;
input n_4275;
input n_1748;
input n_2547;
input n_2415;
input n_4283;
input n_900;
input n_3504;
input n_4194;
input n_1449;
input n_531;
input n_827;
input n_2912;
input n_60;
input n_361;
input n_4272;
input n_2659;
input n_2930;
input n_1025;
input n_3409;
input n_2419;
input n_3111;
input n_2116;
input n_336;
input n_2320;
input n_12;
input n_1885;
input n_2677;
input n_1013;
input n_3182;
input n_1259;
input n_3054;
input n_3283;
input n_192;
input n_2183;
input n_3002;
input n_1538;
input n_51;
input n_649;
input n_4030;
input n_1612;
input n_1240;

output n_16688;

wire n_5643;
wire n_12335;
wire n_12949;
wire n_14428;
wire n_13611;
wire n_15214;
wire n_4452;
wire n_6566;
wire n_13045;
wire n_5172;
wire n_11173;
wire n_15268;
wire n_16218;
wire n_4649;
wire n_5315;
wire n_10487;
wire n_6872;
wire n_16664;
wire n_13998;
wire n_5254;
wire n_11926;
wire n_6441;
wire n_8668;
wire n_6806;
wire n_5362;
wire n_13146;
wire n_13235;
wire n_15125;
wire n_10587;
wire n_5019;
wire n_8713;
wire n_15450;
wire n_7111;
wire n_6141;
wire n_10960;
wire n_11111;
wire n_7933;
wire n_7967;
wire n_5138;
wire n_13522;
wire n_10931;
wire n_4388;
wire n_4395;
wire n_6960;
wire n_15609;
wire n_8169;
wire n_12265;
wire n_9002;
wire n_16423;
wire n_16335;
wire n_14670;
wire n_9130;
wire n_7180;
wire n_5653;
wire n_11574;
wire n_4978;
wire n_13530;
wire n_8604;
wire n_15049;
wire n_16362;
wire n_5409;
wire n_5301;
wire n_7263;
wire n_13125;
wire n_15181;
wire n_8168;
wire n_4829;
wire n_7190;
wire n_7504;
wire n_8186;
wire n_5393;
wire n_6725;
wire n_6126;
wire n_4699;
wire n_4686;
wire n_12322;
wire n_14318;
wire n_8899;
wire n_14196;
wire n_15971;
wire n_5524;
wire n_10236;
wire n_5345;
wire n_11205;
wire n_11776;
wire n_11678;
wire n_8023;
wire n_11802;
wire n_12251;
wire n_10053;
wire n_11650;
wire n_5818;
wire n_16307;
wire n_8005;
wire n_8130;
wire n_8534;
wire n_5963;
wire n_12179;
wire n_13942;
wire n_5055;
wire n_15294;
wire n_14439;
wire n_12570;
wire n_9896;
wire n_11856;
wire n_11905;
wire n_4868;
wire n_10020;
wire n_14825;
wire n_16288;
wire n_7116;
wire n_5267;
wire n_10202;
wire n_11536;
wire n_5950;
wire n_15295;
wire n_9104;
wire n_14914;
wire n_6999;
wire n_14741;
wire n_15665;
wire n_11046;
wire n_11079;
wire n_10283;
wire n_5548;
wire n_5057;
wire n_15581;
wire n_11065;
wire n_15445;
wire n_8339;
wire n_8272;
wire n_14215;
wire n_13997;
wire n_14402;
wire n_7161;
wire n_7868;
wire n_14882;
wire n_5838;
wire n_15764;
wire n_5725;
wire n_6324;
wire n_13437;
wire n_15623;
wire n_5229;
wire n_5325;
wire n_11051;
wire n_11214;
wire n_5101;
wire n_7000;
wire n_8561;
wire n_14998;
wire n_14944;
wire n_11954;
wire n_7398;
wire n_14232;
wire n_10392;
wire n_14341;
wire n_12882;
wire n_5900;
wire n_15074;
wire n_5545;
wire n_12617;
wire n_8411;
wire n_8499;
wire n_8236;
wire n_5102;
wire n_15253;
wire n_15356;
wire n_13137;
wire n_13221;
wire n_6882;
wire n_4501;
wire n_9626;
wire n_10775;
wire n_11163;
wire n_15933;
wire n_9526;
wire n_13657;
wire n_15571;
wire n_6325;
wire n_4724;
wire n_9840;
wire n_14099;
wire n_5598;
wire n_15632;
wire n_7983;
wire n_10348;
wire n_10863;
wire n_12495;
wire n_9581;
wire n_15898;
wire n_16245;
wire n_7389;
wire n_4997;
wire n_10719;
wire n_9018;
wire n_4843;
wire n_11419;
wire n_8070;
wire n_12095;
wire n_13663;
wire n_13990;
wire n_16302;
wire n_4696;
wire n_6660;
wire n_13298;
wire n_9055;
wire n_4347;
wire n_14939;
wire n_11740;
wire n_5259;
wire n_6913;
wire n_8444;
wire n_10015;
wire n_13993;
wire n_10986;
wire n_7802;
wire n_6948;
wire n_5819;
wire n_7008;
wire n_12392;
wire n_15353;
wire n_8366;
wire n_8102;
wire n_9362;
wire n_11979;
wire n_7401;
wire n_7516;
wire n_7596;
wire n_6280;
wire n_6629;
wire n_12767;
wire n_5279;
wire n_15993;
wire n_5894;
wire n_16095;
wire n_10759;
wire n_8022;
wire n_5930;
wire n_9036;
wire n_9551;
wire n_13210;
wire n_10262;
wire n_8175;
wire n_8977;
wire n_9658;
wire n_5239;
wire n_8953;
wire n_8426;
wire n_5354;
wire n_10239;
wire n_14577;
wire n_5332;
wire n_14984;
wire n_15797;
wire n_9962;
wire n_5908;
wire n_4814;
wire n_10373;
wire n_11104;
wire n_8913;
wire n_9525;
wire n_10816;
wire n_9725;
wire n_4956;
wire n_11537;
wire n_14699;
wire n_13814;
wire n_12707;
wire n_14861;
wire n_7686;
wire n_6914;
wire n_10335;
wire n_5337;
wire n_15194;
wire n_15362;
wire n_5129;
wire n_11301;
wire n_12424;
wire n_13681;
wire n_14121;
wire n_15101;
wire n_5420;
wire n_15572;
wire n_5070;
wire n_10381;
wire n_6243;
wire n_4414;
wire n_6585;
wire n_11703;
wire n_16553;
wire n_11699;
wire n_6374;
wire n_4646;
wire n_7651;
wire n_11543;
wire n_10947;
wire n_6628;
wire n_8125;
wire n_13483;
wire n_6015;
wire n_14662;
wire n_11261;
wire n_14811;
wire n_10226;
wire n_16012;
wire n_13247;
wire n_16286;
wire n_6526;
wire n_13929;
wire n_16551;
wire n_7956;
wire n_7369;
wire n_6570;
wire n_16549;
wire n_8556;
wire n_7196;
wire n_15421;
wire n_10767;
wire n_5136;
wire n_8040;
wire n_14646;
wire n_15964;
wire n_11821;
wire n_14095;
wire n_5638;
wire n_13121;
wire n_13989;
wire n_9100;
wire n_14864;
wire n_15069;
wire n_6784;
wire n_16643;
wire n_12107;
wire n_14520;
wire n_10755;
wire n_4950;
wire n_14780;
wire n_10868;
wire n_9067;
wire n_10161;
wire n_9842;
wire n_4729;
wire n_11447;
wire n_6323;
wire n_9614;
wire n_14431;
wire n_15200;
wire n_13515;
wire n_10682;
wire n_6110;
wire n_11684;
wire n_12652;
wire n_16024;
wire n_16324;
wire n_6371;
wire n_14410;
wire n_8079;
wire n_10699;
wire n_15507;
wire n_4751;
wire n_7846;
wire n_8595;
wire n_15800;
wire n_9400;
wire n_5151;
wire n_8142;
wire n_11627;
wire n_5684;
wire n_8598;
wire n_13139;
wire n_15887;
wire n_10022;
wire n_5729;
wire n_7256;
wire n_13803;
wire n_6404;
wire n_12209;
wire n_7331;
wire n_16078;
wire n_14066;
wire n_7774;
wire n_7856;
wire n_15600;
wire n_16267;
wire n_6674;
wire n_5680;
wire n_13606;
wire n_6148;
wire n_6951;
wire n_11659;
wire n_15899;
wire n_7625;
wire n_13501;
wire n_9106;
wire n_13509;
wire n_12775;
wire n_13729;
wire n_4662;
wire n_8869;
wire n_6989;
wire n_4671;
wire n_7863;
wire n_8381;
wire n_5504;
wire n_5522;
wire n_5828;
wire n_7342;
wire n_14813;
wire n_9520;
wire n_14791;
wire n_8958;
wire n_14485;
wire n_14931;
wire n_12833;
wire n_5099;
wire n_12090;
wire n_6896;
wire n_14628;
wire n_7770;
wire n_10606;
wire n_8421;
wire n_11164;
wire n_13687;
wire n_7623;
wire n_6968;
wire n_7217;
wire n_16268;
wire n_12371;
wire n_10114;
wire n_12203;
wire n_10357;
wire n_14540;
wire n_15762;
wire n_7147;
wire n_8115;
wire n_4507;
wire n_16351;
wire n_15883;
wire n_8389;
wire n_9398;
wire n_5902;
wire n_11497;
wire n_14900;
wire n_15320;
wire n_12359;
wire n_4677;
wire n_12915;
wire n_5063;
wire n_6196;
wire n_9037;
wire n_15983;
wire n_13149;
wire n_13711;
wire n_15846;
wire n_13454;
wire n_5275;
wire n_5306;
wire n_12548;
wire n_15874;
wire n_12742;
wire n_16662;
wire n_14091;
wire n_9042;
wire n_15755;
wire n_11768;
wire n_8412;
wire n_9267;
wire n_6485;
wire n_14478;
wire n_8987;
wire n_11805;
wire n_14461;
wire n_10177;
wire n_6107;
wire n_9652;
wire n_5493;
wire n_8849;
wire n_11944;
wire n_9059;
wire n_13958;
wire n_14935;
wire n_15332;
wire n_5346;
wire n_4366;
wire n_5252;
wire n_5309;
wire n_7796;
wire n_6282;
wire n_6863;
wire n_6994;
wire n_12770;
wire n_10012;
wire n_14570;
wire n_15986;
wire n_16068;
wire n_13754;
wire n_12985;
wire n_4698;
wire n_13797;
wire n_4445;
wire n_13013;
wire n_13238;
wire n_4810;
wire n_7564;
wire n_11635;
wire n_16254;
wire n_14989;
wire n_15434;
wire n_16530;
wire n_9446;
wire n_11129;
wire n_12951;
wire n_14171;
wire n_16191;
wire n_10204;
wire n_6768;
wire n_9453;
wire n_6383;
wire n_7234;
wire n_4456;
wire n_8119;
wire n_10296;
wire n_8641;
wire n_11637;
wire n_12988;
wire n_15212;
wire n_15977;
wire n_8151;
wire n_8118;
wire n_12393;
wire n_16442;
wire n_9718;
wire n_9128;
wire n_10281;
wire n_13344;
wire n_9038;
wire n_9872;
wire n_10310;
wire n_11139;
wire n_14380;
wire n_16004;
wire n_8748;
wire n_13984;
wire n_8436;
wire n_5452;
wire n_12685;
wire n_14239;
wire n_6794;
wire n_6151;
wire n_15896;
wire n_8718;
wire n_7110;
wire n_5476;
wire n_12831;
wire n_13920;
wire n_9935;
wire n_6431;
wire n_6990;
wire n_8659;
wire n_14045;
wire n_14288;
wire n_14824;
wire n_10097;
wire n_8223;
wire n_4856;
wire n_15767;
wire n_4369;
wire n_9135;
wire n_7849;
wire n_8915;
wire n_12667;
wire n_15635;
wire n_4331;
wire n_7297;
wire n_10018;
wire n_9866;
wire n_15183;
wire n_16509;
wire n_4972;
wire n_7298;
wire n_4993;
wire n_15118;
wire n_5536;
wire n_9129;
wire n_9858;
wire n_10141;
wire n_12427;
wire n_7533;
wire n_14162;
wire n_13771;
wire n_7221;
wire n_4375;
wire n_13977;
wire n_10656;
wire n_15159;
wire n_16026;
wire n_6575;
wire n_6055;
wire n_8727;
wire n_8224;
wire n_11295;
wire n_5130;
wire n_16538;
wire n_11662;
wire n_13960;
wire n_8246;
wire n_5532;
wire n_5897;
wire n_8952;
wire n_4613;
wire n_15679;
wire n_13014;
wire n_9070;
wire n_11708;
wire n_10266;
wire n_15629;
wire n_14401;
wire n_5609;
wire n_4717;
wire n_10897;
wire n_10827;
wire n_4877;
wire n_5922;
wire n_15154;
wire n_14922;
wire n_10449;
wire n_7569;
wire n_7823;
wire n_7734;
wire n_7062;
wire n_7861;
wire n_8955;
wire n_9477;
wire n_5658;
wire n_4731;
wire n_9680;
wire n_12172;
wire n_12147;
wire n_12923;
wire n_14769;
wire n_7039;
wire n_8577;
wire n_12384;
wire n_14961;
wire n_11349;
wire n_8594;
wire n_5046;
wire n_13227;
wire n_8428;
wire n_9829;
wire n_15438;
wire n_11260;
wire n_8848;
wire n_12825;
wire n_13341;
wire n_5058;
wire n_10685;
wire n_11351;
wire n_4467;
wire n_15185;
wire n_12083;
wire n_7077;
wire n_12014;
wire n_14803;
wire n_5667;
wire n_8259;
wire n_12540;
wire n_15611;
wire n_10607;
wire n_14388;
wire n_15490;
wire n_5865;
wire n_15182;
wire n_12249;
wire n_8349;
wire n_16035;
wire n_6836;
wire n_5305;
wire n_5042;
wire n_14977;
wire n_11998;
wire n_4681;
wire n_8164;
wire n_13239;
wire n_10628;
wire n_4752;
wire n_13429;
wire n_15942;
wire n_7905;
wire n_5281;
wire n_8776;
wire n_11775;
wire n_15100;
wire n_9143;
wire n_8287;
wire n_10769;
wire n_10256;
wire n_7753;
wire n_10368;
wire n_6771;
wire n_14732;
wire n_7950;
wire n_9947;
wire n_16659;
wire n_13999;
wire n_9088;
wire n_8607;
wire n_14037;
wire n_10138;
wire n_12117;
wire n_11706;
wire n_6248;
wire n_11800;
wire n_16134;
wire n_10183;
wire n_10375;
wire n_6952;
wire n_14535;
wire n_6795;
wire n_5314;
wire n_10452;
wire n_11464;
wire n_7806;
wire n_12960;
wire n_14878;
wire n_14094;
wire n_15928;
wire n_13033;
wire n_11642;
wire n_15046;
wire n_4381;
wire n_11143;
wire n_15703;
wire n_16092;
wire n_7595;
wire n_5144;
wire n_7648;
wire n_10383;
wire n_4466;
wire n_4418;
wire n_8066;
wire n_6831;
wire n_11074;
wire n_16352;
wire n_12131;
wire n_4510;
wire n_6776;
wire n_12851;
wire n_5795;
wire n_11934;
wire n_12349;
wire n_4473;
wire n_6043;
wire n_5552;
wire n_7452;
wire n_14282;
wire n_5226;
wire n_9269;
wire n_10320;
wire n_6715;
wire n_6714;
wire n_15518;
wire n_11308;
wire n_13550;
wire n_16266;
wire n_14217;
wire n_7677;
wire n_10903;
wire n_5457;
wire n_13348;
wire n_8416;
wire n_10396;
wire n_13919;
wire n_4518;
wire n_10724;
wire n_13642;
wire n_16398;
wire n_8404;
wire n_8997;
wire n_6584;
wire n_15574;
wire n_11084;
wire n_14062;
wire n_9988;
wire n_7009;
wire n_8453;
wire n_10693;
wire n_14167;
wire n_12740;
wire n_9113;
wire n_7149;
wire n_5291;
wire n_10363;
wire n_15872;
wire n_13240;
wire n_8949;
wire n_10831;
wire n_9131;
wire n_11553;
wire n_12578;
wire n_12795;
wire n_10517;
wire n_4589;
wire n_10323;
wire n_12194;
wire n_13623;
wire n_10842;
wire n_7519;
wire n_16465;
wire n_7400;
wire n_10876;
wire n_11511;
wire n_15833;
wire n_9137;
wire n_15649;
wire n_11180;
wire n_14043;
wire n_9724;
wire n_11146;
wire n_16046;
wire n_9281;
wire n_10883;
wire n_8995;
wire n_10101;
wire n_15863;
wire n_9393;
wire n_15974;
wire n_4394;
wire n_6581;
wire n_13845;
wire n_12709;
wire n_6010;
wire n_13432;
wire n_8711;
wire n_7013;
wire n_12771;
wire n_14150;
wire n_5343;
wire n_12125;
wire n_12505;
wire n_7290;
wire n_12278;
wire n_13721;
wire n_10820;
wire n_13514;
wire n_4921;
wire n_9687;
wire n_14787;
wire n_4329;
wire n_5135;
wire n_7303;
wire n_6616;
wire n_8306;
wire n_10123;
wire n_10781;
wire n_7488;
wire n_7315;
wire n_13194;
wire n_9886;
wire n_10651;
wire n_8887;
wire n_9426;
wire n_4697;
wire n_13244;
wire n_16183;
wire n_11866;
wire n_6185;
wire n_11450;
wire n_13575;
wire n_12522;
wire n_5529;
wire n_15659;
wire n_7889;
wire n_10943;
wire n_12344;
wire n_6042;
wire n_13843;
wire n_9102;
wire n_11526;
wire n_13404;
wire n_9578;
wire n_16115;
wire n_5183;
wire n_13109;
wire n_8500;
wire n_14785;
wire n_7438;
wire n_16631;
wire n_14355;
wire n_14128;
wire n_7268;
wire n_7337;
wire n_11851;
wire n_4964;
wire n_9489;
wire n_12804;
wire n_14123;
wire n_5957;
wire n_6965;
wire n_12116;
wire n_10728;
wire n_6357;
wire n_9144;
wire n_10094;
wire n_6800;
wire n_10084;
wire n_4636;
wire n_10468;
wire n_14126;
wire n_14105;
wire n_7461;
wire n_8285;
wire n_13870;
wire n_4322;
wire n_10655;
wire n_13791;
wire n_9797;
wire n_15133;
wire n_6955;
wire n_8483;
wire n_4946;
wire n_4767;
wire n_9521;
wire n_15288;
wire n_8332;
wire n_9478;
wire n_9932;
wire n_13040;
wire n_7278;
wire n_11370;
wire n_6509;
wire n_13900;
wire n_16224;
wire n_4576;
wire n_7454;
wire n_11253;
wire n_14652;
wire n_11379;
wire n_15527;
wire n_16627;
wire n_10670;
wire n_5929;
wire n_12861;
wire n_9020;
wire n_4615;
wire n_5787;
wire n_11981;
wire n_16146;
wire n_16654;
wire n_9895;
wire n_8741;
wire n_12918;
wire n_16452;
wire n_9351;
wire n_11585;
wire n_5445;
wire n_13140;
wire n_13962;
wire n_14556;
wire n_5501;
wire n_4389;
wire n_5342;
wire n_7232;
wire n_6839;
wire n_7377;
wire n_4345;
wire n_13753;
wire n_16132;
wire n_6646;
wire n_13353;
wire n_8648;
wire n_12388;
wire n_12102;
wire n_9189;
wire n_15149;
wire n_16528;
wire n_15365;
wire n_4664;
wire n_13716;
wire n_14844;
wire n_14701;
wire n_7098;
wire n_7069;
wire n_12560;
wire n_14391;
wire n_7904;
wire n_11691;
wire n_16587;
wire n_6033;
wire n_11541;
wire n_15495;
wire n_13610;
wire n_8851;
wire n_8921;
wire n_4873;
wire n_9410;
wire n_9801;
wire n_13332;
wire n_5748;
wire n_14408;
wire n_15293;
wire n_9356;
wire n_15880;
wire n_12865;
wire n_16499;
wire n_8773;
wire n_6097;
wire n_6369;
wire n_10712;
wire n_8394;
wire n_11155;
wire n_5076;
wire n_5870;
wire n_4713;
wire n_9175;
wire n_7168;
wire n_6508;
wire n_7093;
wire n_4476;
wire n_5026;
wire n_12013;
wire n_11835;
wire n_4995;
wire n_7542;
wire n_7970;
wire n_7091;
wire n_10959;
wire n_6809;
wire n_11233;
wire n_5636;
wire n_7840;
wire n_10972;
wire n_6359;
wire n_7782;
wire n_13213;
wire n_12231;
wire n_5212;
wire n_10024;
wire n_10945;
wire n_8800;
wire n_16386;
wire n_13385;
wire n_15695;
wire n_10845;
wire n_7080;
wire n_6636;
wire n_5286;
wire n_8229;
wire n_16339;
wire n_8410;
wire n_4528;
wire n_14756;
wire n_14863;
wire n_5811;
wire n_14156;
wire n_13992;
wire n_10711;
wire n_7739;
wire n_6766;
wire n_7624;
wire n_4914;
wire n_7629;
wire n_4939;
wire n_13790;
wire n_14384;
wire n_9735;
wire n_16185;
wire n_9186;
wire n_10818;
wire n_5530;
wire n_15905;
wire n_5397;
wire n_10624;
wire n_4634;
wire n_12552;
wire n_13304;
wire n_14633;
wire n_11069;
wire n_5595;
wire n_9941;
wire n_11951;
wire n_12222;
wire n_7003;
wire n_15178;
wire n_11900;
wire n_15699;
wire n_14711;
wire n_13604;
wire n_5427;
wire n_10788;
wire n_11369;
wire n_4379;
wire n_10563;
wire n_14210;
wire n_8810;
wire n_5388;
wire n_4718;
wire n_9802;
wire n_15788;
wire n_5901;
wire n_13362;
wire n_6538;
wire n_14373;
wire n_5962;
wire n_5599;
wire n_7010;
wire n_8107;
wire n_11108;
wire n_12883;
wire n_9728;
wire n_12992;
wire n_11004;
wire n_5324;
wire n_6519;
wire n_15752;
wire n_8983;
wire n_10422;
wire n_11686;
wire n_9818;
wire n_6530;
wire n_7219;
wire n_9662;
wire n_14154;
wire n_12896;
wire n_4440;
wire n_15694;
wire n_8774;
wire n_4402;
wire n_14518;
wire n_16310;
wire n_10566;
wire n_16503;
wire n_16477;
wire n_13397;
wire n_16568;
wire n_10178;
wire n_7299;
wire n_5052;
wire n_12367;
wire n_4541;
wire n_12104;
wire n_5009;
wire n_15360;
wire n_4872;
wire n_6402;
wire n_12469;
wire n_13526;
wire n_9936;
wire n_12563;
wire n_4551;
wire n_15829;
wire n_6195;
wire n_13132;
wire n_7243;
wire n_6609;
wire n_7326;
wire n_9530;
wire n_10115;
wire n_13321;
wire n_14692;
wire n_15042;
wire n_7471;
wire n_5326;
wire n_7067;
wire n_10455;
wire n_11778;
wire n_12793;
wire n_14722;
wire n_13427;
wire n_15488;
wire n_15519;
wire n_4627;
wire n_14835;
wire n_5300;
wire n_15391;
wire n_9909;
wire n_11393;
wire n_14871;
wire n_16226;
wire n_8691;
wire n_8620;
wire n_12406;
wire n_14907;
wire n_6748;
wire n_15264;
wire n_7741;
wire n_5035;
wire n_9466;
wire n_13270;
wire n_16525;
wire n_7790;
wire n_11719;
wire n_16315;
wire n_6149;
wire n_16685;
wire n_10052;
wire n_10109;
wire n_7484;
wire n_7002;
wire n_16639;
wire n_10448;
wire n_6414;
wire n_11196;
wire n_16239;
wire n_15358;
wire n_11963;
wire n_12428;
wire n_14636;
wire n_8424;
wire n_9571;
wire n_16334;
wire n_15814;
wire n_8026;
wire n_7528;
wire n_9470;
wire n_9638;
wire n_4798;
wire n_16003;
wire n_16069;
wire n_15516;
wire n_10265;
wire n_8174;
wire n_12655;
wire n_16676;
wire n_7941;
wire n_13524;
wire n_16096;
wire n_11175;
wire n_13792;
wire n_5010;
wire n_15756;
wire n_11483;
wire n_5352;
wire n_15067;
wire n_11995;
wire n_14378;
wire n_5089;
wire n_13356;
wire n_11371;
wire n_14912;
wire n_10040;
wire n_5394;
wire n_4592;
wire n_9405;
wire n_6264;
wire n_14191;
wire n_16546;
wire n_8861;
wire n_5359;
wire n_13480;
wire n_8644;
wire n_8907;
wire n_16144;
wire n_16669;
wire n_12304;
wire n_13571;
wire n_15156;
wire n_11080;
wire n_10984;
wire n_5137;
wire n_6902;
wire n_5104;
wire n_14079;
wire n_15168;
wire n_10100;
wire n_7117;
wire n_13138;
wire n_9894;
wire n_5741;
wire n_8324;
wire n_15411;
wire n_15743;
wire n_6205;
wire n_9441;
wire n_6380;
wire n_10906;
wire n_7478;
wire n_7913;
wire n_12001;
wire n_5405;
wire n_7136;
wire n_6754;
wire n_7883;
wire n_7456;
wire n_5288;
wire n_15144;
wire n_12692;
wire n_13715;
wire n_13600;
wire n_7939;
wire n_13602;
wire n_14224;
wire n_8503;
wire n_16675;
wire n_9612;
wire n_4756;
wire n_8196;
wire n_10380;
wire n_10790;
wire n_16062;
wire n_14919;
wire n_6449;
wire n_6723;
wire n_7458;
wire n_9108;
wire n_16653;
wire n_9787;
wire n_6440;
wire n_7436;
wire n_10846;
wire n_4746;
wire n_13363;
wire n_15186;
wire n_14101;
wire n_6461;
wire n_4970;
wire n_9376;
wire n_8446;
wire n_5194;
wire n_9786;
wire n_14682;
wire n_14908;
wire n_9033;
wire n_13810;
wire n_14403;
wire n_12933;
wire n_7435;
wire n_12908;
wire n_15031;
wire n_15718;
wire n_9537;
wire n_11297;
wire n_14635;
wire n_6997;
wire n_10509;
wire n_5952;
wire n_13893;
wire n_12996;
wire n_15171;
wire n_14201;
wire n_5947;
wire n_8923;
wire n_13625;
wire n_12643;
wire n_13315;
wire n_13473;
wire n_6124;
wire n_6736;
wire n_7685;
wire n_7363;
wire n_8192;
wire n_14597;
wire n_5985;
wire n_8197;
wire n_15663;
wire n_14353;
wire n_15963;
wire n_16589;
wire n_6622;
wire n_11946;
wire n_9443;
wire n_11521;
wire n_9996;
wire n_11742;
wire n_14950;
wire n_4633;
wire n_6891;
wire n_7800;
wire n_10031;
wire n_12827;
wire n_12678;
wire n_13795;
wire n_9115;
wire n_12235;
wire n_14547;
wire n_4584;
wire n_15416;
wire n_5232;
wire n_11833;
wire n_7663;
wire n_11897;
wire n_12204;
wire n_10898;
wire n_5116;
wire n_14386;
wire n_5001;
wire n_15868;
wire n_7443;
wire n_5176;
wire n_7747;
wire n_9779;
wire n_16472;
wire n_9938;
wire n_11285;
wire n_8082;
wire n_12098;
wire n_4428;
wire n_8730;
wire n_7917;
wire n_7261;
wire n_15533;
wire n_9023;
wire n_12579;
wire n_6528;
wire n_9203;
wire n_14415;
wire n_9977;
wire n_15073;
wire n_7532;
wire n_8051;
wire n_9613;
wire n_11818;
wire n_15165;
wire n_5761;
wire n_13982;
wire n_13475;
wire n_16298;
wire n_9242;
wire n_15079;
wire n_6773;
wire n_4618;
wire n_12611;
wire n_13859;
wire n_13269;
wire n_7375;
wire n_13369;
wire n_4679;
wire n_13569;
wire n_11262;
wire n_4496;
wire n_7968;
wire n_6382;
wire n_7455;
wire n_12713;
wire n_12880;
wire n_13144;
wire n_15930;
wire n_4805;
wire n_8651;
wire n_13959;
wire n_9141;
wire n_15867;
wire n_5760;
wire n_6885;
wire n_9201;
wire n_10732;
wire n_6531;
wire n_10952;
wire n_10851;
wire n_11027;
wire n_13628;
wire n_11852;
wire n_10660;
wire n_7430;
wire n_5472;
wire n_10221;
wire n_9559;
wire n_8377;
wire n_9299;
wire n_11803;
wire n_15738;
wire n_9937;
wire n_5679;
wire n_11162;
wire n_7912;
wire n_9913;
wire n_13685;
wire n_5100;
wire n_9286;
wire n_16301;
wire n_8015;
wire n_5973;
wire n_7921;
wire n_10044;
wire n_7728;
wire n_4410;
wire n_8281;
wire n_10819;
wire n_14693;
wire n_4807;
wire n_15613;
wire n_8842;
wire n_14786;
wire n_4411;
wire n_14521;
wire n_9184;
wire n_9704;
wire n_13585;
wire n_5166;
wire n_9046;
wire n_16576;
wire n_6339;
wire n_14486;
wire n_8024;
wire n_7730;
wire n_12562;
wire n_8814;
wire n_8530;
wire n_11428;
wire n_11592;
wire n_15090;
wire n_16531;
wire n_9193;
wire n_8467;
wire n_11677;
wire n_7281;
wire n_15385;
wire n_9717;
wire n_13577;
wire n_7711;
wire n_16094;
wire n_16181;
wire n_11090;
wire n_15948;
wire n_8984;
wire n_6417;
wire n_5688;
wire n_9290;
wire n_13281;
wire n_5740;
wire n_5820;
wire n_13769;
wire n_5648;
wire n_14870;
wire n_13266;
wire n_13957;
wire n_14580;
wire n_15627;
wire n_5745;
wire n_4707;
wire n_4676;
wire n_9403;
wire n_10996;
wire n_13672;
wire n_14028;
wire n_9875;
wire n_5180;
wire n_6763;
wire n_8956;
wire n_5182;
wire n_7858;
wire n_11561;
wire n_14772;
wire n_8676;
wire n_8003;
wire n_5534;
wire n_4880;
wire n_13827;
wire n_8785;
wire n_9853;
wire n_13192;
wire n_7448;
wire n_6542;
wire n_15681;
wire n_14542;
wire n_6556;
wire n_15048;
wire n_8692;
wire n_7230;
wire n_6889;
wire n_9183;
wire n_16142;
wire n_7989;
wire n_9778;
wire n_14326;
wire n_5196;
wire n_6199;
wire n_9823;
wire n_5171;
wire n_12937;
wire n_10698;
wire n_15739;
wire n_16381;
wire n_10852;
wire n_15003;
wire n_4470;
wire n_14665;
wire n_6726;
wire n_12374;
wire n_13200;
wire n_9529;
wire n_4813;
wire n_5542;
wire n_7011;
wire n_8998;
wire n_10538;
wire n_5261;
wire n_12848;
wire n_11425;
wire n_12158;
wire n_10870;
wire n_13342;
wire n_4704;
wire n_11066;
wire n_10315;
wire n_13886;
wire n_9123;
wire n_6576;
wire n_6471;
wire n_8906;
wire n_5949;
wire n_11455;
wire n_15545;
wire n_4596;
wire n_14924;
wire n_12368;
wire n_4444;
wire n_5255;
wire n_8482;
wire n_6478;
wire n_7952;
wire n_11867;
wire n_13193;
wire n_6100;
wire n_12796;
wire n_16242;
wire n_6516;
wire n_14489;
wire n_16053;
wire n_8462;
wire n_13774;
wire n_6977;
wire n_9380;
wire n_13847;
wire n_10062;
wire n_7660;
wire n_6915;
wire n_12529;
wire n_15708;
wire n_12103;
wire n_7834;
wire n_11716;
wire n_5185;
wire n_8409;
wire n_6911;
wire n_6599;
wire n_8979;
wire n_6522;
wire n_14053;
wire n_4952;
wire n_5023;
wire n_5906;
wire n_8429;
wire n_8930;
wire n_10514;
wire n_16564;
wire n_14581;
wire n_5660;
wire n_7890;
wire n_12785;
wire n_11950;
wire n_7245;
wire n_5334;
wire n_6024;
wire n_9347;
wire n_4761;
wire n_15312;
wire n_6675;
wire n_6270;
wire n_14155;
wire n_12461;
wire n_6808;
wire n_13603;
wire n_16091;
wire n_16395;
wire n_7620;
wire n_11415;
wire n_11886;
wire n_7265;
wire n_7986;
wire n_5783;
wire n_6207;
wire n_7006;
wire n_6931;
wire n_5821;
wire n_14160;
wire n_6245;
wire n_14932;
wire n_6079;
wire n_15818;
wire n_16481;
wire n_7948;
wire n_9082;
wire n_10925;
wire n_4770;
wire n_9879;
wire n_11158;
wire n_9861;
wire n_11390;
wire n_6963;
wire n_8685;
wire n_15878;
wire n_16430;
wire n_4690;
wire n_11669;
wire n_16252;
wire n_14390;
wire n_8264;
wire n_14712;
wire n_15717;
wire n_5556;
wire n_4932;
wire n_8250;
wire n_8492;
wire n_7381;
wire n_16160;
wire n_12078;
wire n_16565;
wire n_10601;
wire n_5456;
wire n_9158;
wire n_10618;
wire n_8135;
wire n_15647;
wire n_9594;
wire n_7837;
wire n_9832;
wire n_16620;
wire n_7717;
wire n_8445;
wire n_9518;
wire n_6427;
wire n_6580;
wire n_5143;
wire n_9898;
wire n_11739;
wire n_5500;
wire n_6412;
wire n_10497;
wire n_14561;
wire n_9445;
wire n_14978;
wire n_7627;
wire n_13301;
wire n_9803;
wire n_13293;
wire n_7601;
wire n_6437;
wire n_8298;
wire n_6346;
wire n_14381;
wire n_7860;
wire n_5215;
wire n_15709;
wire n_15729;
wire n_8408;
wire n_12639;
wire n_14212;
wire n_5386;
wire n_10661;
wire n_7335;
wire n_9815;
wire n_8895;
wire n_9495;
wire n_10028;
wire n_13878;
wire n_15000;
wire n_7811;
wire n_13158;
wire n_14649;
wire n_11676;
wire n_11044;
wire n_14737;
wire n_11771;
wire n_15967;
wire n_12266;
wire n_15940;
wire n_12175;
wire n_5003;
wire n_15530;
wire n_13536;
wire n_10512;
wire n_13833;
wire n_14714;
wire n_11384;
wire n_4827;
wire n_16518;
wire n_12287;
wire n_11679;
wire n_8450;
wire n_8273;
wire n_9867;
wire n_6059;
wire n_7499;
wire n_12353;
wire n_14441;
wire n_14129;
wire n_6065;
wire n_9688;
wire n_9761;
wire n_7292;
wire n_12398;
wire n_5094;
wire n_4610;
wire n_10967;
wire n_13485;
wire n_9087;
wire n_4472;
wire n_7870;
wire n_5433;
wire n_9043;
wire n_6075;
wire n_12991;
wire n_16264;
wire n_7397;
wire n_10789;
wire n_11134;
wire n_12705;
wire n_13735;
wire n_15333;
wire n_6117;
wire n_7977;
wire n_8886;
wire n_12847;
wire n_10434;
wire n_7211;
wire n_12869;
wire n_13047;
wire n_10933;
wire n_5618;
wire n_6861;
wire n_8312;
wire n_6781;
wire n_11828;
wire n_14470;
wire n_12326;
wire n_15497;
wire n_14264;
wire n_7847;
wire n_8506;
wire n_14115;
wire n_15952;
wire n_16635;
wire n_6494;
wire n_13830;
wire n_13178;
wire n_6133;
wire n_16365;
wire n_11548;
wire n_13041;
wire n_13154;
wire n_8963;
wire n_12404;
wire n_14184;
wire n_7822;
wire n_6453;
wire n_4380;
wire n_5978;
wire n_11606;
wire n_11889;
wire n_9307;
wire n_6127;
wire n_4990;
wire n_4996;
wire n_5247;
wire n_14183;
wire n_10762;
wire n_11342;
wire n_4398;
wire n_11452;
wire n_11362;
wire n_15734;
wire n_8078;
wire n_7785;
wire n_6217;
wire n_4515;
wire n_14200;
wire n_5031;
wire n_6006;
wire n_11266;
wire n_10797;
wire n_7289;
wire n_14110;
wire n_16558;
wire n_12309;
wire n_7926;
wire n_14806;
wire n_5082;
wire n_6598;
wire n_7399;
wire n_5338;
wire n_12479;
wire n_7354;
wire n_15568;
wire n_8352;
wire n_12502;
wire n_13824;
wire n_10360;
wire n_7960;
wire n_15620;
wire n_9450;
wire n_5689;
wire n_13953;
wire n_7482;
wire n_12912;
wire n_14847;
wire n_10312;
wire n_12211;
wire n_16665;
wire n_6115;
wire n_13377;
wire n_12454;
wire n_8143;
wire n_10480;
wire n_4626;
wire n_9223;
wire n_13191;
wire n_16493;
wire n_6048;
wire n_6416;
wire n_10131;
wire n_12537;
wire n_6838;
wire n_15464;
wire n_10068;
wire n_6867;
wire n_9693;
wire n_11988;
wire n_12600;
wire n_12921;
wire n_14536;
wire n_13226;
wire n_6139;
wire n_5931;
wire n_13567;
wire n_11957;
wire n_10633;
wire n_12133;
wire n_13686;
wire n_6256;
wire n_7965;
wire n_13645;
wire n_15645;
wire n_16433;
wire n_6613;
wire n_11438;
wire n_11244;
wire n_12919;
wire n_14432;
wire n_15965;
wire n_5221;
wire n_10273;
wire n_5641;
wire n_12215;
wire n_11416;
wire n_10209;
wire n_6361;
wire n_9880;
wire n_13253;
wire n_4689;
wire n_14321;
wire n_8183;
wire n_14981;
wire n_11348;
wire n_16098;
wire n_4547;
wire n_11245;
wire n_9685;
wire n_6085;
wire n_7474;
wire n_11169;
wire n_11685;
wire n_5731;
wire n_12467;
wire n_6329;
wire n_11607;
wire n_8650;
wire n_12422;
wire n_6678;
wire n_11546;
wire n_15259;
wire n_14654;
wire n_15460;
wire n_8662;
wire n_10503;
wire n_14422;
wire n_15058;
wire n_9694;
wire n_16598;
wire n_7158;
wire n_4905;
wire n_14664;
wire n_16539;
wire n_16636;
wire n_13215;
wire n_13400;
wire n_4601;
wire n_14971;
wire n_9905;
wire n_9948;
wire n_10465;
wire n_14630;
wire n_16073;
wire n_12429;
wire n_10590;
wire n_13782;
wire n_14734;
wire n_15476;
wire n_14494;
wire n_8526;
wire n_13331;
wire n_14956;
wire n_4623;
wire n_7325;
wire n_13751;
wire n_10887;
wire n_14866;
wire n_9456;
wire n_5007;
wire n_7044;
wire n_14019;
wire n_9710;
wire n_6370;
wire n_8623;
wire n_11113;
wire n_9923;
wire n_5883;
wire n_13743;
wire n_7166;
wire n_13812;
wire n_14970;
wire n_6554;
wire n_12146;
wire n_7356;
wire n_5754;
wire n_6759;
wire n_10786;
wire n_13378;
wire n_6560;
wire n_14055;
wire n_11319;
wire n_7028;
wire n_7838;
wire n_4842;
wire n_9890;
wire n_11492;
wire n_5629;
wire n_7873;
wire n_6535;
wire n_16418;
wire n_12731;
wire n_16138;
wire n_12399;
wire n_16644;
wire n_7518;
wire n_12342;
wire n_12640;
wire n_7414;
wire n_9744;
wire n_9817;
wire n_6147;
wire n_10063;
wire n_9199;
wire n_13092;
wire n_14292;
wire n_9548;
wire n_8973;
wire n_11160;
wire n_6448;
wire n_13544;
wire n_7791;
wire n_12378;
wire n_8419;
wire n_9782;
wire n_12533;
wire n_9862;
wire n_5934;
wire n_7431;
wire n_5434;
wire n_12616;
wire n_11385;
wire n_12319;
wire n_10805;
wire n_11355;
wire n_11674;
wire n_12535;
wire n_12178;
wire n_14375;
wire n_12653;
wire n_6643;
wire n_12327;
wire n_7146;
wire n_9471;
wire n_4608;
wire n_16580;
wire n_11346;
wire n_10091;
wire n_11638;
wire n_6157;
wire n_14896;
wire n_4859;
wire n_9363;
wire n_12047;
wire n_12930;
wire n_12587;
wire n_5880;
wire n_8351;
wire n_8430;
wire n_10747;
wire n_12058;
wire n_14810;
wire n_9069;
wire n_13110;
wire n_15719;
wire n_14879;
wire n_16628;
wire n_16143;
wire n_5852;
wire n_14030;
wire n_8603;
wire n_9422;
wire n_5218;
wire n_15164;
wire n_8249;
wire n_16660;
wire n_7052;
wire n_11343;
wire n_12348;
wire n_16099;
wire n_10496;
wire n_12257;
wire n_15590;
wire n_15770;
wire n_12575;
wire n_5960;
wire n_11451;
wire n_14149;
wire n_13394;
wire n_4571;
wire n_10843;
wire n_13391;
wire n_7888;
wire n_11823;
wire n_6397;
wire n_5358;
wire n_13384;
wire n_14680;
wire n_8234;
wire n_16048;
wire n_5321;
wire n_9960;
wire n_10997;
wire n_16262;
wire n_9010;
wire n_13707;
wire n_15241;
wire n_10998;
wire n_15422;
wire n_9003;
wire n_9280;
wire n_6073;
wire n_7502;
wire n_12418;
wire n_14216;
wire n_6331;
wire n_5290;
wire n_16380;
wire n_14837;
wire n_13498;
wire n_7312;
wire n_13263;
wire n_7919;
wire n_14877;
wire n_5145;
wire n_15203;
wire n_11269;
wire n_10800;
wire n_7085;
wire n_11491;
wire n_12065;
wire n_13950;
wire n_9341;
wire n_6939;
wire n_7848;
wire n_11408;
wire n_14048;
wire n_11772;
wire n_16063;
wire n_16237;
wire n_14103;
wire n_4774;
wire n_16112;
wire n_5210;
wire n_13183;
wire n_6689;
wire n_13732;
wire n_14968;
wire n_16422;
wire n_10993;
wire n_15891;
wire n_7632;
wire n_12519;
wire n_5109;
wire n_14985;
wire n_15542;
wire n_9172;
wire n_12769;
wire n_15910;
wire n_14653;
wire n_4902;
wire n_6405;
wire n_7580;
wire n_14077;
wire n_5149;
wire n_8980;
wire n_12641;
wire n_13007;
wire n_5571;
wire n_11311;
wire n_10112;
wire n_14443;
wire n_10765;
wire n_16136;
wire n_6698;
wire n_15263;
wire n_11792;
wire n_14285;
wire n_7304;
wire n_9734;
wire n_7288;
wire n_8558;
wire n_13242;
wire n_10489;
wire n_7707;
wire n_16325;
wire n_7223;
wire n_12421;
wire n_13282;
wire n_14436;
wire n_7833;
wire n_12113;
wire n_14868;
wire n_4987;
wire n_14599;
wire n_7274;
wire n_5512;
wire n_16087;
wire n_9297;
wire n_10495;
wire n_10159;
wire n_9004;
wire n_4736;
wire n_14351;
wire n_6206;
wire n_9068;
wire n_13352;
wire n_8136;
wire n_5033;
wire n_9808;
wire n_6610;
wire n_7445;
wire n_14812;
wire n_10612;
wire n_11086;
wire n_7466;
wire n_6529;
wire n_10260;
wire n_11293;
wire n_14728;
wire n_4516;
wire n_6363;
wire n_6750;
wire n_12285;
wire n_13310;
wire n_11710;
wire n_8619;
wire n_11568;
wire n_6290;
wire n_10253;
wire n_7429;
wire n_11766;
wire n_6025;
wire n_11038;
wire n_9150;
wire n_10134;
wire n_14508;
wire n_15122;
wire n_11603;
wire n_13798;
wire n_7277;
wire n_6455;
wire n_15277;
wire n_15092;
wire n_13804;
wire n_12683;
wire n_11271;
wire n_12455;
wire n_14778;
wire n_15714;
wire n_15842;
wire n_13099;
wire n_12015;
wire n_8146;
wire n_4492;
wire n_13690;
wire n_14822;
wire n_8813;
wire n_5607;
wire n_11562;
wire n_7695;
wire n_10194;
wire n_14566;
wire n_7179;
wire n_10356;
wire n_7122;
wire n_10173;
wire n_12157;
wire n_7165;
wire n_7869;
wire n_4789;
wire n_5999;
wire n_13386;
wire n_13846;
wire n_8910;
wire n_12311;
wire n_4376;
wire n_6203;
wire n_6408;
wire n_14374;
wire n_15806;
wire n_6555;
wire n_9448;
wire n_7683;
wire n_10739;
wire n_13064;
wire n_14815;
wire n_6150;
wire n_7630;
wire n_10077;
wire n_16246;
wire n_4708;
wire n_13619;
wire n_16437;
wire n_8470;
wire n_4657;
wire n_9587;
wire n_12031;
wire n_5341;
wire n_16480;
wire n_8643;
wire n_15660;
wire n_4512;
wire n_9278;
wire n_10671;
wire n_15357;
wire n_10889;
wire n_10010;
wire n_10193;
wire n_11718;
wire n_8565;
wire n_10821;
wire n_13648;
wire n_14831;
wire n_14996;
wire n_11170;
wire n_11758;
wire n_12126;
wire n_14383;
wire n_8550;
wire n_14543;
wire n_9396;
wire n_4542;
wire n_6892;
wire n_11094;
wire n_4462;
wire n_14450;
wire n_14747;
wire n_7061;
wire n_11680;
wire n_12480;
wire n_15722;
wire n_14683;
wire n_10599;
wire n_9667;
wire n_14192;
wire n_14181;
wire n_6401;
wire n_7322;
wire n_15278;
wire n_9053;
wire n_11658;
wire n_15504;
wire n_11893;
wire n_13338;
wire n_6685;
wire n_11639;
wire n_12226;
wire n_4931;
wire n_9739;
wire n_10573;
wire n_13492;
wire n_14358;
wire n_4536;
wire n_9480;
wire n_14001;
wire n_14213;
wire n_5562;
wire n_15397;
wire n_4324;
wire n_7051;
wire n_10850;
wire n_9185;
wire n_8477;
wire n_15840;
wire n_7880;
wire n_9793;
wire n_11692;
wire n_15054;
wire n_4382;
wire n_12195;
wire n_13376;
wire n_14842;
wire n_13115;
wire n_11759;
wire n_8230;
wire n_12549;
wire n_6679;
wire n_8092;
wire n_13864;
wire n_5911;
wire n_11601;
wire n_13289;
wire n_15279;
wire n_11971;
wire n_13182;
wire n_11456;
wire n_12314;
wire n_10546;
wire n_16265;
wire n_5622;
wire n_9919;
wire n_12135;
wire n_16466;
wire n_6574;
wire n_11116;
wire n_13324;
wire n_12604;
wire n_6571;
wire n_13305;
wire n_5577;
wire n_9541;
wire n_11286;
wire n_8876;
wire n_15215;
wire n_5124;
wire n_9151;
wire n_8829;
wire n_16379;
wire n_9359;
wire n_7824;
wire n_13381;
wire n_13236;
wire n_14189;
wire n_14299;
wire n_7094;
wire n_15761;
wire n_5123;
wire n_7097;
wire n_16320;
wire n_4639;
wire n_8140;
wire n_5413;
wire n_8971;
wire n_15111;
wire n_8060;
wire n_16667;
wire n_10558;
wire n_7036;
wire n_9579;
wire n_9475;
wire n_11124;
wire n_15273;
wire n_6392;
wire n_5915;
wire n_8527;
wire n_12899;
wire n_13777;
wire n_15301;
wire n_9049;
wire n_7351;
wire n_13718;
wire n_4480;
wire n_9352;
wire n_14775;
wire n_7608;
wire n_5779;
wire n_6260;
wire n_15567;
wire n_6832;
wire n_7394;
wire n_11045;
wire n_13202;
wire n_7909;
wire n_15350;
wire n_7413;
wire n_13638;
wire n_6303;
wire n_8935;
wire n_14392;
wire n_11340;
wire n_15759;
wire n_10734;
wire n_6286;
wire n_16441;
wire n_7675;
wire n_8267;
wire n_15383;
wire n_11903;
wire n_7027;
wire n_7992;
wire n_13279;
wire n_13644;
wire n_6912;
wire n_11560;
wire n_10330;
wire n_7175;
wire n_8276;
wire n_10395;
wire n_13291;
wire n_6019;
wire n_10174;
wire n_11435;
wire n_14966;
wire n_11465;
wire n_7524;
wire n_15255;
wire n_4344;
wire n_8027;
wire n_15897;
wire n_4705;
wire n_11564;
wire n_14015;
wire n_8925;
wire n_6214;
wire n_12946;
wire n_9978;
wire n_11914;
wire n_11265;
wire n_9370;
wire n_11125;
wire n_9670;
wire n_13136;
wire n_13513;
wire n_12916;
wire n_9334;
wire n_7783;
wire n_13220;
wire n_15131;
wire n_6692;
wire n_10276;
wire n_14322;
wire n_12331;
wire n_8978;
wire n_10594;
wire n_8093;
wire n_12531;
wire n_8245;
wire n_15072;
wire n_6036;
wire n_8471;
wire n_4391;
wire n_12521;
wire n_11302;
wire n_12910;
wire n_13349;
wire n_9956;
wire n_9800;
wire n_8454;
wire n_6552;
wire n_8327;
wire n_11382;
wire n_13096;
wire n_9413;
wire n_12727;
wire n_15314;
wire n_10991;
wire n_14173;
wire n_15509;
wire n_10098;
wire n_11745;
wire n_8891;
wire n_15240;
wire n_4947;
wire n_11690;
wire n_16194;
wire n_9487;
wire n_11707;
wire n_5591;
wire n_11373;
wire n_7697;
wire n_14608;
wire n_6403;
wire n_15564;
wire n_7306;
wire n_13835;
wire n_16153;
wire n_16260;
wire n_7947;
wire n_10118;
wire n_14350;
wire n_7470;
wire n_7547;
wire n_6013;
wire n_7733;
wire n_13815;
wire n_13800;
wire n_7693;
wire n_9557;
wire n_15957;
wire n_6491;
wire n_16319;
wire n_4740;
wire n_4631;
wire n_16321;
wire n_14039;
wire n_14072;
wire n_15662;
wire n_11412;
wire n_6348;
wire n_6744;
wire n_13039;
wire n_13773;
wire n_13130;
wire n_14109;
wire n_8582;
wire n_10441;
wire n_6982;
wire n_5518;
wire n_10002;
wire n_6293;
wire n_5068;
wire n_9124;
wire n_6661;
wire n_15671;
wire n_5847;
wire n_13719;
wire n_7345;
wire n_6049;
wire n_9762;
wire n_8847;
wire n_11242;
wire n_8957;
wire n_14136;
wire n_7385;
wire n_10923;
wire n_14548;
wire n_5159;
wire n_15793;
wire n_15923;
wire n_6558;
wire n_14176;
wire n_4625;
wire n_11149;
wire n_10841;
wire n_16076;
wire n_12635;
wire n_12227;
wire n_12258;
wire n_14117;
wire n_13694;
wire n_12313;
wire n_4766;
wire n_8488;
wire n_9271;
wire n_4863;
wire n_9543;
wire n_13688;
wire n_14661;
wire n_11396;
wire n_8356;
wire n_6136;
wire n_9660;
wire n_15196;
wire n_16176;
wire n_16384;
wire n_16416;
wire n_11443;
wire n_9483;
wire n_15765;
wire n_6855;
wire n_15305;
wire n_15588;
wire n_14754;
wire n_10665;
wire n_4744;
wire n_12906;
wire n_8888;
wire n_11810;
wire n_14267;
wire n_15020;
wire n_16233;
wire n_13467;
wire n_5357;
wire n_6091;
wire n_13093;
wire n_13062;
wire n_9328;
wire n_14252;
wire n_7857;
wire n_7481;
wire n_16511;
wire n_14130;
wire n_15830;
wire n_12583;
wire n_6551;
wire n_7691;
wire n_14930;
wire n_7907;
wire n_5541;
wire n_5568;
wire n_10576;
wire n_16596;
wire n_6312;
wire n_8747;
wire n_11532;
wire n_9539;
wire n_6668;
wire n_4817;
wire n_9415;
wire n_15274;
wire n_14343;
wire n_15548;
wire n_16410;
wire n_9385;
wire n_9147;
wire n_11209;
wire n_7653;
wire n_13462;
wire n_8354;
wire n_5381;
wire n_15918;
wire n_9785;
wire n_5723;
wire n_6859;
wire n_14276;
wire n_5918;
wire n_6959;
wire n_16212;
wire n_8353;
wire n_13752;
wire n_8922;
wire n_6388;
wire n_5045;
wire n_10237;
wire n_11053;
wire n_11790;
wire n_13185;
wire n_9027;
wire n_12159;
wire n_9434;
wire n_12750;
wire n_4383;
wire n_13596;
wire n_6995;
wire n_10902;
wire n_4491;
wire n_12889;
wire n_13855;
wire n_5696;
wire n_8348;
wire n_7032;
wire n_8211;
wire n_12050;
wire n_12922;
wire n_12250;
wire n_4486;
wire n_16313;
wire n_9515;
wire n_10420;
wire n_6971;
wire n_11304;
wire n_9642;
wire n_16363;
wire n_9233;
wire n_6131;
wire n_9681;
wire n_5848;
wire n_15232;
wire n_7475;
wire n_10485;
wire n_14231;
wire n_12105;
wire n_4612;
wire n_12385;
wire n_6435;
wire n_10536;
wire n_13219;
wire n_14329;
wire n_5673;
wire n_5443;
wire n_6351;
wire n_9079;
wire n_15544;
wire n_15721;
wire n_9382;
wire n_16392;
wire n_10282;
wire n_5163;
wire n_6212;
wire n_7668;
wire n_16145;
wire n_9775;
wire n_10444;
wire n_4529;
wire n_11377;
wire n_8653;
wire n_8018;
wire n_13295;
wire n_15142;
wire n_8920;
wire n_10913;
wire n_7937;
wire n_9176;
wire n_6829;
wire n_10950;
wire n_5485;
wire n_7819;
wire n_10631;
wire n_15991;
wire n_5823;
wire n_7305;
wire n_13388;
wire n_13160;
wire n_13731;
wire n_11071;
wire n_5473;
wire n_10072;
wire n_15249;
wire n_6682;
wire n_6334;
wire n_6823;
wire n_14550;
wire n_10708;
wire n_10703;
wire n_9089;
wire n_9666;
wire n_14503;
wire n_4390;
wire n_12248;
wire n_13818;
wire n_15024;
wire n_8678;
wire n_10565;
wire n_10011;
wire n_15346;
wire n_13477;
wire n_8884;
wire n_8803;
wire n_14886;
wire n_8942;
wire n_7993;
wire n_7181;
wire n_9865;
wire n_10978;
wire n_5537;
wire n_8222;
wire n_13808;
wire n_14644;
wire n_6822;
wire n_11715;
wire n_4396;
wire n_8553;
wire n_7071;
wire n_9706;
wire n_15174;
wire n_15454;
wire n_10642;
wire n_15213;
wire n_12181;
wire n_10187;
wire n_10387;
wire n_11014;
wire n_13764;
wire n_14560;
wire n_15033;
wire n_8751;
wire n_11864;
wire n_14829;
wire n_11007;
wire n_11224;
wire n_15473;
wire n_11006;
wire n_15584;
wire n_9564;
wire n_15018;
wire n_7391;
wire n_8790;
wire n_15569;
wire n_9230;
wire n_6617;
wire n_10219;
wire n_7511;
wire n_6533;
wire n_11924;
wire n_10768;
wire n_10316;
wire n_9795;
wire n_15193;
wire n_4684;
wire n_14067;
wire n_9591;
wire n_6429;
wire n_6407;
wire n_16515;
wire n_14108;
wire n_6389;
wire n_6137;
wire n_5027;
wire n_15903;
wire n_14833;
wire n_10364;
wire n_15439;
wire n_10479;
wire n_11422;
wire n_16049;
wire n_8338;
wire n_6983;
wire n_10494;
wire n_13660;
wire n_8398;
wire n_4412;
wire n_14480;
wire n_8178;
wire n_13970;
wire n_6801;
wire n_15247;
wire n_16656;
wire n_12489;
wire n_8491;
wire n_14000;
wire n_14372;
wire n_4580;
wire n_5630;
wire n_4758;
wire n_10065;
wire n_4781;
wire n_12046;
wire n_10212;
wire n_16610;
wire n_9283;
wire n_8700;
wire n_12030;
wire n_12738;
wire n_13408;
wire n_15062;
wire n_15248;
wire n_13727;
wire n_5379;
wire n_13025;
wire n_5335;
wire n_11599;
wire n_12565;
wire n_10268;
wire n_15236;
wire n_14801;
wire n_14098;
wire n_6113;
wire n_9468;
wire n_10070;
wire n_12601;
wire n_14482;
wire n_15399;
wire n_16178;
wire n_9425;
wire n_12917;
wire n_14629;
wire n_13641;
wire n_14223;
wire n_15962;
wire n_11172;
wire n_10089;
wire n_5424;
wire n_12415;
wire n_8750;
wire n_14947;
wire n_5505;
wire n_5868;
wire n_10305;
wire n_8560;
wire n_14983;
wire n_14748;
wire n_10559;
wire n_13173;
wire n_8439;
wire n_9641;
wire n_12755;
wire n_10004;
wire n_12807;
wire n_15355;
wire n_15669;
wire n_12059;
wire n_12488;
wire n_15945;
wire n_7321;
wire n_14848;
wire n_5289;
wire n_8200;
wire n_15845;
wire n_11110;
wire n_7154;
wire n_6129;
wire n_5018;
wire n_16055;
wire n_16232;
wire n_6518;
wire n_16211;
wire n_15001;
wire n_8304;
wire n_11418;
wire n_6655;
wire n_8674;
wire n_12981;
wire n_5274;
wire n_9138;
wire n_5401;
wire n_12977;
wire n_7584;
wire n_9958;
wire n_14544;
wire n_4457;
wire n_13328;
wire n_7537;
wire n_10516;
wire n_8675;
wire n_10892;
wire n_6254;
wire n_5989;
wire n_15924;
wire n_10493;
wire n_13542;
wire n_12567;
wire n_9367;
wire n_7320;
wire n_4928;
wire n_5769;
wire n_10405;
wire n_15037;
wire n_4794;
wire n_15130;
wire n_16122;
wire n_5613;
wire n_8212;
wire n_5612;
wire n_14604;
wire n_14735;
wire n_7964;
wire n_4482;
wire n_9016;
wire n_14426;
wire n_13101;
wire n_11887;
wire n_15456;
wire n_14349;
wire n_6278;
wire n_6786;
wire n_7022;
wire n_10026;
wire n_11545;
wire n_9729;
wire n_5073;
wire n_12691;
wire n_8846;
wire n_8315;
wire n_16446;
wire n_12471;
wire n_11033;
wire n_15885;
wire n_12451;
wire n_4834;
wire n_11040;
wire n_12665;
wire n_16367;
wire n_16526;
wire n_16397;
wire n_11754;
wire n_11850;
wire n_14916;
wire n_15740;
wire n_9194;
wire n_8760;
wire n_9756;
wire n_12592;
wire n_14356;
wire n_4762;
wire n_5581;
wire n_13748;
wire n_9029;
wire n_9411;
wire n_11672;
wire n_10353;
wire n_6837;
wire n_16006;
wire n_10847;
wire n_12651;
wire n_10451;
wire n_11043;
wire n_15801;
wire n_5303;
wire n_16476;
wire n_12507;
wire n_7486;
wire n_12240;
wire n_6756;
wire n_16373;
wire n_9414;
wire n_7023;
wire n_12003;
wire n_9615;
wire n_14205;
wire n_14564;
wire n_7496;
wire n_11277;
wire n_12165;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_10866;
wire n_14190;
wire n_7410;
wire n_9940;
wire n_10779;
wire n_8563;
wire n_6200;
wire n_4504;
wire n_14600;
wire n_8777;
wire n_4975;
wire n_11061;
wire n_11763;
wire n_16495;
wire n_15546;
wire n_15010;
wire n_8465;
wire n_6670;
wire n_8535;
wire n_10653;
wire n_11534;
wire n_6373;
wire n_5375;
wire n_11587;
wire n_12280;
wire n_9221;
wire n_12492;
wire n_13581;
wire n_13461;
wire n_14344;
wire n_15742;
wire n_16686;
wire n_12972;
wire n_16282;
wire n_16347;
wire n_5370;
wire n_13789;
wire n_4898;
wire n_4815;
wire n_5601;
wire n_5784;
wire n_9811;
wire n_7899;
wire n_8631;
wire n_13188;
wire n_4819;
wire n_14511;
wire n_7906;
wire n_16385;
wire n_13286;
wire n_5248;
wire n_9951;
wire n_7131;
wire n_14723;
wire n_6411;
wire n_9424;
wire n_9586;
wire n_10285;
wire n_4370;
wire n_8909;
wire n_14488;
wire n_11032;
wire n_5112;
wire n_13582;
wire n_10507;
wire n_16356;
wire n_10520;
wire n_7302;
wire n_11968;
wire n_11843;
wire n_10045;
wire n_11174;
wire n_4645;
wire n_14614;
wire n_13531;
wire n_7797;
wire n_11335;
wire n_11629;
wire n_15147;
wire n_6381;
wire n_7030;
wire n_6656;
wire n_9730;
wire n_13880;
wire n_7687;
wire n_9554;
wire n_10294;
wire n_4755;
wire n_13988;
wire n_4359;
wire n_4960;
wire n_10106;
wire n_5635;
wire n_7582;
wire n_15272;
wire n_9934;
wire n_4933;
wire n_10541;
wire n_5091;
wire n_13609;
wire n_14587;
wire n_4591;
wire n_6546;
wire n_5528;
wire n_9234;
wire n_10674;
wire n_5111;
wire n_8959;
wire n_6534;
wire n_13679;
wire n_10614;
wire n_5227;
wire n_7809;
wire n_11785;
wire n_10417;
wire n_15927;
wire n_16011;
wire n_12841;
wire n_6265;
wire n_12855;
wire n_5778;
wire n_8425;
wire n_11257;
wire n_15176;
wire n_8087;
wire n_15834;
wire n_13276;
wire n_9910;
wire n_7060;
wire n_7607;
wire n_10217;
wire n_14458;
wire n_8938;
wire n_4474;
wire n_5665;
wire n_16058;
wire n_11801;
wire n_13217;
wire n_16519;
wire n_12073;
wire n_13655;
wire n_6898;
wire n_6596;
wire n_5363;
wire n_10743;
wire n_5165;
wire n_13424;
wire n_16332;
wire n_14658;
wire n_15066;
wire n_4884;
wire n_14830;
wire n_14397;
wire n_10853;
wire n_7867;
wire n_9651;
wire n_13565;
wire n_14281;
wire n_13755;
wire n_14643;
wire n_10249;
wire n_8361;
wire n_6135;
wire n_13802;
wire n_14594;
wire n_15474;
wire n_7761;
wire n_10705;
wire n_8007;
wire n_9246;
wire n_10338;
wire n_15316;
wire n_10270;
wire n_6814;
wire n_11115;
wire n_10557;
wire n_8669;
wire n_12978;
wire n_13784;
wire n_8001;
wire n_7525;
wire n_13468;
wire n_7257;
wire n_12363;
wire n_9372;
wire n_7553;
wire n_7529;
wire n_15668;
wire n_4692;
wire n_6791;
wire n_15137;
wire n_14233;
wire n_8496;
wire n_11915;
wire n_13704;
wire n_6824;
wire n_5788;
wire n_11016;
wire n_9326;
wire n_14976;
wire n_11788;
wire n_12544;
wire n_13036;
wire n_14146;
wire n_7650;
wire n_12476;
wire n_13199;
wire n_8568;
wire n_6903;
wire n_13009;
wire n_13043;
wire n_8852;
wire n_12023;
wire n_8637;
wire n_6168;
wire n_16225;
wire n_6881;
wire n_16677;
wire n_4722;
wire n_4606;
wire n_10339;
wire n_9908;
wire n_10908;
wire n_13413;
wire n_9486;
wire n_6450;
wire n_9544;
wire n_13002;
wire n_15153;
wire n_12632;
wire n_12620;
wire n_7520;
wire n_9831;
wire n_13203;
wire n_13868;
wire n_6309;
wire n_7903;
wire n_9697;
wire n_11303;
wire n_11877;
wire n_6733;
wire n_14462;
wire n_8864;
wire n_7384;
wire n_8456;
wire n_5317;
wire n_13285;
wire n_5430;
wire n_8610;
wire n_5942;
wire n_7894;
wire n_7137;
wire n_4563;
wire n_4962;
wire n_9902;
wire n_14933;
wire n_5056;
wire n_8362;
wire n_4820;
wire n_5540;
wire n_11750;
wire n_9900;
wire n_6300;
wire n_8256;
wire n_15521;
wire n_9920;
wire n_7055;
wire n_7202;
wire n_5716;
wire n_8520;
wire n_9310;
wire n_10132;
wire n_12598;
wire n_9039;
wire n_13374;
wire n_11854;
wire n_12416;
wire n_16458;
wire n_8573;
wire n_12055;
wire n_12091;
wire n_8704;
wire n_8265;
wire n_4619;
wire n_7639;
wire n_16520;
wire n_5762;
wire n_6132;
wire n_4327;
wire n_11609;
wire n_5211;
wire n_5336;
wire n_5447;
wire n_16464;
wire n_7743;
wire n_13230;
wire n_9294;
wire n_5036;
wire n_12811;
wire n_12186;
wire n_11747;
wire n_6179;
wire n_6395;
wire n_10327;
wire n_12494;
wire n_13032;
wire n_13826;
wire n_7054;
wire n_7605;
wire n_11556;
wire n_15140;
wire n_11529;
wire n_9512;
wire n_10437;
wire n_11001;
wire n_10021;
wire n_5327;
wire n_13684;
wire n_14199;
wire n_16673;
wire n_9146;
wire n_9125;
wire n_4392;
wire n_9170;
wire n_9139;
wire n_11858;
wire n_14027;
wire n_15108;
wire n_15753;
wire n_7433;
wire n_9616;
wire n_8131;
wire n_8941;
wire n_5014;
wire n_16316;
wire n_5747;
wire n_9073;
wire n_10075;
wire n_16357;
wire n_12733;
wire n_10423;
wire n_12897;
wire n_12623;
wire n_11444;
wire n_5192;
wire n_4334;
wire n_6171;
wire n_13750;
wire n_8775;
wire n_14104;
wire n_12272;
wire n_9302;
wire n_5519;
wire n_13948;
wire n_11798;
wire n_9062;
wire n_14684;
wire n_11895;
wire n_13458;
wire n_6269;
wire n_5753;
wire n_7092;
wire n_6980;
wire n_11213;
wire n_12245;
wire n_15713;
wire n_9171;
wire n_10886;
wire n_5233;
wire n_8279;
wire n_12213;
wire n_6654;
wire n_9358;
wire n_12191;
wire n_9580;
wire n_8019;
wire n_14572;
wire n_13963;
wire n_9972;
wire n_13003;
wire n_6083;
wire n_13091;
wire n_12909;
wire n_4575;
wire n_6434;
wire n_6387;
wire n_9565;
wire n_9157;
wire n_8257;
wire n_13072;
wire n_10192;
wire n_7832;
wire n_9465;
wire n_16417;
wire n_9540;
wire n_9324;
wire n_5808;
wire n_8390;
wire n_11137;
wire n_8898;
wire n_13811;
wire n_14316;
wire n_7726;
wire n_8807;
wire n_5436;
wire n_5139;
wire n_13839;
wire n_6120;
wire n_5231;
wire n_8613;
wire n_6068;
wire n_6933;
wire n_8521;
wire n_14011;
wire n_13954;
wire n_10436;
wire n_8464;
wire n_15701;
wire n_6547;
wire n_8799;
wire n_12794;
wire n_5193;
wire n_6423;
wire n_15496;
wire n_9442;
wire n_6342;
wire n_6641;
wire n_15260;
wire n_6984;
wire n_15612;
wire n_5789;
wire n_15104;
wire n_10763;
wire n_7441;
wire n_9957;
wire n_10124;
wire n_12483;
wire n_12759;
wire n_11793;
wire n_16374;
wire n_7106;
wire n_7213;
wire n_12112;
wire n_13060;
wire n_14689;
wire n_16187;
wire n_10245;
wire n_5961;
wire n_10905;
wire n_14132;
wire n_11235;
wire n_9449;
wire n_14817;
wire n_5866;
wire n_9050;
wire n_6507;
wire n_6399;
wire n_4499;
wire n_9313;
wire n_6687;
wire n_5822;
wire n_9173;
wire n_5195;
wire n_6690;
wire n_6121;
wire n_7412;
wire n_9959;
wire n_12144;
wire n_15055;
wire n_5726;
wire n_11015;
wire n_9563;
wire n_14087;
wire n_9160;
wire n_5364;
wire n_9974;
wire n_12129;
wire n_14753;
wire n_11166;
wire n_15980;
wire n_7031;
wire n_9285;
wire n_13658;
wire n_5533;
wire n_16595;
wire n_7763;
wire n_9631;
wire n_14671;
wire n_8033;
wire n_15172;
wire n_14751;
wire n_4458;
wire n_6194;
wire n_14438;
wire n_16454;
wire n_5103;
wire n_4641;
wire n_8393;
wire n_16253;
wire n_7133;
wire n_16561;
wire n_13572;
wire n_15547;
wire n_12032;
wire n_4720;
wire n_10784;
wire n_12202;
wire n_4893;
wire n_14674;
wire n_13836;
wire n_8463;
wire n_8153;
wire n_12815;
wire n_15913;
wire n_6524;
wire n_10944;
wire n_10211;
wire n_12835;
wire n_10129;
wire n_10431;
wire n_9945;
wire n_8661;
wire n_16089;
wire n_12431;
wire n_7424;
wire n_7523;
wire n_8654;
wire n_5039;
wire n_16314;
wire n_11855;
wire n_4772;
wire n_14229;
wire n_15060;
wire n_6790;
wire n_8746;
wire n_11241;
wire n_15115;
wire n_16671;
wire n_15520;
wire n_5953;
wire n_12870;
wire n_11183;
wire n_10019;
wire n_11156;
wire n_8531;
wire n_14188;
wire n_11508;
wire n_10611;
wire n_12093;
wire n_7141;
wire n_5198;
wire n_11581;
wire n_10715;
wire n_4468;
wire n_13799;
wire n_5718;
wire n_6459;
wire n_6505;
wire n_16139;
wire n_12333;
wire n_12636;
wire n_8379;
wire n_8609;
wire n_13854;
wire n_11227;
wire n_7626;
wire n_13576;
wire n_15380;
wire n_13100;
wire n_4961;
wire n_7310;
wire n_4454;
wire n_16154;
wire n_12334;
wire n_6686;
wire n_15956;
wire n_6001;
wire n_7311;
wire n_9209;
wire n_7669;
wire n_11218;
wire n_4502;
wire n_12119;
wire n_11787;
wire n_12618;
wire n_5958;
wire n_8793;
wire n_16059;
wire n_12355;
wire n_8103;
wire n_15052;
wire n_9767;
wire n_9838;
wire n_10195;
wire n_13722;
wire n_4526;
wire n_9300;
wire n_11500;
wire n_16093;
wire n_4849;
wire n_12943;
wire n_15129;
wire n_7327;
wire n_14306;
wire n_12938;
wire n_13057;
wire n_8873;
wire n_8367;
wire n_11891;
wire n_16276;
wire n_7367;
wire n_14752;
wire n_5792;
wire n_11021;
wire n_12401;
wire n_16439;
wire n_8543;
wire n_16502;
wire n_6183;
wire n_6023;
wire n_13055;
wire n_7323;
wire n_11544;
wire n_7189;
wire n_14897;
wire n_15447;
wire n_7301;
wire n_12173;
wire n_13067;
wire n_10730;
wire n_6258;
wire n_6905;
wire n_10243;
wire n_9700;
wire n_10564;
wire n_8682;
wire n_13829;
wire n_16533;
wire n_8089;
wire n_9218;
wire n_6704;
wire n_14657;
wire n_8533;
wire n_15483;
wire n_9118;
wire n_11122;
wire n_6657;
wire n_7655;
wire n_5554;
wire n_7244;
wire n_15925;
wire n_10745;
wire n_7368;
wire n_10596;
wire n_5553;
wire n_4485;
wire n_8011;
wire n_7633;
wire n_13937;
wire n_5711;
wire n_12140;
wire n_9437;
wire n_10263;
wire n_4340;
wire n_5790;
wire n_11509;
wire n_8640;
wire n_14359;
wire n_8063;
wire n_15141;
wire n_11960;
wire n_4855;
wire n_12599;
wire n_6186;
wire n_7878;
wire n_6803;
wire n_9514;
wire n_12411;
wire n_6210;
wire n_8437;
wire n_6500;
wire n_8427;
wire n_8032;
wire n_10280;
wire n_12465;
wire n_7427;
wire n_10605;
wire n_13532;
wire n_11029;
wire n_14013;
wire n_14419;
wire n_13250;
wire n_13118;
wire n_5404;
wire n_9933;
wire n_11449;
wire n_11190;
wire n_5739;
wire n_10951;
wire n_12152;
wire n_9892;
wire n_15251;
wire n_8570;
wire n_6163;
wire n_11794;
wire n_7628;
wire n_9462;
wire n_9074;
wire n_5972;
wire n_10519;
wire n_5549;
wire n_9408;
wire n_6785;
wire n_6553;
wire n_15854;
wire n_10454;
wire n_10163;
wire n_15401;
wire n_13339;
wire n_4940;
wire n_5444;
wire n_12568;
wire n_16163;
wire n_13478;
wire n_8039;
wire n_12501;
wire n_5757;
wire n_12970;
wire n_8902;
wire n_8916;
wire n_14295;
wire n_7557;
wire n_10087;
wire n_4356;
wire n_16544;
wire n_8843;
wire n_9891;
wire n_10146;
wire n_7128;
wire n_9946;
wire n_12959;
wire n_15810;
wire n_14367;
wire n_9885;
wire n_6849;
wire n_12330;
wire n_7594;
wire n_13915;
wire n_8129;
wire n_8162;
wire n_14819;
wire n_14890;
wire n_15057;
wire n_15871;
wire n_13906;
wire n_7457;
wire n_10643;
wire n_16300;
wire n_8744;
wire n_10504;
wire n_5824;
wire n_7788;
wire n_4361;
wire n_10872;
wire n_5488;
wire n_13783;
wire n_6760;
wire n_10701;
wire n_14265;
wire n_5154;
wire n_13664;
wire n_13987;
wire n_10658;
wire n_11590;
wire n_11238;
wire n_7752;
wire n_13566;
wire n_15626;
wire n_12591;
wire n_12466;
wire n_15775;
wire n_9509;
wire n_8286;
wire n_13416;
wire n_12798;
wire n_14885;
wire n_5329;
wire n_9015;
wire n_9925;
wire n_4367;
wire n_9757;
wire n_5637;
wire n_16066;
wire n_10874;
wire n_6825;
wire n_7586;
wire n_10008;
wire n_6452;
wire n_11831;
wire n_13726;
wire n_9628;
wire n_14399;
wire n_7767;
wire n_14412;
wire n_16213;
wire n_16408;
wire n_8294;
wire n_12279;
wire n_9419;
wire n_12243;
wire n_16402;
wire n_6611;
wire n_8562;
wire n_13705;
wire n_4560;
wire n_12614;
wire n_11378;
wire n_4899;
wire n_10250;
wire n_14631;
wire n_5728;
wire n_5471;
wire n_10032;
wire n_10592;
wire n_11433;
wire n_5164;
wire n_9277;
wire n_9257;
wire n_14063;
wire n_7207;
wire n_8218;
wire n_9806;
wire n_13425;
wire n_16657;
wire n_5843;
wire n_8170;
wire n_9159;
wire n_11558;
wire n_7744;
wire n_7021;
wire n_10595;
wire n_13591;
wire n_7748;
wire n_8537;
wire n_10126;
wire n_6827;
wire n_14421;
wire n_12041;
wire n_15890;
wire n_4663;
wire n_11713;
wire n_13653;
wire n_11073;
wire n_15586;
wire n_5484;
wire n_6355;
wire n_12566;
wire n_12931;
wire n_15525;
wire n_6227;
wire n_13680;
wire n_7215;
wire n_15157;
wire n_7485;
wire n_13074;
wire n_16077;
wire n_9066;
wire n_4802;
wire n_5523;
wire n_14332;
wire n_10302;
wire n_11974;
wire n_12881;
wire n_15736;
wire n_14986;
wire n_14920;
wire n_8016;
wire n_8671;
wire n_5423;
wire n_12546;
wire n_14716;
wire n_10645;
wire n_13058;
wire n_15313;
wire n_10604;
wire n_5074;
wire n_11096;
wire n_12036;
wire n_12876;
wire n_15286;
wire n_6564;
wire n_11161;
wire n_9671;
wire n_8782;
wire n_8709;
wire n_14698;
wire n_12911;
wire n_15715;
wire n_6468;
wire n_12491;
wire n_14994;
wire n_10080;
wire n_16505;
wire n_11216;
wire n_14368;
wire n_12228;
wire n_10570;
wire n_16120;
wire n_9857;
wire n_4701;
wire n_10966;
wire n_12781;
wire n_10057;
wire n_14323;
wire n_12929;
wire n_10882;
wire n_16065;
wire n_9338;
wire n_13071;
wire n_6857;
wire n_8144;
wire n_15075;
wire n_12261;
wire n_10435;
wire n_9542;
wire n_12536;
wire n_10795;
wire n_10921;
wire n_7171;
wire n_16333;
wire n_6442;
wire n_4851;
wire n_12106;
wire n_12061;
wire n_15116;
wire n_16200;
wire n_14585;
wire n_11085;
wire n_8049;
wire n_16041;
wire n_7762;
wire n_5204;
wire n_5333;
wire n_9467;
wire n_16541;
wire n_7068;
wire n_7925;
wire n_7186;
wire n_10609;
wire n_11157;
wire n_13739;
wire n_13649;
wire n_4991;
wire n_14804;
wire n_5594;
wire n_15126;
wire n_12291;
wire n_14510;
wire n_9097;
wire n_5422;
wire n_6871;
wire n_12124;
wire n_11755;
wire n_16497;
wire n_9783;
wire n_13806;
wire n_14364;
wire n_9510;
wire n_15472;
wire n_9389;
wire n_12074;
wire n_4934;
wire n_13497;
wire n_9404;
wire n_15406;
wire n_8357;
wire n_6904;
wire n_10912;
wire n_5087;
wire n_14396;
wire n_9916;
wire n_12645;
wire n_5526;
wire n_13234;
wire n_5292;
wire n_9314;
wire n_11918;
wire n_16198;
wire n_7017;
wire n_11748;
wire n_12433;
wire n_12745;
wire n_14466;
wire n_7777;
wire n_9752;
wire n_12138;
wire n_5000;
wire n_5403;
wire n_14473;
wire n_12887;
wire n_5551;
wire n_7652;
wire n_10220;
wire n_10341;
wire n_8701;
wire n_11347;
wire n_4479;
wire n_6499;
wire n_10550;
wire n_7830;
wire n_14673;
wire n_15816;
wire n_5131;
wire n_12217;
wire n_12365;
wire n_7138;
wire n_12097;
wire n_5257;
wire n_15922;
wire n_8097;
wire n_13738;
wire n_13851;
wire n_9679;
wire n_14972;
wire n_8084;
wire n_9306;
wire n_8645;
wire n_14138;
wire n_13272;
wire n_4753;
wire n_4688;
wire n_8712;
wire n_10232;
wire n_14113;
wire n_10461;
wire n_14586;
wire n_8289;
wire n_11178;
wire n_7966;
wire n_4848;
wire n_8591;
wire n_5059;
wire n_16411;
wire n_8837;
wire n_5887;
wire n_8811;
wire n_16428;
wire n_8824;
wire n_11673;
wire n_14938;
wire n_14784;
wire n_11432;
wire n_14641;
wire n_14179;
wire n_14031;
wire n_7191;
wire n_16506;
wire n_14979;
wire n_7712;
wire n_10412;
wire n_4475;
wire n_5242;
wire n_15433;
wire n_10326;
wire n_12650;
wire n_15953;
wire n_5219;
wire n_8417;
wire n_6276;
wire n_9721;
wire n_11344;
wire n_5631;
wire n_10499;
wire n_8340;
wire n_4443;
wire n_6008;
wire n_12487;
wire n_12658;
wire n_14324;
wire n_9197;
wire n_7997;
wire n_6420;
wire n_5854;
wire n_11387;
wire n_11333;
wire n_5460;
wire n_4587;
wire n_8455;
wire n_7208;
wire n_12288;
wire n_12859;
wire n_13613;
wire n_14740;
wire n_9210;
wire n_12185;
wire n_7961;
wire n_12130;
wire n_9770;
wire n_13120;
wire n_5686;
wire n_5899;
wire n_6893;
wire n_7406;
wire n_8681;
wire n_11417;
wire n_8905;
wire n_13008;
wire n_16044;
wire n_16299;
wire n_10617;
wire n_12271;
wire n_12704;
wire n_7807;
wire n_4749;
wire n_9592;
wire n_5155;
wire n_14198;
wire n_7680;
wire n_9180;
wire n_14846;
wire n_15190;
wire n_10922;
wire n_10544;
wire n_16524;
wire n_12958;
wire n_13030;
wire n_8172;
wire n_9917;
wire n_10718;
wire n_12056;
wire n_14539;
wire n_15094;
wire n_8106;
wire n_9502;
wire n_13821;
wire n_6447;
wire n_13712;
wire n_12238;
wire n_11952;
wire n_5981;
wire n_9625;
wire n_4891;
wire n_5937;
wire n_6422;
wire n_13896;
wire n_14761;
wire n_6751;
wire n_5339;
wire n_12976;
wire n_15243;
wire n_16473;
wire n_14420;
wire n_11087;
wire n_15041;
wire n_11477;
wire n_9873;
wire n_6040;
wire n_11888;
wire n_8375;
wire n_13299;
wire n_15393;
wire n_13243;
wire n_4464;
wire n_14314;
wire n_8612;
wire n_13042;
wire n_14144;
wire n_4624;
wire n_4818;
wire n_6851;
wire n_6460;
wire n_8345;
wire n_16642;
wire n_15658;
wire n_10095;
wire n_14227;
wire n_4659;
wire n_13725;
wire n_10309;
wire n_15873;
wire n_6741;
wire n_8459;
wire n_11773;
wire n_12608;
wire n_5217;
wire n_5465;
wire n_11099;
wire n_5015;
wire n_8974;
wire n_4339;
wire n_8268;
wire n_14164;
wire n_6160;
wire n_9871;
wire n_10050;
wire n_6650;
wire n_8221;
wire n_11682;
wire n_7066;
wire n_15595;
wire n_9164;
wire n_8255;
wire n_7183;
wire n_7789;
wire n_13197;
wire n_10306;
wire n_15081;
wire n_10878;
wire n_7606;
wire n_8461;
wire n_6192;
wire n_6368;
wire n_10056;
wire n_7140;
wire n_16597;
wire n_7193;
wire n_6039;
wire n_16474;
wire n_4487;
wire n_11919;
wire n_14860;
wire n_6583;
wire n_4889;
wire n_4866;
wire n_10450;
wire n_5721;
wire n_11414;
wire n_11472;
wire n_9114;
wire n_11978;
wire n_4816;
wire n_12520;
wire n_8515;
wire n_10529;
wire n_13632;
wire n_5719;
wire n_14685;
wire n_5773;
wire n_5482;
wire n_14892;
wire n_8812;
wire n_14505;
wire n_13020;
wire n_6012;
wire n_12254;
wire n_9392;
wire n_13148;
wire n_10429;
wire n_4937;
wire n_11459;
wire n_10904;
wire n_11317;
wire n_5277;
wire n_8792;
wire n_12436;
wire n_14531;
wire n_7344;
wire n_9888;
wire n_11470;
wire n_11538;
wire n_16344;
wire n_10037;
wire n_12808;
wire n_13871;
wire n_6707;
wire n_9698;
wire n_4874;
wire n_13435;
wire n_4401;
wire n_15408;
wire n_12744;
wire n_6064;
wire n_15173;
wire n_11136;
wire n_9903;
wire n_13801;
wire n_5793;
wire n_9644;
wire n_11353;
wire n_6787;
wire n_11102;
wire n_11620;
wire n_8523;
wire n_15480;
wire n_10179;
wire n_4709;
wire n_9228;
wire n_11539;
wire n_7710;
wire n_4976;
wire n_12143;
wire n_9499;
wire n_16166;
wire n_11899;
wire n_7892;
wire n_13168;
wire n_13879;
wire n_6647;
wire n_6275;
wire n_14038;
wire n_14771;
wire n_9522;
wire n_5578;
wire n_15617;
wire n_15463;
wire n_11215;
wire n_4658;
wire n_5296;
wire n_11076;
wire n_9366;
wire n_11890;
wire n_14339;
wire n_14253;
wire n_7915;
wire n_5893;
wire n_7750;
wire n_9077;
wire n_6769;
wire n_11597;
wire n_16005;
wire n_9148;
wire n_11806;
wire n_11054;
wire n_15902;
wire n_8406;
wire n_6277;
wire n_15919;
wire n_10754;
wire n_5742;
wire n_11050;
wire n_5207;
wire n_16652;
wire n_12443;
wire n_6463;
wire n_11683;
wire n_5676;
wire n_8554;
wire n_10920;
wire n_9275;
wire n_10223;
wire n_6051;
wire n_8896;
wire n_14398;
wire n_4665;
wire n_11484;
wire n_7206;
wire n_11126;
wire n_7538;
wire n_5674;
wire n_12934;
wire n_15758;
wire n_5539;
wire n_6895;
wire n_13598;
wire n_5282;
wire n_10295;
wire n_9409;
wire n_5464;
wire n_6799;
wire n_10336;
wire n_10228;
wire n_12555;
wire n_4362;
wire n_11646;
wire n_7716;
wire n_6487;
wire n_5121;
wire n_8758;
wire n_9768;
wire n_6026;
wire n_6070;
wire n_8818;
wire n_16648;
wire n_4430;
wire n_8617;
wire n_4348;
wire n_12980;
wire n_13966;
wire n_9881;
wire n_12530;
wire n_5013;
wire n_8954;
wire n_6807;
wire n_9463;
wire n_7251;
wire n_4489;
wire n_7254;
wire n_4839;
wire n_12212;
wire n_10466;
wire n_12973;
wire n_7540;
wire n_11953;
wire n_4404;
wire n_13123;
wire n_14669;
wire n_5589;
wire n_13077;
wire n_6563;
wire n_12234;
wire n_10776;
wire n_13231;
wire n_12624;
wire n_7882;
wire n_16309;
wire n_8552;
wire n_16348;
wire n_16514;
wire n_10425;
wire n_7554;
wire n_8069;
wire n_7558;
wire n_8373;
wire n_10848;
wire n_13165;
wire n_6481;
wire n_15926;
wire n_5628;
wire n_4825;
wire n_7765;
wire n_11482;
wire n_5006;
wire n_4513;
wire n_7816;
wire n_12151;
wire n_15201;
wire n_11089;
wire n_9997;
wire n_6341;
wire n_10164;
wire n_13422;
wire n_15809;
wire n_15204;
wire n_6384;
wire n_7421;
wire n_15579;
wire n_13828;
wire n_10166;
wire n_7489;
wire n_4747;
wire n_6906;
wire n_7541;
wire n_14702;
wire n_13179;
wire n_14562;
wire n_15585;
wire n_5251;
wire n_15844;
wire n_12033;
wire n_11839;
wire n_9844;
wire n_12826;
wire n_8318;
wire n_4801;
wire n_14376;
wire n_13834;
wire n_10366;
wire n_8341;
wire n_9970;
wire n_11193;
wire n_11365;
wire n_9595;
wire n_7188;
wire n_15015;
wire n_16081;
wire n_5475;
wire n_11217;
wire n_15651;
wire n_15555;
wire n_15341;
wire n_7334;
wire n_6923;
wire n_5807;
wire n_4448;
wire n_13923;
wire n_9287;
wire n_7991;
wire n_15477;
wire n_13051;
wire n_16376;
wire n_6233;
wire n_10877;
wire n_6377;
wire n_11524;
wire n_9265;
wire n_12402;
wire n_5216;
wire n_14991;
wire n_14686;
wire n_12214;
wire n_10225;
wire n_4869;
wire n_8239;
wire n_16114;
wire n_13330;
wire n_16259;
wire n_8926;
wire n_6257;
wire n_4386;
wire n_10361;
wire n_11228;
wire n_5273;
wire n_7898;
wire n_10766;
wire n_4438;
wire n_4844;
wire n_8383;
wire n_10086;
wire n_4836;
wire n_5439;
wire n_7143;
wire n_9789;
wire n_10424;
wire n_12621;
wire n_13924;
wire n_4955;
wire n_8965;
wire n_11290;
wire n_5936;
wire n_12518;
wire n_9608;
wire n_4355;
wire n_7646;
wire n_9052;
wire n_13476;
wire n_14047;
wire n_8817;
wire n_8190;
wire n_11488;
wire n_13671;
wire n_16033;
wire n_12162;
wire n_6587;
wire n_14627;
wire n_14876;
wire n_6987;
wire n_7781;
wire n_7360;
wire n_11037;
wire n_14568;
wire n_11702;
wire n_6069;
wire n_13699;
wire n_14319;
wire n_7497;
wire n_4655;
wire n_11372;
wire n_5706;
wire n_7665;
wire n_9354;
wire n_10501;
wire n_10817;
wire n_11829;
wire n_14026;
wire n_15324;
wire n_11517;
wire n_7793;
wire n_16102;
wire n_16274;
wire n_8355;
wire n_6991;
wire n_10556;
wire n_15287;
wire n_12741;
wire n_7101;
wire n_7671;
wire n_9436;
wire n_7530;
wire n_8489;
wire n_13150;
wire n_15006;
wire n_13776;
wire n_5431;
wire n_15103;
wire n_15619;
wire n_7248;
wire n_4357;
wire n_10350;
wire n_12541;
wire n_7204;
wire n_12730;
wire n_9860;
wire n_8649;
wire n_12510;
wire n_15835;
wire n_12852;
wire n_6887;
wire n_11756;
wire n_10567;
wire n_7578;
wire n_14818;
wire n_13343;
wire n_7654;
wire n_16123;
wire n_13152;
wire n_8303;
wire n_6153;
wire n_4374;
wire n_5132;
wire n_6637;
wire n_8369;
wire n_9022;
wire n_9238;
wire n_16512;
wire n_13809;
wire n_8059;
wire n_6633;
wire n_10230;
wire n_12675;
wire n_5627;
wire n_9103;
wire n_11031;
wire n_5774;
wire n_6579;
wire n_11665;
wire n_13590;
wire n_13907;
wire n_4400;
wire n_4846;
wire n_5798;
wire n_11138;
wire n_11731;
wire n_16103;
wire n_5875;
wire n_5187;
wire n_9839;
wire n_12821;
wire n_14782;
wire n_16257;
wire n_8831;
wire n_5621;
wire n_5608;
wire n_7900;
wire n_15704;
wire n_6569;
wire n_6335;
wire n_7120;
wire n_8728;
wire n_10807;
wire n_12478;
wire n_12837;
wire n_12233;
wire n_6789;
wire n_8386;
wire n_12100;
wire n_8853;
wire n_14070;
wire n_4582;
wire n_14330;
wire n_15327;
wire n_13491;
wire n_6252;
wire n_13545;
wire n_13471;
wire n_13760;
wire n_13883;
wire n_4860;
wire n_6211;
wire n_15716;
wire n_10511;
wire n_5844;
wire n_8862;
wire n_15748;
wire n_16161;
wire n_10580;
wire n_14235;
wire n_4870;
wire n_6164;
wire n_13261;
wire n_7576;
wire n_6173;
wire n_8081;
wire n_9675;
wire n_14851;
wire n_16608;
wire n_7786;
wire n_11023;
wire n_7313;
wire n_10058;
wire n_16471;
wire n_10873;
wire n_14484;
wire n_4989;
wire n_7676;
wire n_7609;
wire n_7757;
wire n_11454;
wire n_13442;
wire n_8900;
wire n_12523;
wire n_14444;
wire n_6630;
wire n_6934;
wire n_9017;
wire n_10484;
wire n_4558;
wire n_6737;
wire n_11744;
wire n_4488;
wire n_15726;
wire n_8396;
wire n_16560;
wire n_6612;
wire n_14307;
wire n_8478;
wire n_6606;
wire n_13450;
wire n_6695;
wire n_12395;
wire n_8865;
wire n_10288;
wire n_10337;
wire n_15302;
wire n_7779;
wire n_8999;
wire n_6189;
wire n_10388;
wire n_14178;
wire n_11626;
wire n_12148;
wire n_11072;
wire n_15299;
wire n_5867;
wire n_5508;
wire n_6479;
wire n_4656;
wire n_10791;
wire n_10506;
wire n_12907;
wire n_16312;
wire n_15500;
wire n_8497;
wire n_10770;
wire n_16204;
wire n_8820;
wire n_6410;
wire n_14891;
wire n_9318;
wire n_6158;
wire n_11917;
wire n_5597;
wire n_9028;
wire n_13944;
wire n_4915;
wire n_4328;
wire n_9492;
wire n_15592;
wire n_6413;
wire n_6090;
wire n_8020;
wire n_16064;
wire n_16443;
wire n_9374;
wire n_7419;
wire n_15319;
wire n_6506;
wire n_5515;
wire n_5662;
wire n_13634;
wire n_12132;
wire n_6935;
wire n_9727;
wire n_10413;
wire n_10593;
wire n_13019;
wire n_14452;
wire n_5862;
wire n_12703;
wire n_13079;
wire n_13464;
wire n_4397;
wire n_12182;
wire n_12670;
wire n_5050;
wire n_10636;
wire n_12043;
wire n_4808;
wire n_7667;
wire n_16478;
wire n_5697;
wire n_10203;
wire n_10980;
wire n_9174;
wire n_5767;
wire n_15369;
wire n_8992;
wire n_15134;
wire n_12708;
wire n_16110;
wire n_4712;
wire n_8880;
wire n_10369;
wire n_8690;
wire n_6234;
wire n_6821;
wire n_5462;
wire n_9983;
wire n_9375;
wire n_10082;
wire n_6688;
wire n_5980;
wire n_8580;
wire n_7818;
wire n_9993;
wire n_8770;
wire n_11721;
wire n_7182;
wire n_15453;
wire n_5318;
wire n_7365;
wire n_13573;
wire n_6608;
wire n_10467;
wire n_9109;
wire n_9849;
wire n_13622;
wire n_6105;
wire n_4725;
wire n_6022;
wire n_11207;
wire n_9856;
wire n_10964;
wire n_4406;
wire n_5498;
wire n_12493;
wire n_13135;
wire n_8075;
wire n_6798;
wire n_10838;
wire n_10530;
wire n_5053;
wire n_7896;
wire n_7841;
wire n_9458;
wire n_12482;
wire n_14794;
wire n_9237;
wire n_13931;
wire n_11668;
wire n_7885;
wire n_15208;
wire n_15684;
wire n_6860;
wire n_6557;
wire n_14404;
wire n_8466;
wire n_6753;
wire n_12137;
wire n_6527;
wire n_7341;
wire n_11328;
wire n_9349;
wire n_12306;
wire n_15275;
wire n_4908;
wire n_11200;
wire n_12088;
wire n_14442;
wire n_15210;
wire n_15423;
wire n_11091;
wire n_8094;
wire n_10940;
wire n_14377;
wire n_16463;
wire n_15976;
wire n_16536;
wire n_6639;
wire n_4824;
wire n_12508;
wire n_4567;
wire n_12096;
wire n_6430;
wire n_5150;
wire n_13418;
wire n_8832;
wire n_10987;
wire n_4778;
wire n_5477;
wire n_12684;
wire n_5175;
wire n_8839;
wire n_7996;
wire n_4595;
wire n_12891;
wire n_11098;
wire n_15815;
wire n_11615;
wire n_10533;
wire n_11059;
wire n_5987;
wire n_16403;
wire n_5179;
wire n_7957;
wire n_14616;
wire n_11965;
wire n_4904;
wire n_10938;
wire n_16681;
wire n_10176;
wire n_7517;
wire n_6627;
wire n_8080;
wire n_14696;
wire n_5988;
wire n_5585;
wire n_15093;
wire n_12324;
wire n_12345;
wire n_6058;
wire n_7745;
wire n_12941;
wire n_13551;
wire n_14006;
wire n_6666;
wire n_10927;
wire n_14258;
wire n_12200;
wire n_4616;
wire n_8321;
wire n_16060;
wire n_14024;
wire n_8772;
wire n_8735;
wire n_9954;
wire n_4982;
wire n_11722;
wire n_8786;
wire n_8592;
wire n_15597;
wire n_11204;
wire n_8684;
wire n_6190;
wire n_4643;
wire n_13682;
wire n_6249;
wire n_12694;
wire n_12701;
wire n_8083;
wire n_12310;
wire n_5348;
wire n_11060;
wire n_10578;
wire n_6594;
wire n_9805;
wire n_10155;
wire n_5480;
wire n_4323;
wire n_16199;
wire n_13593;
wire n_8157;
wire n_4831;
wire n_7095;
wire n_11461;
wire n_13902;
wire n_10714;
wire n_11701;
wire n_16672;
wire n_6969;
wire n_6615;
wire n_7459;
wire n_6161;
wire n_8206;
wire n_7294;
wire n_4896;
wire n_4916;
wire n_9110;
wire n_11811;
wire n_13745;
wire n_10569;
wire n_8622;
wire n_5904;
wire n_13917;
wire n_4739;
wire n_15367;
wire n_7184;
wire n_9617;
wire n_6607;
wire n_9335;
wire n_13546;
wire n_14595;
wire n_14468;
wire n_6062;
wire n_7908;
wire n_12550;
wire n_9452;
wire n_7974;
wire n_7551;
wire n_11427;
wire n_11980;
wire n_13350;
wire n_13861;
wire n_10051;
wire n_8104;
wire n_10414;
wire n_11255;
wire n_8344;
wire n_13592;
wire n_5284;
wire n_11720;
wire n_12673;
wire n_14694;
wire n_8120;
wire n_8513;
wire n_10120;
wire n_9474;
wire n_5461;
wire n_9075;
wire n_12961;
wire n_13874;
wire n_6482;
wire n_9427;
wire n_11496;
wire n_10746;
wire n_12225;
wire n_9188;
wire n_6294;
wire n_16407;
wire n_5147;
wire n_9611;
wire n_15506;
wire n_4644;
wire n_9021;
wire n_8779;
wire n_9810;
wire n_14469;
wire n_16269;
wire n_8621;
wire n_5503;
wire n_5845;
wire n_9250;
wire n_5945;
wire n_9550;
wire n_11212;
wire n_12884;
wire n_13145;
wire n_16591;
wire n_10697;
wire n_11714;
wire n_16201;
wire n_16179;
wire n_11263;
wire n_10641;
wire n_6246;
wire n_8868;
wire n_15070;
wire n_8134;
wire n_4716;
wire n_12207;
wire n_9975;
wire n_7250;
wire n_5755;
wire n_5600;
wire n_16566;
wire n_8762;
wire n_12011;
wire n_13195;
wire n_8043;
wire n_8694;
wire n_16377;
wire n_14492;
wire n_13965;
wire n_6053;
wire n_5048;
wire n_11994;
wire n_7252;
wire n_13419;
wire n_9207;
wire n_13358;
wire n_14134;
wire n_4944;
wire n_11860;
wire n_11990;
wire n_10103;
wire n_5245;
wire n_4343;
wire n_6843;
wire n_10926;
wire n_14519;
wire n_4715;
wire n_6123;
wire n_8897;
wire n_11000;
wire n_16125;
wire n_10626;
wire n_15457;
wire n_6901;
wire n_14345;
wire n_4935;
wire n_13273;
wire n_4694;
wire n_11503;
wire n_8191;
wire n_10325;
wire n_6841;
wire n_4672;
wire n_10153;
wire n_16354;
wire n_8101;
wire n_5054;
wire n_10298;
wire n_8376;
wire n_8171;
wire n_5448;
wire n_6922;
wire n_9006;
wire n_7698;
wire n_5749;
wire n_6774;
wire n_12854;
wire n_15640;
wire n_6271;
wire n_6489;
wire n_8600;
wire n_16427;
wire n_4407;
wire n_7402;
wire n_8431;
wire n_14816;
wire n_8710;
wire n_15683;
wire n_12806;
wire n_16336;
wire n_4598;
wire n_16202;
wire n_16248;
wire n_14302;
wire n_8599;
wire n_8549;
wire n_13460;
wire n_15451;
wire n_10172;
wire n_5993;
wire n_8054;
wire n_11273;
wire n_13904;
wire n_16614;
wire n_10400;
wire n_15233;
wire n_6716;
wire n_9637;
wire n_11636;
wire n_9418;
wire n_8616;
wire n_4524;
wire n_6020;
wire n_12472;
wire n_9177;
wire n_9060;
wire n_13105;
wire n_11947;
wire n_14035;
wire n_14496;
wire n_14467;
wire n_13218;
wire n_9096;
wire n_9081;
wire n_13952;
wire n_11697;
wire n_14789;
wire n_15784;
wire n_13076;
wire n_15526;
wire n_9236;
wire n_6844;
wire n_11762;
wire n_11969;
wire n_12950;
wire n_7914;
wire n_8628;
wire n_16388;
wire n_6521;
wire n_7891;
wire n_15150;
wire n_13028;
wire n_14413;
wire n_8857;
wire n_8517;
wire n_4850;
wire n_14243;
wire n_8547;
wire n_10156;
wire n_4424;
wire n_9040;
wire n_7113;
wire n_9607;
wire n_6162;
wire n_10433;
wire n_6779;
wire n_8010;
wire n_6432;
wire n_4776;
wire n_9116;
wire n_14096;
wire n_10774;
wire n_12332;
wire n_10901;
wire n_11034;
wire n_11983;
wire n_10549;
wire n_10839;
wire n_12115;
wire n_11813;
wire n_7216;
wire n_12762;
wire n_13574;
wire n_11499;
wire n_15990;
wire n_15364;
wire n_10825;
wire n_14583;
wire n_14893;
wire n_8275;
wire n_6198;
wire n_4723;
wire n_5418;
wire n_6543;
wire n_9830;
wire n_6762;
wire n_6178;
wire n_9621;
wire n_5685;
wire n_10761;
wire n_14777;
wire n_14057;
wire n_5459;
wire n_9035;
wire n_11579;
wire n_16117;
wire n_10398;
wire n_15303;
wire n_8291;
wire n_16459;
wire n_11535;
wire n_15661;
wire n_16406;
wire n_12558;
wire n_14915;
wire n_4650;
wire n_11984;
wire n_11948;
wire n_7706;
wire n_4719;
wire n_5173;
wire n_7477;
wire n_5016;
wire n_15654;
wire n_12975;
wire n_11402;
wire n_6458;
wire n_7642;
wire n_4967;
wire n_9678;
wire n_11401;
wire n_8247;
wire n_6577;
wire n_12506;
wire n_16291;
wire n_13850;
wire n_6740;
wire n_12718;
wire n_12956;
wire n_11510;
wire n_6315;
wire n_10581;
wire n_12638;
wire n_14116;
wire n_14856;
wire n_14949;
wire n_4912;
wire n_15235;
wire n_4799;
wire n_9284;
wire n_12736;
wire n_4423;
wire n_5086;
wire n_5283;
wire n_9111;
wire n_7156;
wire n_4735;
wire n_9163;
wire n_15461;
wire n_12086;
wire n_15711;
wire n_16453;
wire n_16645;
wire n_5170;
wire n_6910;
wire n_7604;
wire n_6262;
wire n_14800;
wire n_7703;
wire n_9606;
wire n_6319;
wire n_13459;
wire n_10470;
wire n_16449;
wire n_14268;
wire n_11589;
wire n_10297;
wire n_11246;
wire n_12553;
wire n_14888;
wire n_15034;
wire n_12350;
wire n_12542;
wire n_13860;
wire n_5839;
wire n_5028;
wire n_14240;
wire n_14504;
wire n_13449;
wire n_14127;
wire n_6536;
wire n_12747;
wire n_6175;
wire n_16209;
wire n_7040;
wire n_8827;
wire n_10625;
wire n_8280;
wire n_12561;
wire n_16606;
wire n_12390;
wire n_14460;
wire n_5514;
wire n_13216;
wire n_8388;
wire n_12849;
wire n_14730;
wire n_10235;
wire n_11312;
wire n_6978;
wire n_13786;
wire n_9589;
wire n_5351;
wire n_5909;
wire n_9344;
wire n_12805;
wire n_10865;
wire n_9549;
wire n_6093;
wire n_11649;
wire n_4543;
wire n_10445;
wire n_15110;
wire n_16306;
wire n_7378;
wire n_10738;
wire n_14894;
wire n_12866;
wire n_8988;
wire n_6845;
wire n_9798;
wire n_15491;
wire n_15025;
wire n_9190;
wire n_14925;
wire n_6947;
wire n_11612;
wire n_14918;
wire n_9482;
wire n_5293;
wire n_12447;
wire n_13417;
wire n_12296;
wire n_8203;
wire n_6099;
wire n_12900;
wire n_13414;
wire n_8569;
wire n_5400;
wire n_14598;
wire n_4892;
wire n_6140;
wire n_8877;
wire n_15489;
wire n_9412;
wire n_7498;
wire n_10679;
wire n_11323;
wire n_10799;
wire n_15561;
wire n_6321;
wire n_12914;
wire n_11916;
wire n_6819;
wire n_7501;
wire n_5201;
wire n_9506;
wire n_10136;
wire n_10421;
wire n_5890;
wire n_6415;
wire n_10976;
wire n_6465;
wire n_9447;
wire n_4439;
wire n_10585;
wire n_12764;
wire n_13696;
wire n_15148;
wire n_15325;
wire n_4783;
wire n_11356;
wire n_16457;
wire n_16542;
wire n_15955;
wire n_12948;
wire n_7931;
wire n_8688;
wire n_10828;
wire n_13322;
wire n_15158;
wire n_14238;
wire n_9092;
wire n_10034;
wire n_9451;
wire n_4910;
wire n_11148;
wire n_12409;
wire n_11625;
wire n_12300;
wire n_13934;
wire n_6899;
wire n_15389;
wire n_7549;
wire n_10692;
wire n_7373;
wire n_7895;
wire n_11281;
wire n_13056;
wire n_14826;
wire n_15331;
wire n_15776;
wire n_16019;
wire n_16421;
wire n_6592;
wire n_11280;
wire n_12337;
wire n_13254;
wire n_14987;
wire n_13466;
wire n_15082;
wire n_15191;
wire n_8686;
wire n_12239;
wire n_8871;
wire n_9712;
wire n_6626;
wire n_8585;
wire n_8951;
wire n_5389;
wire n_5142;
wire n_11114;
wire n_15676;
wire n_9011;
wire n_16023;
wire n_8418;
wire n_7740;
wire n_8403;
wire n_5891;
wire n_13050;
wire n_14042;
wire n_7613;
wire n_11493;
wire n_6101;
wire n_9220;
wire n_14440;
wire n_7556;
wire n_5935;
wire n_10528;
wire n_10860;
wire n_12763;
wire n_4930;
wire n_16208;
wire n_8588;
wire n_15229;
wire n_11339;
wire n_15804;
wire n_5623;
wire n_15209;
wire n_15269;
wire n_12273;
wire n_13875;
wire n_16394;
wire n_8564;
wire n_11943;
wire n_6944;
wire n_9121;
wire n_10471;
wire n_15310;
wire n_12712;
wire n_14076;
wire n_11220;
wire n_9012;
wire n_15078;
wire n_4557;
wire n_13012;
wire n_4917;
wire n_8698;
wire n_8924;
wire n_12584;
wire n_14435;
wire n_4432;
wire n_14638;
wire n_14946;
wire n_10376;
wire n_15510;
wire n_12752;
wire n_15674;
wire n_4352;
wire n_7515;
wire n_6928;
wire n_4416;
wire n_10880;
wire n_15511;
wire n_4593;
wire n_7238;
wire n_9994;
wire n_4465;
wire n_14226;
wire n_8780;
wire n_7309;
wire n_15811;
wire n_14936;
wire n_5114;
wire n_7958;
wire n_16469;
wire n_4980;
wire n_8047;
wire n_11596;
wire n_8559;
wire n_5693;
wire n_4495;
wire n_6273;
wire n_14278;
wire n_11885;
wire n_5117;
wire n_15618;
wire n_7572;
wire n_5663;
wire n_11955;
wire n_8214;
wire n_10224;
wire n_12777;
wire n_14706;
wire n_15849;
wire n_5990;
wire n_7043;
wire n_10777;
wire n_11462;
wire n_11732;
wire n_16156;
wire n_16490;
wire n_5024;
wire n_9391;
wire n_7760;
wire n_4559;
wire n_16105;
wire n_8514;
wire n_9134;
wire n_9753;
wire n_13306;
wire n_12819;
wire n_14159;
wire n_14515;
wire n_8722;
wire n_16489;
wire n_11654;
wire n_12268;
wire n_10214;
wire n_8241;
wire n_8589;
wire n_12077;
wire n_12982;
wire n_7573;
wire n_8442;
wire n_15321;
wire n_6281;
wire n_11619;
wire n_10649;
wire n_7364;
wire n_5647;
wire n_13133;
wire n_14757;
wire n_4938;
wire n_5396;
wire n_9572;
wire n_8608;
wire n_5203;
wire n_12874;
wire n_12534;
wire n_6846;
wire n_6311;
wire n_10469;
wire n_9229;
wire n_11480;
wire n_11194;
wire n_15282;
wire n_16038;
wire n_7590;
wire n_9342;
wire n_12237;
wire n_13271;
wire n_5162;
wire n_6134;
wire n_9329;
wire n_5426;
wire n_10175;
wire n_5803;
wire n_11481;
wire n_13372;
wire n_15812;
wire n_16292;
wire n_9868;
wire n_11375;
wire n_5285;
wire n_11267;
wire n_9602;
wire n_7048;
wire n_6886;
wire n_4335;
wire n_9311;
wire n_12275;
wire n_6593;
wire n_13742;
wire n_8630;
wire n_15177;
wire n_16491;
wire n_12376;
wire n_9884;
wire n_5365;
wire n_13114;
wire n_9876;
wire n_8583;
wire n_4521;
wire n_8145;
wire n_8405;
wire n_10447;
wire n_9260;
wire n_15063;
wire n_7176;
wire n_14534;
wire n_8928;
wire n_13630;
wire n_7682;
wire n_15223;
wire n_9353;
wire n_11350;
wire n_13054;
wire n_16535;
wire n_11925;
wire n_13700;
wire n_6231;
wire n_8948;
wire n_8672;
wire n_10406;
wire n_5715;
wire n_12509;
wire n_14902;
wire n_4920;
wire n_8295;
wire n_6932;
wire n_6746;
wire n_11985;
wire n_13527;
wire n_8447;
wire n_7901;
wire n_5395;
wire n_10522;
wire n_6443;
wire n_5709;
wire n_7658;
wire n_13793;
wire n_11782;
wire n_16532;
wire n_6446;
wire n_16618;
wire n_10278;
wire n_14290;
wire n_10055;
wire n_10979;
wire n_7980;
wire n_6996;
wire n_7218;
wire n_8828;
wire n_9430;
wire n_15935;
wire n_15384;
wire n_11407;
wire n_13882;
wire n_9750;
wire n_9749;
wire n_14139;
wire n_12710;
wire n_15686;
wire n_6749;
wire n_9263;
wire n_11082;
wire n_8440;
wire n_7005;
wire n_15950;
wire n_10408;
wire n_16180;
wire n_8572;
wire n_10965;
wire n_10798;
wire n_7732;
wire n_13325;
wire n_6337;
wire n_14850;
wire n_6181;
wire n_15135;
wire n_16196;
wire n_7447;
wire n_9776;
wire n_11911;
wire n_6777;
wire n_11987;
wire n_11442;
wire n_8227;
wire n_12936;
wire n_12721;
wire n_5634;
wire n_5672;
wire n_16008;
wire n_8475;
wire n_11730;
wire n_10482;
wire n_6924;
wire n_8029;
wire n_9804;
wire n_14064;
wire n_14524;
wire n_4861;
wire n_9304;
wire n_5799;
wire n_8859;
wire n_8380;
wire n_7405;
wire n_12039;
wire n_4926;
wire n_11388;
wire n_11651;
wire n_14151;
wire n_8314;
wire n_9386;
wire n_15120;
wire n_10154;
wire n_5617;
wire n_7922;
wire n_13089;
wire n_15826;
wire n_15459;
wire n_15192;
wire n_10377;
wire n_5266;
wire n_5580;
wire n_4828;
wire n_10033;
wire n_9926;
wire n_11121;
wire n_13167;
wire n_11270;
wire n_12329;
wire n_6310;
wire n_15161;
wire n_11689;
wire n_10003;
wire n_15601;
wire n_15936;
wire n_8311;
wire n_10858;
wire n_10321;
wire n_5450;
wire n_12253;
wire n_15005;
wire n_11147;
wire n_12928;
wire n_5310;
wire n_9661;
wire n_16303;
wire n_9843;
wire n_15013;
wire n_9877;
wire n_8764;
wire n_14284;
wire n_6953;
wire n_14945;
wire n_16559;
wire n_5722;
wire n_4640;
wire n_5122;
wire n_13001;
wire n_5390;
wire n_13232;
wire n_9901;
wire n_16167;
wire n_13320;
wire n_5593;
wire n_12990;
wire n_14246;
wire n_6683;
wire n_4769;
wire n_10683;
wire n_5764;
wire n_9834;
wire n_8934;
wire n_13059;
wire n_16353;
wire n_6365;
wire n_4628;
wire n_6920;
wire n_9921;
wire n_12318;
wire n_8407;
wire n_6229;
wire n_8567;
wire n_5385;
wire n_11817;
wire n_13278;
wire n_15455;
wire n_8729;
wire n_11288;
wire n_12772;
wire n_10359;
wire n_5237;
wire n_13597;
wire n_14957;
wire n_5133;
wire n_13488;
wire n_11042;
wire n_6907;
wire n_5322;
wire n_10726;
wire n_13447;
wire n_15907;
wire n_7089;
wire n_7144;
wire n_16534;
wire n_7286;
wire n_16579;
wire n_11479;
wire n_11737;
wire n_4460;
wire n_8048;
wire n_14681;
wire n_12028;
wire n_13668;
wire n_13016;
wire n_7072;
wire n_11272;
wire n_14230;
wire n_13095;
wire n_8253;
wire n_6177;
wire n_14708;
wire n_6332;
wire n_5853;
wire n_12048;
wire n_15032;
wire n_8283;
wire n_5982;
wire n_10930;
wire n_11600;
wire n_16607;
wire n_15085;
wire n_16390;
wire n_8749;
wire n_8088;
wire n_7403;
wire n_10722;
wire n_5011;
wire n_10666;
wire n_7338;
wire n_5917;
wire n_14546;
wire n_7129;
wire n_4909;
wire n_13938;
wire n_12057;
wire n_6696;
wire n_15440;
wire n_13251;
wire n_9882;
wire n_9527;
wire n_16484;
wire n_8566;
wire n_16450;
wire n_7343;
wire n_12766;
wire n_14875;
wire n_8516;
wire n_10637;
wire n_8302;
wire n_15056;
wire n_8317;
wire n_15860;
wire n_5376;
wire n_15610;
wire n_12229;
wire n_14003;
wire n_16197;
wire n_5106;
wire n_9205;
wire n_6116;
wire n_9511;
wire n_8167;
wire n_15329;
wire n_7859;
wire n_14315;
wire n_6730;
wire n_7492;
wire n_7872;
wire n_13670;
wire n_7972;
wire n_11254;
wire n_13319;
wire n_15023;
wire n_4768;
wire n_11617;
wire n_13858;
wire n_13512;
wire n_9071;
wire n_7916;
wire n_9368;
wire n_7480;
wire n_7694;
wire n_5561;
wire n_10415;
wire n_13069;
wire n_11711;
wire n_5410;
wire n_12362;
wire n_8944;
wire n_6167;
wire n_15666;
wire n_16255;
wire n_13233;
wire n_11931;
wire n_8008;
wire n_10023;
wire n_10999;
wire n_6170;
wire n_8109;
wire n_13297;
wire n_9459;
wire n_14185;
wire n_5156;
wire n_12780;
wire n_13267;
wire n_14017;
wire n_6307;
wire n_10410;
wire n_6094;
wire n_9098;
wire n_7987;
wire n_7483;
wire n_4447;
wire n_14953;
wire n_9133;
wire n_16054;
wire n_12664;
wire n_14942;
wire n_14873;
wire n_15604;
wire n_7434;
wire n_4826;
wire n_9009;
wire n_6155;
wire n_7269;
wire n_9777;
wire n_9504;
wire n_15359;
wire n_14840;
wire n_8975;
wire n_16556;
wire n_6267;
wire n_16000;
wire n_9063;
wire n_7787;
wire n_12360;
wire n_5998;
wire n_9268;
wire n_15431;
wire n_5304;
wire n_6568;
wire n_15035;
wire n_8673;
wire n_7507;
wire n_7159;
wire n_11305;
wire n_5378;
wire n_6028;
wire n_9101;
wire n_10456;
wire n_15631;
wire n_16072;
wire n_6261;
wire n_14083;
wire n_13186;
wire n_5916;
wire n_11907;
wire n_15655;
wire n_4648;
wire n_10096;
wire n_13617;
wire n_10025;
wire n_10627;
wire n_10475;
wire n_10189;
wire n_8697;
wire n_14755;
wire n_6299;
wire n_6813;
wire n_8825;
wire n_12969;
wire n_15430;
wire n_11753;
wire n_7425;
wire n_12260;
wire n_12016;
wire n_6669;
wire n_8581;
wire n_15732;
wire n_8266;
wire n_5691;
wire n_12457;
wire n_16070;
wire n_16045;
wire n_4951;
wire n_8981;
wire n_8420;
wire n_4957;
wire n_8297;
wire n_11150;
wire n_4360;
wire n_8771;
wire n_10881;
wire n_13519;
wire n_16111;
wire n_15750;
wire n_14170;
wire n_16583;
wire n_15641;
wire n_13496;
wire n_4566;
wire n_16007;
wire n_12939;
wire n_6316;
wire n_15038;
wire n_6292;
wire n_4853;
wire n_9726;
wire n_13884;
wire n_10404;
wire n_8639;
wire n_8138;
wire n_8058;
wire n_9308;
wire n_6638;
wire n_12779;
wire n_11838;
wire n_10508;
wire n_16510;
wire n_7719;
wire n_15892;
wire n_10811;
wire n_14049;
wire n_8333;
wire n_5615;
wire n_6220;
wire n_7562;
wire n_15531;
wire n_13547;
wire n_12816;
wire n_7619;
wire n_6985;
wire n_12783;
wire n_7170;
wire n_13853;
wire n_9211;
wire n_12019;
wire n_8176;
wire n_8124;
wire n_14529;
wire n_8823;
wire n_7366;
wire n_9395;
wire n_16106;
wire n_5269;
wire n_10891;
wire n_11457;
wire n_12751;
wire n_9026;
wire n_15284;
wire n_10803;
wire n_8147;
wire n_13190;
wire n_5468;
wire n_6188;
wire n_4730;
wire n_5399;
wire n_8127;
wire n_9402;
wire n_14014;
wire n_14195;
wire n_5262;
wire n_10700;
wire n_7938;
wire n_4670;
wire n_10968;
wire n_4882;
wire n_11695;
wire n_4620;
wire n_7935;
wire n_4738;
wire n_8458;
wire n_5421;
wire n_14247;
wire n_6772;
wire n_8113;
wire n_9716;
wire n_16646;
wire n_15877;
wire n_14300;
wire n_11453;
wire n_16155;
wire n_15443;
wire n_5206;
wire n_6077;
wire n_5713;
wire n_11512;
wire n_5256;
wire n_6318;
wire n_15418;
wire n_16445;
wire n_11970;
wire n_14678;
wire n_7918;
wire n_13599;
wire n_4517;
wire n_13354;
wire n_14690;
wire n_15008;
wire n_5188;
wire n_13647;
wire n_6916;
wire n_15524;
wire n_4490;
wire n_13683;
wire n_6651;
wire n_12308;
wire n_10290;
wire n_10783;
wire n_11862;
wire n_10147;
wire n_12163;
wire n_14839;
wire n_10725;
wire n_11523;
wire n_7845;
wire n_12688;
wire n_5550;
wire n_12944;
wire n_15409;
wire n_8290;
wire n_7536;
wire n_7472;
wire n_16207;
wire n_9433;
wire n_9737;
wire n_9298;
wire n_11660;
wire n_10812;
wire n_14709;
wire n_12297;
wire n_13848;
wire n_6366;
wire n_14249;
wire n_6230;
wire n_14241;
wire n_6604;
wire n_14497;
wire n_16108;
wire n_5161;
wire n_5373;
wire n_10001;
wire n_16101;
wire n_11107;
wire n_14280;
wire n_13724;
wire n_13280;
wire n_9301;
wire n_12145;
wire n_11088;
wire n_5573;
wire n_5939;
wire n_5509;
wire n_8160;
wire n_6391;
wire n_5382;
wire n_10284;
wire n_12757;
wire n_12054;
wire n_15827;
wire n_14379;
wire n_5659;
wire n_8099;
wire n_14446;
wire n_11595;
wire n_8840;
wire n_16284;
wire n_11405;
wire n_14719;
wire n_16001;
wire n_15575;
wire n_13768;
wire n_13189;
wire n_5881;
wire n_8522;
wire n_12971;
wire n_7222;
wire n_7942;
wire n_8578;
wire n_6473;
wire n_13103;
wire n_13838;
wire n_15630;
wire n_16599;
wire n_10046;
wire n_15696;
wire n_12328;
wire n_14558;
wire n_11318;
wire n_9083;
wire n_7725;
wire n_10977;
wire n_11299;
wire n_10397;
wire n_6483;
wire n_10615;
wire n_10994;
wire n_11542;
wire n_14004;
wire n_5863;
wire n_7647;
wire n_8626;
wire n_10936;
wire n_12442;
wire n_16221;
wire n_8611;
wire n_8036;
wire n_8819;
wire n_11485;
wire n_12426;
wire n_16222;
wire n_15123;
wire n_9835;
wire n_15068;
wire n_15442;
wire n_7300;
wire n_15021;
wire n_12839;
wire n_6697;
wire n_9054;
wire n_7875;
wire n_13153;
wire n_6975;
wire n_4446;
wire n_14666;
wire n_13605;
wire n_10532;
wire n_4417;
wire n_5466;
wire n_13995;
wire n_7643;
wire n_13073;
wire n_11048;
wire n_4733;
wire n_13441;
wire n_6729;
wire n_6728;
wire n_4764;
wire n_14237;
wire n_16082;
wire n_15095;
wire n_11240;
wire n_4743;
wire n_10207;
wire n_13857;
wire n_13841;
wire n_16029;
wire n_13556;
wire n_10401;
wire n_11634;
wire n_12580;
wire n_13367;
wire n_5955;
wire n_7242;
wire n_10013;
wire n_10771;
wire n_13816;
wire n_11487;
wire n_11441;
wire n_8441;
wire n_16119;
wire n_14203;
wire n_6076;
wire n_8933;
wire n_15876;
wire n_7778;
wire n_15231;
wire n_12844;
wire n_5851;
wire n_14736;
wire n_7073;
wire n_9755;
wire n_11287;
wire n_5110;
wire n_9774;
wire n_8397;
wire n_6390;
wire n_4879;
wire n_10139;
wire n_13246;
wire n_13409;
wire n_14061;
wire n_5796;
wire n_10104;
wire n_8726;
wire n_12986;
wire n_11381;
wire n_6665;
wire n_16378;
wire n_16109;
wire n_8797;
wire n_10723;
wire n_7224;
wire n_12441;
wire n_15789;
wire n_9117;
wire n_16172;
wire n_9720;
wire n_16611;
wire n_7746;
wire n_9381;
wire n_10169;
wire n_6958;
wire n_15727;
wire n_16277;
wire n_12049;
wire n_12690;
wire n_14498;
wire n_15417;
wire n_7563;
wire n_12475;
wire n_4556;
wire n_12516;
wire n_11765;
wire n_6549;
wire n_8414;
wire n_13921;
wire n_6297;
wire n_16615;
wire n_14667;
wire n_6523;
wire n_6653;
wire n_8434;
wire n_13405;
wire n_12302;
wire n_10477;
wire n_6096;
wire n_14713;
wire n_15512;
wire n_7853;
wire n_12526;
wire n_4687;
wire n_14414;
wire n_15565;
wire n_7531;
wire n_12377;
wire n_8890;
wire n_5492;
wire n_5995;
wire n_9965;
wire n_13214;
wire n_8615;
wire n_15975;
wire n_11062;
wire n_16575;
wire n_13650;
wire n_7721;
wire n_7192;
wire n_14202;
wire n_15636;
wire n_15859;
wire n_5905;
wire n_11933;
wire n_11206;
wire n_14554;
wire n_9887;
wire n_9149;
wire n_15946;
wire n_4600;
wire n_11593;
wire n_7035;
wire n_6193;
wire n_6501;
wire n_15807;
wire n_13211;
wire n_8316;
wire n_9990;
wire n_5829;
wire n_10005;
wire n_11786;
wire n_12737;
wire n_8057;
wire n_12905;
wire n_11426;
wire n_4954;
wire n_5191;
wire n_14874;
wire n_15311;
wire n_8505;
wire n_15113;
wire n_9273;
wire n_7884;
wire n_9345;
wire n_11258;
wire n_11550;
wire n_15498;
wire n_8970;
wire n_7527;
wire n_7417;
wire n_13061;
wire n_9682;
wire n_4881;
wire n_12513;
wire n_10640;
wire n_6582;
wire n_5734;
wire n_15098;
wire n_13395;
wire n_12545;
wire n_10729;
wire n_14656;
wire n_7388;
wire n_16052;
wire n_11657;
wire n_9924;
wire n_14745;
wire n_8717;
wire n_14744;
wire n_13336;
wire n_5770;
wire n_5705;
wire n_16074;
wire n_4605;
wire n_15091;
wire n_9064;
wire n_7635;
wire n_5525;
wire n_13102;
wire n_11268;
wire n_12753;
wire n_14760;
wire n_4691;
wire n_7090;
wire n_9254;
wire n_12894;
wire n_14135;
wire n_8571;
wire n_11641;
wire n_11501;
wire n_7227;
wire n_10492;
wire n_16482;
wire n_7415;
wire n_11211;
wire n_13375;
wire n_13390;
wire n_13691;
wire n_15769;
wire n_6745;
wire n_6972;
wire n_12514;
wire n_10048;
wire n_8030;
wire n_9247;
wire n_6052;
wire n_8378;
wire n_8687;
wire n_13264;
wire n_5374;
wire n_14194;
wire n_10526;
wire n_5575;
wire n_8725;
wire n_12010;
wire n_9570;
wire n_5675;
wire n_9738;
wire n_12026;
wire n_16663;
wire n_12356;
wire n_11857;
wire n_13825;
wire n_11077;
wire n_6240;
wire n_8243;
wire n_6347;
wire n_8633;
wire n_5020;
wire n_9593;
wire n_7689;
wire n_9846;
wire n_13262;
wire n_13482;
wire n_6511;
wire n_5297;
wire n_15778;
wire n_7121;
wire n_9469;
wire n_10764;
wire n_15869;
wire n_13398;
wire n_9677;
wire n_15598;
wire n_4415;
wire n_15988;
wire n_16593;
wire n_6515;
wire n_7099;
wire n_6804;
wire n_14676;
wire n_8449;
wire n_6358;
wire n_13204;
wire n_14331;
wire n_6603;
wire n_4765;
wire n_16604;
wire n_13873;
wire n_15805;
wire n_4364;
wire n_7534;
wire n_9406;
wire n_11313;
wire n_8201;
wire n_8967;
wire n_4354;
wire n_6986;
wire n_4732;
wire n_8801;
wire n_9322;
wire n_10438;
wire n_15017;
wire n_5959;
wire n_11201;
wire n_16485;
wire n_10531;
wire n_14964;
wire n_8031;
wire n_8918;
wire n_12878;
wire n_15591;
wire n_9348;
wire n_14262;
wire n_16438;
wire n_12188;
wire n_8219;
wire n_15373;
wire n_16609;
wire n_8696;
wire n_4745;
wire n_6396;
wire n_8932;
wire n_5642;
wire n_9232;
wire n_10575;
wire n_15167;
wire n_12630;
wire n_4581;
wire n_6890;
wire n_11028;
wire n_12171;
wire n_4377;
wire n_12299;
wire n_16603;
wire n_15706;
wire n_12022;
wire n_9249;
wire n_14193;
wire n_12935;
wire n_7827;
wire n_14906;
wire n_8180;
wire n_10741;
wire n_15211;
wire n_6109;
wire n_14727;
wire n_10760;
wire n_4792;
wire n_15580;
wire n_12425;
wire n_14762;
wire n_9444;
wire n_15334;
wire n_7731;
wire n_10772;
wire n_11527;
wire n_7114;
wire n_4878;
wire n_13507;
wire n_16486;
wire n_11327;
wire n_10915;
wire n_4979;
wire n_9535;
wire n_15984;
wire n_6770;
wire n_7943;
wire n_11743;
wire n_8892;
wire n_15900;
wire n_12199;
wire n_5302;
wire n_12000;
wire n_15410;
wire n_4511;
wire n_9707;
wire n_12490;
wire n_15151;
wire n_16002;
wire n_16626;
wire n_16258;
wire n_13594;
wire n_5639;
wire n_5781;
wire n_14182;
wire n_8943;
wire n_8486;
wire n_14767;
wire n_10279;
wire n_15853;
wire n_4520;
wire n_5299;
wire n_12829;
wire n_4503;
wire n_14352;
wire n_13889;
wire n_14773;
wire n_10680;
wire n_10127;
wire n_5543;
wire n_13654;
wire n_5361;
wire n_11814;
wire n_7132;
wire n_7081;
wire n_11610;
wire n_12255;
wire n_12739;
wire n_13015;
wire n_5885;
wire n_6663;
wire n_14228;
wire n_9723;
wire n_5356;
wire n_12609;
wire n_4441;
wire n_7319;
wire n_15831;
wire n_5458;
wire n_7644;
wire n_11176;
wire n_16131;
wire n_11473;
wire n_9883;
wire n_11135;
wire n_8155;
wire n_11360;
wire n_5668;
wire n_11275;
wire n_11868;
wire n_5038;
wire n_5330;
wire n_4585;
wire n_7199;
wire n_10039;
wire n_11726;
wire n_11358;
wire n_10854;
wire n_5463;
wire n_15944;
wire n_13366;
wire n_8098;
wire n_12574;
wire n_12700;
wire n_12904;
wire n_8833;
wire n_9191;
wire n_5489;
wire n_5892;
wire n_7828;
wire n_10142;
wire n_4773;
wire n_14623;
wire n_7940;
wire n_9918;
wire n_15932;
wire n_7910;
wire n_5654;
wire n_6782;
wire n_16467;
wire n_6009;
wire n_9034;
wire n_16345;
wire n_6503;
wire n_6376;
wire n_4427;
wire n_7084;
wire n_5923;
wire n_14073;
wire n_9390;
wire n_5113;
wire n_12017;
wire n_12888;
wire n_10069;
wire n_5479;
wire n_5714;
wire n_8541;
wire n_8074;
wire n_15381;
wire n_8485;
wire n_13639;
wire n_14852;
wire n_8860;
wire n_15989;
wire n_5510;
wire n_11958;
wire n_6621;
wire n_15624;
wire n_7001;
wire n_9650;
wire n_4822;
wire n_13070;
wire n_8271;
wire n_15514;
wire n_5692;
wire n_16460;
wire n_8473;
wire n_13640;
wire n_14147;
wire n_4800;
wire n_9266;
wire n_14491;
wire n_12728;
wire n_5555;
wire n_15011;
wire n_10027;
wire n_16210;
wire n_12784;
wire n_16651;
wire n_4958;
wire n_5441;
wire n_6783;
wire n_9664;
wire n_13678;
wire n_12458;
wire n_12259;
wire n_6066;
wire n_12877;
wire n_14582;
wire n_8699;
wire n_16305;
wire n_14261;
wire n_14677;
wire n_6897;
wire n_13523;
wire n_10616;
wire n_8587;
wire n_9619;
wire n_11171;
wire n_15117;
wire n_5366;
wire n_14928;
wire n_15550;
wire n_16016;
wire n_15528;
wire n_6925;
wire n_6878;
wire n_15861;
wire n_8225;
wire n_9078;
wire n_9536;
wire n_16297;
wire n_13778;
wire n_14250;
wire n_16171;
wire n_16573;
wire n_4886;
wire n_9931;
wire n_13198;
wire n_16419;
wire n_16470;
wire n_16562;
wire n_15914;
wire n_6296;
wire n_9187;
wire n_7708;
wire n_13741;
wire n_13819;
wire n_16621;
wire n_15777;
wire n_12610;
wire n_14634;
wire n_11671;
wire n_10328;
wire n_14416;
wire n_5968;
wire n_11251;
wire n_14424;
wire n_14523;
wire n_12293;
wire n_11063;
wire n_10753;
wire n_6497;
wire n_8319;
wire n_9989;
wire n_13174;
wire n_15705;
wire n_7108;
wire n_14455;
wire n_12853;
wire n_6470;
wire n_12942;
wire n_11598;
wire n_8368;
wire n_15691;
wire n_9259;
wire n_8322;
wire n_7333;
wire n_11879;
wire n_16127;
wire n_6187;
wire n_7876;
wire n_12397;
wire n_15376;
wire n_16555;
wire n_8546;
wire n_10963;
wire n_16358;
wire n_8300;
wire n_15336;
wire n_7371;
wire n_9378;
wire n_8152;
wire n_15050;
wire n_10826;
wire n_7463;
wire n_12206;
wire n_8525;
wire n_14161;
wire n_6573;
wire n_9656;
wire n_7634;
wire n_5078;
wire n_8148;
wire n_11400;
wire n_13290;
wire n_8150;
wire n_13500;
wire n_11440;
wire n_12596;
wire n_6693;
wire n_15848;
wire n_15398;
wire n_10483;
wire n_15593;
wire n_12160;
wire n_4737;
wire n_11563;
wire n_4925;
wire n_9620;
wire n_16424;
wire n_5415;
wire n_13945;
wire n_8986;
wire n_7285;
wire n_11337;
wire n_12444;
wire n_12005;
wire n_16409;
wire n_5419;
wire n_11243;
wire n_8929;
wire n_9360;
wire n_12697;
wire n_14513;
wire n_7260;
wire n_5205;
wire n_12778;
wire n_12485;
wire n_6409;
wire n_11939;
wire n_7954;
wire n_11119;
wire n_9824;
wire n_14347;
wire n_15089;
wire n_7951;
wire n_7552;
wire n_8096;
wire n_14602;
wire n_11468;
wire n_15995;
wire n_16150;
wire n_13901;
wire n_12166;
wire n_8233;
wire n_6130;
wire n_4603;
wire n_7273;
wire n_9683;
wire n_10646;
wire n_14750;
wire n_7231;
wire n_15725;
wire n_5080;
wire n_5976;
wire n_11704;
wire n_14074;
wire n_15252;
wire n_15132;
wire n_5732;
wire n_5372;
wire n_16238;
wire n_14050;
wire n_11878;
wire n_15843;
wire n_15763;
wire n_16666;
wire n_4471;
wire n_15749;
wire n_15317;
wire n_7449;
wire n_7772;
wire n_8763;
wire n_12800;
wire n_5208;
wire n_14197;
wire n_8679;
wire n_15638;
wire n_16547;
wire n_7239;
wire n_14289;
wire n_15582;
wire n_16415;
wire n_9848;
wire n_14447;
wire n_16479;
wire n_16574;
wire n_11962;
wire n_15145;
wire n_5690;
wire n_9227;
wire n_8187;
wire n_10751;
wire n_7050;
wire n_10240;
wire n_9399;
wire n_8996;
wire n_10691;
wire n_15838;
wire n_15297;
wire n_6623;
wire n_9561;
wire n_13951;
wire n_13968;
wire n_10378;
wire n_13979;
wire n_12070;
wire n_16104;
wire n_9714;
wire n_9740;
wire n_9773;
wire n_13316;
wire n_14898;
wire n_10313;
wire n_15672;
wire n_12947;
wire n_5371;
wire n_4651;
wire n_9745;
wire n_13689;
wire n_15413;
wire n_10216;
wire n_15628;
wire n_15920;
wire n_11928;
wire n_8139;
wire n_9764;
wire n_4854;
wire n_5071;
wire n_15160;
wire n_7597;
wire n_5801;
wire n_10150;
wire n_12354;
wire n_12666;
wire n_14297;
wire n_14395;
wire n_13528;
wire n_6047;
wire n_12581;
wire n_8292;
wire n_16368;
wire n_12631;
wire n_14969;
wire n_14820;
wire n_10133;
wire n_8601;
wire n_10773;
wire n_6652;
wire n_4994;
wire n_9377;
wire n_11932;
wire n_10971;
wire n_8830;
wire n_4483;
wire n_6921;
wire n_6970;
wire n_5347;
wire n_5168;
wire n_14836;
wire n_4661;
wire n_13027;
wire n_12867;
wire n_4988;
wire n_7674;
wire n_14675;
wire n_9826;
wire n_12607;
wire n_14516;
wire n_15960;
wire n_7568;
wire n_15343;
wire n_6354;
wire n_7272;
wire n_15782;
wire n_12075;
wire n_4540;
wire n_11942;
wire n_15998;
wire n_6344;
wire n_12305;
wire n_13489;
wire n_12123;
wire n_9772;
wire n_12170;
wire n_15370;
wire n_6021;
wire n_7949;
wire n_7724;
wire n_6624;
wire n_9630;
wire n_6956;
wire n_13313;
wire n_13927;
wire n_12966;
wire n_13877;
wire n_15851;
wire n_15308;
wire n_6305;
wire n_9255;
wire n_6209;
wire n_8310;
wire n_10231;
wire n_12547;
wire n_9758;
wire n_16148;
wire n_15577;
wire n_16500;
wire n_16550;
wire n_15884;
wire n_11922;
wire n_4971;
wire n_14020;
wire n_15175;
wire n_8936;
wire n_5656;
wire n_7126;
wire n_5125;
wire n_5857;
wire n_12358;
wire n_7329;
wire n_14502;
wire n_15206;
wire n_8646;
wire n_7408;
wire n_13415;
wire n_9691;
wire n_12997;
wire n_14533;
wire n_10259;
wire n_14005;
wire n_7107;
wire n_14293;
wire n_5652;
wire n_6457;
wire n_8597;
wire n_10488;
wire n_14334;
wire n_7690;
wire n_8969;
wire n_14187;
wire n_15245;
wire n_7123;
wire n_10752;
wire n_11577;
wire n_15225;
wire n_5499;
wire n_8117;
wire n_10067;
wire n_15169;
wire n_10399;
wire n_11223;
wire n_10213;
wire n_13562;
wire n_14537;
wire n_12498;
wire n_13888;
wire n_16592;
wire n_11475;
wire n_6950;
wire n_8208;
wire n_10038;
wire n_9048;
wire n_5228;
wire n_11010;
wire n_10274;
wire n_15614;
wire n_9590;
wire n_16017;
wire n_11588;
wire n_16346;
wire n_6694;
wire n_13956;
wire n_15318;
wire n_6880;
wire n_5066;
wire n_7418;
wire n_9168;
wire n_14220;
wire n_11221;
wire n_13837;
wire n_12387;
wire n_9497;
wire n_15772;
wire n_8536;
wire n_13255;
wire n_15911;
wire n_9435;
wire n_7229;
wire n_14245;
wire n_8350;
wire n_16475;
wire n_11448;
wire n_9219;
wire n_5507;
wire n_5569;
wire n_8028;
wire n_8328;
wire n_15502;
wire n_8914;
wire n_15076;
wire n_12576;
wire n_15559;
wire n_7258;
wire n_15276;
wire n_5190;
wire n_13892;
wire n_8391;
wire n_16361;
wire n_14221;
wire n_16343;
wire n_10579;
wire n_10832;
wire n_13345;
wire n_13964;
wire n_13749;
wire n_8336;
wire n_6856;
wire n_6466;
wire n_14559;
wire n_16039;
wire n_7864;
wire n_15552;
wire n_16228;
wire n_6727;
wire n_14360;
wire n_10584;
wire n_5392;
wire n_12862;
wire n_11445;
wire n_13151;
wire n_13621;
wire n_13601;
wire n_14052;
wire n_14311;
wire n_8216;
wire n_11552;
wire n_13765;
wire n_10332;
wire n_7709;
wire n_15290;
wire n_15102;
wire n_14733;
wire n_11874;
wire n_13926;
wire n_9982;
wire n_10171;
wire n_15184;
wire n_14157;
wire n_5455;
wire n_5442;
wire n_6386;
wire n_14317;
wire n_12803;
wire n_5948;
wire n_7804;
wire n_4459;
wire n_4545;
wire n_12656;
wire n_16220;
wire n_9852;
wire n_6820;
wire n_11623;
wire n_8313;
wire n_14828;
wire n_7656;
wire n_5511;
wire n_6208;
wire n_5295;
wire n_6739;
wire n_15779;
wire n_14131;
wire n_8041;
wire n_10676;
wire n_8202;
wire n_8263;
wire n_10299;
wire n_6438;
wire n_5490;
wire n_10540;
wire n_11936;
wire n_15366;
wire n_12845;
wire n_10374;
wire n_11645;
wire n_4771;
wire n_10200;
wire n_13392;
wire n_7332;
wire n_12734;
wire n_10382;
wire n_13164;
wire n_5836;
wire n_7185;
wire n_6291;
wire n_11489;
wire n_13662;
wire n_10269;
wire n_4455;
wire n_8374;
wire n_12262;
wire n_13223;
wire n_16275;
wire n_13340;
wire n_9169;
wire n_14910;
wire n_13451;
wire n_4514;
wire n_13939;
wire n_5834;
wire n_10229;
wire n_5584;
wire n_13728;
wire n_7512;
wire n_14385;
wire n_4806;
wire n_7386;
wire n_9939;
wire n_7766;
wire n_10981;
wire n_8738;
wire n_11018;
wire n_14499;
wire n_9126;
wire n_6469;
wire n_6700;
wire n_15368;
wire n_16014;
wire n_12797;
wire n_6223;
wire n_11376;
wire n_6758;
wire n_9438;
wire n_11398;
wire n_5160;
wire n_7808;
wire n_6544;
wire n_8798;
wire n_9481;
wire n_13379;
wire n_9600;
wire n_13781;
wire n_9122;
wire n_14731;
wire n_8085;
wire n_11274;
wire n_5098;
wire n_8123;
wire n_10344;
wire n_7955;
wire n_5707;
wire n_12012;
wire n_5140;
wire n_4992;
wire n_12512;
wire n_5197;
wire n_7287;
wire n_16337;
wire n_9927;
wire n_14613;
wire n_5497;
wire n_10076;
wire n_11515;
wire n_8721;
wire n_12820;
wire n_6464;
wire n_9912;
wire n_6356;
wire n_13558;
wire n_11554;
wire n_15657;
wire n_15881;
wire n_7637;
wire n_10148;
wire n_16577;
wire n_10318;
wire n_4796;
wire n_4442;
wire n_7127;
wire n_4533;
wire n_9635;
wire n_13890;
wire n_5481;
wire n_12890;
wire n_8666;
wire n_15513;
wire n_5344;
wire n_9264;
wire n_13994;
wire n_14483;
wire n_4419;
wire n_8326;
wire n_8670;
wire n_5308;
wire n_5184;
wire n_5794;
wire n_15179;
wire n_7638;
wire n_11972;
wire n_12284;
wire n_15724;
wire n_14308;
wire n_7801;
wire n_5408;
wire n_13484;
wire n_9155;
wire n_10234;
wire n_8460;
wire n_10416;
wire n_15837;
wire n_14370;
wire n_14593;
wire n_8836;
wire n_7959;
wire n_13430;
wire n_7019;
wire n_8181;
wire n_11325;
wire n_14838;
wire n_15207;
wire n_8254;
wire n_13452;
wire n_13521;
wire n_8071;
wire n_14525;
wire n_7735;
wire n_8004;
wire n_16013;
wire n_6667;
wire n_14926;
wire n_7409;
wire n_5271;
wire n_10731;
wire n_10735;
wire n_10583;
wire n_9878;
wire n_5964;
wire n_6004;
wire n_10806;
wire n_13807;
wire n_14591;
wire n_14363;
wire n_9825;
wire n_5494;
wire n_7444;
wire n_11628;
wire n_14576;
wire n_7546;
wire n_4431;
wire n_5234;
wire n_6272;
wire n_4387;
wire n_14274;
wire n_6588;
wire n_11549;
wire n_5128;
wire n_14033;
wire n_12286;
wire n_9001;
wire n_10393;
wire n_15403;
wire n_11498;
wire n_13081;
wire n_15221;
wire n_16107;
wire n_15602;
wire n_10513;
wire n_12252;
wire n_5467;
wire n_10439;
wire n_7296;
wire n_8013;
wire n_14545;
wire n_12627;
wire n_16090;
wire n_4890;
wire n_7575;
wire n_9045;
wire n_7083;
wire n_12281;
wire n_15637;
wire n_14272;
wire n_11237;
wire n_7720;
wire n_6222;
wire n_11643;
wire n_9373;
wire n_15012;
wire n_14337;
wire n_6268;
wire n_16683;
wire n_5827;
wire n_5199;
wire n_12347;
wire n_14551;
wire n_6456;
wire n_11103;
wire n_11809;
wire n_15720;
wire n_11181;
wire n_13651;
wire n_9967;
wire n_13553;
wire n_7521;
wire n_14088;
wire n_5992;
wire n_12968;
wire n_5313;
wire n_10663;
wire n_13817;
wire n_9971;
wire n_7187;
wire n_15517;
wire n_10894;
wire n_14118;
wire n_13974;
wire n_9524;
wire n_12277;
wire n_14917;
wire n_12698;
wire n_5312;
wire n_6467;
wire n_9182;
wire n_9243;
wire n_9282;
wire n_16075;
wire n_5079;
wire n_9365;
wire n_6540;
wire n_6625;
wire n_10909;
wire n_15680;
wire n_6336;
wire n_10083;
wire n_6796;
wire n_9224;
wire n_10347;
wire n_16086;
wire n_5513;
wire n_5614;
wire n_12417;
wire n_11871;
wire n_6541;
wire n_12410;
wire n_4830;
wire n_4706;
wire n_13225;
wire n_14855;
wire n_16327;
wire n_5225;
wire n_4570;
wire n_14707;
wire n_15326;
wire n_16043;
wire n_10208;
wire n_7722;
wire n_8487;
wire n_9240;
wire n_10804;
wire n_8293;
wire n_6486;
wire n_4622;
wire n_14726;
wire n_8141;
wire n_14612;
wire n_12294;
wire n_14180;
wire n_7603;
wire n_10667;
wire n_4887;
wire n_14058;
wire n_8438;
wire n_10548;
wire n_11020;
wire n_13355;
wire n_12957;
wire n_4693;
wire n_13141;
wire n_11616;
wire n_16461;
wire n_14065;
wire n_8791;
wire n_11920;
wire n_10793;
wire n_8288;
wire n_14672;
wire n_14366;
wire n_15127;
wire n_5835;
wire n_10481;
wire n_6732;
wire n_7979;
wire n_6876;
wire n_12786;
wire n_16022;
wire n_5049;
wire n_13382;
wire n_12711;
wire n_11675;
wire n_12219;
wire n_10678;
wire n_6757;
wire n_9573;
wire n_15543;
wire n_5846;
wire n_8323;
wire n_8657;
wire n_8006;
wire n_8296;
wire n_10391;
wire n_7636;
wire n_9695;
wire n_9799;
wire n_11306;
wire n_5592;
wire n_6954;
wire n_6938;
wire n_7866;
wire n_4609;
wire n_11083;
wire n_13176;
wire n_15143;
wire n_9784;
wire n_11198;
wire n_7205;
wire n_8757;
wire n_7990;
wire n_7020;
wire n_13035;
wire n_10036;
wire n_13021;
wire n_5278;
wire n_11728;
wire n_12893;
wire n_14905;
wire n_8596;
wire n_15128;
wire n_5157;
wire n_11840;
wire n_4754;
wire n_11698;
wire n_4647;
wire n_9556;
wire n_11292;
wire n_13157;
wire n_8590;
wire n_8720;
wire n_10261;
wire n_16682;
wire n_5708;
wire n_13502;
wire n_5223;
wire n_6298;
wire n_12205;
wire n_11989;
wire n_4894;
wire n_5474;
wire n_14084;
wire n_15798;
wire n_12289;
wire n_10813;
wire n_10757;
wire n_4760;
wire n_5649;
wire n_11326;
wire n_13046;
wire n_6421;
wire n_13935;
wire n_11870;
wire n_16215;
wire n_7407;
wire n_9827;
wire n_14009;
wire n_16670;
wire n_13334;
wire n_10907;
wire n_5704;
wire n_15787;
wire n_11431;
wire n_4983;
wire n_7148;
wire n_14002;
wire n_6328;
wire n_5956;
wire n_11283;
wire n_5287;
wire n_13646;
wire n_6236;
wire n_9417;
wire n_11834;
wire n_13361;
wire n_12020;
wire n_5083;
wire n_7214;
wire n_4509;
wire n_15061;
wire n_6007;
wire n_6144;
wire n_11506;
wire n_16205;
wire n_10135;
wire n_13161;
wire n_6197;
wire n_6658;
wire n_6835;
wire n_4906;
wire n_8834;
wire n_11624;
wire n_13399;
wire n_14010;
wire n_8826;
wire n_15083;
wire n_11352;
wire n_15262;
wire n_16429;
wire n_16413;
wire n_5516;
wire n_6247;
wire n_7075;
wire n_4897;
wire n_11234;
wire n_10822;
wire n_14697;
wire n_15030;
wire n_10919;
wire n_7104;
wire n_9152;
wire n_7124;
wire n_13967;
wire n_12099;
wire n_12858;
wire n_7467;
wire n_4399;
wire n_14609;
wire n_16451;
wire n_15351;
wire n_7799;
wire n_8364;
wire n_5698;
wire n_11092;
wire n_9534;
wire n_14310;
wire n_15228;
wire n_13380;
wire n_5084;
wire n_5771;
wire n_7544;
wire n_15832;
wire n_13053;
wire n_9792;
wire n_7513;
wire n_10720;
wire n_9336;
wire n_10535;
wire n_11836;
wire n_6602;
wire n_10924;
wire n_15281;
wire n_15792;
wire n_6708;
wire n_8854;
wire n_11186;
wire n_8917;
wire n_15675;
wire n_9647;
wire n_15515;
wire n_6645;
wire n_9742;
wire n_11236;
wire n_10727;
wire n_16177;
wire n_10885;
wire n_15106;
wire n_6484;
wire n_4710;
wire n_4420;
wire n_13201;
wire n_6242;
wire n_12527;
wire n_4574;
wire n_14759;
wire n_13274;
wire n_12379;
wire n_9312;
wire n_9019;
wire n_13891;
wire n_8985;
wire n_7692;
wire n_12067;
wire n_9214;
wire n_12932;
wire n_5174;
wire n_12477;
wire n_14325;
wire n_7469;
wire n_5538;
wire n_15503;
wire n_14078;
wire n_7776;
wire n_5017;
wire n_10418;
wire n_14309;
wire n_10895;
wire n_10875;
wire n_11977;
wire n_11736;
wire n_7560;
wire n_16270;
wire n_14729;
wire n_9864;
wire n_8548;
wire n_10672;
wire n_7645;
wire n_11846;
wire n_15576;
wire n_16256;
wire n_14222;
wire n_11696;
wire n_12400;
wire n_5096;
wire n_11734;
wire n_12114;
wire n_4660;
wire n_9533;
wire n_9494;
wire n_5241;
wire n_11770;
wire n_10308;
wire n_11608;
wire n_11507;
wire n_14430;
wire n_9145;
wire n_15337;
wire n_13996;
wire n_7082;
wire n_12092;
wire n_14749;
wire n_12295;
wire n_10623;
wire n_9754;
wire n_4797;
wire n_6285;
wire n_9315;
wire n_11320;
wire n_11837;
wire n_5428;
wire n_16545;
wire n_13709;
wire n_7451;
wire n_4945;
wire n_8260;
wire n_13898;
wire n_9000;
wire n_16507;
wire n_5677;
wire n_9454;
wire n_6734;
wire n_7476;
wire n_10864;
wire n_10586;
wire n_16543;
wire n_5570;
wire n_11938;
wire n_6418;
wire n_8742;
wire n_12626;
wire n_14704;
wire n_8307;
wire n_5153;
wire n_11967;
wire n_9383;
wire n_9253;
wire n_15084;
wire n_13559;
wire n_10571;
wire n_4611;
wire n_8874;
wire n_15258;
wire n_5927;
wire n_15071;
wire n_7392;
wire n_7495;
wire n_9566;
wire n_11338;
wire n_11996;
wire n_5435;
wire n_13426;
wire n_12174;
wire n_9765;
wire n_16322;
wire n_9807;
wire n_4333;
wire n_9057;
wire n_5200;
wire n_8706;
wire n_15220;
wire n_6400;
wire n_7666;
wire n_7945;
wire n_8894;
wire n_16304;
wire n_6941;
wire n_5115;
wire n_12053;
wire n_15947;
wire n_5566;
wire n_12619;
wire n_11250;
wire n_7829;
wire n_7543;
wire n_13504;
wire n_15328;
wire n_8680;
wire n_11289;
wire n_13169;
wire n_7877;
wire n_7963;
wire n_13555;
wire n_9672;
wire n_12582;
wire n_16522;
wire n_5487;
wire n_15291;
wire n_8855;
wire n_6398;
wire n_8885;
wire n_10394;
wire n_8329;
wire n_5486;
wire n_9503;
wire n_15345;
wire n_12423;
wire n_11391;
wire n_15426;
wire n_15462;
wire n_5244;
wire n_5092;
wire n_14721;
wire n_14137;
wire n_13265;
wire n_8270;
wire n_4832;
wire n_12714;
wire n_16051;
wire n_12153;
wire n_5889;
wire n_11738;
wire n_7284;
wire n_7264;
wire n_5391;
wire n_11522;
wire n_9763;
wire n_14163;
wire n_7737;
wire n_13666;
wire n_15523;
wire n_6537;
wire n_16569;
wire n_8614;
wire n_11070;
wire n_7328;
wire n_10702;
wire n_13337;
wire n_10958;
wire n_15682;
wire n_15112;
wire n_9479;
wire n_15556;
wire n_9162;
wire n_9568;
wire n_13730;
wire n_14849;
wire n_15621;
wire n_12405;
wire n_8816;
wire n_14041;
wire n_9119;
wire n_10319;
wire n_5849;
wire n_16661;
wire n_9654;
wire n_9181;
wire n_11648;
wire n_4554;
wire n_10322;
wire n_7135;
wire n_13529;
wire n_6224;
wire n_6578;
wire n_8802;
wire n_9859;
wire n_14763;
wire n_8555;
wire n_5240;
wire n_10695;
wire n_8636;
wire n_7024;
wire n_6092;
wire n_15912;
wire n_10879;
wire n_16206;
wire n_5951;
wire n_6241;
wire n_6589;
wire n_8508;
wire n_6614;
wire n_5912;
wire n_8667;
wire n_10639;
wire n_16359;
wire n_16037;
wire n_16529;
wire n_8121;
wire n_8207;
wire n_9645;
wire n_9276;
wire n_8035;
wire n_12554;
wire n_13351;
wire n_11653;
wire n_12722;
wire n_6735;
wire n_7754;
wire n_4680;
wire n_15549;
wire n_10491;
wire n_12037;
wire n_15371;
wire n_13453;
wire n_5152;
wire n_15080;
wire n_5265;
wire n_12792;
wire n_15937;
wire n_11717;
wire n_9943;
wire n_16141;
wire n_4927;
wire n_5574;
wire n_12391;
wire n_14242;
wire n_15622;
wire n_9821;
wire n_11112;
wire n_7152;
wire n_11723;
wire n_15246;
wire n_9575;
wire n_16647;
wire n_14940;
wire n_6165;
wire n_8320;
wire n_9796;
wire n_10409;
wire n_4548;
wire n_11822;
wire n_4862;
wire n_10521;
wire n_9610;
wire n_15889;
wire n_11830;
wire n_12438;
wire n_15395;
wire n_5469;
wire n_14393;
wire n_8766;
wire n_12364;
wire n_12420;
wire n_12838;
wire n_6567;
wire n_9165;
wire n_16173;
wire n_16483;
wire n_13505;
wire n_14016;
wire n_12323;
wire n_5910;
wire n_15566;
wire n_5895;
wire n_5804;
wire n_9508;
wire n_12539;
wire n_12776;
wire n_10527;
wire n_5965;
wire n_9596;
wire n_13652;
wire n_13703;
wire n_16231;
wire n_14369;
wire n_7240;
wire n_7570;
wire n_4553;
wire n_7033;
wire n_15354;
wire n_10476;
wire n_4875;
wire n_9966;
wire n_13156;
wire n_7817;
wire n_5682;
wire n_15529;
wire n_10710;
wire n_5387;
wire n_5557;
wire n_11394;
wire n_8850;
wire n_11906;
wire n_9928;
wire n_11820;
wire n_14647;
wire n_14298;
wire n_8002;
wire n_9741;
wire n_13897;
wire n_11486;
wire n_14792;
wire n_15280;
wire n_15999;
wire n_12677;
wire n_16290;
wire n_10180;
wire n_14248;
wire n_14112;
wire n_8370;
wire n_7237;
wire n_13300;
wire n_16296;
wire n_5681;
wire n_10650;
wire n_12120;
wire n_9090;
wire n_16412;
wire n_16456;
wire n_12021;
wire n_10157;
wire n_6877;
wire n_7423;
wire n_12873;
wire n_12008;
wire n_10402;
wire n_12515;
wire n_16364;
wire n_6949;
wire n_7566;
wire n_6119;
wire n_11940;
wire n_4901;
wire n_4821;
wire n_9217;
wire n_9261;
wire n_9166;
wire n_12901;
wire n_10518;
wire n_8301;
wire n_12895;
wire n_7617;
wire n_12223;
wire n_12045;
wire n_15170;
wire n_9771;
wire n_13401;
wire n_15774;
wire n_7718;
wire n_5316;
wire n_6940;
wire n_9893;
wire n_12276;
wire n_13844;
wire n_14122;
wire n_7396;
wire n_10942;
wire n_12726;
wire n_12668;
wire n_5703;
wire n_7835;
wire n_11430;
wire n_15437;
wire n_13010;
wire n_6320;
wire n_8126;
wire n_11239;
wire n_15819;
wire n_7998;
wire n_10362;
wire n_9239;
wire n_12432;
wire n_4943;
wire n_10953;
wire n_4757;
wire n_7561;
wire n_15603;
wire n_6810;
wire n_7842;
wire n_12352;
wire n_6202;
wire n_9969;
wire n_10099;
wire n_11437;
wire n_12898;
wire n_4682;
wire n_9961;
wire n_14068;
wire n_16130;
wire n_12879;
wire n_14853;
wire n_5564;
wire n_11869;
wire n_13746;
wire n_14895;
wire n_12559;
wire n_13508;
wire n_5620;
wire n_14660;
wire n_15540;
wire n_7163;
wire n_4530;
wire n_16582;
wire n_10343;
wire n_10836;
wire n_4942;
wire n_15270;
wire n_9899;
wire n_9258;
wire n_16375;
wire n_13004;
wire n_10181;
wire n_15670;
wire n_10286;
wire n_5406;
wire n_8072;
wire n_10371;
wire n_13479;
wire n_14990;
wire n_8277;
wire n_7236;
wire n_16295;
wire n_4604;
wire n_13117;
wire n_10257;
wire n_7130;
wire n_5724;
wire n_14437;
wire n_7201;
wire n_11219;
wire n_4841;
wire n_10047;
wire n_14541;
wire n_13759;
wire n_16186;
wire n_5806;
wire n_10949;
wire n_4338;
wire n_13766;
wire n_10486;
wire n_11226;
wire n_11282;
wire n_8724;
wire n_16613;
wire n_5738;
wire n_15938;
wire n_11413;
wire n_14700;
wire n_15146;
wire n_4840;
wire n_4519;
wire n_5355;
wire n_16617;
wire n_5320;
wire n_16382;
wire n_7491;
wire n_13969;
wire n_5353;
wire n_9995;
wire n_13710;
wire n_16548;
wire n_5710;
wire n_5186;
wire n_9076;
wire n_11232;
wire n_12351;
wire n_12693;
wire n_9105;
wire n_6792;
wire n_16360;
wire n_12080;
wire n_16261;
wire n_5093;
wire n_9316;
wire n_5979;
wire n_9636;
wire n_13359;
wire n_9668;
wire n_10372;
wire n_14867;
wire n_7559;
wire n_6044;
wire n_5438;
wire n_8867;
wire n_9491;
wire n_13335;
wire n_4326;
wire n_13259;
wire n_14022;
wire n_12702;
wire n_15188;
wire n_13175;
wire n_5517;
wire n_11276;
wire n_5605;
wire n_12439;
wire n_14954;
wire n_10744;
wire n_12648;
wire n_11008;
wire n_9870;
wire n_9833;
wire n_6125;
wire n_7314;
wire n_9095;
wire n_4726;
wire n_7678;
wire n_5907;
wire n_11334;
wire n_15757;
wire n_15979;
wire n_6045;
wire n_13075;
wire n_13129;
wire n_13736;
wire n_9914;
wire n_8132;
wire n_6731;
wire n_9178;
wire n_14186;
wire n_7526;
wire n_5040;
wire n_14023;
wire n_6063;
wire n_16118;
wire n_10736;
wire n_10917;
wire n_16050;
wire n_6504;
wire n_11575;
wire n_7004;
wire n_7821;
wire n_14418;
wire n_12407;
wire n_13586;
wire n_8308;
wire n_6154;
wire n_15813;
wire n_11284;
wire n_6943;
wire n_10597;
wire n_14668;
wire n_16281;
wire n_11827;
wire n_13049;
wire n_8165;
wire n_13961;
wire n_14283;
wire n_12038;
wire n_14776;
wire n_4788;
wire n_8400;
wire n_10458;
wire n_15745;
wire n_8210;
wire n_11656;
wire n_12644;
wire n_5977;
wire n_10446;
wire n_13134;
wire n_11826;
wire n_7879;
wire n_10271;
wire n_16372;
wire n_10888;
wire n_15958;
wire n_10116;
wire n_15415;
wire n_14808;
wire n_7696;
wire n_11570;
wire n_16567;
wire n_6003;
wire n_12952;
wire n_6684;
wire n_5746;
wire n_6600;
wire n_11764;
wire n_13063;
wire n_14795;
wire n_5451;
wire n_9323;
wire n_14140;
wire n_5402;
wire n_6673;
wire n_10696;
wire n_7355;
wire n_6961;
wire n_9331;
wire n_10170;
wire n_6031;
wire n_9922;
wire n_13252;
wire n_14479;
wire n_12024;
wire n_8331;
wire n_11909;
wire n_13084;
wire n_16425;
wire n_8217;
wire n_10603;
wire n_6962;
wire n_12004;
wire n_15374;
wire n_16622;
wire n_12830;
wire n_12637;
wire n_8858;
wire n_7887;
wire n_7246;
wire n_4365;
wire n_6060;
wire n_15414;
wire n_15783;
wire n_7929;
wire n_10255;
wire n_16440;
wire n_10572;
wire n_14172;
wire n_16431;
wire n_12009;
wire n_13612;
wire n_7270;
wire n_13985;
wire n_11490;
wire n_8689;
wire n_10648;
wire n_5417;
wire n_6967;
wire n_14124;
wire n_10113;
wire n_7550;
wire n_15077;
wire n_15086;
wire n_12414;
wire n_9760;
wire n_10690;
wire n_6853;
wire n_6742;
wire n_10188;
wire n_13525;
wire n_4923;
wire n_5864;
wire n_10686;
wire n_15733;
wire n_15864;
wire n_9841;
wire n_14997;
wire n_15931;
wire n_13552;
wire n_6691;
wire n_8743;
wire n_7087;
wire n_12681;
wire n_14207;
wire n_8753;
wire n_14799;
wire n_6191;
wire n_4741;
wire n_10689;
wire n_13909;
wire n_6172;
wire n_12634;
wire n_10974;
wire n_13022;
wire n_11067;
wire n_13863;
wire n_8627;
wire n_14305;
wire n_9513;
wire n_16447;
wire n_14774;
wire n_9863;
wire n_12680;
wire n_15330;
wire n_11613;
wire n_4885;
wire n_13659;
wire n_16124;
wire n_10233;
wire n_12034;
wire n_10500;
wire n_16586;
wire n_15446;
wire n_10555;
wire n_5432;
wire n_15261;
wire n_15492;
wire n_10314;
wire n_4550;
wire n_6988;
wire n_4652;
wire n_11929;
wire n_10810;
wire n_11075;
wire n_16056;
wire n_7851;
wire n_6894;
wire n_13303;
wire n_13346;
wire n_12176;
wire n_9791;
wire n_13702;
wire n_16605;
wire n_10311;
wire n_9179;
wire n_15894;
wire n_5453;
wire n_13656;
wire n_9140;
wire n_8752;
wire n_6834;
wire n_4900;
wire n_11177;
wire n_13667;
wire n_4408;
wire n_4577;
wire n_6817;
wire n_4748;
wire n_5842;
wire n_10937;
wire n_13126;
wire n_6927;
wire n_12134;
wire n_12449;
wire n_5814;
wire n_7798;
wire n_5253;
wire n_5209;
wire n_10857;
wire n_15470;
wire n_11310;
wire n_13275;
wire n_12094;
wire n_6215;
wire n_16399;
wire n_11165;
wire n_9736;
wire n_5699;
wire n_5531;
wire n_14411;
wire n_5765;
wire n_12823;
wire n_15412;
wire n_12517;
wire n_6517;
wire n_15754;
wire n_6284;
wire n_5943;
wire n_15441;
wire n_10167;
wire n_7862;
wire n_12193;
wire n_9225;
wire n_12524;
wire n_11923;
wire n_12071;
wire n_13832;
wire n_10630;
wire n_8105;
wire n_6088;
wire n_9031;
wire n_5777;
wire n_6883;
wire n_8808;
wire n_10061;
wire n_15257;
wire n_12963;
wire n_10428;
wire n_13087;
wire n_13972;
wire n_15599;
wire n_11865;
wire n_15436;
wire n_12366;
wire n_15633;
wire n_8528;
wire n_8204;
wire n_13024;
wire n_11733;
wire n_11068;
wire n_11035;
wire n_14951;
wire n_5495;
wire n_10694;
wire n_15646;
wire n_12339;
wire n_10602;
wire n_16630;
wire n_7100;
wire n_12729;
wire n_13292;
wire n_12198;
wire n_11041;
wire n_14632;
wire n_9420;
wire n_14490;
wire n_5655;
wire n_6393;
wire n_15969;
wire n_9708;
wire n_14336;
wire n_5064;
wire n_7825;
wire n_10079;
wire n_12242;
wire n_14738;
wire n_15479;
wire n_7119;
wire n_8154;
wire n_7212;
wire n_5610;
wire n_6966;
wire n_8889;
wire n_13986;
wire n_9790;
wire n_13849;
wire n_13796;
wire n_10502;
wire n_11973;
wire n_11131;
wire n_15522;
wire n_5002;
wire n_5759;
wire n_10778;
wire n_6722;
wire n_13258;
wire n_6035;
wire n_7874;
wire n_13329;
wire n_8490;
wire n_7622;
wire n_9014;
wire n_10329;
wire n_9979;
wire n_13166;
wire n_15435;
wire n_8509;
wire n_8767;
wire n_11123;
wire n_8512;
wire n_13946;
wire n_9505;
wire n_8634;
wire n_9531;
wire n_6364;
wire n_14464;
wire n_15028;
wire n_8635;
wire n_7102;
wire n_7420;
wire n_15482;
wire n_4342;
wire n_12605;
wire n_13618;
wire n_10855;
wire n_7995;
wire n_6114;
wire n_16217;
wire n_4568;
wire n_11003;
wire n_6061;
wire n_10662;
wire n_5559;
wire n_15535;
wire n_16633;
wire n_7831;
wire n_6253;
wire n_12828;
wire n_12723;
wire n_10258;
wire n_5786;
wire n_14960;
wire n_8532;
wire n_14993;
wire n_14327;
wire n_12661;
wire n_10227;
wire n_10588;
wire n_8624;
wire n_8991;
wire n_11022;
wire n_14097;
wire n_10574;
wire n_8065;
wire n_10247;
wire n_11140;
wire n_16323;
wire n_5377;
wire n_6201;
wire n_8796;
wire n_12218;
wire n_5737;
wire n_12343;
wire n_10733;
wire n_4373;
wire n_8518;
wire n_8919;
wire n_10472;
wire n_12597;
wire n_12316;
wire n_14937;
wire n_14454;
wire n_4711;
wire n_13744;
wire n_11478;
wire n_12834;
wire n_16067;
wire n_15650;
wire n_10066;
wire n_13017;
wire n_12236;
wire n_14335;
wire n_12902;
wire n_6419;
wire n_8372;
wire n_7784;
wire n_9272;
wire n_5768;
wire n_16230;
wire n_10088;
wire n_14887;
wire n_13038;
wire n_7225;
wire n_15199;
wire n_15087;
wire n_8077;
wire n_12892;
wire n_11294;
wire n_15667;
wire n_6244;
wire n_9812;
wire n_6900;
wire n_9337;
wire n_15419;
wire n_15219;
wire n_6755;
wire n_7361;
wire n_6565;
wire n_9432;
wire n_9949;
wire n_10289;
wire n_7705;
wire n_6942;
wire n_11819;
wire n_14889;
wire n_7228;
wire n_13762;
wire n_5350;
wire n_13037;
wire n_5470;
wire n_7932;
wire n_4812;
wire n_11573;
wire n_4409;
wire n_9576;
wire n_7509;
wire n_10145;
wire n_13420;
wire n_5872;
wire n_6862;
wire n_14225;
wire n_7058;
wire n_11005;
wire n_5858;
wire n_15053;
wire n_4629;
wire n_6255;
wire n_6840;
wire n_4638;
wire n_13005;
wire n_6338;
wire n_14805;
wire n_15267;
wire n_15009;
wire n_8262;
wire n_8423;
wire n_5700;
wire n_6037;
wire n_7981;
wire n_9874;
wire n_9577;
wire n_12588;
wire n_15648;
wire n_4913;
wire n_12589;
wire n_5874;
wire n_6266;
wire n_14796;
wire n_14143;
wire n_6488;
wire n_8337;
wire n_9231;
wire n_7164;
wire n_11844;
wire n_15390;
wire n_14044;
wire n_6635;
wire n_7973;
wire n_6815;
wire n_11364;
wire n_9569;
wire n_13184;
wire n_14823;
wire n_15634;
wire n_12790;
wire n_8632;
wire n_14691;
wire n_13535;
wire n_14982;
wire n_7018;
wire n_5873;
wire n_12247;
wire n_7975;
wire n_12699;
wire n_9719;
wire n_16508;
wire n_8358;
wire n_10009;
wire n_14770;
wire n_9552;
wire n_12927;
wire n_11100;
wire n_9279;
wire n_13822;
wire n_14948;
wire n_11902;
wire n_16588;
wire n_6317;
wire n_8199;
wire n_5588;
wire n_11993;
wire n_10443;
wire n_8656;
wire n_7167;
wire n_10756;
wire n_12813;
wire n_14909;
wire n_6480;
wire n_15105;
wire n_14387;
wire n_10918;
wire n_13122;
wire n_13534;
wire n_16572;
wire n_5075;
wire n_11797;
wire n_4968;
wire n_12765;
wire n_14106;
wire n_7865;
wire n_15553;
wire n_13616;
wire n_15690;
wire n_12663;
wire n_10384;
wire n_9289;
wire n_5085;
wire n_11315;
wire n_16349;
wire n_5736;
wire n_15841;
wire n_6561;
wire n_7978;
wire n_7820;
wire n_12706;
wire n_11127;
wire n_10293;
wire n_8881;
wire n_7844;
wire n_14301;
wire n_7134;
wire n_9633;
wire n_15468;
wire n_11153;
wire n_12312;
wire n_10074;
wire n_4572;
wire n_4845;
wire n_9547;
wire n_13097;
wire n_6875;
wire n_13627;
wire n_10934;
wire n_10197;
wire n_15786;
wire n_16350;
wire n_8346;
wire n_5120;
wire n_8761;
wire n_13112;
wire n_15458;
wire n_9085;
wire n_9632;
wire n_10042;
wire n_13734;
wire n_8226;
wire n_11949;
wire n_8402;
wire n_10478;
wire n_7079;
wire n_9690;
wire n_16581;
wire n_9084;
wire n_5928;
wire n_12256;
wire n_5478;
wire n_6016;
wire n_11746;
wire n_11812;
wire n_9371;
wire n_14051;
wire n_13163;
wire n_9711;
wire n_8754;
wire n_9431;
wire n_9847;
wire n_4779;
wire n_14650;
wire n_7267;
wire n_10367;
wire n_14610;
wire n_4599;
wire n_12315;
wire n_11505;
wire n_4437;
wire n_5222;
wire n_9889;
wire n_7316;
wire n_7850;
wire n_10867;
wire n_14100;
wire n_12556;
wire n_12375;
wire n_12998;
wire n_7812;
wire n_7103;
wire n_13723;
wire n_13143;
wire n_9080;
wire n_14601;
wire n_14549;
wire n_8133;
wire n_10168;
wire n_7460;
wire n_6176;
wire n_9519;
wire n_14717;
wire n_14814;
wire n_6367;
wire n_11363;
wire n_15794;
wire n_12156;
wire n_13564;
wire n_14459;
wire n_16426;
wire n_13128;
wire n_4508;
wire n_13490;
wire n_4727;
wire n_4594;
wire n_11530;
wire n_12671;
wire n_10621;
wire n_14913;
wire n_13411;
wire n_7056;
wire n_14645;
wire n_9731;
wire n_8193;
wire n_6572;
wire n_8714;
wire n_12445;
wire n_4429;
wire n_9604;
wire n_7962;
wire n_12856;
wire n_13260;
wire n_4642;
wire n_10085;
wire n_7813;
wire n_15382;
wire n_7755;
wire n_7514;
wire n_7649;
wire n_11151;
wire n_16031;
wire n_6080;
wire n_4865;
wire n_8182;
wire n_8387;
wire n_12525;
wire n_16116;
wire n_6078;
wire n_10613;
wire n_10716;
wire n_12076;
wire n_14090;
wire n_15825;
wire n_6056;
wire n_6717;
wire n_15823;
wire n_5832;
wire n_10664;
wire n_7473;
wire n_13758;
wire n_7200;
wire n_11359;
wire n_7688;
wire n_4562;
wire n_15997;
wire n_8707;
wire n_12357;
wire n_15424;
wire n_4903;
wire n_10561;
wire n_11434;
wire n_9208;
wire n_11791;
wire n_14695;
wire n_15554;
wire n_7611;
wire n_15836;
wire n_6873;
wire n_15966;
wire n_16251;
wire n_16009;
wire n_15309;
wire n_13212;
wire n_14463;
wire n_8494;
wire n_15166;
wire n_5812;
wire n_5743;
wire n_12468;
wire n_9429;
wire n_15216;
wire n_8544;
wire n_11848;
wire n_13503;
wire n_11152;
wire n_15138;
wire n_4998;
wire n_10749;
wire n_16516;
wire n_16318;
wire n_11632;
wire n_15352;
wire n_7795;
wire n_14166;
wire n_12180;
wire n_8788;
wire n_15608;
wire n_14405;
wire n_4522;
wire n_10122;
wire n_10935;
wire n_7038;
wire n_10992;
wire n_14081;
wire n_7723;
wire n_4341;
wire n_11621;
wire n_10560;
wire n_10160;
wire n_9327;
wire n_7404;
wire n_16175;
wire n_12857;
wire n_13171;
wire n_5368;
wire n_8177;
wire n_9854;
wire n_14271;
wire n_7059;
wire n_7450;
wire n_11667;
wire n_12025;
wire n_14854;
wire n_8962;
wire n_9538;
wire n_14254;
wire n_14425;
wire n_5971;
wire n_6327;
wire n_7362;
wire n_16137;
wire n_12208;
wire n_6145;
wire n_11964;
wire n_6539;
wire n_6926;
wire n_15266;
wire n_13421;
wire n_7271;
wire n_7826;
wire n_9713;
wire n_14565;
wire n_11298;
wire n_15796;
wire n_5933;
wire n_13495;
wire n_16501;
wire n_8993;
wire n_6204;
wire n_7076;
wire n_13474;
wire n_4780;
wire n_10300;
wire n_13949;
wire n_13314;
wire n_9588;
wire n_11403;
wire n_14903;
wire n_14218;
wire n_11741;
wire n_15107;
wire n_12383;
wire n_11912;
wire n_4973;
wire n_15537;
wire n_6842;
wire n_12773;
wire n_6866;
wire n_13876;
wire n_14967;
wire n_9044;
wire n_4803;
wire n_9423;
wire n_16619;
wire n_12381;
wire n_9387;
wire n_6030;
wire n_14487;
wire n_4750;
wire n_14883;
wire n_12962;
wire n_6451;
wire n_9813;
wire n_9127;
wire n_14596;
wire n_6514;
wire n_16263;
wire n_9794;
wire n_5996;
wire n_11666;
wire n_12459;
wire n_7105;
wire n_14500;
wire n_13568;
wire n_10140;
wire n_12612;
wire n_9244;
wire n_16387;
wire n_9869;
wire n_11142;
wire n_16369;
wire n_15304;
wire n_7049;
wire n_5903;
wire n_14449;
wire n_15271;
wire n_5986;
wire n_6710;
wire n_4984;
wire n_8278;
wire n_12885;
wire n_14865;
wire n_11644;
wire n_6345;
wire n_15539;
wire n_16165;
wire n_9715;
wire n_15893;
wire n_8618;
wire n_12108;
wire n_9094;
wire n_15432;
wire n_13108;
wire n_5782;
wire n_7535;
wire n_5041;
wire n_13170;
wire n_10862;
wire n_11531;
wire n_4959;
wire n_8248;
wire n_8911;
wire n_9056;
wire n_11357;
wire n_14471;
wire n_4426;
wire n_9407;
wire n_11476;
wire n_15906;
wire n_14476;
wire n_4425;
wire n_13633;
wire n_9985;
wire n_15244;
wire n_4449;
wire n_12089;
wire n_12496;
wire n_14538;
wire n_11824;
wire n_12814;
wire n_7057;
wire n_11959;
wire n_11367;
wire n_15478;
wire n_6957;
wire n_9361;
wire n_15943;
wire n_11921;
wire n_4809;
wire n_8495;
wire n_14532;
wire n_12676;
wire n_13976;
wire n_16578;
wire n_8783;
wire n_12987;
wire n_13579;
wire n_14557;
wire n_11566;
wire n_16650;
wire n_13913;
wire n_8529;
wire n_8733;
wire n_14639;
wire n_12603;
wire n_8990;
wire n_6050;
wire n_7976;
wire n_6444;
wire n_15392;
wire n_10254;
wire n_14340;
wire n_14032;
wire n_14715;
wire n_7944;
wire n_15970;
wire n_13080;
wire n_11208;
wire n_15702;
wire n_7262;
wire n_8647;
wire n_11374;
wire n_12967;
wire n_12452;
wire n_13403;
wire n_15978;
wire n_15857;
wire n_14899;
wire n_15961;
wire n_8574;
wire n_7016;
wire n_10782;
wire n_12292;
wire n_13557;
wire n_12232;
wire n_14952;
wire n_11859;
wire n_12818;
wire n_15616;
wire n_15773;
wire n_10386;
wire n_12128;
wire n_6379;
wire n_14060;
wire n_15589;
wire n_14018;
wire n_11420;
wire n_12754;
wire n_12500;
wire n_15959;
wire n_5563;
wire n_15307;
wire n_13583;
wire n_11026;
wire n_14111;
wire n_8044;
wire n_13309;
wire n_16330;
wire n_5840;
wire n_6719;
wire n_13580;
wire n_7178;
wire n_9439;
wire n_9553;
wire n_11633;
wire n_15292;
wire n_11467;
wire n_15239;
wire n_7506;
wire n_12672;
wire n_8551;
wire n_12063;
wire n_11630;
wire n_14361;
wire n_8330;
wire n_12760;
wire n_16658;
wire n_15444;
wire n_13455;
wire n_15560;
wire n_15065;
wire n_6232;
wire n_15289;
wire n_9132;
wire n_13172;
wire n_5717;
wire n_16234;
wire n_6017;
wire n_9696;
wire n_14943;
wire n_10861;
wire n_9120;
wire n_8879;
wire n_15771;
wire n_15508;
wire n_11203;
wire n_16157;
wire n_11159;
wire n_8052;
wire n_12168;
wire n_4578;
wire n_6362;
wire n_4777;
wire n_11956;
wire n_11975;
wire n_12121;
wire n_5720;
wire n_9332;
wire n_14148;
wire n_16496;
wire n_8903;
wire n_11030;
wire n_4702;
wire n_12590;
wire n_4895;
wire n_5871;
wire n_12924;
wire n_15605;
wire n_7142;
wire n_12577;
wire n_16331;
wire n_10182;
wire n_12732;
wire n_13928;
wire n_6326;
wire n_12649;
wire n_5898;
wire n_16057;
wire n_7125;
wire n_16401;
wire n_6858;
wire n_9252;
wire n_9464;
wire n_6649;
wire n_6283;
wire n_10073;
wire n_4531;
wire n_14619;
wire n_11655;
wire n_15781;
wire n_5072;
wire n_11017;
wire n_12843;
wire n_7241;
wire n_7247;
wire n_14279;
wire n_14448;
wire n_12069;
wire n_10419;
wire n_7172;
wire n_15656;
wire n_15427;
wire n_14622;
wire n_10333;
wire n_12430;
wire n_10317;
wire n_4666;
wire n_7893;
wire n_6213;
wire n_14739;
wire n_16649;
wire n_15687;
wire n_7235;
wire n_8540;
wire n_11248;
wire n_12613;
wire n_6239;
wire n_12270;
wire n_14365;
wire n_9915;
wire n_4617;
wire n_9325;
wire n_16021;
wire n_9196;
wire n_16448;
wire n_13407;
wire n_5896;
wire n_5882;
wire n_4555;
wire n_5940;
wire n_6089;
wire n_7588;
wire n_5650;
wire n_13676;
wire n_9384;
wire n_4969;
wire n_6057;
wire n_6216;
wire n_10017;
wire n_7340;
wire n_12557;
wire n_6974;
wire n_13788;
wire n_14555;
wire n_11141;
wire n_5105;
wire n_12695;
wire n_15467;
wire n_10893;
wire n_11093;
wire n_16537;
wire n_5021;
wire n_14219;
wire n_9251;
wire n_11576;
wire n_8939;
wire n_13584;
wire n_9973;
wire n_5263;
wire n_11117;
wire n_15471;
wire n_6713;
wire n_12139;
wire n_8064;
wire n_9030;
wire n_7657;
wire n_8468;
wire n_4325;
wire n_15968;
wire n_4602;
wire n_5044;
wire n_9665;
wire n_10201;
wire n_13181;
wire n_5134;
wire n_7096;
wire n_12210;
wire n_13327;
wire n_8778;
wire n_11197;
wire n_16487;
wire n_7442;
wire n_15047;
wire n_10093;
wire n_5567;
wire n_8343;
wire n_15014;
wire n_6174;
wire n_15428;
wire n_12006;
wire n_7999;
wire n_10128;
wire n_10675;
wire n_14168;
wire n_6087;
wire n_7593;
wire n_16311;
wire n_12246;
wire n_5249;
wire n_14085;
wire n_8068;
wire n_15342;
wire n_9955;
wire n_15534;
wire n_10539;
wire n_14080;
wire n_5625;
wire n_9007;
wire n_10143;
wire n_7764;
wire n_11777;
wire n_4919;
wire n_10107;
wire n_13975;
wire n_5969;
wire n_10196;
wire n_10121;
wire n_8198;
wire n_14573;
wire n_13085;
wire n_15536;
wire n_7780;
wire n_6828;
wire n_5158;
wire n_7255;
wire n_8693;
wire n_12189;
wire n_13224;
wire n_11469;
wire n_6454;
wire n_5022;
wire n_12625;
wire n_9270;
wire n_14046;
wire n_8452;
wire n_7041;
wire n_7307;
wire n_11518;
wire n_12177;
wire n_14142;
wire n_10742;
wire n_5670;
wire n_10829;
wire n_14512;
wire n_8557;
wire n_6041;
wire n_6918;
wire n_9099;
wire n_12389;
wire n_16214;
wire n_13761;
wire n_9309;
wire n_7350;
wire n_10620;
wire n_10303;
wire n_16189;
wire n_15097;
wire n_10814;
wire n_5276;
wire n_16034;
wire n_9627;
wire n_16219;
wire n_13971;
wire n_11252;
wire n_16563;
wire n_8012;
wire n_14456;
wire n_13364;
wire n_7672;
wire n_11494;
wire n_6664;
wire n_5047;
wire n_14743;
wire n_7318;
wire n_6472;
wire n_10218;
wire n_8114;
wire n_13131;
wire n_14941;
wire n_12995;
wire n_14406;
wire n_13209;
wire n_4791;
wire n_11154;
wire n_11700;
wire n_14859;
wire n_16227;
wire n_5879;
wire n_14563;
wire n_8062;
wire n_4403;
wire n_11883;
wire n_5238;
wire n_16329;
wire n_11256;
wire n_11832;
wire n_14959;
wire n_6166;
wire n_5855;
wire n_12370;
wire n_9136;
wire n_6375;
wire n_12860;
wire n_15387;
wire n_16128;
wire n_16278;
wire n_10975;
wire n_11901;
wire n_6352;
wire n_12974;
wire n_9460;
wire n_15973;
wire n_8542;
wire n_12136;
wire n_10859;
wire n_13078;
wire n_7063;
wire n_7047;
wire n_11652;
wire n_14768;
wire n_14320;
wire n_6632;
wire n_4549;
wire n_11056;
wire n_8576;
wire n_14807;
wire n_13885;
wire n_6238;
wire n_15795;
wire n_10542;
wire n_8038;
wire n_13631;
wire n_13932;
wire n_4349;
wire n_10681;
wire n_15162;
wire n_15606;
wire n_6081;
wire n_9732;
wire n_10459;
wire n_16494;
wire n_11572;
wire n_13370;
wire n_5141;
wire n_11894;
wire n_15929;
wire n_14493;
wire n_10222;
wire n_6724;
wire n_13113;
wire n_13387;
wire n_10524;
wire n_5429;
wire n_6545;
wire n_11583;
wire n_8716;
wire n_11336;
wire n_6705;
wire n_15866;
wire n_9766;
wire n_12758;
wire n_8629;
wire n_9517;
wire n_10463;
wire n_5535;
wire n_14764;
wire n_7074;
wire n_8734;
wire n_9204;
wire n_9689;
wire n_9476;
wire n_11849;
wire n_12142;
wire n_15237;
wire n_15862;
wire n_10659;
wire n_6591;
wire n_7585;
wire n_4948;
wire n_12564;
wire n_5268;
wire n_13643;
wire n_9780;
wire n_6946;
wire n_6002;
wire n_13433;
wire n_15505;
wire n_10403;
wire n_13607;
wire n_12983;
wire n_15538;
wire n_6289;
wire n_7037;
wire n_13697;
wire n_11784;
wire n_6424;
wire n_4941;
wire n_5506;
wire n_5298;
wire n_11399;
wire n_9025;
wire n_8524;
wire n_14244;
wire n_11210;
wire n_7599;
wire n_7928;
wire n_16271;
wire n_15541;
wire n_8768;
wire n_4393;
wire n_10884;
wire n_12886;
wire n_14114;
wire n_15870;
wire n_13980;
wire n_6532;
wire n_4372;
wire n_7293;
wire n_13000;
wire n_16366;
wire n_12035;
wire n_14362;
wire n_13006;
wire n_5640;
wire n_11191;
wire n_12791;
wire n_7600;
wire n_10547;
wire n_14742;
wire n_15996;
wire n_6778;
wire n_14904;
wire n_6721;
wire n_5560;
wire n_13205;
wire n_6644;
wire n_6512;
wire n_4795;
wire n_5544;
wire n_12810;
wire n_6108;
wire n_8258;
wire n_10370;
wire n_4918;
wire n_9597;
wire n_5067;
wire n_13820;
wire n_13947;
wire n_11322;
wire n_5744;
wire n_11892;
wire n_6703;
wire n_12122;
wire n_5384;
wire n_4544;
wire n_15283;
wire n_13428;
wire n_5841;
wire n_12396;
wire n_12241;
wire n_15407;
wire n_7614;
wire n_9343;
wire n_15731;
wire n_15895;
wire n_16554;
wire n_7839;
wire n_5108;
wire n_8299;
wire n_12473;
wire n_7347;
wire n_6086;
wire n_9837;
wire n_11421;
wire n_11057;
wire n_16668;
wire n_10896;
wire n_10969;
wire n_4477;
wire n_11966;
wire n_14474;
wire n_12748;
wire n_7383;
wire n_6805;
wire n_4337;
wire n_8863;
wire n_10562;
wire n_16042;
wire n_5941;
wire n_7759;
wire n_12184;
wire n_10210;
wire n_14417;
wire n_6340;
wire n_5611;
wire n_10054;
wire n_10355;
wire n_6219;
wire n_11551;
wire n_7479;
wire n_6706;
wire n_12571;
wire n_11853;
wire n_9692;
wire n_7395;
wire n_13402;
wire n_10598;
wire n_13034;
wire n_8947;
wire n_4742;
wire n_15494;
wire n_9609;
wire n_10717;
wire n_11118;
wire n_10029;
wire n_7078;
wire n_8188;
wire n_13831;
wire n_6761;
wire n_10007;
wire n_8972;
wire n_11751;
wire n_11423;
wire n_11725;
wire n_5701;
wire n_13635;
wire n_6067;
wire n_10801;
wire n_9206;
wire n_12674;
wire n_8510;
wire n_11410;
wire n_12230;
wire n_15698;
wire n_9567;
wire n_14637;
wire n_6811;
wire n_9061;
wire n_11495;
wire n_9942;
wire n_11712;
wire n_9703;
wire n_4478;
wire n_7372;
wire n_5367;
wire n_12220;
wire n_6868;
wire n_8664;
wire n_10704;
wire n_11520;
wire n_11622;
wire n_4838;
wire n_16552;
wire n_5970;
wire n_16133;
wire n_12169;
wire n_12283;
wire n_12336;
wire n_16638;
wire n_7174;
wire n_14783;
wire n_13268;
wire n_9421;
wire n_5202;
wire n_10740;
wire n_16338;
wire n_13383;
wire n_10457;
wire n_12543;
wire n_15088;
wire n_16129;
wire n_4965;
wire n_16383;
wire n_8021;
wire n_9705;
wire n_16585;
wire n_7803;
wire n_15124;
wire n_11012;
wire n_6111;
wire n_14158;
wire n_12595;
wire n_9624;
wire n_9701;
wire n_11502;
wire n_14236;
wire n_15348;
wire n_11429;
wire n_15802;
wire n_15163;
wire n_10389;
wire n_11631;
wire n_13588;
wire n_13510;
wire n_13570;
wire n_14640;
wire n_6659;
wire n_15688;
wire n_4523;
wire n_9709;
wire n_13677;
wire n_13983;
wire n_6011;
wire n_9416;
wire n_9295;
wire n_13757;
wire n_14036;
wire n_4371;
wire n_6225;
wire n_11842;
wire n_14710;
wire n_12463;
wire n_10990;
wire n_11640;
wire n_12263;
wire n_5502;
wire n_4552;
wire n_6218;
wire n_8982;
wire n_16678;
wire n_9929;
wire n_12920;
wire n_10264;
wire n_5850;
wire n_13317;
wire n_4673;
wire n_13910;
wire n_15029;
wire n_9953;
wire n_13737;
wire n_7086;
wire n_16590;
wire n_6648;
wire n_4607;
wire n_14286;
wire n_15578;
wire n_16640;
wire n_12528;
wire n_10955;
wire n_11389;
wire n_7226;
wire n_6182;
wire n_7927;
wire n_9013;
wire n_12717;
wire n_6520;
wire n_12660;
wire n_9634;
wire n_9532;
wire n_11011;
wire n_5876;
wire n_9998;
wire n_11795;
wire n_5521;
wire n_4837;
wire n_9850;
wire n_6601;
wire n_10916;
wire n_16247;
wire n_12141;
wire n_8584;
wire n_11547;
wire n_11557;
wire n_9346;
wire n_7920;
wire n_13196;
wire n_13520;
wire n_15363;
wire n_12774;
wire n_7810;
wire n_8501;
wire n_14687;
wire n_11904;
wire n_8480;
wire n_10301;
wire n_5088;
wire n_14955;
wire n_8034;
wire n_13018;
wire n_7025;
wire n_9364;
wire n_15886;
wire n_8228;
wire n_15139;
wire n_8076;
wire n_10440;
wire n_6826;
wire n_15856;
wire n_16015;
wire n_15824;
wire n_5856;
wire n_11395;
wire n_8484;
wire n_9472;
wire n_14304;
wire n_15642;
wire n_9836;
wire n_10929;
wire n_14357;
wire n_9107;
wire n_11279;
wire n_11724;
wire n_16393;
wire n_13044;
wire n_11789;
wire n_14152;
wire n_13228;
wire n_11525;
wire n_13518;
wire n_13862;
wire n_8100;
wire n_11999;
wire n_13446;
wire n_13086;
wire n_10837;
wire n_14869;
wire n_14008;
wire n_10554;
wire n_8014;
wire n_8994;
wire n_8091;
wire n_8413;
wire n_4685;
wire n_12746;
wire n_5837;
wire n_4675;
wire n_10149;
wire n_16162;
wire n_10970;
wire n_7768;
wire n_8638;
wire n_16294;
wire n_5825;
wire n_14651;
wire n_16285;
wire n_5491;
wire n_5496;
wire n_5802;
wire n_14965;
wire n_13887;
wire n_7982;
wire n_15791;
wire n_12190;
wire n_14927;
wire n_12787;
wire n_8804;
wire n_13881;
wire n_15484;
wire n_15152;
wire n_11383;
wire n_12799;
wire n_11847;
wire n_11976;
wire n_5178;
wire n_9317;
wire n_12657;
wire n_9769;
wire n_5547;
wire n_15205;
wire n_15882;
wire n_13747;
wire n_8158;
wire n_12511;
wire n_11167;
wire n_6879;
wire n_12532;
wire n_8469;
wire n_7567;
wire n_10238;
wire n_8765;
wire n_8433;
wire n_10102;
wire n_8931;
wire n_5596;
wire n_6074;
wire n_5983;
wire n_8213;
wire n_14472;
wire n_4588;
wire n_10534;
wire n_11825;
wire n_4653;
wire n_4435;
wire n_10932;
wire n_10619;
wire n_7684;
wire n_11049;
wire n_14354;
wire n_14974;
wire n_15532;
wire n_8451;
wire n_5604;
wire n_5411;
wire n_8334;
wire n_12743;
wire n_16523;
wire n_16083;
wire n_8731;
wire n_10589;
wire n_11681;
wire n_11611;
wire n_8385;
wire n_10890;
wire n_9156;
wire n_16113;
wire n_11202;
wire n_4728;
wire n_4999;
wire n_15587;
wire n_4385;
wire n_6642;
wire n_6847;
wire n_10707;
wire n_4922;
wire n_10552;
wire n_10248;
wire n_5815;
wire n_7370;
wire n_9748;
wire n_13365;
wire n_15254;
wire n_6595;
wire n_7771;
wire n_15322;
wire n_13539;
wire n_9350;
wire n_12408;
wire n_11780;
wire n_16287;
wire n_16169;
wire n_5695;
wire n_6027;
wire n_8539;
wire n_16289;
wire n_10205;
wire n_7026;
wire n_7701;
wire n_7053;
wire n_14618;
wire n_16342;
wire n_15747;
wire n_9226;
wire n_5235;
wire n_10110;
wire n_13899;
wire n_6306;
wire n_11230;
wire n_6720;
wire n_11930;
wire n_10608;
wire n_16355;
wire n_11688;
wire n_6888;
wire n_7173;
wire n_4350;
wire n_7042;
wire n_12715;
wire n_11709;
wire n_12434;
wire n_14328;
wire n_12628;
wire n_8122;
wire n_6095;
wire n_13444;
wire n_16235;
wire n_8432;
wire n_11663;
wire n_5331;
wire n_16504;
wire n_4330;
wire n_7592;
wire n_16540;
wire n_14209;
wire n_11331;
wire n_14429;
wire n_5311;
wire n_12979;
wire n_16436;
wire n_9528;
wire n_6590;
wire n_14348;
wire n_10638;
wire n_7583;
wire n_12201;
wire n_14086;
wire n_12499;
wire n_6559;
wire n_9112;
wire n_15799;
wire n_12448;
wire n_4621;
wire n_11876;
wire n_5797;
wire n_9235;
wire n_16570;
wire n_10610;
wire n_11187;
wire n_12761;
wire n_5572;
wire n_13852;
wire n_16455;
wire n_9333;
wire n_7151;
wire n_15004;
wire n_5565;
wire n_14270;
wire n_15238;
wire n_8950;
wire n_14089;
wire n_10758;
wire n_16625;
wire n_13431;
wire n_10190;
wire n_16025;
wire n_5520;
wire n_11804;
wire n_14234;
wire n_14125;
wire n_5800;
wire n_6562;
wire n_5984;
wire n_6287;
wire n_12809;
wire n_13614;
wire n_4785;
wire n_8347;
wire n_4683;
wire n_14552;
wire n_7353;
wire n_9330;
wire n_12538;
wire n_14208;
wire n_14025;
wire n_7758;
wire n_13779;
wire n_12446;
wire n_9490;
wire n_15693;
wire n_12029;
wire n_9355;
wire n_11052;
wire n_15954;
wire n_5060;
wire n_9523;
wire n_14584;
wire n_15386;
wire n_4986;
wire n_14620;
wire n_5888;
wire n_5669;
wire n_14575;
wire n_9024;
wire n_9574;
wire n_11694;
wire n_5772;
wire n_15349;
wire n_7571;
wire n_9582;
wire n_4775;
wire n_5884;
wire n_10060;
wire n_6671;
wire n_13470;
wire n_16249;
wire n_11009;
wire n_6812;
wire n_12361;
wire n_4864;
wire n_9288;
wire n_9686;
wire n_16435;
wire n_9488;
wire n_5758;
wire n_10748;
wire n_4674;
wire n_13068;
wire n_4481;
wire n_6308;
wire n_7897;
wire n_11446;
wire n_10910;
wire n_10162;
wire n_8242;
wire n_4669;
wire n_7118;
wire n_15002;
wire n_8284;
wire n_9964;
wire n_11540;
wire n_13248;
wire n_7792;
wire n_15985;
wire n_13842;
wire n_8161;
wire n_9702;
wire n_7510;
wire n_9819;
wire n_15338;
wire n_15378;
wire n_6662;
wire n_11291;
wire n_8184;
wire n_5603;
wire n_9154;
wire n_6525;
wire n_7422;
wire n_13107;
wire n_14501;
wire n_6738;
wire n_12307;
wire n_13119;
wire n_5763;
wire n_8703;
wire n_10014;
wire n_15723;
wire n_7109;
wire n_12642;
wire n_15839;
wire n_12484;
wire n_6128;
wire n_16135;
wire n_13549;
wire n_8822;
wire n_6029;
wire n_14790;
wire n_14999;
wire n_10677;
wire n_12187;
wire n_5751;
wire n_15852;
wire n_5264;
wire n_16080;
wire n_4525;
wire n_12321;
wire n_5924;
wire n_9992;
wire n_11247;
wire n_15180;
wire n_15692;
wire n_7253;
wire n_8384;
wire n_5712;
wire n_6445;
wire n_12669;
wire n_13106;
wire n_8476;
wire n_14296;
wire n_14294;
wire n_6702;
wire n_11927;
wire n_16674;
wire n_13720;
wire n_11179;
wire n_16326;
wire n_6701;
wire n_16571;
wire n_7339;
wire n_14862;
wire n_13706;
wire n_8359;
wire n_7380;
wire n_4484;
wire n_13903;
wire n_15808;
wire n_9051;
wire n_8736;
wire n_8545;
wire n_10385;
wire n_4497;
wire n_7749;
wire n_10078;
wire n_10105;
wire n_11514;
wire n_12470;
wire n_12994;
wire n_11321;
wire n_14313;
wire n_15785;
wire n_9500;
wire n_8705;
wire n_14574;
wire n_10215;
wire n_14451;
wire n_11779;
wire n_14059;
wire n_7508;
wire n_5694;
wire n_9455;
wire n_10251;
wire n_4871;
wire n_8708;
wire n_14211;
wire n_15234;
wire n_10834;
wire n_7574;
wire n_14092;
wire n_4700;
wire n_4883;
wire n_9980;
wire n_14509;
wire n_14394;
wire n_11882;
wire n_13516;
wire n_11647;
wire n_12064;
wire n_15027;
wire n_14273;
wire n_15404;
wire n_10706;
wire n_12462;
wire n_6005;
wire n_8872;
wire n_12696;
wire n_4453;
wire n_9555;
wire n_15735;
wire n_11133;
wire n_5449;
wire n_16462;
wire n_14845;
wire n_6169;
wire n_8238;
wire n_15230;
wire n_12735;
wire n_7713;
wire n_15465;
wire n_4564;
wire n_15372;
wire n_13560;
wire n_15700;
wire n_11222;
wire n_9200;
wire n_16279;
wire n_16182;
wire n_5146;
wire n_10709;
wire n_12646;
wire n_10871;
wire n_15858;
wire n_15875;
wire n_7352;
wire n_16405;
wire n_5926;
wire n_10304;
wire n_5398;
wire n_4573;
wire n_5860;
wire n_6936;
wire n_4535;
wire n_14624;
wire n_10244;
wire n_15934;
wire n_16600;
wire n_15036;
wire n_14765;
wire n_16121;
wire n_7704;
wire n_11571;
wire n_7487;
wire n_9986;
wire n_16170;
wire n_14120;
wire n_14995;
wire n_8844;
wire n_13147;
wire n_6302;
wire n_7641;
wire n_13794;
wire n_6106;
wire n_7203;
wire n_12999;
wire n_13537;
wire n_14260;
wire n_14407;
wire n_9397;
wire n_7169;
wire n_10407;
wire n_11259;
wire n_7670;
wire n_12682;
wire n_16010;
wire n_14802;
wire n_9673;
wire n_14434;
wire n_14175;
wire n_4695;
wire n_6848;
wire n_8642;
wire n_10043;
wire n_9855;
wire n_10568;
wire n_11875;
wire n_11941;
wire n_5919;
wire n_4368;
wire n_8159;
wire n_14834;
wire n_12111;
wire n_15780;
wire n_8912;
wire n_14346;
wire n_7439;
wire n_13463;
wire n_9496;
wire n_16241;
wire n_15189;
wire n_8110;
wire n_14275;
wire n_5319;
wire n_10796;
wire n_14506;
wire n_10016;
wire n_9008;
wire n_12903;
wire n_12079;
wire n_15335;
wire n_6343;
wire n_12593;
wire n_16018;
wire n_14615;
wire n_5270;
wire n_10030;
wire n_15222;
wire n_15227;
wire n_8805;
wire n_6850;
wire n_12864;
wire n_15285;
wire n_5005;
wire n_9653;
wire n_11602;
wire n_10272;
wire n_8989;
wire n_13294;
wire n_15689;
wire n_9640;
wire n_6098;
wire n_12413;
wire n_6014;
wire n_7209;
wire n_7112;
wire n_15026;
wire n_13895;
wire n_11307;
wire n_5181;
wire n_13936;
wire n_13933;
wire n_6979;
wire n_7815;
wire n_13222;
wire n_7934;
wire n_9545;
wire n_13813;
wire n_8111;
wire n_16190;
wire n_9629;
wire n_9603;
wire n_11578;
wire n_6865;
wire n_10432;
wire n_12719;
wire n_7276;
wire n_10342;
wire n_8056;
wire n_15361;
wire n_5043;
wire n_8739;
wire n_6747;
wire n_9674;
wire n_13714;
wire n_16244;
wire n_5583;
wire n_4654;
wire n_13438;
wire n_6433;
wire n_15987;
wire n_10462;
wire n_12725;
wire n_6640;
wire n_16030;
wire n_15850;
wire n_15469;
wire n_11769;
wire n_8856;
wire n_6142;
wire n_9930;
wire n_16079;
wire n_11908;
wire n_14371;
wire n_12925;
wire n_5775;
wire n_14901;
wire n_6462;
wire n_7769;
wire n_14988;
wire n_6034;
wire n_9781;
wire n_10291;
wire n_13159;
wire n_4597;
wire n_9659;
wire n_14333;
wire n_16293;
wire n_7233;
wire n_8732;
wire n_13636;
wire n_13506;
wire n_13287;
wire n_11913;
wire n_14788;
wire n_7602;
wire n_9296;
wire n_7034;
wire n_9897;
wire n_5220;
wire n_9241;
wire n_14590;
wire n_11341;
wire n_7390;
wire n_10787;
wire n_4867;
wire n_13256;
wire n_10669;
wire n_13389;
wire n_14567;
wire n_6870;
wire n_6221;
wire n_14603;
wire n_8231;
wire n_16308;
wire n_8185;
wire n_11466;
wire n_6279;
wire n_5061;
wire n_15265;
wire n_15040;
wire n_6775;
wire n_13905;
wire n_9291;
wire n_7881;
wire n_12290;
wire n_9906;
wire n_9369;
wire n_11982;
wire n_13717;
wire n_5029;
wire n_5127;
wire n_12317;
wire n_13302;
wire n_6071;
wire n_11873;
wire n_7598;
wire n_9583;
wire n_12440;
wire n_15119;
wire n_15821;
wire n_8908;
wire n_10185;
wire n_11182;
wire n_10092;
wire n_16085;
wire n_16250;
wire n_15768;
wire n_8220;
wire n_6833;
wire n_12150;
wire n_6793;
wire n_6767;
wire n_11815;
wire n_6295;
wire n_12782;
wire n_4721;
wire n_15256;
wire n_11231;
wire n_14145;
wire n_8090;
wire n_13740;
wire n_8053;
wire n_10184;
wire n_10111;
wire n_11991;
wire n_12875;
wire n_15982;
wire n_15064;
wire n_15300;
wire n_6385;
wire n_11354;
wire n_11807;
wire n_9262;
wire n_7426;
wire n_13918;
wire n_8137;
wire n_7045;
wire n_13775;
wire n_12027;
wire n_9851;
wire n_11799;
wire n_8740;
wire n_8009;
wire n_7852;
wire n_10983;
wire n_9987;
wire n_15218;
wire n_15452;
wire n_7984;
wire n_11727;
wire n_13615;
wire n_15625;
wire n_6788;
wire n_7014;
wire n_12192;
wire n_12633;
wire n_10430;
wire n_14779;
wire n_15114;
wire n_8305;
wire n_4614;
wire n_14973;
wire n_10277;
wire n_8163;
wire n_7220;
wire n_6709;
wire n_16632;
wire n_14465;
wire n_13412;
wire n_16028;
wire n_4422;
wire n_10948;
wire n_11749;
wire n_6712;
wire n_6550;
wire n_10525;
wire n_9507;
wire n_14287;
wire n_11528;
wire n_7416;
wire n_11300;
wire n_6143;
wire n_15296;
wire n_15828;
wire n_8841;
wire n_14553;
wire n_16126;
wire n_13457;
wire n_5177;
wire n_9657;
wire n_12551;
wire n_12196;
wire n_5483;
wire n_16594;
wire n_16370;
wire n_15136;
wire n_6743;
wire n_12497;
wire n_4632;
wire n_15043;
wire n_10354;
wire n_16223;
wire n_12412;
wire n_16168;
wire n_11880;
wire n_5785;
wire n_16602;
wire n_15915;
wire n_7465;
wire n_14528;
wire n_13177;
wire n_5967;
wire n_4546;
wire n_10049;
wire n_12724;
wire n_4583;
wire n_4963;
wire n_14958;
wire n_15551;
wire n_6672;
wire n_9457;
wire n_4966;
wire n_9485;
wire n_5780;
wire n_4714;
wire n_7679;
wire n_5037;
wire n_13940;
wire n_7936;
wire n_8966;
wire n_6084;
wire n_11249;
wire n_15449;
wire n_4847;
wire n_10287;
wire n_15992;
wire n_8538;
wire n_11039;
wire n_7738;
wire n_14342;
wire n_12101;
wire n_10119;
wire n_13693;
wire n_11145;
wire n_12606;
wire n_11986;
wire n_16684;
wire n_8395;
wire n_10900;
wire n_14798;
wire n_5966;
wire n_10349;
wire n_6634;
wire n_14107;
wire n_14758;
wire n_4668;
wire n_5213;
wire n_8961;
wire n_14781;
wire n_10849;
wire n_7462;
wire n_13333;
wire n_4635;
wire n_13229;
wire n_5735;
wire n_12118;
wire n_13311;
wire n_14409;
wire n_14724;
wire n_16340;
wire n_7490;
wire n_11380;
wire n_15737;
wire n_14291;
wire n_7545;
wire n_10792;
wire n_15573;
wire n_11513;
wire n_8625;
wire n_13296;
wire n_16020;
wire n_7160;
wire n_7464;
wire n_8937;
wire n_9809;
wire n_6919;
wire n_14611;
wire n_10750;
wire n_13756;
wire n_7805;
wire n_10995;
wire n_7115;
wire n_7295;
wire n_12087;
wire n_13675;
wire n_9192;
wire n_15022;
wire n_14338;
wire n_7348;
wire n_5752;
wire n_11618;
wire n_14266;
wire n_12594;
wire n_5360;
wire n_10673;
wire n_12460;
wire n_6681;
wire n_6104;
wire n_16071;
wire n_8179;
wire n_10537;
wire n_11861;
wire n_15051;
wire n_6548;
wire n_15394;
wire n_6082;
wire n_6993;
wire n_8511;
wire n_15916;
wire n_6973;
wire n_12081;
wire n_15941;
wire n_10426;
wire n_4405;
wire n_4413;
wire n_9558;
wire n_11594;
wire n_7453;
wire n_16468;
wire n_9167;
wire n_12082;
wire n_8715;
wire n_9655;
wire n_10241;
wire n_12474;
wire n_15639;
wire n_10684;
wire n_4759;
wire n_7162;
wire n_11436;
wire n_12346;
wire n_16655;
wire n_4667;
wire n_5081;
wire n_11729;
wire n_15039;
wire n_8371;
wire n_8702;
wire n_13916;
wire n_15195;
wire n_8116;
wire n_7946;
wire n_8195;
wire n_8806;
wire n_11458;
wire n_12989;
wire n_14069;
wire n_12244;
wire n_5877;
wire n_9991;
wire n_16188;
wire n_15644;
wire n_14255;
wire n_11670;
wire n_11366;
wire n_11872;
wire n_7681;
wire n_8845;
wire n_15198;
wire n_11504;
wire n_6018;
wire n_6619;
wire n_13620;
wire n_16434;
wire n_5189;
wire n_13930;
wire n_7702;
wire n_6676;
wire n_13981;
wire n_8149;
wire n_10823;
wire n_4637;
wire n_9976;
wire n_8042;
wire n_11516;
wire n_14766;
wire n_10390;
wire n_12464;
wire n_11106;
wire n_8392;
wire n_9560;
wire n_14592;
wire n_8095;
wire n_7210;
wire n_5869;
wire n_14659;
wire n_10830;
wire n_15109;
wire n_11132;
wire n_6718;
wire n_15007;
wire n_5118;
wire n_7503;
wire n_10824;
wire n_6854;
wire n_15400;
wire n_15197;
wire n_16216;
wire n_15485;
wire n_4977;
wire n_14841;
wire n_13624;
wire n_5632;
wire n_8519;
wire n_5582;
wire n_14277;
wire n_5425;
wire n_5886;
wire n_8269;
wire n_13493;
wire n_6032;
wire n_9047;
wire n_13805;
wire n_16389;
wire n_12953;
wire n_12842;
wire n_15224;
wire n_8968;
wire n_12481;
wire n_16243;
wire n_9319;
wire n_9215;
wire n_11406;
wire n_5446;
wire n_11316;
wire n_7855;
wire n_14029;
wire n_11047;
wire n_14963;
wire n_8050;
wire n_12450;
wire n_5224;
wire n_12817;
wire n_4590;
wire n_8399;
wire n_5090;
wire n_14648;
wire n_11767;
wire n_9599;
wire n_14056;
wire n_10985;
wire n_11559;
wire n_9072;
wire n_13866;
wire n_4929;
wire n_9401;
wire n_5678;
wire n_13695;
wire n_12435;
wire n_9428;
wire n_10340;
wire n_10946;
wire n_11586;
wire n_6981;
wire n_15817;
wire n_15344;
wire n_13288;
wire n_7065;
wire n_12149;
wire n_13669;
wire n_9216;
wire n_12002;
wire n_12836;
wire n_4835;
wire n_11519;
wire n_11109;
wire n_13065;
wire n_13840;
wire n_11229;
wire n_13548;
wire n_15710;
wire n_16601;
wire n_16159;
wire n_11591;
wire n_11961;
wire n_11195;
wire n_14251;
wire n_6122;
wire n_11397;
wire n_11225;
wire n_16240;
wire n_7911;
wire n_6765;
wire n_9747;
wire n_4565;
wire n_5414;
wire n_14526;
wire n_13487;
wire n_12840;
wire n_7330;
wire n_14605;
wire n_5437;
wire n_8883;
wire n_10634;
wire n_8586;
wire n_12846;
wire n_9202;
wire n_4586;
wire n_11058;
wire n_9058;
wire n_15888;
wire n_7336;
wire n_11471;
wire n_14705;
wire n_7446;
wire n_13543;
wire n_8401;
wire n_7854;
wire n_10577;
wire n_5454;
wire n_10351;
wire n_13772;
wire n_14679;
wire n_4734;
wire n_7493;
wire n_10961;
wire n_12940;
wire n_10460;
wire n_10780;
wire n_15487;
wire n_7357;
wire n_8756;
wire n_11324;
wire n_8737;
wire n_13925;
wire n_10334;
wire n_4434;
wire n_12945;
wire n_13406;
wire n_16371;
wire n_7923;
wire n_5307;
wire n_10379;
wire n_10151;
wire n_6439;
wire n_11614;
wire n_14040;
wire n_8602;
wire n_14054;
wire n_13368;
wire n_8240;
wire n_12850;
wire n_13469;
wire n_14507;
wire n_7714;
wire n_5407;
wire n_10411;
wire n_15242;
wire n_13249;
wire n_9484;
wire n_12984;
wire n_16193;
wire n_10989;
wire n_8422;
wire n_10939;
wire n_13587;
wire n_12224;
wire n_5913;
wire n_7088;
wire n_9305;
wire n_9394;
wire n_9999;
wire n_8878;
wire n_11361;
wire n_10090;
wire n_6406;
wire n_7440;
wire n_11144;
wire n_14857;
wire n_6945;
wire n_14872;
wire n_8112;
wire n_14034;
wire n_11567;
wire n_10962;
wire n_7029;
wire n_14797;
wire n_11128;
wire n_9292;
wire n_9622;
wire n_15677;
wire n_10721;
wire n_8593;
wire n_12197;
wire n_14177;
wire n_14093;
wire n_10186;
wire n_14607;
wire n_4833;
wire n_11580;
wire n_11841;
wire n_11025;
wire n_12007;
wire n_5062;
wire n_6618;
wire n_13326;
wire n_15901;
wire n_6474;
wire n_13082;
wire n_14453;
wire n_10191;
wire n_5230;
wire n_5944;
wire n_6226;
wire n_4888;
wire n_13094;
wire n_7317;
wire n_10856;
wire n_12403;
wire n_6000;
wire n_12679;
wire n_13481;
wire n_9584;
wire n_13692;
wire n_8194;
wire n_9461;
wire n_8055;
wire n_11168;
wire n_14921;
wire n_8579;
wire n_6816;
wire n_10914;
wire n_10911;
wire n_10928;
wire n_12756;
wire n_8360;
wire n_12018;
wire n_5008;
wire n_6425;
wire n_14457;
wire n_5004;
wire n_5294;
wire n_6493;
wire n_16097;
wire n_9845;
wire n_16147;
wire n_6502;
wire n_6250;
wire n_7374;
wire n_6288;
wire n_5974;
wire n_14382;
wire n_14389;
wire n_11937;
wire n_12872;
wire n_13396;
wire n_7522;
wire n_6492;
wire n_10071;
wire n_8755;
wire n_4527;
wire n_6046;
wire n_11460;
wire n_14517;
wire n_8251;
wire n_13713;
wire n_5323;
wire n_11565;
wire n_4790;
wire n_14621;
wire n_12372;
wire n_9618;
wire n_14911;
wire n_6118;
wire n_13608;
wire n_5810;
wire n_4561;
wire n_15405;
wire n_4461;
wire n_7046;
wire n_11192;
wire n_11808;
wire n_15643;
wire n_13257;
wire n_10956;
wire n_4949;
wire n_6852;
wire n_15420;
wire n_8677;
wire n_13052;
wire n_7468;
wire n_9091;
wire n_11013;
wire n_5991;
wire n_14934;
wire n_13914;
wire n_16634;
wire n_5069;
wire n_12453;
wire n_12572;
wire n_14663;
wire n_10035;
wire n_5702;
wire n_13393;
wire n_6251;
wire n_9828;
wire n_14962;
wire n_15652;
wire n_13922;
wire n_9699;
wire n_13277;
wire n_12340;
wire n_13423;
wire n_8108;
wire n_14578;
wire n_15653;
wire n_5914;
wire n_5243;
wire n_12955;
wire n_12068;
wire n_10252;
wire n_5250;
wire n_16641;
wire n_11555;
wire n_13494;
wire n_6869;
wire n_10041;
wire n_9321;
wire n_15499;
wire n_14625;
wire n_5590;
wire n_10345;
wire n_14514;
wire n_10059;
wire n_5260;
wire n_8325;
wire n_9751;
wire n_7621;
wire n_7359;
wire n_8498;
wire n_5809;
wire n_14256;
wire n_15016;
wire n_10543;
wire n_7924;
wire n_4782;
wire n_12394;
wire n_13578;
wire n_7659;
wire n_9005;
wire n_9161;
wire n_14204;
wire n_16203;
wire n_8875;
wire n_4378;
wire n_5349;
wire n_8274;
wire n_9585;
wire n_15855;
wire n_7153;
wire n_11101;
wire n_12954;
wire n_7836;
wire n_10737;
wire n_12662;
wire n_15697;
wire n_4876;
wire n_14082;
wire n_6146;
wire n_8504;
wire n_10464;
wire n_7280;
wire n_10644;
wire n_12801;
wire n_13448;
wire n_14688;
wire n_15865;
wire n_5813;
wire n_9293;
wire n_12503;
wire n_13708;
wire n_10365;
wire n_13767;
wire n_5833;
wire n_11781;
wire n_11055;
wire n_7886;
wire n_4358;
wire n_15728;
wire n_16616;
wire n_14832;
wire n_15202;
wire n_10982;
wire n_5805;
wire n_5616;
wire n_9648;
wire n_12871;
wire n_6884;
wire n_7664;
wire n_7012;
wire n_12965;
wire n_13029;
wire n_10591;
wire n_11845;
wire n_12486;
wire n_14571;
wire n_16400;
wire n_6631;
wire n_12788;
wire n_12369;
wire n_4469;
wire n_9498;
wire n_7376;
wire n_7577;
wire n_7308;
wire n_5169;
wire n_15707;
wire n_16328;
wire n_5816;
wire n_10809;
wire n_15396;
wire n_8927;
wire n_10899;
wire n_15347;
wire n_15909;
wire n_16396;
wire n_9639;
wire n_15155;
wire n_11898;
wire n_10137;
wire n_12084;
wire n_12686;
wire n_15250;
wire n_6228;
wire n_6711;
wire n_11997;
wire n_11884;
wire n_5416;
wire n_8946;
wire n_14881;
wire n_16517;
wire n_13090;
wire n_14527;
wire n_12822;
wire n_13541;
wire n_13307;
wire n_13371;
wire n_11863;
wire n_4493;
wire n_4924;
wire n_7279;
wire n_7971;
wire n_13908;
wire n_9646;
wire n_8017;
wire n_12264;
wire n_13312;
wire n_11761;
wire n_8474;
wire n_9984;
wire n_16174;
wire n_8232;
wire n_7275;
wire n_8795;
wire n_7195;
wire n_10600;
wire n_10794;
wire n_6102;
wire n_9649;
wire n_14703;
wire n_8904;
wire n_11199;
wire n_13533;
wire n_6274;
wire n_10833;
wire n_8838;
wire n_11264;
wire n_12109;
wire n_16283;
wire n_10629;
wire n_9562;
wire n_7007;
wire n_7070;
wire n_4539;
wire n_8382;
wire n_4421;
wire n_13023;
wire n_16088;
wire n_6072;
wire n_7610;
wire n_12303;
wire n_9501;
wire n_11896;
wire n_4793;
wire n_13856;
wire n_16229;
wire n_15607;
wire n_4498;
wire n_10006;
wire n_7259;
wire n_11757;
wire n_12274;
wire n_12320;
wire n_14588;
wire n_15879;
wire n_15315;
wire n_9759;
wire n_6353;
wire n_4953;
wire n_12622;
wire n_6992;
wire n_11185;
wire n_8128;
wire n_12659;
wire n_13440;
wire n_6818;
wire n_15226;
wire n_15746;
wire n_13436;
wire n_10206;
wire n_15921;
wire n_6322;
wire n_5167;
wire n_15425;
wire n_5661;
wire n_5830;
wire n_5932;
wire n_11345;
wire n_12380;
wire n_13245;
wire n_12629;
wire n_7539;
wire n_12586;
wire n_8794;
wire n_11760;
wire n_7616;
wire n_9733;
wire n_12868;
wire n_12282;
wire n_8189;
wire n_6498;
wire n_11081;
wire n_8481;
wire n_10275;
wire n_7775;
wire n_13011;
wire n_16687;
wire n_4505;
wire n_11392;
wire n_9981;
wire n_14858;
wire n_7930;
wire n_5558;
wire n_8787;
wire n_5687;
wire n_7661;
wire n_16513;
wire n_6378;
wire n_13911;
wire n_5383;
wire n_14495;
wire n_16498;
wire n_5126;
wire n_8205;
wire n_14165;
wire n_5051;
wire n_9907;
wire n_13088;
wire n_6976;
wire n_5587;
wire n_10941;
wire n_11024;
wire n_6304;
wire n_5236;
wire n_12269;
wire n_13538;
wire n_7640;
wire n_14617;
wire n_13701;
wire n_9816;
wire n_13787;
wire n_10498;
wire n_11424;
wire n_13486;
wire n_12585;
wire n_5012;
wire n_14021;
wire n_13674;
wire n_14263;
wire n_11463;
wire n_13912;
wire n_14303;
wire n_10292;
wire n_7969;
wire n_6864;
wire n_8605;
wire n_11278;
wire n_14445;
wire n_10358;
wire n_7548;
wire n_10635;
wire n_13626;
wire n_9944;
wire n_4450;
wire n_5954;
wire n_6156;
wire n_12832;
wire n_12913;
wire n_6998;
wire n_5025;
wire n_8067;
wire n_7587;
wire n_7064;
wire n_16158;
wire n_12301;
wire n_12338;
wire n_9643;
wire n_7615;
wire n_5651;
wire n_6930;
wire n_4630;
wire n_9605;
wire n_12802;
wire n_12154;
wire n_8000;
wire n_11569;
wire n_10064;
wire n_14427;
wire n_7197;
wire n_9676;
wire n_5645;
wire n_15822;
wire n_11881;
wire n_7393;
wire n_11332;
wire n_6917;
wire n_13629;
wire n_6937;
wire n_7591;
wire n_13207;
wire n_14980;
wire n_9963;
wire n_5766;
wire n_11404;
wire n_7727;
wire n_7358;
wire n_16488;
wire n_15994;
wire n_7324;
wire n_9950;
wire n_5878;
wire n_5671;
wire n_10152;
wire n_11935;
wire n_13589;
wire n_15730;
wire n_4534;
wire n_15685;
wire n_6301;
wire n_9788;
wire n_6929;
wire n_15570;
wire n_15562;
wire n_11309;
wire n_16273;
wire n_8719;
wire n_16140;
wire n_8045;
wire n_10785;
wire n_16032;
wire n_7729;
wire n_13872;
wire n_15493;
wire n_12341;
wire n_12615;
wire n_4494;
wire n_6436;
wire n_5412;
wire n_14475;
wire n_8209;
wire n_13357;
wire n_10802;
wire n_14477;
wire n_4786;
wire n_10815;
wire n_7565;
wire n_6699;
wire n_12926;
wire n_16624;
wire n_14809;
wire n_9213;
wire n_4579;
wire n_7291;
wire n_14725;
wire n_7631;
wire n_14522;
wire n_8784;
wire n_7382;
wire n_4811;
wire n_13869;
wire n_13955;
wire n_6874;
wire n_7387;
wire n_6259;
wire n_9212;
wire n_9340;
wire n_16527;
wire n_13561;
wire n_12167;
wire n_14720;
wire n_9473;
wire n_14400;
wire n_4857;
wire n_13026;
wire n_10490;
wire n_7437;
wire n_15019;
wire n_6677;
wire n_12161;
wire n_16432;
wire n_13499;
wire n_12085;
wire n_14843;
wire n_11735;
wire n_7618;
wire n_10647;
wire n_16084;
wire n_9320;
wire n_10523;
wire n_8769;
wire n_6764;
wire n_8575;
wire n_13554;
wire n_12298;
wire n_10081;
wire n_5733;
wire n_10324;
wire n_11189;
wire n_6780;
wire n_12569;
wire n_8815;
wire n_11582;
wire n_14929;
wire n_6620;
wire n_6597;
wire n_12044;
wire n_9303;
wire n_11105;
wire n_11705;
wire n_5148;
wire n_8261;
wire n_7673;
wire n_13698;
wire n_6830;
wire n_13894;
wire n_12456;
wire n_13104;
wire n_8655;
wire n_7282;
wire n_6586;
wire n_9968;
wire n_11474;
wire n_10808;
wire n_6333;
wire n_10474;
wire n_7139;
wire n_8745;
wire n_12689;
wire n_5791;
wire n_5727;
wire n_10657;
wire n_8086;
wire n_16612;
wire n_15466;
wire n_13595;
wire n_5946;
wire n_8789;
wire n_5997;
wire n_13943;
wire n_7953;
wire n_13540;
wire n_6428;
wire n_5328;
wire n_7379;
wire n_10687;
wire n_14642;
wire n_9722;
wire n_13283;
wire n_12042;
wire n_12155;
wire n_14827;
wire n_5657;
wire n_15481;
wire n_8901;
wire n_11078;
wire n_11130;
wire n_13465;
wire n_8695;
wire n_4974;
wire n_12373;
wire n_15615;
wire n_5975;
wire n_15664;
wire n_16149;
wire n_4911;
wire n_8173;
wire n_11664;
wire n_12072;
wire n_12110;
wire n_4436;
wire n_14579;
wire n_8363;
wire n_15388;
wire n_5119;
wire n_10652;
wire n_4569;
wire n_10545;
wire n_9669;
wire n_8665;
wire n_13098;
wire n_13733;
wire n_16557;
wire n_6510;
wire n_8282;
wire n_15847;
wire n_9388;
wire n_5938;
wire n_15972;
wire n_6237;
wire n_12216;
wire n_11752;
wire n_12040;
wire n_12654;
wire n_14141;
wire n_5602;
wire n_9379;
wire n_11992;
wire n_5097;
wire n_15790;
wire n_4985;
wire n_7751;
wire n_10869;
wire n_14880;
wire n_14718;
wire n_4384;
wire n_14975;
wire n_13142;
wire n_7581;
wire n_13180;
wire n_13116;
wire n_11783;
wire n_6360;
wire n_15217;
wire n_14589;
wire n_5246;
wire n_10453;
wire n_12386;
wire n_14257;
wire n_4858;
wire n_4678;
wire n_13308;
wire n_9952;
wire n_16492;
wire n_15323;
wire n_9911;
wire n_12183;
wire n_5579;
wire n_8835;
wire n_16317;
wire n_15187;
wire n_9256;
wire n_10668;
wire n_10346;
wire n_12419;
wire n_13763;
wire n_5750;
wire n_10688;
wire n_4823;
wire n_13785;
wire n_5831;
wire n_4363;
wire n_7742;
wire n_9274;
wire n_12964;
wire n_10473;
wire n_15712;
wire n_16404;
wire n_14007;
wire n_5107;
wire n_5095;
wire n_15099;
wire n_8493;
wire n_7346;
wire n_10331;
wire n_11439;
wire n_14655;
wire n_10957;
wire n_13373;
wire n_7579;
wire n_13517;
wire n_12863;
wire n_10352;
wire n_11188;
wire n_7428;
wire n_12221;
wire n_5666;
wire n_9195;
wire n_10442;
wire n_16236;
wire n_11687;
wire n_8870;
wire n_13973;
wire n_7150;
wire n_7155;
wire n_8252;
wire n_11774;
wire n_7283;
wire n_6475;
wire n_7015;
wire n_8507;
wire n_7699;
wire n_6314;
wire n_8415;
wire n_10632;
wire n_13206;
wire n_9623;
wire n_6103;
wire n_15951;
wire n_7249;
wire n_5546;
wire n_10713;
wire n_6394;
wire n_8781;
wire n_6964;
wire n_15939;
wire n_14102;
wire n_6680;
wire n_10954;
wire n_7985;
wire n_13637;
wire n_12267;
wire n_15803;
wire n_7432;
wire n_8365;
wire n_16036;
wire n_13978;
wire n_13941;
wire n_4532;
wire n_15339;
wire n_13439;
wire n_13780;
wire n_8893;
wire n_16152;
wire n_6372;
wire n_14133;
wire n_14433;
wire n_11329;
wire n_15904;
wire n_5994;
wire n_6495;
wire n_7194;
wire n_9516;
wire n_13241;
wire n_16027;
wire n_13187;
wire n_13162;
wire n_6752;
wire n_12768;
wire n_8976;
wire n_6426;
wire n_7505;
wire n_5626;
wire n_16047;
wire n_8025;
wire n_8502;
wire n_10165;
wire n_15059;
wire n_8244;
wire n_10130;
wire n_7612;
wire n_8156;
wire n_11661;
wire n_7494;
wire n_4353;
wire n_11120;
wire n_14923;
wire n_9222;
wire n_13031;
wire n_8435;
wire n_6350;
wire n_8882;
wire n_16391;
wire n_4787;
wire n_7736;
wire n_15949;
wire n_16040;
wire n_10622;
wire n_5633;
wire n_13661;
wire n_13155;
wire n_9546;
wire n_5664;
wire n_7589;
wire n_14259;
wire n_5921;
wire n_6797;
wire n_15673;
wire n_13410;
wire n_4537;
wire n_14012;
wire n_4346;
wire n_8759;
wire n_4351;
wire n_6159;
wire n_7177;
wire n_7814;
wire n_13066;
wire n_8660;
wire n_13360;
wire n_11296;
wire n_13665;
wire n_8479;
wire n_14214;
wire n_15558;
wire n_13770;
wire n_12993;
wire n_13124;
wire n_6054;
wire n_11095;
wire n_11314;
wire n_8723;
wire n_13511;
wire n_11019;
wire n_8606;
wire n_9663;
wire n_7843;
wire n_6235;
wire n_15678;
wire n_8235;
wire n_13083;
wire n_12647;
wire n_7662;
wire n_16164;
wire n_4784;
wire n_16584;
wire n_6152;
wire n_16444;
wire n_15340;
wire n_16061;
wire n_9820;
wire n_14569;
wire n_7773;
wire n_7902;
wire n_5340;
wire n_14071;
wire n_9743;
wire n_6496;
wire n_15744;
wire n_7756;
wire n_12749;
wire n_15557;
wire n_8342;
wire n_8940;
wire n_13048;
wire n_11584;
wire n_5280;
wire n_8448;
wire n_13563;
wire n_8472;
wire n_7700;
wire n_4451;
wire n_14169;
wire n_4332;
wire n_7555;
wire n_10000;
wire n_4538;
wire n_4506;
wire n_10158;
wire n_12812;
wire n_10582;
wire n_12066;
wire n_16151;
wire n_10427;
wire n_11816;
wire n_12060;
wire n_10199;
wire n_7988;
wire n_8658;
wire n_14174;
wire n_6513;
wire n_7500;
wire n_10246;
wire n_11910;
wire n_15377;
wire n_16420;
wire n_11693;
wire n_15583;
wire n_15429;
wire n_13347;
wire n_15908;
wire n_14269;
wire n_5925;
wire n_9248;
wire n_6138;
wire n_5369;
wire n_8061;
wire n_8866;
wire n_9822;
wire n_10835;
wire n_5730;
wire n_11411;
wire n_5576;
wire n_11184;
wire n_13991;
wire n_13823;
wire n_11386;
wire n_11945;
wire n_11604;
wire n_14821;
wire n_13323;
wire n_12164;
wire n_15096;
wire n_16623;
wire n_5272;
wire n_11368;
wire n_14992;
wire n_10125;
wire n_12824;
wire n_13111;
wire n_13434;
wire n_6330;
wire n_15563;
wire n_16680;
wire n_10117;
wire n_9065;
wire n_12716;
wire n_10844;
wire n_16341;
wire n_16679;
wire n_16637;
wire n_14153;
wire n_8457;
wire n_6802;
wire n_13456;
wire n_10654;
wire n_9153;
wire n_9086;
wire n_10505;
wire n_9339;
wire n_10198;
wire n_6909;
wire n_7157;
wire n_11064;
wire n_13237;
wire n_6908;
wire n_14312;
wire n_8237;
wire n_13445;
wire n_15448;
wire n_7411;
wire n_9601;
wire n_9093;
wire n_15045;
wire n_11409;
wire n_4336;
wire n_7266;
wire n_15760;
wire n_8046;
wire n_14746;
wire n_7871;
wire n_5646;
wire n_12051;
wire n_11097;
wire n_13284;
wire n_12437;
wire n_5624;
wire n_4852;
wire n_4981;
wire n_10840;
wire n_12052;
wire n_6477;
wire n_9746;
wire n_14606;
wire n_6263;
wire n_10515;
wire n_8073;
wire n_15501;
wire n_5440;
wire n_6490;
wire n_15751;
wire n_16521;
wire n_15298;
wire n_11533;
wire n_11605;
wire n_8652;
wire n_9198;
wire n_8821;
wire n_7198;
wire n_8335;
wire n_9904;
wire n_10242;
wire n_9142;
wire n_9440;
wire n_10144;
wire n_9684;
wire n_15741;
wire n_16195;
wire n_6184;
wire n_14793;
wire n_5817;
wire n_15820;
wire n_5214;
wire n_15486;
wire n_10973;
wire n_13472;
wire n_4936;
wire n_15596;
wire n_9493;
wire n_4763;
wire n_15475;
wire n_5586;
wire n_11036;
wire n_8663;
wire n_11330;
wire n_12720;
wire n_4463;
wire n_7794;
wire n_10267;
wire n_6038;
wire n_10551;
wire n_13318;
wire n_15379;
wire n_5861;
wire n_10553;
wire n_16272;
wire n_15917;
wire n_13127;
wire n_14884;
wire n_8309;
wire n_5258;
wire n_8945;
wire n_11002;
wire n_6605;
wire n_15121;
wire n_12687;
wire n_5032;
wire n_8964;
wire n_10988;
wire n_14075;
wire n_9032;
wire n_9814;
wire n_16629;
wire n_6313;
wire n_16184;
wire n_4804;
wire n_6112;
wire n_5619;
wire n_16192;
wire n_13208;
wire n_7145;
wire n_9041;
wire n_13867;
wire n_15594;
wire n_5859;
wire n_12325;
wire n_14423;
wire n_16280;
wire n_16414;
wire n_5380;
wire n_4500;
wire n_9245;
wire n_5065;
wire n_13443;
wire n_5776;
wire n_8166;
wire n_4433;
wire n_5606;
wire n_9357;
wire n_5644;
wire n_11796;
wire n_14626;
wire n_5826;
wire n_15766;
wire n_10108;
wire n_8960;
wire n_13865;
wire n_12789;
wire n_5920;
wire n_10307;
wire n_5030;
wire n_14530;
wire n_15402;
wire n_7994;
wire n_14206;
wire n_4703;
wire n_8443;
wire n_7349;
wire n_9598;
wire n_8215;
wire n_7715;
wire n_6180;
wire n_8683;
wire n_14481;
wire n_8809;
wire n_5683;
wire n_6349;
wire n_10510;
wire n_15044;
wire n_12127;
wire n_12504;
wire n_12382;
wire n_5756;
wire n_15306;
wire n_12602;
wire n_5527;
wire n_6476;
wire n_8037;
wire n_13673;
wire n_12062;
wire n_14119;
wire n_15981;
wire n_15375;
wire n_12573;
wire n_16100;

CKINVDCx5p33_ASAP7_75t_R g4322 ( 
.A(n_220),
.Y(n_4322)
);

BUFx10_ASAP7_75t_L g4323 ( 
.A(n_4221),
.Y(n_4323)
);

CKINVDCx5p33_ASAP7_75t_R g4324 ( 
.A(n_4172),
.Y(n_4324)
);

CKINVDCx5p33_ASAP7_75t_R g4325 ( 
.A(n_1399),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4294),
.Y(n_4326)
);

CKINVDCx20_ASAP7_75t_R g4327 ( 
.A(n_4213),
.Y(n_4327)
);

CKINVDCx5p33_ASAP7_75t_R g4328 ( 
.A(n_1507),
.Y(n_4328)
);

HB1xp67_ASAP7_75t_L g4329 ( 
.A(n_2699),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_222),
.Y(n_4330)
);

BUFx10_ASAP7_75t_L g4331 ( 
.A(n_603),
.Y(n_4331)
);

CKINVDCx5p33_ASAP7_75t_R g4332 ( 
.A(n_731),
.Y(n_4332)
);

CKINVDCx5p33_ASAP7_75t_R g4333 ( 
.A(n_1531),
.Y(n_4333)
);

CKINVDCx5p33_ASAP7_75t_R g4334 ( 
.A(n_4059),
.Y(n_4334)
);

HB1xp67_ASAP7_75t_L g4335 ( 
.A(n_214),
.Y(n_4335)
);

INVx1_ASAP7_75t_L g4336 ( 
.A(n_1326),
.Y(n_4336)
);

CKINVDCx5p33_ASAP7_75t_R g4337 ( 
.A(n_1274),
.Y(n_4337)
);

CKINVDCx5p33_ASAP7_75t_R g4338 ( 
.A(n_1088),
.Y(n_4338)
);

CKINVDCx5p33_ASAP7_75t_R g4339 ( 
.A(n_2664),
.Y(n_4339)
);

CKINVDCx5p33_ASAP7_75t_R g4340 ( 
.A(n_3796),
.Y(n_4340)
);

INVx1_ASAP7_75t_SL g4341 ( 
.A(n_4115),
.Y(n_4341)
);

CKINVDCx5p33_ASAP7_75t_R g4342 ( 
.A(n_1407),
.Y(n_4342)
);

CKINVDCx5p33_ASAP7_75t_R g4343 ( 
.A(n_1704),
.Y(n_4343)
);

CKINVDCx5p33_ASAP7_75t_R g4344 ( 
.A(n_2650),
.Y(n_4344)
);

BUFx10_ASAP7_75t_L g4345 ( 
.A(n_2239),
.Y(n_4345)
);

CKINVDCx5p33_ASAP7_75t_R g4346 ( 
.A(n_4217),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_4150),
.Y(n_4347)
);

CKINVDCx5p33_ASAP7_75t_R g4348 ( 
.A(n_917),
.Y(n_4348)
);

CKINVDCx5p33_ASAP7_75t_R g4349 ( 
.A(n_1930),
.Y(n_4349)
);

INVx1_ASAP7_75t_L g4350 ( 
.A(n_3526),
.Y(n_4350)
);

CKINVDCx5p33_ASAP7_75t_R g4351 ( 
.A(n_1156),
.Y(n_4351)
);

INVx1_ASAP7_75t_L g4352 ( 
.A(n_3807),
.Y(n_4352)
);

CKINVDCx20_ASAP7_75t_R g4353 ( 
.A(n_3101),
.Y(n_4353)
);

CKINVDCx5p33_ASAP7_75t_R g4354 ( 
.A(n_734),
.Y(n_4354)
);

CKINVDCx5p33_ASAP7_75t_R g4355 ( 
.A(n_2673),
.Y(n_4355)
);

CKINVDCx5p33_ASAP7_75t_R g4356 ( 
.A(n_2194),
.Y(n_4356)
);

BUFx3_ASAP7_75t_L g4357 ( 
.A(n_4158),
.Y(n_4357)
);

INVx2_ASAP7_75t_L g4358 ( 
.A(n_3265),
.Y(n_4358)
);

CKINVDCx5p33_ASAP7_75t_R g4359 ( 
.A(n_649),
.Y(n_4359)
);

CKINVDCx5p33_ASAP7_75t_R g4360 ( 
.A(n_1418),
.Y(n_4360)
);

CKINVDCx5p33_ASAP7_75t_R g4361 ( 
.A(n_1287),
.Y(n_4361)
);

INVx1_ASAP7_75t_SL g4362 ( 
.A(n_3950),
.Y(n_4362)
);

INVx2_ASAP7_75t_L g4363 ( 
.A(n_1702),
.Y(n_4363)
);

CKINVDCx5p33_ASAP7_75t_R g4364 ( 
.A(n_2680),
.Y(n_4364)
);

CKINVDCx5p33_ASAP7_75t_R g4365 ( 
.A(n_2695),
.Y(n_4365)
);

CKINVDCx5p33_ASAP7_75t_R g4366 ( 
.A(n_2291),
.Y(n_4366)
);

CKINVDCx5p33_ASAP7_75t_R g4367 ( 
.A(n_3398),
.Y(n_4367)
);

INVx2_ASAP7_75t_L g4368 ( 
.A(n_189),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_1139),
.Y(n_4369)
);

CKINVDCx5p33_ASAP7_75t_R g4370 ( 
.A(n_508),
.Y(n_4370)
);

CKINVDCx5p33_ASAP7_75t_R g4371 ( 
.A(n_3480),
.Y(n_4371)
);

CKINVDCx5p33_ASAP7_75t_R g4372 ( 
.A(n_3252),
.Y(n_4372)
);

CKINVDCx5p33_ASAP7_75t_R g4373 ( 
.A(n_3796),
.Y(n_4373)
);

CKINVDCx5p33_ASAP7_75t_R g4374 ( 
.A(n_4170),
.Y(n_4374)
);

CKINVDCx5p33_ASAP7_75t_R g4375 ( 
.A(n_373),
.Y(n_4375)
);

CKINVDCx20_ASAP7_75t_R g4376 ( 
.A(n_1813),
.Y(n_4376)
);

HB1xp67_ASAP7_75t_L g4377 ( 
.A(n_3826),
.Y(n_4377)
);

CKINVDCx20_ASAP7_75t_R g4378 ( 
.A(n_2192),
.Y(n_4378)
);

CKINVDCx5p33_ASAP7_75t_R g4379 ( 
.A(n_3173),
.Y(n_4379)
);

CKINVDCx5p33_ASAP7_75t_R g4380 ( 
.A(n_527),
.Y(n_4380)
);

INVx1_ASAP7_75t_L g4381 ( 
.A(n_3369),
.Y(n_4381)
);

BUFx10_ASAP7_75t_L g4382 ( 
.A(n_2360),
.Y(n_4382)
);

CKINVDCx5p33_ASAP7_75t_R g4383 ( 
.A(n_4174),
.Y(n_4383)
);

CKINVDCx20_ASAP7_75t_R g4384 ( 
.A(n_1982),
.Y(n_4384)
);

INVx1_ASAP7_75t_L g4385 ( 
.A(n_4145),
.Y(n_4385)
);

CKINVDCx5p33_ASAP7_75t_R g4386 ( 
.A(n_804),
.Y(n_4386)
);

CKINVDCx5p33_ASAP7_75t_R g4387 ( 
.A(n_701),
.Y(n_4387)
);

CKINVDCx5p33_ASAP7_75t_R g4388 ( 
.A(n_4051),
.Y(n_4388)
);

INVx1_ASAP7_75t_L g4389 ( 
.A(n_4216),
.Y(n_4389)
);

CKINVDCx16_ASAP7_75t_R g4390 ( 
.A(n_1244),
.Y(n_4390)
);

CKINVDCx5p33_ASAP7_75t_R g4391 ( 
.A(n_3226),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_3148),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_3474),
.Y(n_4393)
);

CKINVDCx5p33_ASAP7_75t_R g4394 ( 
.A(n_652),
.Y(n_4394)
);

CKINVDCx5p33_ASAP7_75t_R g4395 ( 
.A(n_1173),
.Y(n_4395)
);

INVx1_ASAP7_75t_L g4396 ( 
.A(n_1202),
.Y(n_4396)
);

CKINVDCx16_ASAP7_75t_R g4397 ( 
.A(n_3288),
.Y(n_4397)
);

CKINVDCx5p33_ASAP7_75t_R g4398 ( 
.A(n_1462),
.Y(n_4398)
);

CKINVDCx5p33_ASAP7_75t_R g4399 ( 
.A(n_4215),
.Y(n_4399)
);

CKINVDCx5p33_ASAP7_75t_R g4400 ( 
.A(n_1310),
.Y(n_4400)
);

CKINVDCx5p33_ASAP7_75t_R g4401 ( 
.A(n_3533),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_1139),
.Y(n_4402)
);

BUFx6f_ASAP7_75t_L g4403 ( 
.A(n_4127),
.Y(n_4403)
);

CKINVDCx5p33_ASAP7_75t_R g4404 ( 
.A(n_4164),
.Y(n_4404)
);

CKINVDCx5p33_ASAP7_75t_R g4405 ( 
.A(n_105),
.Y(n_4405)
);

INVx1_ASAP7_75t_L g4406 ( 
.A(n_1379),
.Y(n_4406)
);

CKINVDCx5p33_ASAP7_75t_R g4407 ( 
.A(n_2371),
.Y(n_4407)
);

CKINVDCx5p33_ASAP7_75t_R g4408 ( 
.A(n_4),
.Y(n_4408)
);

INVx1_ASAP7_75t_L g4409 ( 
.A(n_2216),
.Y(n_4409)
);

CKINVDCx5p33_ASAP7_75t_R g4410 ( 
.A(n_1176),
.Y(n_4410)
);

CKINVDCx5p33_ASAP7_75t_R g4411 ( 
.A(n_1989),
.Y(n_4411)
);

CKINVDCx5p33_ASAP7_75t_R g4412 ( 
.A(n_1345),
.Y(n_4412)
);

INVx2_ASAP7_75t_L g4413 ( 
.A(n_2164),
.Y(n_4413)
);

CKINVDCx20_ASAP7_75t_R g4414 ( 
.A(n_2918),
.Y(n_4414)
);

CKINVDCx20_ASAP7_75t_R g4415 ( 
.A(n_4243),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_3081),
.Y(n_4416)
);

CKINVDCx20_ASAP7_75t_R g4417 ( 
.A(n_4063),
.Y(n_4417)
);

CKINVDCx16_ASAP7_75t_R g4418 ( 
.A(n_3983),
.Y(n_4418)
);

CKINVDCx5p33_ASAP7_75t_R g4419 ( 
.A(n_3988),
.Y(n_4419)
);

INVx2_ASAP7_75t_SL g4420 ( 
.A(n_1364),
.Y(n_4420)
);

INVx1_ASAP7_75t_L g4421 ( 
.A(n_1663),
.Y(n_4421)
);

CKINVDCx5p33_ASAP7_75t_R g4422 ( 
.A(n_3765),
.Y(n_4422)
);

CKINVDCx5p33_ASAP7_75t_R g4423 ( 
.A(n_822),
.Y(n_4423)
);

INVx1_ASAP7_75t_L g4424 ( 
.A(n_1008),
.Y(n_4424)
);

CKINVDCx5p33_ASAP7_75t_R g4425 ( 
.A(n_2581),
.Y(n_4425)
);

INVx1_ASAP7_75t_L g4426 ( 
.A(n_3005),
.Y(n_4426)
);

INVx1_ASAP7_75t_L g4427 ( 
.A(n_3018),
.Y(n_4427)
);

INVx1_ASAP7_75t_L g4428 ( 
.A(n_1376),
.Y(n_4428)
);

CKINVDCx5p33_ASAP7_75t_R g4429 ( 
.A(n_3940),
.Y(n_4429)
);

CKINVDCx5p33_ASAP7_75t_R g4430 ( 
.A(n_3428),
.Y(n_4430)
);

CKINVDCx5p33_ASAP7_75t_R g4431 ( 
.A(n_2359),
.Y(n_4431)
);

CKINVDCx5p33_ASAP7_75t_R g4432 ( 
.A(n_4075),
.Y(n_4432)
);

INVx1_ASAP7_75t_L g4433 ( 
.A(n_2060),
.Y(n_4433)
);

BUFx10_ASAP7_75t_L g4434 ( 
.A(n_4096),
.Y(n_4434)
);

CKINVDCx5p33_ASAP7_75t_R g4435 ( 
.A(n_3996),
.Y(n_4435)
);

CKINVDCx5p33_ASAP7_75t_R g4436 ( 
.A(n_4102),
.Y(n_4436)
);

INVxp67_ASAP7_75t_L g4437 ( 
.A(n_2748),
.Y(n_4437)
);

INVx1_ASAP7_75t_L g4438 ( 
.A(n_1757),
.Y(n_4438)
);

INVx1_ASAP7_75t_L g4439 ( 
.A(n_3713),
.Y(n_4439)
);

CKINVDCx5p33_ASAP7_75t_R g4440 ( 
.A(n_1088),
.Y(n_4440)
);

CKINVDCx5p33_ASAP7_75t_R g4441 ( 
.A(n_1934),
.Y(n_4441)
);

CKINVDCx5p33_ASAP7_75t_R g4442 ( 
.A(n_3260),
.Y(n_4442)
);

CKINVDCx5p33_ASAP7_75t_R g4443 ( 
.A(n_4311),
.Y(n_4443)
);

INVx1_ASAP7_75t_L g4444 ( 
.A(n_3571),
.Y(n_4444)
);

INVx1_ASAP7_75t_L g4445 ( 
.A(n_3398),
.Y(n_4445)
);

CKINVDCx5p33_ASAP7_75t_R g4446 ( 
.A(n_4176),
.Y(n_4446)
);

INVx2_ASAP7_75t_SL g4447 ( 
.A(n_3123),
.Y(n_4447)
);

INVx1_ASAP7_75t_L g4448 ( 
.A(n_1864),
.Y(n_4448)
);

CKINVDCx5p33_ASAP7_75t_R g4449 ( 
.A(n_4121),
.Y(n_4449)
);

CKINVDCx5p33_ASAP7_75t_R g4450 ( 
.A(n_1227),
.Y(n_4450)
);

CKINVDCx5p33_ASAP7_75t_R g4451 ( 
.A(n_2094),
.Y(n_4451)
);

CKINVDCx5p33_ASAP7_75t_R g4452 ( 
.A(n_4101),
.Y(n_4452)
);

CKINVDCx5p33_ASAP7_75t_R g4453 ( 
.A(n_2077),
.Y(n_4453)
);

INVx1_ASAP7_75t_L g4454 ( 
.A(n_1255),
.Y(n_4454)
);

INVx2_ASAP7_75t_SL g4455 ( 
.A(n_4189),
.Y(n_4455)
);

INVx2_ASAP7_75t_L g4456 ( 
.A(n_1779),
.Y(n_4456)
);

INVx1_ASAP7_75t_L g4457 ( 
.A(n_2037),
.Y(n_4457)
);

INVx1_ASAP7_75t_L g4458 ( 
.A(n_3557),
.Y(n_4458)
);

CKINVDCx5p33_ASAP7_75t_R g4459 ( 
.A(n_2873),
.Y(n_4459)
);

INVx1_ASAP7_75t_L g4460 ( 
.A(n_4111),
.Y(n_4460)
);

INVx1_ASAP7_75t_L g4461 ( 
.A(n_3808),
.Y(n_4461)
);

CKINVDCx5p33_ASAP7_75t_R g4462 ( 
.A(n_1820),
.Y(n_4462)
);

CKINVDCx5p33_ASAP7_75t_R g4463 ( 
.A(n_2820),
.Y(n_4463)
);

CKINVDCx20_ASAP7_75t_R g4464 ( 
.A(n_2914),
.Y(n_4464)
);

CKINVDCx5p33_ASAP7_75t_R g4465 ( 
.A(n_103),
.Y(n_4465)
);

CKINVDCx5p33_ASAP7_75t_R g4466 ( 
.A(n_4018),
.Y(n_4466)
);

CKINVDCx5p33_ASAP7_75t_R g4467 ( 
.A(n_1359),
.Y(n_4467)
);

CKINVDCx5p33_ASAP7_75t_R g4468 ( 
.A(n_1638),
.Y(n_4468)
);

CKINVDCx20_ASAP7_75t_R g4469 ( 
.A(n_1983),
.Y(n_4469)
);

BUFx10_ASAP7_75t_L g4470 ( 
.A(n_30),
.Y(n_4470)
);

CKINVDCx5p33_ASAP7_75t_R g4471 ( 
.A(n_2967),
.Y(n_4471)
);

CKINVDCx5p33_ASAP7_75t_R g4472 ( 
.A(n_1535),
.Y(n_4472)
);

CKINVDCx5p33_ASAP7_75t_R g4473 ( 
.A(n_1558),
.Y(n_4473)
);

CKINVDCx5p33_ASAP7_75t_R g4474 ( 
.A(n_2623),
.Y(n_4474)
);

CKINVDCx5p33_ASAP7_75t_R g4475 ( 
.A(n_1052),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_4105),
.Y(n_4476)
);

CKINVDCx5p33_ASAP7_75t_R g4477 ( 
.A(n_2803),
.Y(n_4477)
);

CKINVDCx5p33_ASAP7_75t_R g4478 ( 
.A(n_514),
.Y(n_4478)
);

INVx2_ASAP7_75t_L g4479 ( 
.A(n_2457),
.Y(n_4479)
);

CKINVDCx5p33_ASAP7_75t_R g4480 ( 
.A(n_689),
.Y(n_4480)
);

CKINVDCx5p33_ASAP7_75t_R g4481 ( 
.A(n_1317),
.Y(n_4481)
);

CKINVDCx5p33_ASAP7_75t_R g4482 ( 
.A(n_4278),
.Y(n_4482)
);

CKINVDCx5p33_ASAP7_75t_R g4483 ( 
.A(n_1435),
.Y(n_4483)
);

BUFx8_ASAP7_75t_SL g4484 ( 
.A(n_3157),
.Y(n_4484)
);

CKINVDCx5p33_ASAP7_75t_R g4485 ( 
.A(n_1172),
.Y(n_4485)
);

BUFx3_ASAP7_75t_L g4486 ( 
.A(n_4198),
.Y(n_4486)
);

CKINVDCx5p33_ASAP7_75t_R g4487 ( 
.A(n_216),
.Y(n_4487)
);

BUFx2_ASAP7_75t_L g4488 ( 
.A(n_1967),
.Y(n_4488)
);

CKINVDCx5p33_ASAP7_75t_R g4489 ( 
.A(n_2529),
.Y(n_4489)
);

INVx1_ASAP7_75t_L g4490 ( 
.A(n_1953),
.Y(n_4490)
);

CKINVDCx5p33_ASAP7_75t_R g4491 ( 
.A(n_501),
.Y(n_4491)
);

CKINVDCx5p33_ASAP7_75t_R g4492 ( 
.A(n_4109),
.Y(n_4492)
);

CKINVDCx20_ASAP7_75t_R g4493 ( 
.A(n_3069),
.Y(n_4493)
);

CKINVDCx5p33_ASAP7_75t_R g4494 ( 
.A(n_909),
.Y(n_4494)
);

INVx1_ASAP7_75t_L g4495 ( 
.A(n_1820),
.Y(n_4495)
);

CKINVDCx5p33_ASAP7_75t_R g4496 ( 
.A(n_294),
.Y(n_4496)
);

INVx2_ASAP7_75t_SL g4497 ( 
.A(n_1076),
.Y(n_4497)
);

INVx1_ASAP7_75t_L g4498 ( 
.A(n_3407),
.Y(n_4498)
);

CKINVDCx5p33_ASAP7_75t_R g4499 ( 
.A(n_4005),
.Y(n_4499)
);

CKINVDCx5p33_ASAP7_75t_R g4500 ( 
.A(n_2671),
.Y(n_4500)
);

CKINVDCx16_ASAP7_75t_R g4501 ( 
.A(n_1320),
.Y(n_4501)
);

INVx3_ASAP7_75t_L g4502 ( 
.A(n_251),
.Y(n_4502)
);

CKINVDCx5p33_ASAP7_75t_R g4503 ( 
.A(n_1729),
.Y(n_4503)
);

CKINVDCx5p33_ASAP7_75t_R g4504 ( 
.A(n_2753),
.Y(n_4504)
);

CKINVDCx5p33_ASAP7_75t_R g4505 ( 
.A(n_1642),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_1441),
.Y(n_4506)
);

CKINVDCx20_ASAP7_75t_R g4507 ( 
.A(n_3087),
.Y(n_4507)
);

INVx2_ASAP7_75t_L g4508 ( 
.A(n_45),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_2311),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_2164),
.Y(n_4510)
);

HB1xp67_ASAP7_75t_L g4511 ( 
.A(n_2541),
.Y(n_4511)
);

CKINVDCx5p33_ASAP7_75t_R g4512 ( 
.A(n_3143),
.Y(n_4512)
);

CKINVDCx5p33_ASAP7_75t_R g4513 ( 
.A(n_1845),
.Y(n_4513)
);

CKINVDCx5p33_ASAP7_75t_R g4514 ( 
.A(n_3835),
.Y(n_4514)
);

BUFx2_ASAP7_75t_L g4515 ( 
.A(n_1242),
.Y(n_4515)
);

INVx1_ASAP7_75t_L g4516 ( 
.A(n_2659),
.Y(n_4516)
);

INVx1_ASAP7_75t_L g4517 ( 
.A(n_1069),
.Y(n_4517)
);

INVx1_ASAP7_75t_L g4518 ( 
.A(n_2338),
.Y(n_4518)
);

INVx1_ASAP7_75t_L g4519 ( 
.A(n_2394),
.Y(n_4519)
);

INVx1_ASAP7_75t_L g4520 ( 
.A(n_1733),
.Y(n_4520)
);

CKINVDCx5p33_ASAP7_75t_R g4521 ( 
.A(n_1485),
.Y(n_4521)
);

CKINVDCx5p33_ASAP7_75t_R g4522 ( 
.A(n_4098),
.Y(n_4522)
);

CKINVDCx5p33_ASAP7_75t_R g4523 ( 
.A(n_1631),
.Y(n_4523)
);

CKINVDCx5p33_ASAP7_75t_R g4524 ( 
.A(n_645),
.Y(n_4524)
);

INVxp67_ASAP7_75t_SL g4525 ( 
.A(n_4116),
.Y(n_4525)
);

CKINVDCx20_ASAP7_75t_R g4526 ( 
.A(n_1172),
.Y(n_4526)
);

INVx1_ASAP7_75t_L g4527 ( 
.A(n_1683),
.Y(n_4527)
);

INVx1_ASAP7_75t_L g4528 ( 
.A(n_3094),
.Y(n_4528)
);

BUFx3_ASAP7_75t_L g4529 ( 
.A(n_1394),
.Y(n_4529)
);

CKINVDCx5p33_ASAP7_75t_R g4530 ( 
.A(n_3093),
.Y(n_4530)
);

CKINVDCx5p33_ASAP7_75t_R g4531 ( 
.A(n_4015),
.Y(n_4531)
);

INVx2_ASAP7_75t_SL g4532 ( 
.A(n_724),
.Y(n_4532)
);

INVx1_ASAP7_75t_L g4533 ( 
.A(n_3310),
.Y(n_4533)
);

CKINVDCx5p33_ASAP7_75t_R g4534 ( 
.A(n_1518),
.Y(n_4534)
);

CKINVDCx5p33_ASAP7_75t_R g4535 ( 
.A(n_4160),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_509),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_2937),
.Y(n_4537)
);

CKINVDCx5p33_ASAP7_75t_R g4538 ( 
.A(n_4193),
.Y(n_4538)
);

INVx1_ASAP7_75t_L g4539 ( 
.A(n_2334),
.Y(n_4539)
);

CKINVDCx5p33_ASAP7_75t_R g4540 ( 
.A(n_435),
.Y(n_4540)
);

CKINVDCx5p33_ASAP7_75t_R g4541 ( 
.A(n_4088),
.Y(n_4541)
);

CKINVDCx5p33_ASAP7_75t_R g4542 ( 
.A(n_1456),
.Y(n_4542)
);

INVx1_ASAP7_75t_L g4543 ( 
.A(n_2039),
.Y(n_4543)
);

CKINVDCx5p33_ASAP7_75t_R g4544 ( 
.A(n_172),
.Y(n_4544)
);

CKINVDCx5p33_ASAP7_75t_R g4545 ( 
.A(n_798),
.Y(n_4545)
);

INVx1_ASAP7_75t_L g4546 ( 
.A(n_4177),
.Y(n_4546)
);

BUFx2_ASAP7_75t_L g4547 ( 
.A(n_321),
.Y(n_4547)
);

BUFx10_ASAP7_75t_L g4548 ( 
.A(n_619),
.Y(n_4548)
);

INVx2_ASAP7_75t_L g4549 ( 
.A(n_227),
.Y(n_4549)
);

CKINVDCx5p33_ASAP7_75t_R g4550 ( 
.A(n_2518),
.Y(n_4550)
);

BUFx6f_ASAP7_75t_L g4551 ( 
.A(n_2723),
.Y(n_4551)
);

CKINVDCx5p33_ASAP7_75t_R g4552 ( 
.A(n_521),
.Y(n_4552)
);

INVx1_ASAP7_75t_L g4553 ( 
.A(n_1671),
.Y(n_4553)
);

CKINVDCx5p33_ASAP7_75t_R g4554 ( 
.A(n_852),
.Y(n_4554)
);

INVx1_ASAP7_75t_L g4555 ( 
.A(n_1057),
.Y(n_4555)
);

INVxp67_ASAP7_75t_L g4556 ( 
.A(n_1159),
.Y(n_4556)
);

CKINVDCx5p33_ASAP7_75t_R g4557 ( 
.A(n_4155),
.Y(n_4557)
);

INVx1_ASAP7_75t_L g4558 ( 
.A(n_2900),
.Y(n_4558)
);

BUFx3_ASAP7_75t_L g4559 ( 
.A(n_2701),
.Y(n_4559)
);

INVx1_ASAP7_75t_L g4560 ( 
.A(n_3882),
.Y(n_4560)
);

CKINVDCx5p33_ASAP7_75t_R g4561 ( 
.A(n_4095),
.Y(n_4561)
);

CKINVDCx5p33_ASAP7_75t_R g4562 ( 
.A(n_2730),
.Y(n_4562)
);

CKINVDCx5p33_ASAP7_75t_R g4563 ( 
.A(n_925),
.Y(n_4563)
);

CKINVDCx5p33_ASAP7_75t_R g4564 ( 
.A(n_4227),
.Y(n_4564)
);

CKINVDCx20_ASAP7_75t_R g4565 ( 
.A(n_4241),
.Y(n_4565)
);

CKINVDCx5p33_ASAP7_75t_R g4566 ( 
.A(n_1738),
.Y(n_4566)
);

BUFx5_ASAP7_75t_L g4567 ( 
.A(n_2897),
.Y(n_4567)
);

CKINVDCx20_ASAP7_75t_R g4568 ( 
.A(n_883),
.Y(n_4568)
);

CKINVDCx5p33_ASAP7_75t_R g4569 ( 
.A(n_3504),
.Y(n_4569)
);

CKINVDCx5p33_ASAP7_75t_R g4570 ( 
.A(n_2155),
.Y(n_4570)
);

CKINVDCx5p33_ASAP7_75t_R g4571 ( 
.A(n_4162),
.Y(n_4571)
);

CKINVDCx20_ASAP7_75t_R g4572 ( 
.A(n_1024),
.Y(n_4572)
);

CKINVDCx5p33_ASAP7_75t_R g4573 ( 
.A(n_428),
.Y(n_4573)
);

CKINVDCx5p33_ASAP7_75t_R g4574 ( 
.A(n_2618),
.Y(n_4574)
);

INVx1_ASAP7_75t_L g4575 ( 
.A(n_1074),
.Y(n_4575)
);

CKINVDCx20_ASAP7_75t_R g4576 ( 
.A(n_3843),
.Y(n_4576)
);

CKINVDCx5p33_ASAP7_75t_R g4577 ( 
.A(n_889),
.Y(n_4577)
);

INVx1_ASAP7_75t_L g4578 ( 
.A(n_1352),
.Y(n_4578)
);

BUFx3_ASAP7_75t_L g4579 ( 
.A(n_2650),
.Y(n_4579)
);

INVx1_ASAP7_75t_L g4580 ( 
.A(n_1785),
.Y(n_4580)
);

CKINVDCx5p33_ASAP7_75t_R g4581 ( 
.A(n_1745),
.Y(n_4581)
);

CKINVDCx5p33_ASAP7_75t_R g4582 ( 
.A(n_2623),
.Y(n_4582)
);

BUFx3_ASAP7_75t_L g4583 ( 
.A(n_947),
.Y(n_4583)
);

CKINVDCx20_ASAP7_75t_R g4584 ( 
.A(n_541),
.Y(n_4584)
);

CKINVDCx5p33_ASAP7_75t_R g4585 ( 
.A(n_4139),
.Y(n_4585)
);

CKINVDCx5p33_ASAP7_75t_R g4586 ( 
.A(n_1730),
.Y(n_4586)
);

CKINVDCx5p33_ASAP7_75t_R g4587 ( 
.A(n_3835),
.Y(n_4587)
);

INVx1_ASAP7_75t_L g4588 ( 
.A(n_54),
.Y(n_4588)
);

CKINVDCx5p33_ASAP7_75t_R g4589 ( 
.A(n_2517),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_1298),
.Y(n_4590)
);

INVx1_ASAP7_75t_L g4591 ( 
.A(n_932),
.Y(n_4591)
);

CKINVDCx5p33_ASAP7_75t_R g4592 ( 
.A(n_2104),
.Y(n_4592)
);

CKINVDCx5p33_ASAP7_75t_R g4593 ( 
.A(n_50),
.Y(n_4593)
);

CKINVDCx5p33_ASAP7_75t_R g4594 ( 
.A(n_2868),
.Y(n_4594)
);

BUFx10_ASAP7_75t_L g4595 ( 
.A(n_4098),
.Y(n_4595)
);

CKINVDCx5p33_ASAP7_75t_R g4596 ( 
.A(n_3880),
.Y(n_4596)
);

CKINVDCx5p33_ASAP7_75t_R g4597 ( 
.A(n_909),
.Y(n_4597)
);

INVx1_ASAP7_75t_L g4598 ( 
.A(n_1957),
.Y(n_4598)
);

CKINVDCx5p33_ASAP7_75t_R g4599 ( 
.A(n_3657),
.Y(n_4599)
);

CKINVDCx5p33_ASAP7_75t_R g4600 ( 
.A(n_4092),
.Y(n_4600)
);

INVx2_ASAP7_75t_L g4601 ( 
.A(n_880),
.Y(n_4601)
);

CKINVDCx5p33_ASAP7_75t_R g4602 ( 
.A(n_396),
.Y(n_4602)
);

INVx1_ASAP7_75t_L g4603 ( 
.A(n_4295),
.Y(n_4603)
);

CKINVDCx5p33_ASAP7_75t_R g4604 ( 
.A(n_1231),
.Y(n_4604)
);

CKINVDCx5p33_ASAP7_75t_R g4605 ( 
.A(n_3064),
.Y(n_4605)
);

CKINVDCx5p33_ASAP7_75t_R g4606 ( 
.A(n_1776),
.Y(n_4606)
);

CKINVDCx5p33_ASAP7_75t_R g4607 ( 
.A(n_2512),
.Y(n_4607)
);

CKINVDCx5p33_ASAP7_75t_R g4608 ( 
.A(n_445),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_1664),
.Y(n_4609)
);

INVx1_ASAP7_75t_L g4610 ( 
.A(n_3070),
.Y(n_4610)
);

CKINVDCx5p33_ASAP7_75t_R g4611 ( 
.A(n_2693),
.Y(n_4611)
);

INVx1_ASAP7_75t_SL g4612 ( 
.A(n_4112),
.Y(n_4612)
);

CKINVDCx5p33_ASAP7_75t_R g4613 ( 
.A(n_2359),
.Y(n_4613)
);

CKINVDCx5p33_ASAP7_75t_R g4614 ( 
.A(n_1599),
.Y(n_4614)
);

CKINVDCx5p33_ASAP7_75t_R g4615 ( 
.A(n_2367),
.Y(n_4615)
);

INVx1_ASAP7_75t_L g4616 ( 
.A(n_2137),
.Y(n_4616)
);

INVx1_ASAP7_75t_L g4617 ( 
.A(n_1904),
.Y(n_4617)
);

CKINVDCx5p33_ASAP7_75t_R g4618 ( 
.A(n_180),
.Y(n_4618)
);

INVx1_ASAP7_75t_SL g4619 ( 
.A(n_3352),
.Y(n_4619)
);

CKINVDCx20_ASAP7_75t_R g4620 ( 
.A(n_2562),
.Y(n_4620)
);

CKINVDCx5p33_ASAP7_75t_R g4621 ( 
.A(n_1288),
.Y(n_4621)
);

CKINVDCx20_ASAP7_75t_R g4622 ( 
.A(n_3576),
.Y(n_4622)
);

INVx1_ASAP7_75t_L g4623 ( 
.A(n_2760),
.Y(n_4623)
);

HB1xp67_ASAP7_75t_L g4624 ( 
.A(n_660),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_3925),
.Y(n_4625)
);

CKINVDCx5p33_ASAP7_75t_R g4626 ( 
.A(n_195),
.Y(n_4626)
);

CKINVDCx5p33_ASAP7_75t_R g4627 ( 
.A(n_3530),
.Y(n_4627)
);

CKINVDCx20_ASAP7_75t_R g4628 ( 
.A(n_3227),
.Y(n_4628)
);

CKINVDCx5p33_ASAP7_75t_R g4629 ( 
.A(n_3355),
.Y(n_4629)
);

INVx2_ASAP7_75t_L g4630 ( 
.A(n_1947),
.Y(n_4630)
);

CKINVDCx5p33_ASAP7_75t_R g4631 ( 
.A(n_3040),
.Y(n_4631)
);

CKINVDCx5p33_ASAP7_75t_R g4632 ( 
.A(n_1),
.Y(n_4632)
);

INVx1_ASAP7_75t_L g4633 ( 
.A(n_2735),
.Y(n_4633)
);

INVx2_ASAP7_75t_L g4634 ( 
.A(n_2248),
.Y(n_4634)
);

INVx1_ASAP7_75t_L g4635 ( 
.A(n_1765),
.Y(n_4635)
);

CKINVDCx5p33_ASAP7_75t_R g4636 ( 
.A(n_314),
.Y(n_4636)
);

INVx1_ASAP7_75t_L g4637 ( 
.A(n_3191),
.Y(n_4637)
);

CKINVDCx5p33_ASAP7_75t_R g4638 ( 
.A(n_4208),
.Y(n_4638)
);

CKINVDCx5p33_ASAP7_75t_R g4639 ( 
.A(n_1153),
.Y(n_4639)
);

CKINVDCx5p33_ASAP7_75t_R g4640 ( 
.A(n_376),
.Y(n_4640)
);

CKINVDCx5p33_ASAP7_75t_R g4641 ( 
.A(n_4185),
.Y(n_4641)
);

INVx1_ASAP7_75t_L g4642 ( 
.A(n_4203),
.Y(n_4642)
);

CKINVDCx5p33_ASAP7_75t_R g4643 ( 
.A(n_4129),
.Y(n_4643)
);

CKINVDCx5p33_ASAP7_75t_R g4644 ( 
.A(n_4177),
.Y(n_4644)
);

INVx1_ASAP7_75t_SL g4645 ( 
.A(n_2610),
.Y(n_4645)
);

CKINVDCx5p33_ASAP7_75t_R g4646 ( 
.A(n_4183),
.Y(n_4646)
);

CKINVDCx5p33_ASAP7_75t_R g4647 ( 
.A(n_4168),
.Y(n_4647)
);

CKINVDCx5p33_ASAP7_75t_R g4648 ( 
.A(n_2554),
.Y(n_4648)
);

INVx1_ASAP7_75t_L g4649 ( 
.A(n_91),
.Y(n_4649)
);

CKINVDCx5p33_ASAP7_75t_R g4650 ( 
.A(n_280),
.Y(n_4650)
);

INVx2_ASAP7_75t_L g4651 ( 
.A(n_517),
.Y(n_4651)
);

CKINVDCx5p33_ASAP7_75t_R g4652 ( 
.A(n_697),
.Y(n_4652)
);

INVx1_ASAP7_75t_L g4653 ( 
.A(n_294),
.Y(n_4653)
);

CKINVDCx5p33_ASAP7_75t_R g4654 ( 
.A(n_1079),
.Y(n_4654)
);

CKINVDCx5p33_ASAP7_75t_R g4655 ( 
.A(n_3857),
.Y(n_4655)
);

CKINVDCx5p33_ASAP7_75t_R g4656 ( 
.A(n_1514),
.Y(n_4656)
);

CKINVDCx5p33_ASAP7_75t_R g4657 ( 
.A(n_3638),
.Y(n_4657)
);

CKINVDCx5p33_ASAP7_75t_R g4658 ( 
.A(n_3097),
.Y(n_4658)
);

INVx1_ASAP7_75t_L g4659 ( 
.A(n_2512),
.Y(n_4659)
);

CKINVDCx5p33_ASAP7_75t_R g4660 ( 
.A(n_1549),
.Y(n_4660)
);

INVx1_ASAP7_75t_L g4661 ( 
.A(n_4103),
.Y(n_4661)
);

CKINVDCx5p33_ASAP7_75t_R g4662 ( 
.A(n_1887),
.Y(n_4662)
);

CKINVDCx5p33_ASAP7_75t_R g4663 ( 
.A(n_2731),
.Y(n_4663)
);

INVx1_ASAP7_75t_L g4664 ( 
.A(n_2184),
.Y(n_4664)
);

CKINVDCx5p33_ASAP7_75t_R g4665 ( 
.A(n_1878),
.Y(n_4665)
);

CKINVDCx5p33_ASAP7_75t_R g4666 ( 
.A(n_992),
.Y(n_4666)
);

CKINVDCx5p33_ASAP7_75t_R g4667 ( 
.A(n_411),
.Y(n_4667)
);

CKINVDCx5p33_ASAP7_75t_R g4668 ( 
.A(n_2183),
.Y(n_4668)
);

HB1xp67_ASAP7_75t_L g4669 ( 
.A(n_3262),
.Y(n_4669)
);

INVx1_ASAP7_75t_L g4670 ( 
.A(n_1124),
.Y(n_4670)
);

CKINVDCx5p33_ASAP7_75t_R g4671 ( 
.A(n_554),
.Y(n_4671)
);

INVxp67_ASAP7_75t_L g4672 ( 
.A(n_266),
.Y(n_4672)
);

INVx1_ASAP7_75t_L g4673 ( 
.A(n_4194),
.Y(n_4673)
);

INVx1_ASAP7_75t_L g4674 ( 
.A(n_3289),
.Y(n_4674)
);

CKINVDCx5p33_ASAP7_75t_R g4675 ( 
.A(n_2398),
.Y(n_4675)
);

CKINVDCx5p33_ASAP7_75t_R g4676 ( 
.A(n_2342),
.Y(n_4676)
);

BUFx6f_ASAP7_75t_L g4677 ( 
.A(n_1890),
.Y(n_4677)
);

CKINVDCx5p33_ASAP7_75t_R g4678 ( 
.A(n_4236),
.Y(n_4678)
);

CKINVDCx5p33_ASAP7_75t_R g4679 ( 
.A(n_3005),
.Y(n_4679)
);

CKINVDCx5p33_ASAP7_75t_R g4680 ( 
.A(n_3863),
.Y(n_4680)
);

CKINVDCx5p33_ASAP7_75t_R g4681 ( 
.A(n_4082),
.Y(n_4681)
);

INVx1_ASAP7_75t_L g4682 ( 
.A(n_3023),
.Y(n_4682)
);

INVx1_ASAP7_75t_L g4683 ( 
.A(n_468),
.Y(n_4683)
);

CKINVDCx5p33_ASAP7_75t_R g4684 ( 
.A(n_3590),
.Y(n_4684)
);

BUFx2_ASAP7_75t_L g4685 ( 
.A(n_2274),
.Y(n_4685)
);

CKINVDCx5p33_ASAP7_75t_R g4686 ( 
.A(n_3096),
.Y(n_4686)
);

CKINVDCx20_ASAP7_75t_R g4687 ( 
.A(n_4071),
.Y(n_4687)
);

CKINVDCx5p33_ASAP7_75t_R g4688 ( 
.A(n_116),
.Y(n_4688)
);

INVx1_ASAP7_75t_L g4689 ( 
.A(n_74),
.Y(n_4689)
);

INVx1_ASAP7_75t_L g4690 ( 
.A(n_2708),
.Y(n_4690)
);

CKINVDCx20_ASAP7_75t_R g4691 ( 
.A(n_919),
.Y(n_4691)
);

CKINVDCx16_ASAP7_75t_R g4692 ( 
.A(n_520),
.Y(n_4692)
);

CKINVDCx5p33_ASAP7_75t_R g4693 ( 
.A(n_244),
.Y(n_4693)
);

INVx1_ASAP7_75t_L g4694 ( 
.A(n_2546),
.Y(n_4694)
);

INVx2_ASAP7_75t_L g4695 ( 
.A(n_4067),
.Y(n_4695)
);

CKINVDCx5p33_ASAP7_75t_R g4696 ( 
.A(n_572),
.Y(n_4696)
);

INVx1_ASAP7_75t_L g4697 ( 
.A(n_3225),
.Y(n_4697)
);

INVx1_ASAP7_75t_SL g4698 ( 
.A(n_4014),
.Y(n_4698)
);

CKINVDCx5p33_ASAP7_75t_R g4699 ( 
.A(n_3690),
.Y(n_4699)
);

CKINVDCx5p33_ASAP7_75t_R g4700 ( 
.A(n_3569),
.Y(n_4700)
);

CKINVDCx5p33_ASAP7_75t_R g4701 ( 
.A(n_3943),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_2966),
.Y(n_4702)
);

CKINVDCx5p33_ASAP7_75t_R g4703 ( 
.A(n_619),
.Y(n_4703)
);

CKINVDCx5p33_ASAP7_75t_R g4704 ( 
.A(n_4135),
.Y(n_4704)
);

CKINVDCx5p33_ASAP7_75t_R g4705 ( 
.A(n_3995),
.Y(n_4705)
);

INVxp67_ASAP7_75t_L g4706 ( 
.A(n_2795),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_1761),
.Y(n_4707)
);

INVx1_ASAP7_75t_L g4708 ( 
.A(n_2699),
.Y(n_4708)
);

CKINVDCx5p33_ASAP7_75t_R g4709 ( 
.A(n_1092),
.Y(n_4709)
);

CKINVDCx16_ASAP7_75t_R g4710 ( 
.A(n_2425),
.Y(n_4710)
);

INVx2_ASAP7_75t_L g4711 ( 
.A(n_3064),
.Y(n_4711)
);

INVx1_ASAP7_75t_L g4712 ( 
.A(n_597),
.Y(n_4712)
);

INVx2_ASAP7_75t_SL g4713 ( 
.A(n_3039),
.Y(n_4713)
);

CKINVDCx5p33_ASAP7_75t_R g4714 ( 
.A(n_3942),
.Y(n_4714)
);

INVx1_ASAP7_75t_L g4715 ( 
.A(n_2817),
.Y(n_4715)
);

CKINVDCx5p33_ASAP7_75t_R g4716 ( 
.A(n_4133),
.Y(n_4716)
);

CKINVDCx5p33_ASAP7_75t_R g4717 ( 
.A(n_3903),
.Y(n_4717)
);

CKINVDCx5p33_ASAP7_75t_R g4718 ( 
.A(n_4195),
.Y(n_4718)
);

CKINVDCx20_ASAP7_75t_R g4719 ( 
.A(n_1430),
.Y(n_4719)
);

BUFx10_ASAP7_75t_L g4720 ( 
.A(n_3336),
.Y(n_4720)
);

CKINVDCx5p33_ASAP7_75t_R g4721 ( 
.A(n_2959),
.Y(n_4721)
);

BUFx3_ASAP7_75t_L g4722 ( 
.A(n_665),
.Y(n_4722)
);

CKINVDCx5p33_ASAP7_75t_R g4723 ( 
.A(n_521),
.Y(n_4723)
);

INVx2_ASAP7_75t_L g4724 ( 
.A(n_4090),
.Y(n_4724)
);

CKINVDCx5p33_ASAP7_75t_R g4725 ( 
.A(n_2477),
.Y(n_4725)
);

CKINVDCx5p33_ASAP7_75t_R g4726 ( 
.A(n_4210),
.Y(n_4726)
);

BUFx8_ASAP7_75t_SL g4727 ( 
.A(n_4191),
.Y(n_4727)
);

INVx2_ASAP7_75t_SL g4728 ( 
.A(n_203),
.Y(n_4728)
);

CKINVDCx14_ASAP7_75t_R g4729 ( 
.A(n_2559),
.Y(n_4729)
);

CKINVDCx5p33_ASAP7_75t_R g4730 ( 
.A(n_2088),
.Y(n_4730)
);

INVx1_ASAP7_75t_L g4731 ( 
.A(n_2255),
.Y(n_4731)
);

CKINVDCx5p33_ASAP7_75t_R g4732 ( 
.A(n_1661),
.Y(n_4732)
);

CKINVDCx5p33_ASAP7_75t_R g4733 ( 
.A(n_4264),
.Y(n_4733)
);

CKINVDCx5p33_ASAP7_75t_R g4734 ( 
.A(n_4228),
.Y(n_4734)
);

CKINVDCx5p33_ASAP7_75t_R g4735 ( 
.A(n_2208),
.Y(n_4735)
);

CKINVDCx5p33_ASAP7_75t_R g4736 ( 
.A(n_4149),
.Y(n_4736)
);

CKINVDCx5p33_ASAP7_75t_R g4737 ( 
.A(n_2351),
.Y(n_4737)
);

INVx1_ASAP7_75t_L g4738 ( 
.A(n_2729),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_2638),
.Y(n_4739)
);

CKINVDCx5p33_ASAP7_75t_R g4740 ( 
.A(n_2144),
.Y(n_4740)
);

CKINVDCx5p33_ASAP7_75t_R g4741 ( 
.A(n_766),
.Y(n_4741)
);

INVx1_ASAP7_75t_L g4742 ( 
.A(n_1525),
.Y(n_4742)
);

CKINVDCx5p33_ASAP7_75t_R g4743 ( 
.A(n_217),
.Y(n_4743)
);

CKINVDCx5p33_ASAP7_75t_R g4744 ( 
.A(n_2826),
.Y(n_4744)
);

INVx2_ASAP7_75t_SL g4745 ( 
.A(n_4159),
.Y(n_4745)
);

INVx1_ASAP7_75t_L g4746 ( 
.A(n_143),
.Y(n_4746)
);

CKINVDCx5p33_ASAP7_75t_R g4747 ( 
.A(n_357),
.Y(n_4747)
);

CKINVDCx5p33_ASAP7_75t_R g4748 ( 
.A(n_3762),
.Y(n_4748)
);

INVx1_ASAP7_75t_L g4749 ( 
.A(n_1490),
.Y(n_4749)
);

BUFx10_ASAP7_75t_L g4750 ( 
.A(n_1062),
.Y(n_4750)
);

CKINVDCx5p33_ASAP7_75t_R g4751 ( 
.A(n_2885),
.Y(n_4751)
);

CKINVDCx14_ASAP7_75t_R g4752 ( 
.A(n_2127),
.Y(n_4752)
);

INVx1_ASAP7_75t_L g4753 ( 
.A(n_4036),
.Y(n_4753)
);

CKINVDCx5p33_ASAP7_75t_R g4754 ( 
.A(n_4192),
.Y(n_4754)
);

CKINVDCx5p33_ASAP7_75t_R g4755 ( 
.A(n_2184),
.Y(n_4755)
);

BUFx10_ASAP7_75t_L g4756 ( 
.A(n_638),
.Y(n_4756)
);

CKINVDCx5p33_ASAP7_75t_R g4757 ( 
.A(n_2475),
.Y(n_4757)
);

INVx1_ASAP7_75t_L g4758 ( 
.A(n_2967),
.Y(n_4758)
);

INVx1_ASAP7_75t_L g4759 ( 
.A(n_2913),
.Y(n_4759)
);

INVx1_ASAP7_75t_L g4760 ( 
.A(n_379),
.Y(n_4760)
);

CKINVDCx5p33_ASAP7_75t_R g4761 ( 
.A(n_2159),
.Y(n_4761)
);

BUFx10_ASAP7_75t_L g4762 ( 
.A(n_1748),
.Y(n_4762)
);

INVx1_ASAP7_75t_L g4763 ( 
.A(n_2442),
.Y(n_4763)
);

INVx2_ASAP7_75t_L g4764 ( 
.A(n_4247),
.Y(n_4764)
);

INVx1_ASAP7_75t_L g4765 ( 
.A(n_4142),
.Y(n_4765)
);

INVx2_ASAP7_75t_L g4766 ( 
.A(n_399),
.Y(n_4766)
);

INVx1_ASAP7_75t_SL g4767 ( 
.A(n_2117),
.Y(n_4767)
);

CKINVDCx5p33_ASAP7_75t_R g4768 ( 
.A(n_3711),
.Y(n_4768)
);

CKINVDCx5p33_ASAP7_75t_R g4769 ( 
.A(n_3057),
.Y(n_4769)
);

CKINVDCx5p33_ASAP7_75t_R g4770 ( 
.A(n_305),
.Y(n_4770)
);

INVx2_ASAP7_75t_L g4771 ( 
.A(n_1996),
.Y(n_4771)
);

INVx2_ASAP7_75t_SL g4772 ( 
.A(n_4052),
.Y(n_4772)
);

INVxp67_ASAP7_75t_L g4773 ( 
.A(n_1748),
.Y(n_4773)
);

CKINVDCx5p33_ASAP7_75t_R g4774 ( 
.A(n_4219),
.Y(n_4774)
);

CKINVDCx5p33_ASAP7_75t_R g4775 ( 
.A(n_390),
.Y(n_4775)
);

INVx1_ASAP7_75t_L g4776 ( 
.A(n_1734),
.Y(n_4776)
);

CKINVDCx5p33_ASAP7_75t_R g4777 ( 
.A(n_1824),
.Y(n_4777)
);

CKINVDCx5p33_ASAP7_75t_R g4778 ( 
.A(n_157),
.Y(n_4778)
);

BUFx6f_ASAP7_75t_L g4779 ( 
.A(n_2975),
.Y(n_4779)
);

CKINVDCx5p33_ASAP7_75t_R g4780 ( 
.A(n_3105),
.Y(n_4780)
);

CKINVDCx5p33_ASAP7_75t_R g4781 ( 
.A(n_3864),
.Y(n_4781)
);

CKINVDCx5p33_ASAP7_75t_R g4782 ( 
.A(n_420),
.Y(n_4782)
);

INVx1_ASAP7_75t_L g4783 ( 
.A(n_3179),
.Y(n_4783)
);

CKINVDCx5p33_ASAP7_75t_R g4784 ( 
.A(n_1729),
.Y(n_4784)
);

CKINVDCx5p33_ASAP7_75t_R g4785 ( 
.A(n_2392),
.Y(n_4785)
);

INVx1_ASAP7_75t_L g4786 ( 
.A(n_4220),
.Y(n_4786)
);

INVx2_ASAP7_75t_SL g4787 ( 
.A(n_249),
.Y(n_4787)
);

CKINVDCx5p33_ASAP7_75t_R g4788 ( 
.A(n_3447),
.Y(n_4788)
);

BUFx3_ASAP7_75t_L g4789 ( 
.A(n_1006),
.Y(n_4789)
);

CKINVDCx20_ASAP7_75t_R g4790 ( 
.A(n_686),
.Y(n_4790)
);

CKINVDCx5p33_ASAP7_75t_R g4791 ( 
.A(n_2278),
.Y(n_4791)
);

INVx1_ASAP7_75t_SL g4792 ( 
.A(n_2887),
.Y(n_4792)
);

CKINVDCx5p33_ASAP7_75t_R g4793 ( 
.A(n_1831),
.Y(n_4793)
);

INVx1_ASAP7_75t_SL g4794 ( 
.A(n_1296),
.Y(n_4794)
);

INVx1_ASAP7_75t_L g4795 ( 
.A(n_4044),
.Y(n_4795)
);

CKINVDCx5p33_ASAP7_75t_R g4796 ( 
.A(n_2047),
.Y(n_4796)
);

INVx1_ASAP7_75t_L g4797 ( 
.A(n_3320),
.Y(n_4797)
);

CKINVDCx5p33_ASAP7_75t_R g4798 ( 
.A(n_3580),
.Y(n_4798)
);

CKINVDCx5p33_ASAP7_75t_R g4799 ( 
.A(n_3236),
.Y(n_4799)
);

CKINVDCx5p33_ASAP7_75t_R g4800 ( 
.A(n_109),
.Y(n_4800)
);

CKINVDCx20_ASAP7_75t_R g4801 ( 
.A(n_1316),
.Y(n_4801)
);

CKINVDCx5p33_ASAP7_75t_R g4802 ( 
.A(n_4171),
.Y(n_4802)
);

INVx1_ASAP7_75t_L g4803 ( 
.A(n_3653),
.Y(n_4803)
);

CKINVDCx5p33_ASAP7_75t_R g4804 ( 
.A(n_2975),
.Y(n_4804)
);

INVx1_ASAP7_75t_L g4805 ( 
.A(n_3155),
.Y(n_4805)
);

CKINVDCx5p33_ASAP7_75t_R g4806 ( 
.A(n_1695),
.Y(n_4806)
);

INVx1_ASAP7_75t_L g4807 ( 
.A(n_2785),
.Y(n_4807)
);

CKINVDCx5p33_ASAP7_75t_R g4808 ( 
.A(n_1837),
.Y(n_4808)
);

INVx1_ASAP7_75t_L g4809 ( 
.A(n_1560),
.Y(n_4809)
);

INVx1_ASAP7_75t_L g4810 ( 
.A(n_1319),
.Y(n_4810)
);

CKINVDCx5p33_ASAP7_75t_R g4811 ( 
.A(n_951),
.Y(n_4811)
);

CKINVDCx5p33_ASAP7_75t_R g4812 ( 
.A(n_4060),
.Y(n_4812)
);

INVx1_ASAP7_75t_L g4813 ( 
.A(n_1929),
.Y(n_4813)
);

BUFx10_ASAP7_75t_L g4814 ( 
.A(n_4136),
.Y(n_4814)
);

INVx1_ASAP7_75t_L g4815 ( 
.A(n_2128),
.Y(n_4815)
);

CKINVDCx16_ASAP7_75t_R g4816 ( 
.A(n_2309),
.Y(n_4816)
);

CKINVDCx5p33_ASAP7_75t_R g4817 ( 
.A(n_4137),
.Y(n_4817)
);

BUFx3_ASAP7_75t_L g4818 ( 
.A(n_3259),
.Y(n_4818)
);

INVx1_ASAP7_75t_L g4819 ( 
.A(n_4077),
.Y(n_4819)
);

CKINVDCx5p33_ASAP7_75t_R g4820 ( 
.A(n_2233),
.Y(n_4820)
);

CKINVDCx20_ASAP7_75t_R g4821 ( 
.A(n_4190),
.Y(n_4821)
);

INVx2_ASAP7_75t_L g4822 ( 
.A(n_1),
.Y(n_4822)
);

CKINVDCx5p33_ASAP7_75t_R g4823 ( 
.A(n_3537),
.Y(n_4823)
);

CKINVDCx5p33_ASAP7_75t_R g4824 ( 
.A(n_908),
.Y(n_4824)
);

CKINVDCx5p33_ASAP7_75t_R g4825 ( 
.A(n_477),
.Y(n_4825)
);

BUFx3_ASAP7_75t_L g4826 ( 
.A(n_455),
.Y(n_4826)
);

CKINVDCx5p33_ASAP7_75t_R g4827 ( 
.A(n_1154),
.Y(n_4827)
);

CKINVDCx5p33_ASAP7_75t_R g4828 ( 
.A(n_3706),
.Y(n_4828)
);

BUFx10_ASAP7_75t_L g4829 ( 
.A(n_87),
.Y(n_4829)
);

CKINVDCx5p33_ASAP7_75t_R g4830 ( 
.A(n_887),
.Y(n_4830)
);

CKINVDCx20_ASAP7_75t_R g4831 ( 
.A(n_3082),
.Y(n_4831)
);

CKINVDCx20_ASAP7_75t_R g4832 ( 
.A(n_3336),
.Y(n_4832)
);

INVx1_ASAP7_75t_SL g4833 ( 
.A(n_3806),
.Y(n_4833)
);

CKINVDCx20_ASAP7_75t_R g4834 ( 
.A(n_4094),
.Y(n_4834)
);

BUFx3_ASAP7_75t_L g4835 ( 
.A(n_2238),
.Y(n_4835)
);

CKINVDCx5p33_ASAP7_75t_R g4836 ( 
.A(n_2564),
.Y(n_4836)
);

CKINVDCx5p33_ASAP7_75t_R g4837 ( 
.A(n_2481),
.Y(n_4837)
);

INVx1_ASAP7_75t_L g4838 ( 
.A(n_2013),
.Y(n_4838)
);

CKINVDCx5p33_ASAP7_75t_R g4839 ( 
.A(n_2231),
.Y(n_4839)
);

INVx1_ASAP7_75t_L g4840 ( 
.A(n_1671),
.Y(n_4840)
);

CKINVDCx20_ASAP7_75t_R g4841 ( 
.A(n_3240),
.Y(n_4841)
);

CKINVDCx5p33_ASAP7_75t_R g4842 ( 
.A(n_2342),
.Y(n_4842)
);

INVx1_ASAP7_75t_L g4843 ( 
.A(n_53),
.Y(n_4843)
);

INVx1_ASAP7_75t_L g4844 ( 
.A(n_2044),
.Y(n_4844)
);

CKINVDCx5p33_ASAP7_75t_R g4845 ( 
.A(n_3775),
.Y(n_4845)
);

CKINVDCx5p33_ASAP7_75t_R g4846 ( 
.A(n_1479),
.Y(n_4846)
);

CKINVDCx5p33_ASAP7_75t_R g4847 ( 
.A(n_18),
.Y(n_4847)
);

CKINVDCx5p33_ASAP7_75t_R g4848 ( 
.A(n_1397),
.Y(n_4848)
);

CKINVDCx5p33_ASAP7_75t_R g4849 ( 
.A(n_4154),
.Y(n_4849)
);

CKINVDCx20_ASAP7_75t_R g4850 ( 
.A(n_3716),
.Y(n_4850)
);

CKINVDCx5p33_ASAP7_75t_R g4851 ( 
.A(n_949),
.Y(n_4851)
);

INVx2_ASAP7_75t_L g4852 ( 
.A(n_4165),
.Y(n_4852)
);

BUFx6f_ASAP7_75t_L g4853 ( 
.A(n_566),
.Y(n_4853)
);

INVx1_ASAP7_75t_L g4854 ( 
.A(n_3669),
.Y(n_4854)
);

INVx1_ASAP7_75t_L g4855 ( 
.A(n_334),
.Y(n_4855)
);

INVx2_ASAP7_75t_SL g4856 ( 
.A(n_862),
.Y(n_4856)
);

CKINVDCx5p33_ASAP7_75t_R g4857 ( 
.A(n_4083),
.Y(n_4857)
);

CKINVDCx5p33_ASAP7_75t_R g4858 ( 
.A(n_4202),
.Y(n_4858)
);

CKINVDCx20_ASAP7_75t_R g4859 ( 
.A(n_4152),
.Y(n_4859)
);

CKINVDCx5p33_ASAP7_75t_R g4860 ( 
.A(n_214),
.Y(n_4860)
);

CKINVDCx5p33_ASAP7_75t_R g4861 ( 
.A(n_4104),
.Y(n_4861)
);

CKINVDCx5p33_ASAP7_75t_R g4862 ( 
.A(n_4298),
.Y(n_4862)
);

INVx2_ASAP7_75t_L g4863 ( 
.A(n_1230),
.Y(n_4863)
);

CKINVDCx5p33_ASAP7_75t_R g4864 ( 
.A(n_857),
.Y(n_4864)
);

BUFx6f_ASAP7_75t_L g4865 ( 
.A(n_3062),
.Y(n_4865)
);

INVx1_ASAP7_75t_L g4866 ( 
.A(n_936),
.Y(n_4866)
);

CKINVDCx5p33_ASAP7_75t_R g4867 ( 
.A(n_787),
.Y(n_4867)
);

INVx1_ASAP7_75t_L g4868 ( 
.A(n_4275),
.Y(n_4868)
);

INVx1_ASAP7_75t_L g4869 ( 
.A(n_406),
.Y(n_4869)
);

CKINVDCx5p33_ASAP7_75t_R g4870 ( 
.A(n_740),
.Y(n_4870)
);

CKINVDCx5p33_ASAP7_75t_R g4871 ( 
.A(n_4318),
.Y(n_4871)
);

INVx1_ASAP7_75t_L g4872 ( 
.A(n_3454),
.Y(n_4872)
);

INVx2_ASAP7_75t_SL g4873 ( 
.A(n_3542),
.Y(n_4873)
);

CKINVDCx5p33_ASAP7_75t_R g4874 ( 
.A(n_4197),
.Y(n_4874)
);

CKINVDCx5p33_ASAP7_75t_R g4875 ( 
.A(n_2807),
.Y(n_4875)
);

CKINVDCx5p33_ASAP7_75t_R g4876 ( 
.A(n_3483),
.Y(n_4876)
);

CKINVDCx5p33_ASAP7_75t_R g4877 ( 
.A(n_600),
.Y(n_4877)
);

INVxp67_ASAP7_75t_L g4878 ( 
.A(n_963),
.Y(n_4878)
);

INVx1_ASAP7_75t_L g4879 ( 
.A(n_3603),
.Y(n_4879)
);

CKINVDCx5p33_ASAP7_75t_R g4880 ( 
.A(n_3483),
.Y(n_4880)
);

INVx1_ASAP7_75t_L g4881 ( 
.A(n_4093),
.Y(n_4881)
);

CKINVDCx5p33_ASAP7_75t_R g4882 ( 
.A(n_1846),
.Y(n_4882)
);

CKINVDCx5p33_ASAP7_75t_R g4883 ( 
.A(n_2466),
.Y(n_4883)
);

CKINVDCx5p33_ASAP7_75t_R g4884 ( 
.A(n_3546),
.Y(n_4884)
);

INVx1_ASAP7_75t_SL g4885 ( 
.A(n_2398),
.Y(n_4885)
);

CKINVDCx5p33_ASAP7_75t_R g4886 ( 
.A(n_3356),
.Y(n_4886)
);

CKINVDCx5p33_ASAP7_75t_R g4887 ( 
.A(n_128),
.Y(n_4887)
);

CKINVDCx20_ASAP7_75t_R g4888 ( 
.A(n_3152),
.Y(n_4888)
);

CKINVDCx16_ASAP7_75t_R g4889 ( 
.A(n_195),
.Y(n_4889)
);

CKINVDCx14_ASAP7_75t_R g4890 ( 
.A(n_609),
.Y(n_4890)
);

CKINVDCx5p33_ASAP7_75t_R g4891 ( 
.A(n_1777),
.Y(n_4891)
);

CKINVDCx5p33_ASAP7_75t_R g4892 ( 
.A(n_400),
.Y(n_4892)
);

INVx1_ASAP7_75t_L g4893 ( 
.A(n_2750),
.Y(n_4893)
);

CKINVDCx14_ASAP7_75t_R g4894 ( 
.A(n_285),
.Y(n_4894)
);

CKINVDCx5p33_ASAP7_75t_R g4895 ( 
.A(n_3499),
.Y(n_4895)
);

INVx1_ASAP7_75t_L g4896 ( 
.A(n_2644),
.Y(n_4896)
);

CKINVDCx5p33_ASAP7_75t_R g4897 ( 
.A(n_2786),
.Y(n_4897)
);

CKINVDCx5p33_ASAP7_75t_R g4898 ( 
.A(n_2680),
.Y(n_4898)
);

CKINVDCx5p33_ASAP7_75t_R g4899 ( 
.A(n_2929),
.Y(n_4899)
);

INVx1_ASAP7_75t_L g4900 ( 
.A(n_2226),
.Y(n_4900)
);

CKINVDCx14_ASAP7_75t_R g4901 ( 
.A(n_4153),
.Y(n_4901)
);

INVx1_ASAP7_75t_SL g4902 ( 
.A(n_4117),
.Y(n_4902)
);

BUFx3_ASAP7_75t_L g4903 ( 
.A(n_2191),
.Y(n_4903)
);

CKINVDCx5p33_ASAP7_75t_R g4904 ( 
.A(n_1968),
.Y(n_4904)
);

CKINVDCx5p33_ASAP7_75t_R g4905 ( 
.A(n_1160),
.Y(n_4905)
);

INVx1_ASAP7_75t_L g4906 ( 
.A(n_966),
.Y(n_4906)
);

INVx1_ASAP7_75t_SL g4907 ( 
.A(n_2380),
.Y(n_4907)
);

INVx1_ASAP7_75t_L g4908 ( 
.A(n_2436),
.Y(n_4908)
);

INVx2_ASAP7_75t_L g4909 ( 
.A(n_3471),
.Y(n_4909)
);

INVx1_ASAP7_75t_L g4910 ( 
.A(n_542),
.Y(n_4910)
);

CKINVDCx20_ASAP7_75t_R g4911 ( 
.A(n_1230),
.Y(n_4911)
);

CKINVDCx20_ASAP7_75t_R g4912 ( 
.A(n_1913),
.Y(n_4912)
);

CKINVDCx5p33_ASAP7_75t_R g4913 ( 
.A(n_4056),
.Y(n_4913)
);

CKINVDCx5p33_ASAP7_75t_R g4914 ( 
.A(n_2265),
.Y(n_4914)
);

CKINVDCx20_ASAP7_75t_R g4915 ( 
.A(n_4187),
.Y(n_4915)
);

INVx1_ASAP7_75t_L g4916 ( 
.A(n_2723),
.Y(n_4916)
);

BUFx10_ASAP7_75t_L g4917 ( 
.A(n_907),
.Y(n_4917)
);

CKINVDCx5p33_ASAP7_75t_R g4918 ( 
.A(n_4126),
.Y(n_4918)
);

INVx2_ASAP7_75t_SL g4919 ( 
.A(n_2462),
.Y(n_4919)
);

INVx2_ASAP7_75t_SL g4920 ( 
.A(n_2313),
.Y(n_4920)
);

CKINVDCx5p33_ASAP7_75t_R g4921 ( 
.A(n_2001),
.Y(n_4921)
);

BUFx3_ASAP7_75t_L g4922 ( 
.A(n_1087),
.Y(n_4922)
);

CKINVDCx5p33_ASAP7_75t_R g4923 ( 
.A(n_3068),
.Y(n_4923)
);

CKINVDCx20_ASAP7_75t_R g4924 ( 
.A(n_747),
.Y(n_4924)
);

INVx2_ASAP7_75t_SL g4925 ( 
.A(n_1913),
.Y(n_4925)
);

CKINVDCx5p33_ASAP7_75t_R g4926 ( 
.A(n_1390),
.Y(n_4926)
);

CKINVDCx5p33_ASAP7_75t_R g4927 ( 
.A(n_4204),
.Y(n_4927)
);

INVx1_ASAP7_75t_L g4928 ( 
.A(n_1191),
.Y(n_4928)
);

HB1xp67_ASAP7_75t_L g4929 ( 
.A(n_3090),
.Y(n_4929)
);

CKINVDCx5p33_ASAP7_75t_R g4930 ( 
.A(n_1123),
.Y(n_4930)
);

CKINVDCx5p33_ASAP7_75t_R g4931 ( 
.A(n_4206),
.Y(n_4931)
);

CKINVDCx5p33_ASAP7_75t_R g4932 ( 
.A(n_3642),
.Y(n_4932)
);

CKINVDCx5p33_ASAP7_75t_R g4933 ( 
.A(n_1852),
.Y(n_4933)
);

CKINVDCx5p33_ASAP7_75t_R g4934 ( 
.A(n_3366),
.Y(n_4934)
);

INVx1_ASAP7_75t_L g4935 ( 
.A(n_3181),
.Y(n_4935)
);

CKINVDCx5p33_ASAP7_75t_R g4936 ( 
.A(n_477),
.Y(n_4936)
);

CKINVDCx5p33_ASAP7_75t_R g4937 ( 
.A(n_2847),
.Y(n_4937)
);

BUFx2_ASAP7_75t_L g4938 ( 
.A(n_3718),
.Y(n_4938)
);

INVx1_ASAP7_75t_L g4939 ( 
.A(n_615),
.Y(n_4939)
);

INVx1_ASAP7_75t_L g4940 ( 
.A(n_4110),
.Y(n_4940)
);

CKINVDCx20_ASAP7_75t_R g4941 ( 
.A(n_693),
.Y(n_4941)
);

CKINVDCx5p33_ASAP7_75t_R g4942 ( 
.A(n_495),
.Y(n_4942)
);

CKINVDCx5p33_ASAP7_75t_R g4943 ( 
.A(n_795),
.Y(n_4943)
);

INVx1_ASAP7_75t_L g4944 ( 
.A(n_638),
.Y(n_4944)
);

INVx1_ASAP7_75t_SL g4945 ( 
.A(n_3583),
.Y(n_4945)
);

BUFx2_ASAP7_75t_SL g4946 ( 
.A(n_3695),
.Y(n_4946)
);

CKINVDCx5p33_ASAP7_75t_R g4947 ( 
.A(n_3044),
.Y(n_4947)
);

CKINVDCx20_ASAP7_75t_R g4948 ( 
.A(n_1417),
.Y(n_4948)
);

INVx1_ASAP7_75t_SL g4949 ( 
.A(n_2245),
.Y(n_4949)
);

INVx2_ASAP7_75t_L g4950 ( 
.A(n_728),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_886),
.Y(n_4951)
);

CKINVDCx5p33_ASAP7_75t_R g4952 ( 
.A(n_2587),
.Y(n_4952)
);

CKINVDCx5p33_ASAP7_75t_R g4953 ( 
.A(n_1634),
.Y(n_4953)
);

INVx1_ASAP7_75t_L g4954 ( 
.A(n_2751),
.Y(n_4954)
);

INVx1_ASAP7_75t_L g4955 ( 
.A(n_2368),
.Y(n_4955)
);

BUFx3_ASAP7_75t_L g4956 ( 
.A(n_2074),
.Y(n_4956)
);

CKINVDCx20_ASAP7_75t_R g4957 ( 
.A(n_2984),
.Y(n_4957)
);

INVx1_ASAP7_75t_L g4958 ( 
.A(n_2858),
.Y(n_4958)
);

CKINVDCx5p33_ASAP7_75t_R g4959 ( 
.A(n_533),
.Y(n_4959)
);

INVx2_ASAP7_75t_L g4960 ( 
.A(n_3313),
.Y(n_4960)
);

CKINVDCx5p33_ASAP7_75t_R g4961 ( 
.A(n_3823),
.Y(n_4961)
);

INVx1_ASAP7_75t_L g4962 ( 
.A(n_3791),
.Y(n_4962)
);

CKINVDCx5p33_ASAP7_75t_R g4963 ( 
.A(n_2738),
.Y(n_4963)
);

INVx1_ASAP7_75t_L g4964 ( 
.A(n_4062),
.Y(n_4964)
);

INVx2_ASAP7_75t_SL g4965 ( 
.A(n_3910),
.Y(n_4965)
);

INVx1_ASAP7_75t_L g4966 ( 
.A(n_4218),
.Y(n_4966)
);

INVx2_ASAP7_75t_L g4967 ( 
.A(n_4068),
.Y(n_4967)
);

INVx1_ASAP7_75t_L g4968 ( 
.A(n_1511),
.Y(n_4968)
);

CKINVDCx5p33_ASAP7_75t_R g4969 ( 
.A(n_3268),
.Y(n_4969)
);

INVx1_ASAP7_75t_SL g4970 ( 
.A(n_2617),
.Y(n_4970)
);

CKINVDCx5p33_ASAP7_75t_R g4971 ( 
.A(n_2642),
.Y(n_4971)
);

CKINVDCx5p33_ASAP7_75t_R g4972 ( 
.A(n_4188),
.Y(n_4972)
);

CKINVDCx5p33_ASAP7_75t_R g4973 ( 
.A(n_3251),
.Y(n_4973)
);

BUFx6f_ASAP7_75t_L g4974 ( 
.A(n_1218),
.Y(n_4974)
);

INVx1_ASAP7_75t_L g4975 ( 
.A(n_2080),
.Y(n_4975)
);

CKINVDCx5p33_ASAP7_75t_R g4976 ( 
.A(n_1759),
.Y(n_4976)
);

CKINVDCx5p33_ASAP7_75t_R g4977 ( 
.A(n_2710),
.Y(n_4977)
);

INVx2_ASAP7_75t_SL g4978 ( 
.A(n_4196),
.Y(n_4978)
);

CKINVDCx5p33_ASAP7_75t_R g4979 ( 
.A(n_2256),
.Y(n_4979)
);

INVx1_ASAP7_75t_L g4980 ( 
.A(n_3741),
.Y(n_4980)
);

CKINVDCx5p33_ASAP7_75t_R g4981 ( 
.A(n_2293),
.Y(n_4981)
);

CKINVDCx5p33_ASAP7_75t_R g4982 ( 
.A(n_3352),
.Y(n_4982)
);

CKINVDCx5p33_ASAP7_75t_R g4983 ( 
.A(n_1130),
.Y(n_4983)
);

BUFx3_ASAP7_75t_L g4984 ( 
.A(n_4120),
.Y(n_4984)
);

INVx2_ASAP7_75t_L g4985 ( 
.A(n_2471),
.Y(n_4985)
);

CKINVDCx20_ASAP7_75t_R g4986 ( 
.A(n_3479),
.Y(n_4986)
);

CKINVDCx5p33_ASAP7_75t_R g4987 ( 
.A(n_821),
.Y(n_4987)
);

CKINVDCx5p33_ASAP7_75t_R g4988 ( 
.A(n_2109),
.Y(n_4988)
);

INVx1_ASAP7_75t_L g4989 ( 
.A(n_1281),
.Y(n_4989)
);

INVx2_ASAP7_75t_L g4990 ( 
.A(n_3183),
.Y(n_4990)
);

CKINVDCx5p33_ASAP7_75t_R g4991 ( 
.A(n_2566),
.Y(n_4991)
);

INVx1_ASAP7_75t_L g4992 ( 
.A(n_2008),
.Y(n_4992)
);

CKINVDCx5p33_ASAP7_75t_R g4993 ( 
.A(n_4084),
.Y(n_4993)
);

CKINVDCx5p33_ASAP7_75t_R g4994 ( 
.A(n_1865),
.Y(n_4994)
);

CKINVDCx5p33_ASAP7_75t_R g4995 ( 
.A(n_3035),
.Y(n_4995)
);

CKINVDCx5p33_ASAP7_75t_R g4996 ( 
.A(n_2944),
.Y(n_4996)
);

CKINVDCx5p33_ASAP7_75t_R g4997 ( 
.A(n_2070),
.Y(n_4997)
);

CKINVDCx5p33_ASAP7_75t_R g4998 ( 
.A(n_725),
.Y(n_4998)
);

INVx2_ASAP7_75t_L g4999 ( 
.A(n_881),
.Y(n_4999)
);

CKINVDCx20_ASAP7_75t_R g5000 ( 
.A(n_1336),
.Y(n_5000)
);

CKINVDCx5p33_ASAP7_75t_R g5001 ( 
.A(n_1921),
.Y(n_5001)
);

CKINVDCx5p33_ASAP7_75t_R g5002 ( 
.A(n_1772),
.Y(n_5002)
);

INVx1_ASAP7_75t_L g5003 ( 
.A(n_3),
.Y(n_5003)
);

CKINVDCx5p33_ASAP7_75t_R g5004 ( 
.A(n_4055),
.Y(n_5004)
);

INVx1_ASAP7_75t_L g5005 ( 
.A(n_1062),
.Y(n_5005)
);

CKINVDCx5p33_ASAP7_75t_R g5006 ( 
.A(n_2932),
.Y(n_5006)
);

INVx1_ASAP7_75t_L g5007 ( 
.A(n_557),
.Y(n_5007)
);

BUFx3_ASAP7_75t_L g5008 ( 
.A(n_3875),
.Y(n_5008)
);

CKINVDCx5p33_ASAP7_75t_R g5009 ( 
.A(n_3636),
.Y(n_5009)
);

INVx2_ASAP7_75t_SL g5010 ( 
.A(n_3092),
.Y(n_5010)
);

INVx1_ASAP7_75t_L g5011 ( 
.A(n_2952),
.Y(n_5011)
);

CKINVDCx20_ASAP7_75t_R g5012 ( 
.A(n_4284),
.Y(n_5012)
);

INVx1_ASAP7_75t_L g5013 ( 
.A(n_4169),
.Y(n_5013)
);

INVx1_ASAP7_75t_L g5014 ( 
.A(n_579),
.Y(n_5014)
);

CKINVDCx5p33_ASAP7_75t_R g5015 ( 
.A(n_321),
.Y(n_5015)
);

CKINVDCx20_ASAP7_75t_R g5016 ( 
.A(n_3884),
.Y(n_5016)
);

CKINVDCx5p33_ASAP7_75t_R g5017 ( 
.A(n_729),
.Y(n_5017)
);

CKINVDCx5p33_ASAP7_75t_R g5018 ( 
.A(n_3225),
.Y(n_5018)
);

CKINVDCx5p33_ASAP7_75t_R g5019 ( 
.A(n_1386),
.Y(n_5019)
);

INVx3_ASAP7_75t_L g5020 ( 
.A(n_1003),
.Y(n_5020)
);

INVx1_ASAP7_75t_L g5021 ( 
.A(n_1448),
.Y(n_5021)
);

CKINVDCx5p33_ASAP7_75t_R g5022 ( 
.A(n_1756),
.Y(n_5022)
);

INVx1_ASAP7_75t_L g5023 ( 
.A(n_4195),
.Y(n_5023)
);

BUFx10_ASAP7_75t_L g5024 ( 
.A(n_348),
.Y(n_5024)
);

CKINVDCx5p33_ASAP7_75t_R g5025 ( 
.A(n_3681),
.Y(n_5025)
);

CKINVDCx5p33_ASAP7_75t_R g5026 ( 
.A(n_598),
.Y(n_5026)
);

CKINVDCx20_ASAP7_75t_R g5027 ( 
.A(n_2995),
.Y(n_5027)
);

INVx1_ASAP7_75t_L g5028 ( 
.A(n_3523),
.Y(n_5028)
);

INVx1_ASAP7_75t_L g5029 ( 
.A(n_741),
.Y(n_5029)
);

CKINVDCx5p33_ASAP7_75t_R g5030 ( 
.A(n_3637),
.Y(n_5030)
);

CKINVDCx16_ASAP7_75t_R g5031 ( 
.A(n_2462),
.Y(n_5031)
);

INVx1_ASAP7_75t_L g5032 ( 
.A(n_3439),
.Y(n_5032)
);

CKINVDCx5p33_ASAP7_75t_R g5033 ( 
.A(n_1365),
.Y(n_5033)
);

CKINVDCx5p33_ASAP7_75t_R g5034 ( 
.A(n_4285),
.Y(n_5034)
);

INVx1_ASAP7_75t_L g5035 ( 
.A(n_2874),
.Y(n_5035)
);

CKINVDCx5p33_ASAP7_75t_R g5036 ( 
.A(n_2726),
.Y(n_5036)
);

CKINVDCx5p33_ASAP7_75t_R g5037 ( 
.A(n_540),
.Y(n_5037)
);

CKINVDCx5p33_ASAP7_75t_R g5038 ( 
.A(n_1869),
.Y(n_5038)
);

CKINVDCx5p33_ASAP7_75t_R g5039 ( 
.A(n_4209),
.Y(n_5039)
);

INVx1_ASAP7_75t_SL g5040 ( 
.A(n_1563),
.Y(n_5040)
);

CKINVDCx5p33_ASAP7_75t_R g5041 ( 
.A(n_2685),
.Y(n_5041)
);

INVx1_ASAP7_75t_L g5042 ( 
.A(n_3842),
.Y(n_5042)
);

CKINVDCx5p33_ASAP7_75t_R g5043 ( 
.A(n_349),
.Y(n_5043)
);

CKINVDCx5p33_ASAP7_75t_R g5044 ( 
.A(n_2411),
.Y(n_5044)
);

CKINVDCx5p33_ASAP7_75t_R g5045 ( 
.A(n_2960),
.Y(n_5045)
);

BUFx5_ASAP7_75t_L g5046 ( 
.A(n_3592),
.Y(n_5046)
);

CKINVDCx5p33_ASAP7_75t_R g5047 ( 
.A(n_2483),
.Y(n_5047)
);

CKINVDCx5p33_ASAP7_75t_R g5048 ( 
.A(n_4123),
.Y(n_5048)
);

CKINVDCx16_ASAP7_75t_R g5049 ( 
.A(n_2515),
.Y(n_5049)
);

CKINVDCx5p33_ASAP7_75t_R g5050 ( 
.A(n_3878),
.Y(n_5050)
);

CKINVDCx5p33_ASAP7_75t_R g5051 ( 
.A(n_352),
.Y(n_5051)
);

CKINVDCx5p33_ASAP7_75t_R g5052 ( 
.A(n_639),
.Y(n_5052)
);

INVx2_ASAP7_75t_L g5053 ( 
.A(n_843),
.Y(n_5053)
);

INVx1_ASAP7_75t_L g5054 ( 
.A(n_1418),
.Y(n_5054)
);

CKINVDCx5p33_ASAP7_75t_R g5055 ( 
.A(n_4179),
.Y(n_5055)
);

CKINVDCx20_ASAP7_75t_R g5056 ( 
.A(n_3866),
.Y(n_5056)
);

CKINVDCx5p33_ASAP7_75t_R g5057 ( 
.A(n_982),
.Y(n_5057)
);

INVxp33_ASAP7_75t_SL g5058 ( 
.A(n_4050),
.Y(n_5058)
);

INVx1_ASAP7_75t_L g5059 ( 
.A(n_2334),
.Y(n_5059)
);

CKINVDCx5p33_ASAP7_75t_R g5060 ( 
.A(n_1102),
.Y(n_5060)
);

INVx2_ASAP7_75t_SL g5061 ( 
.A(n_1796),
.Y(n_5061)
);

CKINVDCx20_ASAP7_75t_R g5062 ( 
.A(n_3860),
.Y(n_5062)
);

CKINVDCx5p33_ASAP7_75t_R g5063 ( 
.A(n_3134),
.Y(n_5063)
);

CKINVDCx5p33_ASAP7_75t_R g5064 ( 
.A(n_3364),
.Y(n_5064)
);

CKINVDCx5p33_ASAP7_75t_R g5065 ( 
.A(n_1536),
.Y(n_5065)
);

INVx2_ASAP7_75t_L g5066 ( 
.A(n_2784),
.Y(n_5066)
);

BUFx6f_ASAP7_75t_L g5067 ( 
.A(n_303),
.Y(n_5067)
);

CKINVDCx5p33_ASAP7_75t_R g5068 ( 
.A(n_256),
.Y(n_5068)
);

INVx1_ASAP7_75t_L g5069 ( 
.A(n_3920),
.Y(n_5069)
);

HB1xp67_ASAP7_75t_L g5070 ( 
.A(n_4113),
.Y(n_5070)
);

BUFx6f_ASAP7_75t_L g5071 ( 
.A(n_2537),
.Y(n_5071)
);

INVx1_ASAP7_75t_L g5072 ( 
.A(n_4011),
.Y(n_5072)
);

CKINVDCx5p33_ASAP7_75t_R g5073 ( 
.A(n_2563),
.Y(n_5073)
);

CKINVDCx20_ASAP7_75t_R g5074 ( 
.A(n_52),
.Y(n_5074)
);

CKINVDCx5p33_ASAP7_75t_R g5075 ( 
.A(n_4181),
.Y(n_5075)
);

CKINVDCx5p33_ASAP7_75t_R g5076 ( 
.A(n_382),
.Y(n_5076)
);

CKINVDCx5p33_ASAP7_75t_R g5077 ( 
.A(n_2916),
.Y(n_5077)
);

CKINVDCx5p33_ASAP7_75t_R g5078 ( 
.A(n_18),
.Y(n_5078)
);

CKINVDCx5p33_ASAP7_75t_R g5079 ( 
.A(n_4108),
.Y(n_5079)
);

BUFx10_ASAP7_75t_L g5080 ( 
.A(n_4081),
.Y(n_5080)
);

CKINVDCx5p33_ASAP7_75t_R g5081 ( 
.A(n_2166),
.Y(n_5081)
);

CKINVDCx5p33_ASAP7_75t_R g5082 ( 
.A(n_2187),
.Y(n_5082)
);

CKINVDCx5p33_ASAP7_75t_R g5083 ( 
.A(n_1970),
.Y(n_5083)
);

CKINVDCx5p33_ASAP7_75t_R g5084 ( 
.A(n_3223),
.Y(n_5084)
);

CKINVDCx5p33_ASAP7_75t_R g5085 ( 
.A(n_1504),
.Y(n_5085)
);

CKINVDCx5p33_ASAP7_75t_R g5086 ( 
.A(n_4201),
.Y(n_5086)
);

CKINVDCx5p33_ASAP7_75t_R g5087 ( 
.A(n_2287),
.Y(n_5087)
);

CKINVDCx16_ASAP7_75t_R g5088 ( 
.A(n_3189),
.Y(n_5088)
);

CKINVDCx5p33_ASAP7_75t_R g5089 ( 
.A(n_332),
.Y(n_5089)
);

INVx1_ASAP7_75t_L g5090 ( 
.A(n_2709),
.Y(n_5090)
);

INVx1_ASAP7_75t_L g5091 ( 
.A(n_1565),
.Y(n_5091)
);

CKINVDCx20_ASAP7_75t_R g5092 ( 
.A(n_1714),
.Y(n_5092)
);

CKINVDCx5p33_ASAP7_75t_R g5093 ( 
.A(n_762),
.Y(n_5093)
);

CKINVDCx5p33_ASAP7_75t_R g5094 ( 
.A(n_3320),
.Y(n_5094)
);

CKINVDCx5p33_ASAP7_75t_R g5095 ( 
.A(n_2857),
.Y(n_5095)
);

CKINVDCx5p33_ASAP7_75t_R g5096 ( 
.A(n_2100),
.Y(n_5096)
);

INVx1_ASAP7_75t_L g5097 ( 
.A(n_864),
.Y(n_5097)
);

CKINVDCx5p33_ASAP7_75t_R g5098 ( 
.A(n_2773),
.Y(n_5098)
);

INVx1_ASAP7_75t_L g5099 ( 
.A(n_3187),
.Y(n_5099)
);

CKINVDCx5p33_ASAP7_75t_R g5100 ( 
.A(n_839),
.Y(n_5100)
);

CKINVDCx5p33_ASAP7_75t_R g5101 ( 
.A(n_3620),
.Y(n_5101)
);

BUFx6f_ASAP7_75t_L g5102 ( 
.A(n_4036),
.Y(n_5102)
);

CKINVDCx5p33_ASAP7_75t_R g5103 ( 
.A(n_4119),
.Y(n_5103)
);

INVx2_ASAP7_75t_SL g5104 ( 
.A(n_2376),
.Y(n_5104)
);

CKINVDCx5p33_ASAP7_75t_R g5105 ( 
.A(n_1307),
.Y(n_5105)
);

INVx1_ASAP7_75t_L g5106 ( 
.A(n_4147),
.Y(n_5106)
);

INVx2_ASAP7_75t_L g5107 ( 
.A(n_3586),
.Y(n_5107)
);

INVx1_ASAP7_75t_L g5108 ( 
.A(n_979),
.Y(n_5108)
);

BUFx2_ASAP7_75t_L g5109 ( 
.A(n_2684),
.Y(n_5109)
);

CKINVDCx5p33_ASAP7_75t_R g5110 ( 
.A(n_2361),
.Y(n_5110)
);

INVx1_ASAP7_75t_L g5111 ( 
.A(n_1099),
.Y(n_5111)
);

INVx1_ASAP7_75t_L g5112 ( 
.A(n_4194),
.Y(n_5112)
);

CKINVDCx5p33_ASAP7_75t_R g5113 ( 
.A(n_4207),
.Y(n_5113)
);

INVx1_ASAP7_75t_L g5114 ( 
.A(n_794),
.Y(n_5114)
);

CKINVDCx20_ASAP7_75t_R g5115 ( 
.A(n_3650),
.Y(n_5115)
);

INVx1_ASAP7_75t_L g5116 ( 
.A(n_3272),
.Y(n_5116)
);

BUFx5_ASAP7_75t_L g5117 ( 
.A(n_1519),
.Y(n_5117)
);

BUFx6f_ASAP7_75t_L g5118 ( 
.A(n_2030),
.Y(n_5118)
);

INVx1_ASAP7_75t_L g5119 ( 
.A(n_2984),
.Y(n_5119)
);

CKINVDCx5p33_ASAP7_75t_R g5120 ( 
.A(n_737),
.Y(n_5120)
);

CKINVDCx5p33_ASAP7_75t_R g5121 ( 
.A(n_3839),
.Y(n_5121)
);

INVx1_ASAP7_75t_L g5122 ( 
.A(n_2042),
.Y(n_5122)
);

CKINVDCx5p33_ASAP7_75t_R g5123 ( 
.A(n_944),
.Y(n_5123)
);

CKINVDCx5p33_ASAP7_75t_R g5124 ( 
.A(n_4227),
.Y(n_5124)
);

CKINVDCx16_ASAP7_75t_R g5125 ( 
.A(n_1723),
.Y(n_5125)
);

INVx1_ASAP7_75t_L g5126 ( 
.A(n_4107),
.Y(n_5126)
);

INVx2_ASAP7_75t_SL g5127 ( 
.A(n_3370),
.Y(n_5127)
);

CKINVDCx5p33_ASAP7_75t_R g5128 ( 
.A(n_1955),
.Y(n_5128)
);

INVx1_ASAP7_75t_L g5129 ( 
.A(n_1196),
.Y(n_5129)
);

CKINVDCx5p33_ASAP7_75t_R g5130 ( 
.A(n_1893),
.Y(n_5130)
);

CKINVDCx5p33_ASAP7_75t_R g5131 ( 
.A(n_769),
.Y(n_5131)
);

CKINVDCx5p33_ASAP7_75t_R g5132 ( 
.A(n_2907),
.Y(n_5132)
);

CKINVDCx5p33_ASAP7_75t_R g5133 ( 
.A(n_3764),
.Y(n_5133)
);

INVx2_ASAP7_75t_L g5134 ( 
.A(n_1936),
.Y(n_5134)
);

BUFx3_ASAP7_75t_L g5135 ( 
.A(n_255),
.Y(n_5135)
);

INVx1_ASAP7_75t_L g5136 ( 
.A(n_2821),
.Y(n_5136)
);

CKINVDCx5p33_ASAP7_75t_R g5137 ( 
.A(n_4057),
.Y(n_5137)
);

CKINVDCx5p33_ASAP7_75t_R g5138 ( 
.A(n_2573),
.Y(n_5138)
);

BUFx10_ASAP7_75t_L g5139 ( 
.A(n_2870),
.Y(n_5139)
);

BUFx2_ASAP7_75t_SL g5140 ( 
.A(n_3433),
.Y(n_5140)
);

BUFx6f_ASAP7_75t_L g5141 ( 
.A(n_1420),
.Y(n_5141)
);

INVx1_ASAP7_75t_L g5142 ( 
.A(n_2870),
.Y(n_5142)
);

INVx1_ASAP7_75t_L g5143 ( 
.A(n_1113),
.Y(n_5143)
);

CKINVDCx14_ASAP7_75t_R g5144 ( 
.A(n_4140),
.Y(n_5144)
);

INVx1_ASAP7_75t_L g5145 ( 
.A(n_2073),
.Y(n_5145)
);

INVx1_ASAP7_75t_L g5146 ( 
.A(n_3127),
.Y(n_5146)
);

INVx1_ASAP7_75t_L g5147 ( 
.A(n_4103),
.Y(n_5147)
);

INVx1_ASAP7_75t_L g5148 ( 
.A(n_629),
.Y(n_5148)
);

CKINVDCx5p33_ASAP7_75t_R g5149 ( 
.A(n_104),
.Y(n_5149)
);

CKINVDCx5p33_ASAP7_75t_R g5150 ( 
.A(n_2877),
.Y(n_5150)
);

INVx2_ASAP7_75t_L g5151 ( 
.A(n_3864),
.Y(n_5151)
);

INVx1_ASAP7_75t_L g5152 ( 
.A(n_4218),
.Y(n_5152)
);

INVx1_ASAP7_75t_L g5153 ( 
.A(n_3640),
.Y(n_5153)
);

CKINVDCx5p33_ASAP7_75t_R g5154 ( 
.A(n_4080),
.Y(n_5154)
);

INVx1_ASAP7_75t_L g5155 ( 
.A(n_2751),
.Y(n_5155)
);

CKINVDCx5p33_ASAP7_75t_R g5156 ( 
.A(n_1817),
.Y(n_5156)
);

INVx2_ASAP7_75t_L g5157 ( 
.A(n_2096),
.Y(n_5157)
);

CKINVDCx5p33_ASAP7_75t_R g5158 ( 
.A(n_4154),
.Y(n_5158)
);

INVx1_ASAP7_75t_L g5159 ( 
.A(n_164),
.Y(n_5159)
);

INVx1_ASAP7_75t_L g5160 ( 
.A(n_2744),
.Y(n_5160)
);

INVx2_ASAP7_75t_SL g5161 ( 
.A(n_1048),
.Y(n_5161)
);

CKINVDCx5p33_ASAP7_75t_R g5162 ( 
.A(n_2997),
.Y(n_5162)
);

BUFx2_ASAP7_75t_L g5163 ( 
.A(n_934),
.Y(n_5163)
);

BUFx3_ASAP7_75t_L g5164 ( 
.A(n_1319),
.Y(n_5164)
);

INVx1_ASAP7_75t_SL g5165 ( 
.A(n_4151),
.Y(n_5165)
);

BUFx10_ASAP7_75t_L g5166 ( 
.A(n_1399),
.Y(n_5166)
);

CKINVDCx5p33_ASAP7_75t_R g5167 ( 
.A(n_1052),
.Y(n_5167)
);

INVx2_ASAP7_75t_SL g5168 ( 
.A(n_3871),
.Y(n_5168)
);

BUFx2_ASAP7_75t_L g5169 ( 
.A(n_4111),
.Y(n_5169)
);

CKINVDCx5p33_ASAP7_75t_R g5170 ( 
.A(n_634),
.Y(n_5170)
);

INVx1_ASAP7_75t_L g5171 ( 
.A(n_3959),
.Y(n_5171)
);

CKINVDCx5p33_ASAP7_75t_R g5172 ( 
.A(n_1340),
.Y(n_5172)
);

INVx1_ASAP7_75t_SL g5173 ( 
.A(n_3851),
.Y(n_5173)
);

INVx2_ASAP7_75t_L g5174 ( 
.A(n_2103),
.Y(n_5174)
);

CKINVDCx5p33_ASAP7_75t_R g5175 ( 
.A(n_539),
.Y(n_5175)
);

CKINVDCx5p33_ASAP7_75t_R g5176 ( 
.A(n_4054),
.Y(n_5176)
);

CKINVDCx5p33_ASAP7_75t_R g5177 ( 
.A(n_2804),
.Y(n_5177)
);

CKINVDCx5p33_ASAP7_75t_R g5178 ( 
.A(n_3992),
.Y(n_5178)
);

CKINVDCx5p33_ASAP7_75t_R g5179 ( 
.A(n_2927),
.Y(n_5179)
);

CKINVDCx5p33_ASAP7_75t_R g5180 ( 
.A(n_13),
.Y(n_5180)
);

CKINVDCx5p33_ASAP7_75t_R g5181 ( 
.A(n_206),
.Y(n_5181)
);

INVx1_ASAP7_75t_L g5182 ( 
.A(n_4235),
.Y(n_5182)
);

CKINVDCx20_ASAP7_75t_R g5183 ( 
.A(n_3761),
.Y(n_5183)
);

CKINVDCx5p33_ASAP7_75t_R g5184 ( 
.A(n_158),
.Y(n_5184)
);

CKINVDCx5p33_ASAP7_75t_R g5185 ( 
.A(n_3088),
.Y(n_5185)
);

INVx1_ASAP7_75t_L g5186 ( 
.A(n_3901),
.Y(n_5186)
);

INVx1_ASAP7_75t_L g5187 ( 
.A(n_125),
.Y(n_5187)
);

INVx1_ASAP7_75t_L g5188 ( 
.A(n_4125),
.Y(n_5188)
);

CKINVDCx5p33_ASAP7_75t_R g5189 ( 
.A(n_2508),
.Y(n_5189)
);

CKINVDCx5p33_ASAP7_75t_R g5190 ( 
.A(n_4049),
.Y(n_5190)
);

CKINVDCx5p33_ASAP7_75t_R g5191 ( 
.A(n_1436),
.Y(n_5191)
);

CKINVDCx5p33_ASAP7_75t_R g5192 ( 
.A(n_2873),
.Y(n_5192)
);

INVx1_ASAP7_75t_L g5193 ( 
.A(n_334),
.Y(n_5193)
);

CKINVDCx5p33_ASAP7_75t_R g5194 ( 
.A(n_4070),
.Y(n_5194)
);

INVxp67_ASAP7_75t_L g5195 ( 
.A(n_1347),
.Y(n_5195)
);

CKINVDCx5p33_ASAP7_75t_R g5196 ( 
.A(n_3151),
.Y(n_5196)
);

CKINVDCx5p33_ASAP7_75t_R g5197 ( 
.A(n_3892),
.Y(n_5197)
);

CKINVDCx5p33_ASAP7_75t_R g5198 ( 
.A(n_2773),
.Y(n_5198)
);

CKINVDCx5p33_ASAP7_75t_R g5199 ( 
.A(n_797),
.Y(n_5199)
);

CKINVDCx5p33_ASAP7_75t_R g5200 ( 
.A(n_1558),
.Y(n_5200)
);

CKINVDCx5p33_ASAP7_75t_R g5201 ( 
.A(n_2884),
.Y(n_5201)
);

CKINVDCx5p33_ASAP7_75t_R g5202 ( 
.A(n_493),
.Y(n_5202)
);

CKINVDCx5p33_ASAP7_75t_R g5203 ( 
.A(n_1893),
.Y(n_5203)
);

CKINVDCx5p33_ASAP7_75t_R g5204 ( 
.A(n_3607),
.Y(n_5204)
);

CKINVDCx16_ASAP7_75t_R g5205 ( 
.A(n_273),
.Y(n_5205)
);

BUFx10_ASAP7_75t_L g5206 ( 
.A(n_2560),
.Y(n_5206)
);

INVx1_ASAP7_75t_L g5207 ( 
.A(n_455),
.Y(n_5207)
);

CKINVDCx5p33_ASAP7_75t_R g5208 ( 
.A(n_610),
.Y(n_5208)
);

CKINVDCx5p33_ASAP7_75t_R g5209 ( 
.A(n_4210),
.Y(n_5209)
);

CKINVDCx5p33_ASAP7_75t_R g5210 ( 
.A(n_1432),
.Y(n_5210)
);

CKINVDCx20_ASAP7_75t_R g5211 ( 
.A(n_4258),
.Y(n_5211)
);

INVx1_ASAP7_75t_SL g5212 ( 
.A(n_3058),
.Y(n_5212)
);

CKINVDCx5p33_ASAP7_75t_R g5213 ( 
.A(n_3558),
.Y(n_5213)
);

BUFx2_ASAP7_75t_L g5214 ( 
.A(n_2040),
.Y(n_5214)
);

CKINVDCx5p33_ASAP7_75t_R g5215 ( 
.A(n_3565),
.Y(n_5215)
);

CKINVDCx5p33_ASAP7_75t_R g5216 ( 
.A(n_1731),
.Y(n_5216)
);

INVx1_ASAP7_75t_L g5217 ( 
.A(n_2039),
.Y(n_5217)
);

BUFx10_ASAP7_75t_L g5218 ( 
.A(n_3268),
.Y(n_5218)
);

CKINVDCx5p33_ASAP7_75t_R g5219 ( 
.A(n_557),
.Y(n_5219)
);

BUFx10_ASAP7_75t_L g5220 ( 
.A(n_994),
.Y(n_5220)
);

CKINVDCx5p33_ASAP7_75t_R g5221 ( 
.A(n_2008),
.Y(n_5221)
);

CKINVDCx5p33_ASAP7_75t_R g5222 ( 
.A(n_2142),
.Y(n_5222)
);

CKINVDCx5p33_ASAP7_75t_R g5223 ( 
.A(n_964),
.Y(n_5223)
);

CKINVDCx5p33_ASAP7_75t_R g5224 ( 
.A(n_2012),
.Y(n_5224)
);

CKINVDCx5p33_ASAP7_75t_R g5225 ( 
.A(n_4315),
.Y(n_5225)
);

CKINVDCx5p33_ASAP7_75t_R g5226 ( 
.A(n_4016),
.Y(n_5226)
);

CKINVDCx5p33_ASAP7_75t_R g5227 ( 
.A(n_1130),
.Y(n_5227)
);

INVx1_ASAP7_75t_L g5228 ( 
.A(n_169),
.Y(n_5228)
);

CKINVDCx5p33_ASAP7_75t_R g5229 ( 
.A(n_1536),
.Y(n_5229)
);

INVx1_ASAP7_75t_L g5230 ( 
.A(n_4061),
.Y(n_5230)
);

CKINVDCx5p33_ASAP7_75t_R g5231 ( 
.A(n_4116),
.Y(n_5231)
);

CKINVDCx5p33_ASAP7_75t_R g5232 ( 
.A(n_2520),
.Y(n_5232)
);

INVx1_ASAP7_75t_L g5233 ( 
.A(n_219),
.Y(n_5233)
);

CKINVDCx5p33_ASAP7_75t_R g5234 ( 
.A(n_3858),
.Y(n_5234)
);

BUFx6f_ASAP7_75t_L g5235 ( 
.A(n_2607),
.Y(n_5235)
);

INVx1_ASAP7_75t_L g5236 ( 
.A(n_3079),
.Y(n_5236)
);

CKINVDCx5p33_ASAP7_75t_R g5237 ( 
.A(n_2668),
.Y(n_5237)
);

CKINVDCx5p33_ASAP7_75t_R g5238 ( 
.A(n_1280),
.Y(n_5238)
);

INVx1_ASAP7_75t_L g5239 ( 
.A(n_1212),
.Y(n_5239)
);

INVx2_ASAP7_75t_L g5240 ( 
.A(n_1964),
.Y(n_5240)
);

CKINVDCx5p33_ASAP7_75t_R g5241 ( 
.A(n_1976),
.Y(n_5241)
);

INVx1_ASAP7_75t_L g5242 ( 
.A(n_3788),
.Y(n_5242)
);

INVx1_ASAP7_75t_L g5243 ( 
.A(n_2733),
.Y(n_5243)
);

BUFx8_ASAP7_75t_SL g5244 ( 
.A(n_1355),
.Y(n_5244)
);

INVx2_ASAP7_75t_SL g5245 ( 
.A(n_2855),
.Y(n_5245)
);

CKINVDCx5p33_ASAP7_75t_R g5246 ( 
.A(n_3135),
.Y(n_5246)
);

CKINVDCx5p33_ASAP7_75t_R g5247 ( 
.A(n_2977),
.Y(n_5247)
);

CKINVDCx5p33_ASAP7_75t_R g5248 ( 
.A(n_354),
.Y(n_5248)
);

INVx1_ASAP7_75t_L g5249 ( 
.A(n_401),
.Y(n_5249)
);

INVx1_ASAP7_75t_L g5250 ( 
.A(n_4097),
.Y(n_5250)
);

INVx1_ASAP7_75t_L g5251 ( 
.A(n_1895),
.Y(n_5251)
);

CKINVDCx5p33_ASAP7_75t_R g5252 ( 
.A(n_3259),
.Y(n_5252)
);

INVx1_ASAP7_75t_L g5253 ( 
.A(n_516),
.Y(n_5253)
);

BUFx2_ASAP7_75t_SL g5254 ( 
.A(n_3075),
.Y(n_5254)
);

BUFx6f_ASAP7_75t_L g5255 ( 
.A(n_937),
.Y(n_5255)
);

CKINVDCx5p33_ASAP7_75t_R g5256 ( 
.A(n_627),
.Y(n_5256)
);

CKINVDCx20_ASAP7_75t_R g5257 ( 
.A(n_3513),
.Y(n_5257)
);

CKINVDCx5p33_ASAP7_75t_R g5258 ( 
.A(n_203),
.Y(n_5258)
);

CKINVDCx5p33_ASAP7_75t_R g5259 ( 
.A(n_833),
.Y(n_5259)
);

CKINVDCx5p33_ASAP7_75t_R g5260 ( 
.A(n_1967),
.Y(n_5260)
);

INVx1_ASAP7_75t_L g5261 ( 
.A(n_3046),
.Y(n_5261)
);

INVx1_ASAP7_75t_L g5262 ( 
.A(n_3742),
.Y(n_5262)
);

INVx1_ASAP7_75t_L g5263 ( 
.A(n_1720),
.Y(n_5263)
);

INVx1_ASAP7_75t_L g5264 ( 
.A(n_1942),
.Y(n_5264)
);

INVx1_ASAP7_75t_SL g5265 ( 
.A(n_4222),
.Y(n_5265)
);

CKINVDCx20_ASAP7_75t_R g5266 ( 
.A(n_1830),
.Y(n_5266)
);

INVx1_ASAP7_75t_L g5267 ( 
.A(n_265),
.Y(n_5267)
);

CKINVDCx5p33_ASAP7_75t_R g5268 ( 
.A(n_841),
.Y(n_5268)
);

CKINVDCx5p33_ASAP7_75t_R g5269 ( 
.A(n_3629),
.Y(n_5269)
);

INVx1_ASAP7_75t_L g5270 ( 
.A(n_409),
.Y(n_5270)
);

CKINVDCx5p33_ASAP7_75t_R g5271 ( 
.A(n_4078),
.Y(n_5271)
);

INVx2_ASAP7_75t_L g5272 ( 
.A(n_2655),
.Y(n_5272)
);

CKINVDCx16_ASAP7_75t_R g5273 ( 
.A(n_2709),
.Y(n_5273)
);

CKINVDCx5p33_ASAP7_75t_R g5274 ( 
.A(n_2639),
.Y(n_5274)
);

CKINVDCx5p33_ASAP7_75t_R g5275 ( 
.A(n_1547),
.Y(n_5275)
);

CKINVDCx5p33_ASAP7_75t_R g5276 ( 
.A(n_4131),
.Y(n_5276)
);

CKINVDCx5p33_ASAP7_75t_R g5277 ( 
.A(n_2678),
.Y(n_5277)
);

CKINVDCx5p33_ASAP7_75t_R g5278 ( 
.A(n_3584),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_3157),
.Y(n_5279)
);

CKINVDCx5p33_ASAP7_75t_R g5280 ( 
.A(n_1831),
.Y(n_5280)
);

INVx1_ASAP7_75t_L g5281 ( 
.A(n_1165),
.Y(n_5281)
);

CKINVDCx5p33_ASAP7_75t_R g5282 ( 
.A(n_3690),
.Y(n_5282)
);

CKINVDCx5p33_ASAP7_75t_R g5283 ( 
.A(n_1264),
.Y(n_5283)
);

CKINVDCx5p33_ASAP7_75t_R g5284 ( 
.A(n_3651),
.Y(n_5284)
);

BUFx2_ASAP7_75t_SL g5285 ( 
.A(n_954),
.Y(n_5285)
);

CKINVDCx5p33_ASAP7_75t_R g5286 ( 
.A(n_1420),
.Y(n_5286)
);

CKINVDCx5p33_ASAP7_75t_R g5287 ( 
.A(n_3982),
.Y(n_5287)
);

INVx1_ASAP7_75t_L g5288 ( 
.A(n_3821),
.Y(n_5288)
);

INVx2_ASAP7_75t_L g5289 ( 
.A(n_4205),
.Y(n_5289)
);

INVx1_ASAP7_75t_L g5290 ( 
.A(n_2912),
.Y(n_5290)
);

CKINVDCx16_ASAP7_75t_R g5291 ( 
.A(n_1840),
.Y(n_5291)
);

CKINVDCx5p33_ASAP7_75t_R g5292 ( 
.A(n_239),
.Y(n_5292)
);

BUFx5_ASAP7_75t_L g5293 ( 
.A(n_664),
.Y(n_5293)
);

CKINVDCx5p33_ASAP7_75t_R g5294 ( 
.A(n_3391),
.Y(n_5294)
);

CKINVDCx5p33_ASAP7_75t_R g5295 ( 
.A(n_1753),
.Y(n_5295)
);

CKINVDCx5p33_ASAP7_75t_R g5296 ( 
.A(n_1994),
.Y(n_5296)
);

INVx1_ASAP7_75t_L g5297 ( 
.A(n_1995),
.Y(n_5297)
);

CKINVDCx5p33_ASAP7_75t_R g5298 ( 
.A(n_4262),
.Y(n_5298)
);

CKINVDCx5p33_ASAP7_75t_R g5299 ( 
.A(n_4124),
.Y(n_5299)
);

HB1xp67_ASAP7_75t_L g5300 ( 
.A(n_518),
.Y(n_5300)
);

CKINVDCx5p33_ASAP7_75t_R g5301 ( 
.A(n_3756),
.Y(n_5301)
);

INVx1_ASAP7_75t_L g5302 ( 
.A(n_4048),
.Y(n_5302)
);

INVx1_ASAP7_75t_L g5303 ( 
.A(n_2819),
.Y(n_5303)
);

CKINVDCx5p33_ASAP7_75t_R g5304 ( 
.A(n_1828),
.Y(n_5304)
);

BUFx2_ASAP7_75t_L g5305 ( 
.A(n_512),
.Y(n_5305)
);

CKINVDCx16_ASAP7_75t_R g5306 ( 
.A(n_4058),
.Y(n_5306)
);

INVx1_ASAP7_75t_L g5307 ( 
.A(n_2085),
.Y(n_5307)
);

CKINVDCx5p33_ASAP7_75t_R g5308 ( 
.A(n_1431),
.Y(n_5308)
);

INVx1_ASAP7_75t_SL g5309 ( 
.A(n_4178),
.Y(n_5309)
);

CKINVDCx5p33_ASAP7_75t_R g5310 ( 
.A(n_1760),
.Y(n_5310)
);

INVx1_ASAP7_75t_SL g5311 ( 
.A(n_3615),
.Y(n_5311)
);

INVx1_ASAP7_75t_L g5312 ( 
.A(n_3773),
.Y(n_5312)
);

INVx1_ASAP7_75t_L g5313 ( 
.A(n_1079),
.Y(n_5313)
);

CKINVDCx5p33_ASAP7_75t_R g5314 ( 
.A(n_828),
.Y(n_5314)
);

INVxp67_ASAP7_75t_L g5315 ( 
.A(n_1133),
.Y(n_5315)
);

INVx1_ASAP7_75t_L g5316 ( 
.A(n_2432),
.Y(n_5316)
);

CKINVDCx5p33_ASAP7_75t_R g5317 ( 
.A(n_2109),
.Y(n_5317)
);

INVx2_ASAP7_75t_L g5318 ( 
.A(n_1367),
.Y(n_5318)
);

INVx1_ASAP7_75t_L g5319 ( 
.A(n_2514),
.Y(n_5319)
);

CKINVDCx5p33_ASAP7_75t_R g5320 ( 
.A(n_2775),
.Y(n_5320)
);

BUFx10_ASAP7_75t_L g5321 ( 
.A(n_2214),
.Y(n_5321)
);

INVx1_ASAP7_75t_L g5322 ( 
.A(n_1425),
.Y(n_5322)
);

BUFx6f_ASAP7_75t_L g5323 ( 
.A(n_3314),
.Y(n_5323)
);

BUFx6f_ASAP7_75t_L g5324 ( 
.A(n_1076),
.Y(n_5324)
);

CKINVDCx5p33_ASAP7_75t_R g5325 ( 
.A(n_2095),
.Y(n_5325)
);

CKINVDCx5p33_ASAP7_75t_R g5326 ( 
.A(n_4118),
.Y(n_5326)
);

CKINVDCx5p33_ASAP7_75t_R g5327 ( 
.A(n_2033),
.Y(n_5327)
);

CKINVDCx5p33_ASAP7_75t_R g5328 ( 
.A(n_1433),
.Y(n_5328)
);

INVx1_ASAP7_75t_SL g5329 ( 
.A(n_615),
.Y(n_5329)
);

INVx1_ASAP7_75t_L g5330 ( 
.A(n_754),
.Y(n_5330)
);

CKINVDCx5p33_ASAP7_75t_R g5331 ( 
.A(n_1254),
.Y(n_5331)
);

CKINVDCx5p33_ASAP7_75t_R g5332 ( 
.A(n_2435),
.Y(n_5332)
);

CKINVDCx5p33_ASAP7_75t_R g5333 ( 
.A(n_2287),
.Y(n_5333)
);

CKINVDCx5p33_ASAP7_75t_R g5334 ( 
.A(n_890),
.Y(n_5334)
);

INVx1_ASAP7_75t_L g5335 ( 
.A(n_4066),
.Y(n_5335)
);

INVx1_ASAP7_75t_L g5336 ( 
.A(n_3545),
.Y(n_5336)
);

BUFx2_ASAP7_75t_L g5337 ( 
.A(n_1814),
.Y(n_5337)
);

CKINVDCx20_ASAP7_75t_R g5338 ( 
.A(n_2795),
.Y(n_5338)
);

INVx1_ASAP7_75t_L g5339 ( 
.A(n_2436),
.Y(n_5339)
);

CKINVDCx5p33_ASAP7_75t_R g5340 ( 
.A(n_2603),
.Y(n_5340)
);

INVx1_ASAP7_75t_SL g5341 ( 
.A(n_3165),
.Y(n_5341)
);

HB1xp67_ASAP7_75t_L g5342 ( 
.A(n_1188),
.Y(n_5342)
);

CKINVDCx5p33_ASAP7_75t_R g5343 ( 
.A(n_1548),
.Y(n_5343)
);

INVx1_ASAP7_75t_L g5344 ( 
.A(n_4211),
.Y(n_5344)
);

INVx1_ASAP7_75t_L g5345 ( 
.A(n_3107),
.Y(n_5345)
);

INVx1_ASAP7_75t_L g5346 ( 
.A(n_2079),
.Y(n_5346)
);

INVx1_ASAP7_75t_L g5347 ( 
.A(n_4122),
.Y(n_5347)
);

CKINVDCx20_ASAP7_75t_R g5348 ( 
.A(n_4163),
.Y(n_5348)
);

CKINVDCx5p33_ASAP7_75t_R g5349 ( 
.A(n_2445),
.Y(n_5349)
);

CKINVDCx5p33_ASAP7_75t_R g5350 ( 
.A(n_325),
.Y(n_5350)
);

CKINVDCx5p33_ASAP7_75t_R g5351 ( 
.A(n_729),
.Y(n_5351)
);

CKINVDCx5p33_ASAP7_75t_R g5352 ( 
.A(n_4086),
.Y(n_5352)
);

INVx1_ASAP7_75t_L g5353 ( 
.A(n_3163),
.Y(n_5353)
);

INVx1_ASAP7_75t_L g5354 ( 
.A(n_1529),
.Y(n_5354)
);

CKINVDCx20_ASAP7_75t_R g5355 ( 
.A(n_3518),
.Y(n_5355)
);

CKINVDCx5p33_ASAP7_75t_R g5356 ( 
.A(n_3123),
.Y(n_5356)
);

CKINVDCx5p33_ASAP7_75t_R g5357 ( 
.A(n_4099),
.Y(n_5357)
);

CKINVDCx5p33_ASAP7_75t_R g5358 ( 
.A(n_3411),
.Y(n_5358)
);

CKINVDCx5p33_ASAP7_75t_R g5359 ( 
.A(n_522),
.Y(n_5359)
);

INVx1_ASAP7_75t_L g5360 ( 
.A(n_3350),
.Y(n_5360)
);

CKINVDCx5p33_ASAP7_75t_R g5361 ( 
.A(n_3306),
.Y(n_5361)
);

BUFx3_ASAP7_75t_L g5362 ( 
.A(n_4163),
.Y(n_5362)
);

CKINVDCx5p33_ASAP7_75t_R g5363 ( 
.A(n_977),
.Y(n_5363)
);

INVx1_ASAP7_75t_L g5364 ( 
.A(n_4144),
.Y(n_5364)
);

CKINVDCx5p33_ASAP7_75t_R g5365 ( 
.A(n_1148),
.Y(n_5365)
);

CKINVDCx5p33_ASAP7_75t_R g5366 ( 
.A(n_564),
.Y(n_5366)
);

BUFx2_ASAP7_75t_L g5367 ( 
.A(n_4143),
.Y(n_5367)
);

CKINVDCx5p33_ASAP7_75t_R g5368 ( 
.A(n_2237),
.Y(n_5368)
);

CKINVDCx5p33_ASAP7_75t_R g5369 ( 
.A(n_3503),
.Y(n_5369)
);

CKINVDCx5p33_ASAP7_75t_R g5370 ( 
.A(n_2294),
.Y(n_5370)
);

INVx1_ASAP7_75t_L g5371 ( 
.A(n_3697),
.Y(n_5371)
);

BUFx10_ASAP7_75t_L g5372 ( 
.A(n_1739),
.Y(n_5372)
);

INVx1_ASAP7_75t_L g5373 ( 
.A(n_4224),
.Y(n_5373)
);

INVx1_ASAP7_75t_L g5374 ( 
.A(n_1113),
.Y(n_5374)
);

CKINVDCx5p33_ASAP7_75t_R g5375 ( 
.A(n_204),
.Y(n_5375)
);

CKINVDCx5p33_ASAP7_75t_R g5376 ( 
.A(n_3628),
.Y(n_5376)
);

INVx1_ASAP7_75t_L g5377 ( 
.A(n_2191),
.Y(n_5377)
);

CKINVDCx20_ASAP7_75t_R g5378 ( 
.A(n_3947),
.Y(n_5378)
);

CKINVDCx5p33_ASAP7_75t_R g5379 ( 
.A(n_2947),
.Y(n_5379)
);

CKINVDCx5p33_ASAP7_75t_R g5380 ( 
.A(n_2024),
.Y(n_5380)
);

INVx1_ASAP7_75t_L g5381 ( 
.A(n_3862),
.Y(n_5381)
);

INVx1_ASAP7_75t_L g5382 ( 
.A(n_3325),
.Y(n_5382)
);

CKINVDCx5p33_ASAP7_75t_R g5383 ( 
.A(n_1639),
.Y(n_5383)
);

INVx1_ASAP7_75t_L g5384 ( 
.A(n_3232),
.Y(n_5384)
);

CKINVDCx5p33_ASAP7_75t_R g5385 ( 
.A(n_2114),
.Y(n_5385)
);

CKINVDCx20_ASAP7_75t_R g5386 ( 
.A(n_538),
.Y(n_5386)
);

INVx1_ASAP7_75t_L g5387 ( 
.A(n_3945),
.Y(n_5387)
);

INVx1_ASAP7_75t_L g5388 ( 
.A(n_1239),
.Y(n_5388)
);

CKINVDCx16_ASAP7_75t_R g5389 ( 
.A(n_3206),
.Y(n_5389)
);

HB1xp67_ASAP7_75t_L g5390 ( 
.A(n_4180),
.Y(n_5390)
);

CKINVDCx5p33_ASAP7_75t_R g5391 ( 
.A(n_4050),
.Y(n_5391)
);

CKINVDCx5p33_ASAP7_75t_R g5392 ( 
.A(n_2521),
.Y(n_5392)
);

CKINVDCx5p33_ASAP7_75t_R g5393 ( 
.A(n_461),
.Y(n_5393)
);

INVx2_ASAP7_75t_L g5394 ( 
.A(n_3905),
.Y(n_5394)
);

CKINVDCx5p33_ASAP7_75t_R g5395 ( 
.A(n_3353),
.Y(n_5395)
);

CKINVDCx5p33_ASAP7_75t_R g5396 ( 
.A(n_1373),
.Y(n_5396)
);

CKINVDCx20_ASAP7_75t_R g5397 ( 
.A(n_3032),
.Y(n_5397)
);

CKINVDCx5p33_ASAP7_75t_R g5398 ( 
.A(n_1846),
.Y(n_5398)
);

CKINVDCx5p33_ASAP7_75t_R g5399 ( 
.A(n_4069),
.Y(n_5399)
);

CKINVDCx5p33_ASAP7_75t_R g5400 ( 
.A(n_3815),
.Y(n_5400)
);

CKINVDCx5p33_ASAP7_75t_R g5401 ( 
.A(n_4247),
.Y(n_5401)
);

INVx1_ASAP7_75t_SL g5402 ( 
.A(n_2322),
.Y(n_5402)
);

CKINVDCx5p33_ASAP7_75t_R g5403 ( 
.A(n_2215),
.Y(n_5403)
);

INVx1_ASAP7_75t_L g5404 ( 
.A(n_2763),
.Y(n_5404)
);

CKINVDCx20_ASAP7_75t_R g5405 ( 
.A(n_3880),
.Y(n_5405)
);

BUFx2_ASAP7_75t_L g5406 ( 
.A(n_1785),
.Y(n_5406)
);

HB1xp67_ASAP7_75t_L g5407 ( 
.A(n_2557),
.Y(n_5407)
);

CKINVDCx5p33_ASAP7_75t_R g5408 ( 
.A(n_3761),
.Y(n_5408)
);

CKINVDCx5p33_ASAP7_75t_R g5409 ( 
.A(n_3102),
.Y(n_5409)
);

INVx1_ASAP7_75t_L g5410 ( 
.A(n_1492),
.Y(n_5410)
);

INVx2_ASAP7_75t_L g5411 ( 
.A(n_2797),
.Y(n_5411)
);

BUFx5_ASAP7_75t_L g5412 ( 
.A(n_2760),
.Y(n_5412)
);

CKINVDCx5p33_ASAP7_75t_R g5413 ( 
.A(n_4023),
.Y(n_5413)
);

BUFx6f_ASAP7_75t_L g5414 ( 
.A(n_1768),
.Y(n_5414)
);

CKINVDCx5p33_ASAP7_75t_R g5415 ( 
.A(n_4185),
.Y(n_5415)
);

INVx1_ASAP7_75t_L g5416 ( 
.A(n_1810),
.Y(n_5416)
);

INVx1_ASAP7_75t_L g5417 ( 
.A(n_3832),
.Y(n_5417)
);

INVx2_ASAP7_75t_L g5418 ( 
.A(n_3114),
.Y(n_5418)
);

INVx1_ASAP7_75t_L g5419 ( 
.A(n_2983),
.Y(n_5419)
);

CKINVDCx5p33_ASAP7_75t_R g5420 ( 
.A(n_4128),
.Y(n_5420)
);

CKINVDCx5p33_ASAP7_75t_R g5421 ( 
.A(n_724),
.Y(n_5421)
);

BUFx3_ASAP7_75t_L g5422 ( 
.A(n_4114),
.Y(n_5422)
);

CKINVDCx5p33_ASAP7_75t_R g5423 ( 
.A(n_1801),
.Y(n_5423)
);

CKINVDCx5p33_ASAP7_75t_R g5424 ( 
.A(n_2708),
.Y(n_5424)
);

CKINVDCx5p33_ASAP7_75t_R g5425 ( 
.A(n_690),
.Y(n_5425)
);

CKINVDCx5p33_ASAP7_75t_R g5426 ( 
.A(n_1159),
.Y(n_5426)
);

CKINVDCx5p33_ASAP7_75t_R g5427 ( 
.A(n_3593),
.Y(n_5427)
);

CKINVDCx5p33_ASAP7_75t_R g5428 ( 
.A(n_2253),
.Y(n_5428)
);

CKINVDCx5p33_ASAP7_75t_R g5429 ( 
.A(n_864),
.Y(n_5429)
);

INVx1_ASAP7_75t_L g5430 ( 
.A(n_2275),
.Y(n_5430)
);

CKINVDCx5p33_ASAP7_75t_R g5431 ( 
.A(n_4172),
.Y(n_5431)
);

CKINVDCx5p33_ASAP7_75t_R g5432 ( 
.A(n_930),
.Y(n_5432)
);

INVx1_ASAP7_75t_L g5433 ( 
.A(n_346),
.Y(n_5433)
);

INVx1_ASAP7_75t_L g5434 ( 
.A(n_302),
.Y(n_5434)
);

CKINVDCx20_ASAP7_75t_R g5435 ( 
.A(n_2275),
.Y(n_5435)
);

INVx2_ASAP7_75t_L g5436 ( 
.A(n_4225),
.Y(n_5436)
);

INVx1_ASAP7_75t_L g5437 ( 
.A(n_3691),
.Y(n_5437)
);

INVx2_ASAP7_75t_SL g5438 ( 
.A(n_2062),
.Y(n_5438)
);

CKINVDCx5p33_ASAP7_75t_R g5439 ( 
.A(n_2662),
.Y(n_5439)
);

CKINVDCx20_ASAP7_75t_R g5440 ( 
.A(n_2061),
.Y(n_5440)
);

INVx1_ASAP7_75t_L g5441 ( 
.A(n_734),
.Y(n_5441)
);

CKINVDCx5p33_ASAP7_75t_R g5442 ( 
.A(n_3617),
.Y(n_5442)
);

CKINVDCx5p33_ASAP7_75t_R g5443 ( 
.A(n_3082),
.Y(n_5443)
);

CKINVDCx5p33_ASAP7_75t_R g5444 ( 
.A(n_3443),
.Y(n_5444)
);

CKINVDCx5p33_ASAP7_75t_R g5445 ( 
.A(n_1971),
.Y(n_5445)
);

BUFx6f_ASAP7_75t_L g5446 ( 
.A(n_554),
.Y(n_5446)
);

INVx1_ASAP7_75t_SL g5447 ( 
.A(n_1055),
.Y(n_5447)
);

CKINVDCx5p33_ASAP7_75t_R g5448 ( 
.A(n_2080),
.Y(n_5448)
);

INVx1_ASAP7_75t_L g5449 ( 
.A(n_395),
.Y(n_5449)
);

INVx3_ASAP7_75t_L g5450 ( 
.A(n_3342),
.Y(n_5450)
);

INVx1_ASAP7_75t_L g5451 ( 
.A(n_3510),
.Y(n_5451)
);

INVx1_ASAP7_75t_L g5452 ( 
.A(n_3175),
.Y(n_5452)
);

INVx2_ASAP7_75t_L g5453 ( 
.A(n_2279),
.Y(n_5453)
);

CKINVDCx5p33_ASAP7_75t_R g5454 ( 
.A(n_3565),
.Y(n_5454)
);

INVx1_ASAP7_75t_L g5455 ( 
.A(n_2246),
.Y(n_5455)
);

CKINVDCx20_ASAP7_75t_R g5456 ( 
.A(n_3914),
.Y(n_5456)
);

INVx1_ASAP7_75t_L g5457 ( 
.A(n_4134),
.Y(n_5457)
);

CKINVDCx5p33_ASAP7_75t_R g5458 ( 
.A(n_1251),
.Y(n_5458)
);

CKINVDCx5p33_ASAP7_75t_R g5459 ( 
.A(n_3701),
.Y(n_5459)
);

CKINVDCx5p33_ASAP7_75t_R g5460 ( 
.A(n_2919),
.Y(n_5460)
);

INVx1_ASAP7_75t_L g5461 ( 
.A(n_2774),
.Y(n_5461)
);

INVx1_ASAP7_75t_L g5462 ( 
.A(n_2620),
.Y(n_5462)
);

CKINVDCx5p33_ASAP7_75t_R g5463 ( 
.A(n_720),
.Y(n_5463)
);

CKINVDCx5p33_ASAP7_75t_R g5464 ( 
.A(n_3650),
.Y(n_5464)
);

CKINVDCx20_ASAP7_75t_R g5465 ( 
.A(n_2369),
.Y(n_5465)
);

BUFx2_ASAP7_75t_L g5466 ( 
.A(n_543),
.Y(n_5466)
);

INVx1_ASAP7_75t_SL g5467 ( 
.A(n_2003),
.Y(n_5467)
);

CKINVDCx5p33_ASAP7_75t_R g5468 ( 
.A(n_4232),
.Y(n_5468)
);

CKINVDCx5p33_ASAP7_75t_R g5469 ( 
.A(n_2115),
.Y(n_5469)
);

BUFx6f_ASAP7_75t_L g5470 ( 
.A(n_370),
.Y(n_5470)
);

CKINVDCx5p33_ASAP7_75t_R g5471 ( 
.A(n_4200),
.Y(n_5471)
);

CKINVDCx6p67_ASAP7_75t_R g5472 ( 
.A(n_4277),
.Y(n_5472)
);

CKINVDCx5p33_ASAP7_75t_R g5473 ( 
.A(n_2904),
.Y(n_5473)
);

CKINVDCx5p33_ASAP7_75t_R g5474 ( 
.A(n_3737),
.Y(n_5474)
);

INVx1_ASAP7_75t_L g5475 ( 
.A(n_4215),
.Y(n_5475)
);

BUFx10_ASAP7_75t_L g5476 ( 
.A(n_1912),
.Y(n_5476)
);

CKINVDCx5p33_ASAP7_75t_R g5477 ( 
.A(n_2027),
.Y(n_5477)
);

INVx1_ASAP7_75t_L g5478 ( 
.A(n_3527),
.Y(n_5478)
);

CKINVDCx20_ASAP7_75t_R g5479 ( 
.A(n_3402),
.Y(n_5479)
);

CKINVDCx5p33_ASAP7_75t_R g5480 ( 
.A(n_3957),
.Y(n_5480)
);

INVx2_ASAP7_75t_L g5481 ( 
.A(n_365),
.Y(n_5481)
);

INVx1_ASAP7_75t_L g5482 ( 
.A(n_50),
.Y(n_5482)
);

CKINVDCx5p33_ASAP7_75t_R g5483 ( 
.A(n_1543),
.Y(n_5483)
);

CKINVDCx5p33_ASAP7_75t_R g5484 ( 
.A(n_16),
.Y(n_5484)
);

CKINVDCx20_ASAP7_75t_R g5485 ( 
.A(n_49),
.Y(n_5485)
);

INVx1_ASAP7_75t_L g5486 ( 
.A(n_241),
.Y(n_5486)
);

INVx1_ASAP7_75t_L g5487 ( 
.A(n_4212),
.Y(n_5487)
);

CKINVDCx5p33_ASAP7_75t_R g5488 ( 
.A(n_1495),
.Y(n_5488)
);

CKINVDCx5p33_ASAP7_75t_R g5489 ( 
.A(n_2478),
.Y(n_5489)
);

CKINVDCx5p33_ASAP7_75t_R g5490 ( 
.A(n_976),
.Y(n_5490)
);

CKINVDCx5p33_ASAP7_75t_R g5491 ( 
.A(n_3455),
.Y(n_5491)
);

CKINVDCx5p33_ASAP7_75t_R g5492 ( 
.A(n_2659),
.Y(n_5492)
);

INVx1_ASAP7_75t_L g5493 ( 
.A(n_4091),
.Y(n_5493)
);

CKINVDCx20_ASAP7_75t_R g5494 ( 
.A(n_3141),
.Y(n_5494)
);

CKINVDCx5p33_ASAP7_75t_R g5495 ( 
.A(n_3890),
.Y(n_5495)
);

INVx2_ASAP7_75t_SL g5496 ( 
.A(n_4106),
.Y(n_5496)
);

CKINVDCx5p33_ASAP7_75t_R g5497 ( 
.A(n_4132),
.Y(n_5497)
);

INVx1_ASAP7_75t_L g5498 ( 
.A(n_2188),
.Y(n_5498)
);

CKINVDCx20_ASAP7_75t_R g5499 ( 
.A(n_1538),
.Y(n_5499)
);

INVx1_ASAP7_75t_L g5500 ( 
.A(n_1405),
.Y(n_5500)
);

BUFx3_ASAP7_75t_L g5501 ( 
.A(n_2832),
.Y(n_5501)
);

INVx1_ASAP7_75t_L g5502 ( 
.A(n_1676),
.Y(n_5502)
);

BUFx3_ASAP7_75t_L g5503 ( 
.A(n_3109),
.Y(n_5503)
);

CKINVDCx5p33_ASAP7_75t_R g5504 ( 
.A(n_1690),
.Y(n_5504)
);

INVx1_ASAP7_75t_L g5505 ( 
.A(n_1682),
.Y(n_5505)
);

INVx1_ASAP7_75t_L g5506 ( 
.A(n_492),
.Y(n_5506)
);

INVx1_ASAP7_75t_L g5507 ( 
.A(n_1295),
.Y(n_5507)
);

INVx1_ASAP7_75t_SL g5508 ( 
.A(n_1311),
.Y(n_5508)
);

INVx2_ASAP7_75t_SL g5509 ( 
.A(n_2567),
.Y(n_5509)
);

CKINVDCx5p33_ASAP7_75t_R g5510 ( 
.A(n_1181),
.Y(n_5510)
);

CKINVDCx5p33_ASAP7_75t_R g5511 ( 
.A(n_1317),
.Y(n_5511)
);

CKINVDCx5p33_ASAP7_75t_R g5512 ( 
.A(n_507),
.Y(n_5512)
);

CKINVDCx20_ASAP7_75t_R g5513 ( 
.A(n_1635),
.Y(n_5513)
);

BUFx6f_ASAP7_75t_L g5514 ( 
.A(n_418),
.Y(n_5514)
);

INVx1_ASAP7_75t_L g5515 ( 
.A(n_481),
.Y(n_5515)
);

CKINVDCx20_ASAP7_75t_R g5516 ( 
.A(n_1219),
.Y(n_5516)
);

CKINVDCx5p33_ASAP7_75t_R g5517 ( 
.A(n_4085),
.Y(n_5517)
);

CKINVDCx20_ASAP7_75t_R g5518 ( 
.A(n_2835),
.Y(n_5518)
);

CKINVDCx5p33_ASAP7_75t_R g5519 ( 
.A(n_1932),
.Y(n_5519)
);

INVx1_ASAP7_75t_L g5520 ( 
.A(n_3440),
.Y(n_5520)
);

BUFx6f_ASAP7_75t_L g5521 ( 
.A(n_3236),
.Y(n_5521)
);

INVx1_ASAP7_75t_L g5522 ( 
.A(n_2466),
.Y(n_5522)
);

INVx1_ASAP7_75t_SL g5523 ( 
.A(n_3167),
.Y(n_5523)
);

INVx1_ASAP7_75t_L g5524 ( 
.A(n_4223),
.Y(n_5524)
);

CKINVDCx5p33_ASAP7_75t_R g5525 ( 
.A(n_4079),
.Y(n_5525)
);

CKINVDCx5p33_ASAP7_75t_R g5526 ( 
.A(n_3467),
.Y(n_5526)
);

BUFx6f_ASAP7_75t_L g5527 ( 
.A(n_4160),
.Y(n_5527)
);

HB1xp67_ASAP7_75t_L g5528 ( 
.A(n_2019),
.Y(n_5528)
);

CKINVDCx5p33_ASAP7_75t_R g5529 ( 
.A(n_1645),
.Y(n_5529)
);

INVx1_ASAP7_75t_SL g5530 ( 
.A(n_4093),
.Y(n_5530)
);

CKINVDCx5p33_ASAP7_75t_R g5531 ( 
.A(n_4199),
.Y(n_5531)
);

CKINVDCx5p33_ASAP7_75t_R g5532 ( 
.A(n_1035),
.Y(n_5532)
);

CKINVDCx5p33_ASAP7_75t_R g5533 ( 
.A(n_3707),
.Y(n_5533)
);

CKINVDCx5p33_ASAP7_75t_R g5534 ( 
.A(n_1614),
.Y(n_5534)
);

INVx1_ASAP7_75t_L g5535 ( 
.A(n_2931),
.Y(n_5535)
);

BUFx3_ASAP7_75t_L g5536 ( 
.A(n_2786),
.Y(n_5536)
);

CKINVDCx5p33_ASAP7_75t_R g5537 ( 
.A(n_61),
.Y(n_5537)
);

INVx2_ASAP7_75t_L g5538 ( 
.A(n_2502),
.Y(n_5538)
);

CKINVDCx5p33_ASAP7_75t_R g5539 ( 
.A(n_4236),
.Y(n_5539)
);

CKINVDCx20_ASAP7_75t_R g5540 ( 
.A(n_1442),
.Y(n_5540)
);

CKINVDCx5p33_ASAP7_75t_R g5541 ( 
.A(n_3511),
.Y(n_5541)
);

BUFx3_ASAP7_75t_L g5542 ( 
.A(n_3062),
.Y(n_5542)
);

CKINVDCx5p33_ASAP7_75t_R g5543 ( 
.A(n_1384),
.Y(n_5543)
);

INVx1_ASAP7_75t_L g5544 ( 
.A(n_1105),
.Y(n_5544)
);

CKINVDCx5p33_ASAP7_75t_R g5545 ( 
.A(n_634),
.Y(n_5545)
);

CKINVDCx11_ASAP7_75t_R g5546 ( 
.A(n_470),
.Y(n_5546)
);

INVx2_ASAP7_75t_L g5547 ( 
.A(n_1120),
.Y(n_5547)
);

BUFx2_ASAP7_75t_L g5548 ( 
.A(n_3719),
.Y(n_5548)
);

BUFx10_ASAP7_75t_L g5549 ( 
.A(n_438),
.Y(n_5549)
);

CKINVDCx5p33_ASAP7_75t_R g5550 ( 
.A(n_868),
.Y(n_5550)
);

CKINVDCx5p33_ASAP7_75t_R g5551 ( 
.A(n_1122),
.Y(n_5551)
);

INVx1_ASAP7_75t_L g5552 ( 
.A(n_735),
.Y(n_5552)
);

BUFx2_ASAP7_75t_L g5553 ( 
.A(n_1291),
.Y(n_5553)
);

CKINVDCx5p33_ASAP7_75t_R g5554 ( 
.A(n_237),
.Y(n_5554)
);

INVx1_ASAP7_75t_L g5555 ( 
.A(n_1433),
.Y(n_5555)
);

BUFx3_ASAP7_75t_L g5556 ( 
.A(n_4076),
.Y(n_5556)
);

CKINVDCx5p33_ASAP7_75t_R g5557 ( 
.A(n_1356),
.Y(n_5557)
);

CKINVDCx16_ASAP7_75t_R g5558 ( 
.A(n_808),
.Y(n_5558)
);

CKINVDCx5p33_ASAP7_75t_R g5559 ( 
.A(n_2264),
.Y(n_5559)
);

CKINVDCx5p33_ASAP7_75t_R g5560 ( 
.A(n_3877),
.Y(n_5560)
);

CKINVDCx5p33_ASAP7_75t_R g5561 ( 
.A(n_4141),
.Y(n_5561)
);

CKINVDCx5p33_ASAP7_75t_R g5562 ( 
.A(n_538),
.Y(n_5562)
);

INVx1_ASAP7_75t_L g5563 ( 
.A(n_2928),
.Y(n_5563)
);

CKINVDCx5p33_ASAP7_75t_R g5564 ( 
.A(n_3359),
.Y(n_5564)
);

INVx2_ASAP7_75t_L g5565 ( 
.A(n_571),
.Y(n_5565)
);

INVx2_ASAP7_75t_L g5566 ( 
.A(n_4146),
.Y(n_5566)
);

INVx1_ASAP7_75t_SL g5567 ( 
.A(n_2946),
.Y(n_5567)
);

INVx1_ASAP7_75t_L g5568 ( 
.A(n_3467),
.Y(n_5568)
);

CKINVDCx5p33_ASAP7_75t_R g5569 ( 
.A(n_762),
.Y(n_5569)
);

INVx1_ASAP7_75t_L g5570 ( 
.A(n_3767),
.Y(n_5570)
);

INVxp67_ASAP7_75t_L g5571 ( 
.A(n_77),
.Y(n_5571)
);

INVx1_ASAP7_75t_L g5572 ( 
.A(n_816),
.Y(n_5572)
);

CKINVDCx5p33_ASAP7_75t_R g5573 ( 
.A(n_4182),
.Y(n_5573)
);

CKINVDCx5p33_ASAP7_75t_R g5574 ( 
.A(n_2061),
.Y(n_5574)
);

CKINVDCx20_ASAP7_75t_R g5575 ( 
.A(n_1274),
.Y(n_5575)
);

CKINVDCx5p33_ASAP7_75t_R g5576 ( 
.A(n_4072),
.Y(n_5576)
);

CKINVDCx5p33_ASAP7_75t_R g5577 ( 
.A(n_1154),
.Y(n_5577)
);

BUFx6f_ASAP7_75t_L g5578 ( 
.A(n_1740),
.Y(n_5578)
);

CKINVDCx5p33_ASAP7_75t_R g5579 ( 
.A(n_527),
.Y(n_5579)
);

CKINVDCx5p33_ASAP7_75t_R g5580 ( 
.A(n_1683),
.Y(n_5580)
);

CKINVDCx5p33_ASAP7_75t_R g5581 ( 
.A(n_4157),
.Y(n_5581)
);

CKINVDCx5p33_ASAP7_75t_R g5582 ( 
.A(n_3004),
.Y(n_5582)
);

CKINVDCx5p33_ASAP7_75t_R g5583 ( 
.A(n_4074),
.Y(n_5583)
);

CKINVDCx5p33_ASAP7_75t_R g5584 ( 
.A(n_4186),
.Y(n_5584)
);

INVx2_ASAP7_75t_L g5585 ( 
.A(n_2868),
.Y(n_5585)
);

CKINVDCx5p33_ASAP7_75t_R g5586 ( 
.A(n_3085),
.Y(n_5586)
);

INVx2_ASAP7_75t_L g5587 ( 
.A(n_4173),
.Y(n_5587)
);

BUFx10_ASAP7_75t_L g5588 ( 
.A(n_1990),
.Y(n_5588)
);

INVx2_ASAP7_75t_L g5589 ( 
.A(n_4156),
.Y(n_5589)
);

CKINVDCx5p33_ASAP7_75t_R g5590 ( 
.A(n_2273),
.Y(n_5590)
);

INVx1_ASAP7_75t_L g5591 ( 
.A(n_2951),
.Y(n_5591)
);

CKINVDCx5p33_ASAP7_75t_R g5592 ( 
.A(n_4161),
.Y(n_5592)
);

CKINVDCx5p33_ASAP7_75t_R g5593 ( 
.A(n_2818),
.Y(n_5593)
);

INVx1_ASAP7_75t_L g5594 ( 
.A(n_1872),
.Y(n_5594)
);

INVx1_ASAP7_75t_L g5595 ( 
.A(n_386),
.Y(n_5595)
);

INVx1_ASAP7_75t_L g5596 ( 
.A(n_2000),
.Y(n_5596)
);

CKINVDCx5p33_ASAP7_75t_R g5597 ( 
.A(n_471),
.Y(n_5597)
);

INVx1_ASAP7_75t_L g5598 ( 
.A(n_4053),
.Y(n_5598)
);

BUFx6f_ASAP7_75t_L g5599 ( 
.A(n_2269),
.Y(n_5599)
);

INVx1_ASAP7_75t_SL g5600 ( 
.A(n_4064),
.Y(n_5600)
);

INVx1_ASAP7_75t_L g5601 ( 
.A(n_165),
.Y(n_5601)
);

CKINVDCx5p33_ASAP7_75t_R g5602 ( 
.A(n_4167),
.Y(n_5602)
);

CKINVDCx5p33_ASAP7_75t_R g5603 ( 
.A(n_743),
.Y(n_5603)
);

CKINVDCx5p33_ASAP7_75t_R g5604 ( 
.A(n_4184),
.Y(n_5604)
);

CKINVDCx5p33_ASAP7_75t_R g5605 ( 
.A(n_1301),
.Y(n_5605)
);

CKINVDCx5p33_ASAP7_75t_R g5606 ( 
.A(n_4226),
.Y(n_5606)
);

CKINVDCx20_ASAP7_75t_R g5607 ( 
.A(n_450),
.Y(n_5607)
);

CKINVDCx5p33_ASAP7_75t_R g5608 ( 
.A(n_3613),
.Y(n_5608)
);

CKINVDCx5p33_ASAP7_75t_R g5609 ( 
.A(n_3423),
.Y(n_5609)
);

CKINVDCx5p33_ASAP7_75t_R g5610 ( 
.A(n_415),
.Y(n_5610)
);

CKINVDCx5p33_ASAP7_75t_R g5611 ( 
.A(n_3672),
.Y(n_5611)
);

CKINVDCx5p33_ASAP7_75t_R g5612 ( 
.A(n_899),
.Y(n_5612)
);

INVx2_ASAP7_75t_SL g5613 ( 
.A(n_2171),
.Y(n_5613)
);

INVx1_ASAP7_75t_L g5614 ( 
.A(n_4061),
.Y(n_5614)
);

CKINVDCx5p33_ASAP7_75t_R g5615 ( 
.A(n_3529),
.Y(n_5615)
);

INVx2_ASAP7_75t_L g5616 ( 
.A(n_916),
.Y(n_5616)
);

CKINVDCx5p33_ASAP7_75t_R g5617 ( 
.A(n_496),
.Y(n_5617)
);

CKINVDCx5p33_ASAP7_75t_R g5618 ( 
.A(n_4085),
.Y(n_5618)
);

INVx1_ASAP7_75t_L g5619 ( 
.A(n_4150),
.Y(n_5619)
);

INVx1_ASAP7_75t_L g5620 ( 
.A(n_2662),
.Y(n_5620)
);

INVx2_ASAP7_75t_L g5621 ( 
.A(n_2104),
.Y(n_5621)
);

CKINVDCx5p33_ASAP7_75t_R g5622 ( 
.A(n_2835),
.Y(n_5622)
);

HB1xp67_ASAP7_75t_L g5623 ( 
.A(n_4214),
.Y(n_5623)
);

CKINVDCx5p33_ASAP7_75t_R g5624 ( 
.A(n_2283),
.Y(n_5624)
);

INVx1_ASAP7_75t_L g5625 ( 
.A(n_2520),
.Y(n_5625)
);

CKINVDCx5p33_ASAP7_75t_R g5626 ( 
.A(n_3409),
.Y(n_5626)
);

CKINVDCx5p33_ASAP7_75t_R g5627 ( 
.A(n_922),
.Y(n_5627)
);

INVx1_ASAP7_75t_L g5628 ( 
.A(n_2652),
.Y(n_5628)
);

INVx2_ASAP7_75t_L g5629 ( 
.A(n_2822),
.Y(n_5629)
);

CKINVDCx5p33_ASAP7_75t_R g5630 ( 
.A(n_3056),
.Y(n_5630)
);

CKINVDCx5p33_ASAP7_75t_R g5631 ( 
.A(n_1474),
.Y(n_5631)
);

CKINVDCx5p33_ASAP7_75t_R g5632 ( 
.A(n_1450),
.Y(n_5632)
);

INVx1_ASAP7_75t_L g5633 ( 
.A(n_3326),
.Y(n_5633)
);

CKINVDCx5p33_ASAP7_75t_R g5634 ( 
.A(n_3297),
.Y(n_5634)
);

INVx1_ASAP7_75t_L g5635 ( 
.A(n_2923),
.Y(n_5635)
);

INVx1_ASAP7_75t_SL g5636 ( 
.A(n_2153),
.Y(n_5636)
);

CKINVDCx5p33_ASAP7_75t_R g5637 ( 
.A(n_1153),
.Y(n_5637)
);

CKINVDCx5p33_ASAP7_75t_R g5638 ( 
.A(n_4053),
.Y(n_5638)
);

CKINVDCx5p33_ASAP7_75t_R g5639 ( 
.A(n_28),
.Y(n_5639)
);

INVx1_ASAP7_75t_L g5640 ( 
.A(n_245),
.Y(n_5640)
);

CKINVDCx5p33_ASAP7_75t_R g5641 ( 
.A(n_625),
.Y(n_5641)
);

CKINVDCx5p33_ASAP7_75t_R g5642 ( 
.A(n_1142),
.Y(n_5642)
);

INVx2_ASAP7_75t_L g5643 ( 
.A(n_2454),
.Y(n_5643)
);

BUFx3_ASAP7_75t_L g5644 ( 
.A(n_2685),
.Y(n_5644)
);

CKINVDCx5p33_ASAP7_75t_R g5645 ( 
.A(n_1031),
.Y(n_5645)
);

INVx1_ASAP7_75t_L g5646 ( 
.A(n_4175),
.Y(n_5646)
);

CKINVDCx5p33_ASAP7_75t_R g5647 ( 
.A(n_3891),
.Y(n_5647)
);

CKINVDCx5p33_ASAP7_75t_R g5648 ( 
.A(n_2514),
.Y(n_5648)
);

CKINVDCx16_ASAP7_75t_R g5649 ( 
.A(n_2159),
.Y(n_5649)
);

CKINVDCx5p33_ASAP7_75t_R g5650 ( 
.A(n_3711),
.Y(n_5650)
);

CKINVDCx5p33_ASAP7_75t_R g5651 ( 
.A(n_1855),
.Y(n_5651)
);

INVx2_ASAP7_75t_L g5652 ( 
.A(n_1324),
.Y(n_5652)
);

BUFx10_ASAP7_75t_L g5653 ( 
.A(n_343),
.Y(n_5653)
);

INVx1_ASAP7_75t_L g5654 ( 
.A(n_3319),
.Y(n_5654)
);

CKINVDCx5p33_ASAP7_75t_R g5655 ( 
.A(n_3720),
.Y(n_5655)
);

INVx1_ASAP7_75t_L g5656 ( 
.A(n_971),
.Y(n_5656)
);

CKINVDCx14_ASAP7_75t_R g5657 ( 
.A(n_4073),
.Y(n_5657)
);

CKINVDCx5p33_ASAP7_75t_R g5658 ( 
.A(n_3958),
.Y(n_5658)
);

CKINVDCx5p33_ASAP7_75t_R g5659 ( 
.A(n_3592),
.Y(n_5659)
);

INVx1_ASAP7_75t_L g5660 ( 
.A(n_1826),
.Y(n_5660)
);

INVx1_ASAP7_75t_SL g5661 ( 
.A(n_3256),
.Y(n_5661)
);

CKINVDCx5p33_ASAP7_75t_R g5662 ( 
.A(n_298),
.Y(n_5662)
);

CKINVDCx5p33_ASAP7_75t_R g5663 ( 
.A(n_1772),
.Y(n_5663)
);

CKINVDCx5p33_ASAP7_75t_R g5664 ( 
.A(n_3707),
.Y(n_5664)
);

CKINVDCx5p33_ASAP7_75t_R g5665 ( 
.A(n_2782),
.Y(n_5665)
);

CKINVDCx16_ASAP7_75t_R g5666 ( 
.A(n_2820),
.Y(n_5666)
);

CKINVDCx20_ASAP7_75t_R g5667 ( 
.A(n_4089),
.Y(n_5667)
);

INVx1_ASAP7_75t_L g5668 ( 
.A(n_285),
.Y(n_5668)
);

CKINVDCx5p33_ASAP7_75t_R g5669 ( 
.A(n_1158),
.Y(n_5669)
);

INVx1_ASAP7_75t_L g5670 ( 
.A(n_372),
.Y(n_5670)
);

BUFx6f_ASAP7_75t_L g5671 ( 
.A(n_2644),
.Y(n_5671)
);

INVx1_ASAP7_75t_L g5672 ( 
.A(n_2569),
.Y(n_5672)
);

CKINVDCx16_ASAP7_75t_R g5673 ( 
.A(n_3570),
.Y(n_5673)
);

INVx1_ASAP7_75t_L g5674 ( 
.A(n_1992),
.Y(n_5674)
);

INVx1_ASAP7_75t_L g5675 ( 
.A(n_3009),
.Y(n_5675)
);

CKINVDCx5p33_ASAP7_75t_R g5676 ( 
.A(n_4148),
.Y(n_5676)
);

INVx1_ASAP7_75t_L g5677 ( 
.A(n_1326),
.Y(n_5677)
);

CKINVDCx5p33_ASAP7_75t_R g5678 ( 
.A(n_1273),
.Y(n_5678)
);

INVx1_ASAP7_75t_L g5679 ( 
.A(n_1987),
.Y(n_5679)
);

CKINVDCx5p33_ASAP7_75t_R g5680 ( 
.A(n_1910),
.Y(n_5680)
);

INVx1_ASAP7_75t_L g5681 ( 
.A(n_4019),
.Y(n_5681)
);

CKINVDCx5p33_ASAP7_75t_R g5682 ( 
.A(n_2665),
.Y(n_5682)
);

CKINVDCx5p33_ASAP7_75t_R g5683 ( 
.A(n_1806),
.Y(n_5683)
);

INVx2_ASAP7_75t_SL g5684 ( 
.A(n_2728),
.Y(n_5684)
);

BUFx6f_ASAP7_75t_L g5685 ( 
.A(n_2399),
.Y(n_5685)
);

BUFx6f_ASAP7_75t_L g5686 ( 
.A(n_2748),
.Y(n_5686)
);

CKINVDCx5p33_ASAP7_75t_R g5687 ( 
.A(n_129),
.Y(n_5687)
);

INVx2_ASAP7_75t_L g5688 ( 
.A(n_1688),
.Y(n_5688)
);

INVx1_ASAP7_75t_L g5689 ( 
.A(n_2441),
.Y(n_5689)
);

INVx1_ASAP7_75t_SL g5690 ( 
.A(n_821),
.Y(n_5690)
);

CKINVDCx5p33_ASAP7_75t_R g5691 ( 
.A(n_4062),
.Y(n_5691)
);

CKINVDCx5p33_ASAP7_75t_R g5692 ( 
.A(n_1725),
.Y(n_5692)
);

INVx1_ASAP7_75t_L g5693 ( 
.A(n_844),
.Y(n_5693)
);

INVx1_ASAP7_75t_L g5694 ( 
.A(n_2422),
.Y(n_5694)
);

INVx1_ASAP7_75t_L g5695 ( 
.A(n_3686),
.Y(n_5695)
);

INVx1_ASAP7_75t_L g5696 ( 
.A(n_3022),
.Y(n_5696)
);

CKINVDCx5p33_ASAP7_75t_R g5697 ( 
.A(n_4138),
.Y(n_5697)
);

CKINVDCx5p33_ASAP7_75t_R g5698 ( 
.A(n_1849),
.Y(n_5698)
);

CKINVDCx5p33_ASAP7_75t_R g5699 ( 
.A(n_2268),
.Y(n_5699)
);

CKINVDCx20_ASAP7_75t_R g5700 ( 
.A(n_1505),
.Y(n_5700)
);

CKINVDCx5p33_ASAP7_75t_R g5701 ( 
.A(n_3524),
.Y(n_5701)
);

CKINVDCx5p33_ASAP7_75t_R g5702 ( 
.A(n_2702),
.Y(n_5702)
);

CKINVDCx5p33_ASAP7_75t_R g5703 ( 
.A(n_2494),
.Y(n_5703)
);

HB1xp67_ASAP7_75t_L g5704 ( 
.A(n_1856),
.Y(n_5704)
);

CKINVDCx5p33_ASAP7_75t_R g5705 ( 
.A(n_1503),
.Y(n_5705)
);

INVx1_ASAP7_75t_L g5706 ( 
.A(n_193),
.Y(n_5706)
);

CKINVDCx5p33_ASAP7_75t_R g5707 ( 
.A(n_4087),
.Y(n_5707)
);

CKINVDCx5p33_ASAP7_75t_R g5708 ( 
.A(n_4052),
.Y(n_5708)
);

BUFx8_ASAP7_75t_SL g5709 ( 
.A(n_2085),
.Y(n_5709)
);

INVx1_ASAP7_75t_L g5710 ( 
.A(n_1676),
.Y(n_5710)
);

CKINVDCx5p33_ASAP7_75t_R g5711 ( 
.A(n_2989),
.Y(n_5711)
);

CKINVDCx5p33_ASAP7_75t_R g5712 ( 
.A(n_2727),
.Y(n_5712)
);

INVx2_ASAP7_75t_L g5713 ( 
.A(n_3844),
.Y(n_5713)
);

CKINVDCx5p33_ASAP7_75t_R g5714 ( 
.A(n_4130),
.Y(n_5714)
);

CKINVDCx5p33_ASAP7_75t_R g5715 ( 
.A(n_2917),
.Y(n_5715)
);

INVx1_ASAP7_75t_L g5716 ( 
.A(n_3812),
.Y(n_5716)
);

CKINVDCx5p33_ASAP7_75t_R g5717 ( 
.A(n_3579),
.Y(n_5717)
);

CKINVDCx20_ASAP7_75t_R g5718 ( 
.A(n_66),
.Y(n_5718)
);

CKINVDCx5p33_ASAP7_75t_R g5719 ( 
.A(n_726),
.Y(n_5719)
);

INVx1_ASAP7_75t_L g5720 ( 
.A(n_878),
.Y(n_5720)
);

BUFx6f_ASAP7_75t_L g5721 ( 
.A(n_3224),
.Y(n_5721)
);

INVx2_ASAP7_75t_SL g5722 ( 
.A(n_3000),
.Y(n_5722)
);

INVx2_ASAP7_75t_SL g5723 ( 
.A(n_365),
.Y(n_5723)
);

BUFx10_ASAP7_75t_L g5724 ( 
.A(n_323),
.Y(n_5724)
);

CKINVDCx5p33_ASAP7_75t_R g5725 ( 
.A(n_654),
.Y(n_5725)
);

CKINVDCx5p33_ASAP7_75t_R g5726 ( 
.A(n_3739),
.Y(n_5726)
);

BUFx6f_ASAP7_75t_L g5727 ( 
.A(n_1745),
.Y(n_5727)
);

CKINVDCx5p33_ASAP7_75t_R g5728 ( 
.A(n_1979),
.Y(n_5728)
);

CKINVDCx5p33_ASAP7_75t_R g5729 ( 
.A(n_747),
.Y(n_5729)
);

INVx1_ASAP7_75t_L g5730 ( 
.A(n_163),
.Y(n_5730)
);

CKINVDCx5p33_ASAP7_75t_R g5731 ( 
.A(n_3464),
.Y(n_5731)
);

CKINVDCx5p33_ASAP7_75t_R g5732 ( 
.A(n_4166),
.Y(n_5732)
);

CKINVDCx5p33_ASAP7_75t_R g5733 ( 
.A(n_3738),
.Y(n_5733)
);

CKINVDCx5p33_ASAP7_75t_R g5734 ( 
.A(n_3102),
.Y(n_5734)
);

INVx2_ASAP7_75t_L g5735 ( 
.A(n_172),
.Y(n_5735)
);

CKINVDCx5p33_ASAP7_75t_R g5736 ( 
.A(n_2433),
.Y(n_5736)
);

CKINVDCx5p33_ASAP7_75t_R g5737 ( 
.A(n_3351),
.Y(n_5737)
);

CKINVDCx5p33_ASAP7_75t_R g5738 ( 
.A(n_1594),
.Y(n_5738)
);

CKINVDCx5p33_ASAP7_75t_R g5739 ( 
.A(n_3451),
.Y(n_5739)
);

BUFx3_ASAP7_75t_L g5740 ( 
.A(n_3737),
.Y(n_5740)
);

INVx1_ASAP7_75t_L g5741 ( 
.A(n_2323),
.Y(n_5741)
);

CKINVDCx5p33_ASAP7_75t_R g5742 ( 
.A(n_2588),
.Y(n_5742)
);

INVx1_ASAP7_75t_L g5743 ( 
.A(n_3623),
.Y(n_5743)
);

INVx1_ASAP7_75t_L g5744 ( 
.A(n_1101),
.Y(n_5744)
);

BUFx3_ASAP7_75t_L g5745 ( 
.A(n_979),
.Y(n_5745)
);

CKINVDCx5p33_ASAP7_75t_R g5746 ( 
.A(n_3194),
.Y(n_5746)
);

INVx1_ASAP7_75t_L g5747 ( 
.A(n_1505),
.Y(n_5747)
);

INVx1_ASAP7_75t_L g5748 ( 
.A(n_4100),
.Y(n_5748)
);

CKINVDCx5p33_ASAP7_75t_R g5749 ( 
.A(n_938),
.Y(n_5749)
);

INVx2_ASAP7_75t_L g5750 ( 
.A(n_4065),
.Y(n_5750)
);

CKINVDCx20_ASAP7_75t_R g5751 ( 
.A(n_1183),
.Y(n_5751)
);

CKINVDCx5p33_ASAP7_75t_R g5752 ( 
.A(n_576),
.Y(n_5752)
);

CKINVDCx5p33_ASAP7_75t_R g5753 ( 
.A(n_5546),
.Y(n_5753)
);

INVx1_ASAP7_75t_L g5754 ( 
.A(n_4567),
.Y(n_5754)
);

INVxp67_ASAP7_75t_L g5755 ( 
.A(n_4488),
.Y(n_5755)
);

CKINVDCx20_ASAP7_75t_R g5756 ( 
.A(n_5012),
.Y(n_5756)
);

INVx1_ASAP7_75t_SL g5757 ( 
.A(n_4515),
.Y(n_5757)
);

INVx1_ASAP7_75t_L g5758 ( 
.A(n_4567),
.Y(n_5758)
);

INVx1_ASAP7_75t_L g5759 ( 
.A(n_4567),
.Y(n_5759)
);

INVx1_ASAP7_75t_L g5760 ( 
.A(n_4567),
.Y(n_5760)
);

INVx1_ASAP7_75t_L g5761 ( 
.A(n_4567),
.Y(n_5761)
);

INVx1_ASAP7_75t_L g5762 ( 
.A(n_5046),
.Y(n_5762)
);

CKINVDCx5p33_ASAP7_75t_R g5763 ( 
.A(n_4484),
.Y(n_5763)
);

INVx1_ASAP7_75t_SL g5764 ( 
.A(n_4547),
.Y(n_5764)
);

CKINVDCx5p33_ASAP7_75t_R g5765 ( 
.A(n_4727),
.Y(n_5765)
);

INVx1_ASAP7_75t_L g5766 ( 
.A(n_5046),
.Y(n_5766)
);

NOR2xp67_ASAP7_75t_L g5767 ( 
.A(n_4502),
.B(n_0),
.Y(n_5767)
);

INVx1_ASAP7_75t_L g5768 ( 
.A(n_5046),
.Y(n_5768)
);

INVx1_ASAP7_75t_L g5769 ( 
.A(n_5046),
.Y(n_5769)
);

BUFx2_ASAP7_75t_SL g5770 ( 
.A(n_4326),
.Y(n_5770)
);

CKINVDCx5p33_ASAP7_75t_R g5771 ( 
.A(n_5244),
.Y(n_5771)
);

INVx1_ASAP7_75t_L g5772 ( 
.A(n_5046),
.Y(n_5772)
);

BUFx2_ASAP7_75t_L g5773 ( 
.A(n_5709),
.Y(n_5773)
);

BUFx6f_ASAP7_75t_L g5774 ( 
.A(n_4403),
.Y(n_5774)
);

CKINVDCx5p33_ASAP7_75t_R g5775 ( 
.A(n_4443),
.Y(n_5775)
);

INVx2_ASAP7_75t_L g5776 ( 
.A(n_5117),
.Y(n_5776)
);

INVx2_ASAP7_75t_L g5777 ( 
.A(n_5117),
.Y(n_5777)
);

INVx1_ASAP7_75t_L g5778 ( 
.A(n_5117),
.Y(n_5778)
);

INVx2_ASAP7_75t_L g5779 ( 
.A(n_5117),
.Y(n_5779)
);

INVx2_ASAP7_75t_L g5780 ( 
.A(n_5117),
.Y(n_5780)
);

CKINVDCx5p33_ASAP7_75t_R g5781 ( 
.A(n_4482),
.Y(n_5781)
);

CKINVDCx5p33_ASAP7_75t_R g5782 ( 
.A(n_4862),
.Y(n_5782)
);

INVx1_ASAP7_75t_L g5783 ( 
.A(n_5293),
.Y(n_5783)
);

CKINVDCx5p33_ASAP7_75t_R g5784 ( 
.A(n_4871),
.Y(n_5784)
);

CKINVDCx5p33_ASAP7_75t_R g5785 ( 
.A(n_5034),
.Y(n_5785)
);

BUFx3_ASAP7_75t_L g5786 ( 
.A(n_4357),
.Y(n_5786)
);

CKINVDCx5p33_ASAP7_75t_R g5787 ( 
.A(n_5225),
.Y(n_5787)
);

CKINVDCx20_ASAP7_75t_R g5788 ( 
.A(n_4729),
.Y(n_5788)
);

CKINVDCx14_ASAP7_75t_R g5789 ( 
.A(n_4752),
.Y(n_5789)
);

CKINVDCx5p33_ASAP7_75t_R g5790 ( 
.A(n_4890),
.Y(n_5790)
);

CKINVDCx5p33_ASAP7_75t_R g5791 ( 
.A(n_4894),
.Y(n_5791)
);

CKINVDCx5p33_ASAP7_75t_R g5792 ( 
.A(n_4901),
.Y(n_5792)
);

CKINVDCx20_ASAP7_75t_R g5793 ( 
.A(n_5144),
.Y(n_5793)
);

INVx2_ASAP7_75t_L g5794 ( 
.A(n_5293),
.Y(n_5794)
);

HB1xp67_ASAP7_75t_L g5795 ( 
.A(n_4390),
.Y(n_5795)
);

CKINVDCx5p33_ASAP7_75t_R g5796 ( 
.A(n_5657),
.Y(n_5796)
);

HB1xp67_ASAP7_75t_L g5797 ( 
.A(n_4397),
.Y(n_5797)
);

CKINVDCx5p33_ASAP7_75t_R g5798 ( 
.A(n_4418),
.Y(n_5798)
);

INVx1_ASAP7_75t_L g5799 ( 
.A(n_5293),
.Y(n_5799)
);

CKINVDCx5p33_ASAP7_75t_R g5800 ( 
.A(n_4501),
.Y(n_5800)
);

CKINVDCx5p33_ASAP7_75t_R g5801 ( 
.A(n_4692),
.Y(n_5801)
);

INVx1_ASAP7_75t_L g5802 ( 
.A(n_5293),
.Y(n_5802)
);

INVx2_ASAP7_75t_L g5803 ( 
.A(n_5293),
.Y(n_5803)
);

CKINVDCx5p33_ASAP7_75t_R g5804 ( 
.A(n_4710),
.Y(n_5804)
);

CKINVDCx5p33_ASAP7_75t_R g5805 ( 
.A(n_4816),
.Y(n_5805)
);

CKINVDCx5p33_ASAP7_75t_R g5806 ( 
.A(n_4889),
.Y(n_5806)
);

INVx1_ASAP7_75t_L g5807 ( 
.A(n_5412),
.Y(n_5807)
);

CKINVDCx5p33_ASAP7_75t_R g5808 ( 
.A(n_5031),
.Y(n_5808)
);

CKINVDCx14_ASAP7_75t_R g5809 ( 
.A(n_4685),
.Y(n_5809)
);

CKINVDCx5p33_ASAP7_75t_R g5810 ( 
.A(n_5049),
.Y(n_5810)
);

INVx1_ASAP7_75t_L g5811 ( 
.A(n_5412),
.Y(n_5811)
);

INVx1_ASAP7_75t_L g5812 ( 
.A(n_5412),
.Y(n_5812)
);

CKINVDCx5p33_ASAP7_75t_R g5813 ( 
.A(n_5088),
.Y(n_5813)
);

BUFx10_ASAP7_75t_L g5814 ( 
.A(n_5407),
.Y(n_5814)
);

CKINVDCx5p33_ASAP7_75t_R g5815 ( 
.A(n_5125),
.Y(n_5815)
);

INVx1_ASAP7_75t_L g5816 ( 
.A(n_5412),
.Y(n_5816)
);

INVx2_ASAP7_75t_L g5817 ( 
.A(n_5412),
.Y(n_5817)
);

CKINVDCx5p33_ASAP7_75t_R g5818 ( 
.A(n_5205),
.Y(n_5818)
);

INVxp67_ASAP7_75t_L g5819 ( 
.A(n_4938),
.Y(n_5819)
);

INVx1_ASAP7_75t_L g5820 ( 
.A(n_4502),
.Y(n_5820)
);

INVx1_ASAP7_75t_L g5821 ( 
.A(n_5020),
.Y(n_5821)
);

CKINVDCx5p33_ASAP7_75t_R g5822 ( 
.A(n_5273),
.Y(n_5822)
);

INVx1_ASAP7_75t_L g5823 ( 
.A(n_5020),
.Y(n_5823)
);

INVx1_ASAP7_75t_L g5824 ( 
.A(n_5450),
.Y(n_5824)
);

INVxp67_ASAP7_75t_SL g5825 ( 
.A(n_5450),
.Y(n_5825)
);

INVx1_ASAP7_75t_L g5826 ( 
.A(n_4403),
.Y(n_5826)
);

CKINVDCx5p33_ASAP7_75t_R g5827 ( 
.A(n_5291),
.Y(n_5827)
);

CKINVDCx20_ASAP7_75t_R g5828 ( 
.A(n_5306),
.Y(n_5828)
);

INVx1_ASAP7_75t_L g5829 ( 
.A(n_4403),
.Y(n_5829)
);

CKINVDCx16_ASAP7_75t_R g5830 ( 
.A(n_5389),
.Y(n_5830)
);

INVx1_ASAP7_75t_L g5831 ( 
.A(n_4551),
.Y(n_5831)
);

INVx1_ASAP7_75t_L g5832 ( 
.A(n_4551),
.Y(n_5832)
);

CKINVDCx20_ASAP7_75t_R g5833 ( 
.A(n_5558),
.Y(n_5833)
);

INVx1_ASAP7_75t_L g5834 ( 
.A(n_4551),
.Y(n_5834)
);

INVx1_ASAP7_75t_L g5835 ( 
.A(n_4677),
.Y(n_5835)
);

CKINVDCx5p33_ASAP7_75t_R g5836 ( 
.A(n_5649),
.Y(n_5836)
);

INVx1_ASAP7_75t_L g5837 ( 
.A(n_4677),
.Y(n_5837)
);

CKINVDCx5p33_ASAP7_75t_R g5838 ( 
.A(n_5666),
.Y(n_5838)
);

INVx1_ASAP7_75t_L g5839 ( 
.A(n_4677),
.Y(n_5839)
);

CKINVDCx5p33_ASAP7_75t_R g5840 ( 
.A(n_5673),
.Y(n_5840)
);

CKINVDCx5p33_ASAP7_75t_R g5841 ( 
.A(n_5472),
.Y(n_5841)
);

INVx1_ASAP7_75t_L g5842 ( 
.A(n_4779),
.Y(n_5842)
);

CKINVDCx5p33_ASAP7_75t_R g5843 ( 
.A(n_5742),
.Y(n_5843)
);

CKINVDCx5p33_ASAP7_75t_R g5844 ( 
.A(n_5746),
.Y(n_5844)
);

INVx1_ASAP7_75t_L g5845 ( 
.A(n_4779),
.Y(n_5845)
);

CKINVDCx16_ASAP7_75t_R g5846 ( 
.A(n_4323),
.Y(n_5846)
);

INVx1_ASAP7_75t_L g5847 ( 
.A(n_4779),
.Y(n_5847)
);

CKINVDCx20_ASAP7_75t_R g5848 ( 
.A(n_4327),
.Y(n_5848)
);

INVx1_ASAP7_75t_SL g5849 ( 
.A(n_5109),
.Y(n_5849)
);

INVx1_ASAP7_75t_L g5850 ( 
.A(n_4853),
.Y(n_5850)
);

INVx1_ASAP7_75t_L g5851 ( 
.A(n_4853),
.Y(n_5851)
);

BUFx6f_ASAP7_75t_L g5852 ( 
.A(n_4853),
.Y(n_5852)
);

INVx1_ASAP7_75t_L g5853 ( 
.A(n_4865),
.Y(n_5853)
);

CKINVDCx5p33_ASAP7_75t_R g5854 ( 
.A(n_5749),
.Y(n_5854)
);

NOR2xp67_ASAP7_75t_L g5855 ( 
.A(n_4437),
.B(n_0),
.Y(n_5855)
);

BUFx3_ASAP7_75t_L g5856 ( 
.A(n_4486),
.Y(n_5856)
);

INVx1_ASAP7_75t_L g5857 ( 
.A(n_4865),
.Y(n_5857)
);

CKINVDCx5p33_ASAP7_75t_R g5858 ( 
.A(n_5752),
.Y(n_5858)
);

INVx1_ASAP7_75t_L g5859 ( 
.A(n_4865),
.Y(n_5859)
);

INVx1_ASAP7_75t_L g5860 ( 
.A(n_4974),
.Y(n_5860)
);

CKINVDCx5p33_ASAP7_75t_R g5861 ( 
.A(n_4322),
.Y(n_5861)
);

CKINVDCx5p33_ASAP7_75t_R g5862 ( 
.A(n_5734),
.Y(n_5862)
);

CKINVDCx20_ASAP7_75t_R g5863 ( 
.A(n_4353),
.Y(n_5863)
);

INVx1_ASAP7_75t_L g5864 ( 
.A(n_4974),
.Y(n_5864)
);

CKINVDCx5p33_ASAP7_75t_R g5865 ( 
.A(n_5736),
.Y(n_5865)
);

INVx1_ASAP7_75t_L g5866 ( 
.A(n_4974),
.Y(n_5866)
);

CKINVDCx16_ASAP7_75t_R g5867 ( 
.A(n_4323),
.Y(n_5867)
);

INVx1_ASAP7_75t_L g5868 ( 
.A(n_5067),
.Y(n_5868)
);

CKINVDCx5p33_ASAP7_75t_R g5869 ( 
.A(n_5739),
.Y(n_5869)
);

INVx1_ASAP7_75t_L g5870 ( 
.A(n_5067),
.Y(n_5870)
);

CKINVDCx5p33_ASAP7_75t_R g5871 ( 
.A(n_4324),
.Y(n_5871)
);

INVx1_ASAP7_75t_L g5872 ( 
.A(n_5067),
.Y(n_5872)
);

CKINVDCx20_ASAP7_75t_R g5873 ( 
.A(n_4376),
.Y(n_5873)
);

INVx1_ASAP7_75t_SL g5874 ( 
.A(n_5163),
.Y(n_5874)
);

INVx1_ASAP7_75t_L g5875 ( 
.A(n_5071),
.Y(n_5875)
);

INVx1_ASAP7_75t_L g5876 ( 
.A(n_5071),
.Y(n_5876)
);

INVx1_ASAP7_75t_L g5877 ( 
.A(n_5071),
.Y(n_5877)
);

CKINVDCx5p33_ASAP7_75t_R g5878 ( 
.A(n_4325),
.Y(n_5878)
);

CKINVDCx5p33_ASAP7_75t_R g5879 ( 
.A(n_4328),
.Y(n_5879)
);

CKINVDCx5p33_ASAP7_75t_R g5880 ( 
.A(n_4332),
.Y(n_5880)
);

INVx1_ASAP7_75t_L g5881 ( 
.A(n_5102),
.Y(n_5881)
);

BUFx5_ASAP7_75t_L g5882 ( 
.A(n_4603),
.Y(n_5882)
);

CKINVDCx5p33_ASAP7_75t_R g5883 ( 
.A(n_4333),
.Y(n_5883)
);

INVx2_ASAP7_75t_L g5884 ( 
.A(n_5102),
.Y(n_5884)
);

CKINVDCx16_ASAP7_75t_R g5885 ( 
.A(n_4331),
.Y(n_5885)
);

INVx1_ASAP7_75t_L g5886 ( 
.A(n_5102),
.Y(n_5886)
);

CKINVDCx5p33_ASAP7_75t_R g5887 ( 
.A(n_5732),
.Y(n_5887)
);

INVx2_ASAP7_75t_L g5888 ( 
.A(n_5118),
.Y(n_5888)
);

CKINVDCx5p33_ASAP7_75t_R g5889 ( 
.A(n_5733),
.Y(n_5889)
);

CKINVDCx5p33_ASAP7_75t_R g5890 ( 
.A(n_5737),
.Y(n_5890)
);

INVx1_ASAP7_75t_L g5891 ( 
.A(n_5118),
.Y(n_5891)
);

CKINVDCx5p33_ASAP7_75t_R g5892 ( 
.A(n_5738),
.Y(n_5892)
);

INVx1_ASAP7_75t_L g5893 ( 
.A(n_5118),
.Y(n_5893)
);

BUFx10_ASAP7_75t_L g5894 ( 
.A(n_4329),
.Y(n_5894)
);

INVx2_ASAP7_75t_L g5895 ( 
.A(n_5141),
.Y(n_5895)
);

INVx1_ASAP7_75t_L g5896 ( 
.A(n_5141),
.Y(n_5896)
);

NOR2xp67_ASAP7_75t_L g5897 ( 
.A(n_4556),
.B(n_2),
.Y(n_5897)
);

CKINVDCx5p33_ASAP7_75t_R g5898 ( 
.A(n_4334),
.Y(n_5898)
);

INVx1_ASAP7_75t_L g5899 ( 
.A(n_5141),
.Y(n_5899)
);

CKINVDCx20_ASAP7_75t_R g5900 ( 
.A(n_4378),
.Y(n_5900)
);

BUFx3_ASAP7_75t_L g5901 ( 
.A(n_4529),
.Y(n_5901)
);

BUFx3_ASAP7_75t_L g5902 ( 
.A(n_4559),
.Y(n_5902)
);

INVx1_ASAP7_75t_L g5903 ( 
.A(n_5235),
.Y(n_5903)
);

INVx2_ASAP7_75t_L g5904 ( 
.A(n_5235),
.Y(n_5904)
);

INVx1_ASAP7_75t_L g5905 ( 
.A(n_5235),
.Y(n_5905)
);

CKINVDCx5p33_ASAP7_75t_R g5906 ( 
.A(n_4337),
.Y(n_5906)
);

INVx1_ASAP7_75t_L g5907 ( 
.A(n_5255),
.Y(n_5907)
);

CKINVDCx5p33_ASAP7_75t_R g5908 ( 
.A(n_4338),
.Y(n_5908)
);

INVx1_ASAP7_75t_L g5909 ( 
.A(n_5255),
.Y(n_5909)
);

INVx1_ASAP7_75t_L g5910 ( 
.A(n_5255),
.Y(n_5910)
);

CKINVDCx5p33_ASAP7_75t_R g5911 ( 
.A(n_5728),
.Y(n_5911)
);

BUFx6f_ASAP7_75t_L g5912 ( 
.A(n_5323),
.Y(n_5912)
);

CKINVDCx5p33_ASAP7_75t_R g5913 ( 
.A(n_5729),
.Y(n_5913)
);

INVx1_ASAP7_75t_L g5914 ( 
.A(n_5323),
.Y(n_5914)
);

CKINVDCx5p33_ASAP7_75t_R g5915 ( 
.A(n_5731),
.Y(n_5915)
);

INVx1_ASAP7_75t_L g5916 ( 
.A(n_5323),
.Y(n_5916)
);

BUFx10_ASAP7_75t_L g5917 ( 
.A(n_4511),
.Y(n_5917)
);

CKINVDCx5p33_ASAP7_75t_R g5918 ( 
.A(n_4339),
.Y(n_5918)
);

INVx1_ASAP7_75t_L g5919 ( 
.A(n_5324),
.Y(n_5919)
);

INVx1_ASAP7_75t_L g5920 ( 
.A(n_5324),
.Y(n_5920)
);

CKINVDCx5p33_ASAP7_75t_R g5921 ( 
.A(n_4340),
.Y(n_5921)
);

CKINVDCx5p33_ASAP7_75t_R g5922 ( 
.A(n_4342),
.Y(n_5922)
);

CKINVDCx5p33_ASAP7_75t_R g5923 ( 
.A(n_4343),
.Y(n_5923)
);

CKINVDCx20_ASAP7_75t_R g5924 ( 
.A(n_4384),
.Y(n_5924)
);

INVx1_ASAP7_75t_L g5925 ( 
.A(n_5324),
.Y(n_5925)
);

CKINVDCx5p33_ASAP7_75t_R g5926 ( 
.A(n_4344),
.Y(n_5926)
);

CKINVDCx5p33_ASAP7_75t_R g5927 ( 
.A(n_4346),
.Y(n_5927)
);

INVxp67_ASAP7_75t_L g5928 ( 
.A(n_5169),
.Y(n_5928)
);

CKINVDCx5p33_ASAP7_75t_R g5929 ( 
.A(n_4348),
.Y(n_5929)
);

BUFx2_ASAP7_75t_L g5930 ( 
.A(n_5214),
.Y(n_5930)
);

BUFx3_ASAP7_75t_L g5931 ( 
.A(n_4579),
.Y(n_5931)
);

CKINVDCx5p33_ASAP7_75t_R g5932 ( 
.A(n_5726),
.Y(n_5932)
);

INVx1_ASAP7_75t_L g5933 ( 
.A(n_5414),
.Y(n_5933)
);

CKINVDCx5p33_ASAP7_75t_R g5934 ( 
.A(n_4349),
.Y(n_5934)
);

CKINVDCx5p33_ASAP7_75t_R g5935 ( 
.A(n_4351),
.Y(n_5935)
);

INVx1_ASAP7_75t_L g5936 ( 
.A(n_5414),
.Y(n_5936)
);

NOR2xp33_ASAP7_75t_L g5937 ( 
.A(n_5058),
.B(n_2),
.Y(n_5937)
);

CKINVDCx5p33_ASAP7_75t_R g5938 ( 
.A(n_4354),
.Y(n_5938)
);

BUFx2_ASAP7_75t_SL g5939 ( 
.A(n_4420),
.Y(n_5939)
);

INVx1_ASAP7_75t_L g5940 ( 
.A(n_5414),
.Y(n_5940)
);

INVx1_ASAP7_75t_L g5941 ( 
.A(n_5446),
.Y(n_5941)
);

INVx1_ASAP7_75t_L g5942 ( 
.A(n_5446),
.Y(n_5942)
);

BUFx3_ASAP7_75t_L g5943 ( 
.A(n_4583),
.Y(n_5943)
);

INVx1_ASAP7_75t_L g5944 ( 
.A(n_5446),
.Y(n_5944)
);

INVx1_ASAP7_75t_L g5945 ( 
.A(n_5470),
.Y(n_5945)
);

BUFx6f_ASAP7_75t_L g5946 ( 
.A(n_5470),
.Y(n_5946)
);

INVx1_ASAP7_75t_L g5947 ( 
.A(n_5470),
.Y(n_5947)
);

HB1xp67_ASAP7_75t_L g5948 ( 
.A(n_4335),
.Y(n_5948)
);

CKINVDCx5p33_ASAP7_75t_R g5949 ( 
.A(n_4355),
.Y(n_5949)
);

CKINVDCx5p33_ASAP7_75t_R g5950 ( 
.A(n_4356),
.Y(n_5950)
);

CKINVDCx20_ASAP7_75t_R g5951 ( 
.A(n_4414),
.Y(n_5951)
);

INVx1_ASAP7_75t_L g5952 ( 
.A(n_5514),
.Y(n_5952)
);

CKINVDCx5p33_ASAP7_75t_R g5953 ( 
.A(n_5725),
.Y(n_5953)
);

CKINVDCx5p33_ASAP7_75t_R g5954 ( 
.A(n_4359),
.Y(n_5954)
);

HB1xp67_ASAP7_75t_L g5955 ( 
.A(n_4377),
.Y(n_5955)
);

CKINVDCx16_ASAP7_75t_R g5956 ( 
.A(n_4331),
.Y(n_5956)
);

CKINVDCx5p33_ASAP7_75t_R g5957 ( 
.A(n_4360),
.Y(n_5957)
);

INVx1_ASAP7_75t_L g5958 ( 
.A(n_5514),
.Y(n_5958)
);

INVx1_ASAP7_75t_L g5959 ( 
.A(n_5514),
.Y(n_5959)
);

CKINVDCx5p33_ASAP7_75t_R g5960 ( 
.A(n_4361),
.Y(n_5960)
);

CKINVDCx14_ASAP7_75t_R g5961 ( 
.A(n_5305),
.Y(n_5961)
);

INVx1_ASAP7_75t_L g5962 ( 
.A(n_5521),
.Y(n_5962)
);

INVx2_ASAP7_75t_L g5963 ( 
.A(n_5521),
.Y(n_5963)
);

CKINVDCx5p33_ASAP7_75t_R g5964 ( 
.A(n_4364),
.Y(n_5964)
);

NOR2xp67_ASAP7_75t_L g5965 ( 
.A(n_4672),
.B(n_3),
.Y(n_5965)
);

INVx1_ASAP7_75t_L g5966 ( 
.A(n_5521),
.Y(n_5966)
);

INVx2_ASAP7_75t_L g5967 ( 
.A(n_5527),
.Y(n_5967)
);

CKINVDCx5p33_ASAP7_75t_R g5968 ( 
.A(n_4365),
.Y(n_5968)
);

INVx1_ASAP7_75t_L g5969 ( 
.A(n_5527),
.Y(n_5969)
);

CKINVDCx20_ASAP7_75t_R g5970 ( 
.A(n_4415),
.Y(n_5970)
);

INVx1_ASAP7_75t_L g5971 ( 
.A(n_5527),
.Y(n_5971)
);

CKINVDCx5p33_ASAP7_75t_R g5972 ( 
.A(n_4366),
.Y(n_5972)
);

INVx1_ASAP7_75t_L g5973 ( 
.A(n_5578),
.Y(n_5973)
);

INVx1_ASAP7_75t_L g5974 ( 
.A(n_5578),
.Y(n_5974)
);

INVx2_ASAP7_75t_L g5975 ( 
.A(n_5578),
.Y(n_5975)
);

INVxp67_ASAP7_75t_L g5976 ( 
.A(n_5337),
.Y(n_5976)
);

INVx1_ASAP7_75t_L g5977 ( 
.A(n_5599),
.Y(n_5977)
);

INVx1_ASAP7_75t_L g5978 ( 
.A(n_5599),
.Y(n_5978)
);

INVx1_ASAP7_75t_L g5979 ( 
.A(n_5599),
.Y(n_5979)
);

CKINVDCx5p33_ASAP7_75t_R g5980 ( 
.A(n_4367),
.Y(n_5980)
);

CKINVDCx5p33_ASAP7_75t_R g5981 ( 
.A(n_4370),
.Y(n_5981)
);

CKINVDCx14_ASAP7_75t_R g5982 ( 
.A(n_5367),
.Y(n_5982)
);

CKINVDCx5p33_ASAP7_75t_R g5983 ( 
.A(n_4371),
.Y(n_5983)
);

INVx1_ASAP7_75t_L g5984 ( 
.A(n_5671),
.Y(n_5984)
);

CKINVDCx5p33_ASAP7_75t_R g5985 ( 
.A(n_4372),
.Y(n_5985)
);

INVx1_ASAP7_75t_L g5986 ( 
.A(n_5671),
.Y(n_5986)
);

CKINVDCx20_ASAP7_75t_R g5987 ( 
.A(n_4417),
.Y(n_5987)
);

INVx1_ASAP7_75t_L g5988 ( 
.A(n_5671),
.Y(n_5988)
);

NOR2xp67_ASAP7_75t_L g5989 ( 
.A(n_4706),
.B(n_4),
.Y(n_5989)
);

CKINVDCx5p33_ASAP7_75t_R g5990 ( 
.A(n_4373),
.Y(n_5990)
);

BUFx6f_ASAP7_75t_L g5991 ( 
.A(n_5685),
.Y(n_5991)
);

CKINVDCx5p33_ASAP7_75t_R g5992 ( 
.A(n_4374),
.Y(n_5992)
);

CKINVDCx20_ASAP7_75t_R g5993 ( 
.A(n_4464),
.Y(n_5993)
);

INVx1_ASAP7_75t_L g5994 ( 
.A(n_5685),
.Y(n_5994)
);

CKINVDCx5p33_ASAP7_75t_R g5995 ( 
.A(n_4375),
.Y(n_5995)
);

INVx2_ASAP7_75t_L g5996 ( 
.A(n_5685),
.Y(n_5996)
);

CKINVDCx5p33_ASAP7_75t_R g5997 ( 
.A(n_4379),
.Y(n_5997)
);

CKINVDCx20_ASAP7_75t_R g5998 ( 
.A(n_4469),
.Y(n_5998)
);

CKINVDCx5p33_ASAP7_75t_R g5999 ( 
.A(n_4380),
.Y(n_5999)
);

NOR2xp33_ASAP7_75t_L g6000 ( 
.A(n_5406),
.B(n_5),
.Y(n_6000)
);

INVx1_ASAP7_75t_L g6001 ( 
.A(n_5686),
.Y(n_6001)
);

BUFx5_ASAP7_75t_L g6002 ( 
.A(n_4330),
.Y(n_6002)
);

CKINVDCx5p33_ASAP7_75t_R g6003 ( 
.A(n_4383),
.Y(n_6003)
);

CKINVDCx5p33_ASAP7_75t_R g6004 ( 
.A(n_4386),
.Y(n_6004)
);

CKINVDCx5p33_ASAP7_75t_R g6005 ( 
.A(n_4387),
.Y(n_6005)
);

CKINVDCx5p33_ASAP7_75t_R g6006 ( 
.A(n_4388),
.Y(n_6006)
);

INVx1_ASAP7_75t_L g6007 ( 
.A(n_5686),
.Y(n_6007)
);

OR2x2_ASAP7_75t_L g6008 ( 
.A(n_5466),
.B(n_5),
.Y(n_6008)
);

INVx1_ASAP7_75t_L g6009 ( 
.A(n_5686),
.Y(n_6009)
);

CKINVDCx5p33_ASAP7_75t_R g6010 ( 
.A(n_4391),
.Y(n_6010)
);

BUFx5_ASAP7_75t_L g6011 ( 
.A(n_4336),
.Y(n_6011)
);

INVx2_ASAP7_75t_L g6012 ( 
.A(n_5721),
.Y(n_6012)
);

BUFx3_ASAP7_75t_L g6013 ( 
.A(n_4722),
.Y(n_6013)
);

BUFx3_ASAP7_75t_L g6014 ( 
.A(n_4789),
.Y(n_6014)
);

CKINVDCx5p33_ASAP7_75t_R g6015 ( 
.A(n_4394),
.Y(n_6015)
);

CKINVDCx5p33_ASAP7_75t_R g6016 ( 
.A(n_4395),
.Y(n_6016)
);

CKINVDCx5p33_ASAP7_75t_R g6017 ( 
.A(n_4398),
.Y(n_6017)
);

CKINVDCx5p33_ASAP7_75t_R g6018 ( 
.A(n_4399),
.Y(n_6018)
);

BUFx2_ASAP7_75t_L g6019 ( 
.A(n_5548),
.Y(n_6019)
);

CKINVDCx5p33_ASAP7_75t_R g6020 ( 
.A(n_4400),
.Y(n_6020)
);

BUFx2_ASAP7_75t_L g6021 ( 
.A(n_5553),
.Y(n_6021)
);

CKINVDCx5p33_ASAP7_75t_R g6022 ( 
.A(n_4401),
.Y(n_6022)
);

INVx1_ASAP7_75t_L g6023 ( 
.A(n_5721),
.Y(n_6023)
);

INVxp33_ASAP7_75t_L g6024 ( 
.A(n_4624),
.Y(n_6024)
);

INVx1_ASAP7_75t_L g6025 ( 
.A(n_5721),
.Y(n_6025)
);

CKINVDCx20_ASAP7_75t_R g6026 ( 
.A(n_4493),
.Y(n_6026)
);

CKINVDCx20_ASAP7_75t_R g6027 ( 
.A(n_4507),
.Y(n_6027)
);

CKINVDCx20_ASAP7_75t_R g6028 ( 
.A(n_4526),
.Y(n_6028)
);

INVx2_ASAP7_75t_L g6029 ( 
.A(n_5727),
.Y(n_6029)
);

INVx1_ASAP7_75t_L g6030 ( 
.A(n_5727),
.Y(n_6030)
);

CKINVDCx5p33_ASAP7_75t_R g6031 ( 
.A(n_4404),
.Y(n_6031)
);

CKINVDCx5p33_ASAP7_75t_R g6032 ( 
.A(n_4405),
.Y(n_6032)
);

INVx2_ASAP7_75t_L g6033 ( 
.A(n_5727),
.Y(n_6033)
);

CKINVDCx5p33_ASAP7_75t_R g6034 ( 
.A(n_4407),
.Y(n_6034)
);

INVx1_ASAP7_75t_L g6035 ( 
.A(n_4818),
.Y(n_6035)
);

CKINVDCx5p33_ASAP7_75t_R g6036 ( 
.A(n_4408),
.Y(n_6036)
);

INVx1_ASAP7_75t_L g6037 ( 
.A(n_4826),
.Y(n_6037)
);

INVx1_ASAP7_75t_L g6038 ( 
.A(n_4835),
.Y(n_6038)
);

INVx1_ASAP7_75t_L g6039 ( 
.A(n_4903),
.Y(n_6039)
);

CKINVDCx5p33_ASAP7_75t_R g6040 ( 
.A(n_4410),
.Y(n_6040)
);

INVx1_ASAP7_75t_L g6041 ( 
.A(n_4922),
.Y(n_6041)
);

CKINVDCx5p33_ASAP7_75t_R g6042 ( 
.A(n_4411),
.Y(n_6042)
);

INVx1_ASAP7_75t_L g6043 ( 
.A(n_4956),
.Y(n_6043)
);

INVx1_ASAP7_75t_L g6044 ( 
.A(n_4984),
.Y(n_6044)
);

CKINVDCx5p33_ASAP7_75t_R g6045 ( 
.A(n_4412),
.Y(n_6045)
);

INVx1_ASAP7_75t_L g6046 ( 
.A(n_5008),
.Y(n_6046)
);

CKINVDCx5p33_ASAP7_75t_R g6047 ( 
.A(n_4419),
.Y(n_6047)
);

NOR2xp67_ASAP7_75t_L g6048 ( 
.A(n_4773),
.B(n_6),
.Y(n_6048)
);

BUFx3_ASAP7_75t_L g6049 ( 
.A(n_5135),
.Y(n_6049)
);

CKINVDCx5p33_ASAP7_75t_R g6050 ( 
.A(n_4422),
.Y(n_6050)
);

BUFx2_ASAP7_75t_L g6051 ( 
.A(n_5164),
.Y(n_6051)
);

INVx1_ASAP7_75t_L g6052 ( 
.A(n_5362),
.Y(n_6052)
);

BUFx6f_ASAP7_75t_L g6053 ( 
.A(n_5422),
.Y(n_6053)
);

INVx1_ASAP7_75t_SL g6054 ( 
.A(n_4719),
.Y(n_6054)
);

CKINVDCx5p33_ASAP7_75t_R g6055 ( 
.A(n_4423),
.Y(n_6055)
);

CKINVDCx20_ASAP7_75t_R g6056 ( 
.A(n_4565),
.Y(n_6056)
);

INVx1_ASAP7_75t_L g6057 ( 
.A(n_5501),
.Y(n_6057)
);

CKINVDCx16_ASAP7_75t_R g6058 ( 
.A(n_4345),
.Y(n_6058)
);

BUFx3_ASAP7_75t_L g6059 ( 
.A(n_5503),
.Y(n_6059)
);

CKINVDCx5p33_ASAP7_75t_R g6060 ( 
.A(n_4425),
.Y(n_6060)
);

BUFx6f_ASAP7_75t_L g6061 ( 
.A(n_5536),
.Y(n_6061)
);

CKINVDCx5p33_ASAP7_75t_R g6062 ( 
.A(n_4429),
.Y(n_6062)
);

CKINVDCx5p33_ASAP7_75t_R g6063 ( 
.A(n_4430),
.Y(n_6063)
);

CKINVDCx5p33_ASAP7_75t_R g6064 ( 
.A(n_4431),
.Y(n_6064)
);

INVx1_ASAP7_75t_L g6065 ( 
.A(n_5542),
.Y(n_6065)
);

CKINVDCx5p33_ASAP7_75t_R g6066 ( 
.A(n_4432),
.Y(n_6066)
);

CKINVDCx16_ASAP7_75t_R g6067 ( 
.A(n_4345),
.Y(n_6067)
);

INVx1_ASAP7_75t_L g6068 ( 
.A(n_5556),
.Y(n_6068)
);

INVxp33_ASAP7_75t_SL g6069 ( 
.A(n_4669),
.Y(n_6069)
);

CKINVDCx16_ASAP7_75t_R g6070 ( 
.A(n_5724),
.Y(n_6070)
);

INVx1_ASAP7_75t_L g6071 ( 
.A(n_5644),
.Y(n_6071)
);

INVx1_ASAP7_75t_L g6072 ( 
.A(n_5740),
.Y(n_6072)
);

INVx1_ASAP7_75t_L g6073 ( 
.A(n_5745),
.Y(n_6073)
);

INVx2_ASAP7_75t_L g6074 ( 
.A(n_4347),
.Y(n_6074)
);

CKINVDCx5p33_ASAP7_75t_R g6075 ( 
.A(n_4435),
.Y(n_6075)
);

INVx1_ASAP7_75t_L g6076 ( 
.A(n_5730),
.Y(n_6076)
);

BUFx10_ASAP7_75t_L g6077 ( 
.A(n_4929),
.Y(n_6077)
);

CKINVDCx5p33_ASAP7_75t_R g6078 ( 
.A(n_4436),
.Y(n_6078)
);

INVx1_ASAP7_75t_L g6079 ( 
.A(n_5743),
.Y(n_6079)
);

CKINVDCx5p33_ASAP7_75t_R g6080 ( 
.A(n_4440),
.Y(n_6080)
);

INVx2_ASAP7_75t_L g6081 ( 
.A(n_4350),
.Y(n_6081)
);

CKINVDCx5p33_ASAP7_75t_R g6082 ( 
.A(n_4441),
.Y(n_6082)
);

CKINVDCx5p33_ASAP7_75t_R g6083 ( 
.A(n_4442),
.Y(n_6083)
);

INVx1_ASAP7_75t_L g6084 ( 
.A(n_4352),
.Y(n_6084)
);

INVx2_ASAP7_75t_L g6085 ( 
.A(n_4369),
.Y(n_6085)
);

INVx2_ASAP7_75t_SL g6086 ( 
.A(n_4382),
.Y(n_6086)
);

INVx1_ASAP7_75t_L g6087 ( 
.A(n_5716),
.Y(n_6087)
);

INVx1_ASAP7_75t_L g6088 ( 
.A(n_5720),
.Y(n_6088)
);

INVx1_ASAP7_75t_L g6089 ( 
.A(n_5741),
.Y(n_6089)
);

CKINVDCx5p33_ASAP7_75t_R g6090 ( 
.A(n_5717),
.Y(n_6090)
);

CKINVDCx5p33_ASAP7_75t_R g6091 ( 
.A(n_5719),
.Y(n_6091)
);

INVx1_ASAP7_75t_L g6092 ( 
.A(n_5744),
.Y(n_6092)
);

CKINVDCx5p33_ASAP7_75t_R g6093 ( 
.A(n_4446),
.Y(n_6093)
);

CKINVDCx5p33_ASAP7_75t_R g6094 ( 
.A(n_4449),
.Y(n_6094)
);

BUFx10_ASAP7_75t_L g6095 ( 
.A(n_5070),
.Y(n_6095)
);

INVx1_ASAP7_75t_L g6096 ( 
.A(n_5747),
.Y(n_6096)
);

CKINVDCx5p33_ASAP7_75t_R g6097 ( 
.A(n_4450),
.Y(n_6097)
);

INVx1_ASAP7_75t_L g6098 ( 
.A(n_5748),
.Y(n_6098)
);

CKINVDCx5p33_ASAP7_75t_R g6099 ( 
.A(n_4451),
.Y(n_6099)
);

CKINVDCx5p33_ASAP7_75t_R g6100 ( 
.A(n_4452),
.Y(n_6100)
);

CKINVDCx5p33_ASAP7_75t_R g6101 ( 
.A(n_4453),
.Y(n_6101)
);

CKINVDCx5p33_ASAP7_75t_R g6102 ( 
.A(n_4459),
.Y(n_6102)
);

BUFx3_ASAP7_75t_L g6103 ( 
.A(n_4382),
.Y(n_6103)
);

INVx1_ASAP7_75t_L g6104 ( 
.A(n_5710),
.Y(n_6104)
);

CKINVDCx5p33_ASAP7_75t_R g6105 ( 
.A(n_5708),
.Y(n_6105)
);

CKINVDCx5p33_ASAP7_75t_R g6106 ( 
.A(n_5711),
.Y(n_6106)
);

INVx1_ASAP7_75t_L g6107 ( 
.A(n_4381),
.Y(n_6107)
);

INVx2_ASAP7_75t_L g6108 ( 
.A(n_4385),
.Y(n_6108)
);

BUFx5_ASAP7_75t_L g6109 ( 
.A(n_4389),
.Y(n_6109)
);

INVx1_ASAP7_75t_L g6110 ( 
.A(n_4392),
.Y(n_6110)
);

CKINVDCx20_ASAP7_75t_R g6111 ( 
.A(n_4568),
.Y(n_6111)
);

INVx1_ASAP7_75t_L g6112 ( 
.A(n_4393),
.Y(n_6112)
);

CKINVDCx5p33_ASAP7_75t_R g6113 ( 
.A(n_4462),
.Y(n_6113)
);

INVx1_ASAP7_75t_L g6114 ( 
.A(n_4396),
.Y(n_6114)
);

CKINVDCx5p33_ASAP7_75t_R g6115 ( 
.A(n_4463),
.Y(n_6115)
);

INVx1_ASAP7_75t_L g6116 ( 
.A(n_4402),
.Y(n_6116)
);

INVx1_ASAP7_75t_L g6117 ( 
.A(n_4406),
.Y(n_6117)
);

CKINVDCx5p33_ASAP7_75t_R g6118 ( 
.A(n_4465),
.Y(n_6118)
);

NOR2xp33_ASAP7_75t_L g6119 ( 
.A(n_5300),
.B(n_6),
.Y(n_6119)
);

CKINVDCx5p33_ASAP7_75t_R g6120 ( 
.A(n_5705),
.Y(n_6120)
);

CKINVDCx16_ASAP7_75t_R g6121 ( 
.A(n_5724),
.Y(n_6121)
);

CKINVDCx5p33_ASAP7_75t_R g6122 ( 
.A(n_5707),
.Y(n_6122)
);

CKINVDCx5p33_ASAP7_75t_R g6123 ( 
.A(n_5712),
.Y(n_6123)
);

INVx1_ASAP7_75t_L g6124 ( 
.A(n_5706),
.Y(n_6124)
);

INVx2_ASAP7_75t_SL g6125 ( 
.A(n_4434),
.Y(n_6125)
);

BUFx5_ASAP7_75t_L g6126 ( 
.A(n_4409),
.Y(n_6126)
);

INVxp67_ASAP7_75t_SL g6127 ( 
.A(n_5342),
.Y(n_6127)
);

INVx1_ASAP7_75t_L g6128 ( 
.A(n_4416),
.Y(n_6128)
);

CKINVDCx16_ASAP7_75t_R g6129 ( 
.A(n_4434),
.Y(n_6129)
);

OR2x2_ASAP7_75t_L g6130 ( 
.A(n_5390),
.B(n_7),
.Y(n_6130)
);

BUFx3_ASAP7_75t_L g6131 ( 
.A(n_4470),
.Y(n_6131)
);

CKINVDCx16_ASAP7_75t_R g6132 ( 
.A(n_4470),
.Y(n_6132)
);

CKINVDCx5p33_ASAP7_75t_R g6133 ( 
.A(n_4466),
.Y(n_6133)
);

INVx1_ASAP7_75t_L g6134 ( 
.A(n_4421),
.Y(n_6134)
);

CKINVDCx20_ASAP7_75t_R g6135 ( 
.A(n_4572),
.Y(n_6135)
);

INVx1_ASAP7_75t_SL g6136 ( 
.A(n_4620),
.Y(n_6136)
);

CKINVDCx20_ASAP7_75t_R g6137 ( 
.A(n_4576),
.Y(n_6137)
);

INVx1_ASAP7_75t_L g6138 ( 
.A(n_4424),
.Y(n_6138)
);

INVx1_ASAP7_75t_L g6139 ( 
.A(n_4426),
.Y(n_6139)
);

INVx1_ASAP7_75t_L g6140 ( 
.A(n_4427),
.Y(n_6140)
);

INVx1_ASAP7_75t_L g6141 ( 
.A(n_4428),
.Y(n_6141)
);

CKINVDCx5p33_ASAP7_75t_R g6142 ( 
.A(n_5714),
.Y(n_6142)
);

INVx1_ASAP7_75t_L g6143 ( 
.A(n_4433),
.Y(n_6143)
);

CKINVDCx5p33_ASAP7_75t_R g6144 ( 
.A(n_5715),
.Y(n_6144)
);

INVx2_ASAP7_75t_L g6145 ( 
.A(n_4438),
.Y(n_6145)
);

INVx1_ASAP7_75t_L g6146 ( 
.A(n_4439),
.Y(n_6146)
);

INVx2_ASAP7_75t_L g6147 ( 
.A(n_4444),
.Y(n_6147)
);

CKINVDCx5p33_ASAP7_75t_R g6148 ( 
.A(n_4467),
.Y(n_6148)
);

INVx1_ASAP7_75t_L g6149 ( 
.A(n_4445),
.Y(n_6149)
);

CKINVDCx5p33_ASAP7_75t_R g6150 ( 
.A(n_4468),
.Y(n_6150)
);

INVx1_ASAP7_75t_L g6151 ( 
.A(n_4448),
.Y(n_6151)
);

HB1xp67_ASAP7_75t_L g6152 ( 
.A(n_5528),
.Y(n_6152)
);

INVxp67_ASAP7_75t_L g6153 ( 
.A(n_5623),
.Y(n_6153)
);

INVx1_ASAP7_75t_L g6154 ( 
.A(n_4454),
.Y(n_6154)
);

CKINVDCx5p33_ASAP7_75t_R g6155 ( 
.A(n_5699),
.Y(n_6155)
);

INVx1_ASAP7_75t_L g6156 ( 
.A(n_4457),
.Y(n_6156)
);

CKINVDCx5p33_ASAP7_75t_R g6157 ( 
.A(n_5701),
.Y(n_6157)
);

INVx1_ASAP7_75t_L g6158 ( 
.A(n_4458),
.Y(n_6158)
);

CKINVDCx5p33_ASAP7_75t_R g6159 ( 
.A(n_5703),
.Y(n_6159)
);

CKINVDCx5p33_ASAP7_75t_R g6160 ( 
.A(n_4471),
.Y(n_6160)
);

BUFx3_ASAP7_75t_L g6161 ( 
.A(n_4548),
.Y(n_6161)
);

INVx1_ASAP7_75t_L g6162 ( 
.A(n_4460),
.Y(n_6162)
);

CKINVDCx5p33_ASAP7_75t_R g6163 ( 
.A(n_4472),
.Y(n_6163)
);

CKINVDCx5p33_ASAP7_75t_R g6164 ( 
.A(n_4473),
.Y(n_6164)
);

INVx1_ASAP7_75t_L g6165 ( 
.A(n_4461),
.Y(n_6165)
);

BUFx2_ASAP7_75t_L g6166 ( 
.A(n_5704),
.Y(n_6166)
);

CKINVDCx16_ASAP7_75t_R g6167 ( 
.A(n_4548),
.Y(n_6167)
);

INVx2_ASAP7_75t_L g6168 ( 
.A(n_4476),
.Y(n_6168)
);

INVx1_ASAP7_75t_L g6169 ( 
.A(n_4490),
.Y(n_6169)
);

INVx1_ASAP7_75t_L g6170 ( 
.A(n_5693),
.Y(n_6170)
);

CKINVDCx5p33_ASAP7_75t_R g6171 ( 
.A(n_5697),
.Y(n_6171)
);

INVx1_ASAP7_75t_L g6172 ( 
.A(n_5694),
.Y(n_6172)
);

BUFx6f_ASAP7_75t_L g6173 ( 
.A(n_4358),
.Y(n_6173)
);

INVx1_ASAP7_75t_L g6174 ( 
.A(n_5696),
.Y(n_6174)
);

INVx1_ASAP7_75t_L g6175 ( 
.A(n_4495),
.Y(n_6175)
);

CKINVDCx5p33_ASAP7_75t_R g6176 ( 
.A(n_5702),
.Y(n_6176)
);

CKINVDCx20_ASAP7_75t_R g6177 ( 
.A(n_4584),
.Y(n_6177)
);

INVxp67_ASAP7_75t_L g6178 ( 
.A(n_4595),
.Y(n_6178)
);

INVx1_ASAP7_75t_L g6179 ( 
.A(n_4498),
.Y(n_6179)
);

INVx1_ASAP7_75t_L g6180 ( 
.A(n_4506),
.Y(n_6180)
);

CKINVDCx5p33_ASAP7_75t_R g6181 ( 
.A(n_4474),
.Y(n_6181)
);

CKINVDCx5p33_ASAP7_75t_R g6182 ( 
.A(n_4475),
.Y(n_6182)
);

INVx1_ASAP7_75t_SL g6183 ( 
.A(n_4831),
.Y(n_6183)
);

CKINVDCx20_ASAP7_75t_R g6184 ( 
.A(n_4622),
.Y(n_6184)
);

INVxp67_ASAP7_75t_L g6185 ( 
.A(n_4595),
.Y(n_6185)
);

INVx1_ASAP7_75t_L g6186 ( 
.A(n_4509),
.Y(n_6186)
);

INVx1_ASAP7_75t_L g6187 ( 
.A(n_5689),
.Y(n_6187)
);

CKINVDCx5p33_ASAP7_75t_R g6188 ( 
.A(n_5691),
.Y(n_6188)
);

INVx2_ASAP7_75t_L g6189 ( 
.A(n_4510),
.Y(n_6189)
);

INVx2_ASAP7_75t_SL g6190 ( 
.A(n_4720),
.Y(n_6190)
);

INVx1_ASAP7_75t_L g6191 ( 
.A(n_5695),
.Y(n_6191)
);

INVx1_ASAP7_75t_L g6192 ( 
.A(n_4516),
.Y(n_6192)
);

BUFx6f_ASAP7_75t_L g6193 ( 
.A(n_4363),
.Y(n_6193)
);

INVx1_ASAP7_75t_L g6194 ( 
.A(n_4517),
.Y(n_6194)
);

INVx1_ASAP7_75t_L g6195 ( 
.A(n_4518),
.Y(n_6195)
);

INVx1_ASAP7_75t_SL g6196 ( 
.A(n_4832),
.Y(n_6196)
);

INVxp67_ASAP7_75t_L g6197 ( 
.A(n_4720),
.Y(n_6197)
);

CKINVDCx5p33_ASAP7_75t_R g6198 ( 
.A(n_4477),
.Y(n_6198)
);

CKINVDCx5p33_ASAP7_75t_R g6199 ( 
.A(n_4478),
.Y(n_6199)
);

INVx1_ASAP7_75t_L g6200 ( 
.A(n_5774),
.Y(n_6200)
);

INVx1_ASAP7_75t_L g6201 ( 
.A(n_5774),
.Y(n_6201)
);

INVx1_ASAP7_75t_L g6202 ( 
.A(n_5774),
.Y(n_6202)
);

INVx1_ASAP7_75t_L g6203 ( 
.A(n_5852),
.Y(n_6203)
);

INVxp67_ASAP7_75t_L g6204 ( 
.A(n_5795),
.Y(n_6204)
);

INVx1_ASAP7_75t_L g6205 ( 
.A(n_5852),
.Y(n_6205)
);

CKINVDCx20_ASAP7_75t_R g6206 ( 
.A(n_5756),
.Y(n_6206)
);

CKINVDCx5p33_ASAP7_75t_R g6207 ( 
.A(n_5775),
.Y(n_6207)
);

INVxp33_ASAP7_75t_SL g6208 ( 
.A(n_5763),
.Y(n_6208)
);

INVx1_ASAP7_75t_L g6209 ( 
.A(n_5852),
.Y(n_6209)
);

CKINVDCx14_ASAP7_75t_R g6210 ( 
.A(n_5789),
.Y(n_6210)
);

INVx1_ASAP7_75t_L g6211 ( 
.A(n_5912),
.Y(n_6211)
);

INVxp67_ASAP7_75t_SL g6212 ( 
.A(n_5786),
.Y(n_6212)
);

BUFx2_ASAP7_75t_SL g6213 ( 
.A(n_5788),
.Y(n_6213)
);

CKINVDCx20_ASAP7_75t_R g6214 ( 
.A(n_5848),
.Y(n_6214)
);

INVx1_ASAP7_75t_L g6215 ( 
.A(n_5912),
.Y(n_6215)
);

INVx1_ASAP7_75t_L g6216 ( 
.A(n_5912),
.Y(n_6216)
);

INVx1_ASAP7_75t_L g6217 ( 
.A(n_5946),
.Y(n_6217)
);

INVx1_ASAP7_75t_L g6218 ( 
.A(n_5946),
.Y(n_6218)
);

CKINVDCx5p33_ASAP7_75t_R g6219 ( 
.A(n_5781),
.Y(n_6219)
);

INVxp67_ASAP7_75t_SL g6220 ( 
.A(n_5856),
.Y(n_6220)
);

CKINVDCx5p33_ASAP7_75t_R g6221 ( 
.A(n_5782),
.Y(n_6221)
);

CKINVDCx20_ASAP7_75t_R g6222 ( 
.A(n_5863),
.Y(n_6222)
);

INVxp33_ASAP7_75t_SL g6223 ( 
.A(n_5765),
.Y(n_6223)
);

INVx1_ASAP7_75t_L g6224 ( 
.A(n_5946),
.Y(n_6224)
);

BUFx2_ASAP7_75t_L g6225 ( 
.A(n_5828),
.Y(n_6225)
);

CKINVDCx20_ASAP7_75t_R g6226 ( 
.A(n_5873),
.Y(n_6226)
);

INVx1_ASAP7_75t_L g6227 ( 
.A(n_5991),
.Y(n_6227)
);

INVx1_ASAP7_75t_L g6228 ( 
.A(n_5991),
.Y(n_6228)
);

INVx1_ASAP7_75t_L g6229 ( 
.A(n_5991),
.Y(n_6229)
);

INVx1_ASAP7_75t_L g6230 ( 
.A(n_5884),
.Y(n_6230)
);

INVx1_ASAP7_75t_L g6231 ( 
.A(n_5888),
.Y(n_6231)
);

CKINVDCx20_ASAP7_75t_R g6232 ( 
.A(n_5900),
.Y(n_6232)
);

INVx1_ASAP7_75t_L g6233 ( 
.A(n_5895),
.Y(n_6233)
);

CKINVDCx5p33_ASAP7_75t_R g6234 ( 
.A(n_5784),
.Y(n_6234)
);

INVx2_ASAP7_75t_L g6235 ( 
.A(n_5904),
.Y(n_6235)
);

CKINVDCx20_ASAP7_75t_R g6236 ( 
.A(n_5924),
.Y(n_6236)
);

INVxp33_ASAP7_75t_L g6237 ( 
.A(n_5797),
.Y(n_6237)
);

INVx1_ASAP7_75t_L g6238 ( 
.A(n_5963),
.Y(n_6238)
);

CKINVDCx20_ASAP7_75t_R g6239 ( 
.A(n_5951),
.Y(n_6239)
);

CKINVDCx20_ASAP7_75t_R g6240 ( 
.A(n_5970),
.Y(n_6240)
);

INVx1_ASAP7_75t_L g6241 ( 
.A(n_5967),
.Y(n_6241)
);

INVxp67_ASAP7_75t_SL g6242 ( 
.A(n_5901),
.Y(n_6242)
);

INVx1_ASAP7_75t_L g6243 ( 
.A(n_5975),
.Y(n_6243)
);

INVx1_ASAP7_75t_L g6244 ( 
.A(n_5996),
.Y(n_6244)
);

INVx1_ASAP7_75t_L g6245 ( 
.A(n_6012),
.Y(n_6245)
);

INVx1_ASAP7_75t_L g6246 ( 
.A(n_6029),
.Y(n_6246)
);

CKINVDCx20_ASAP7_75t_R g6247 ( 
.A(n_5987),
.Y(n_6247)
);

INVx2_ASAP7_75t_L g6248 ( 
.A(n_6033),
.Y(n_6248)
);

INVx1_ASAP7_75t_L g6249 ( 
.A(n_5826),
.Y(n_6249)
);

CKINVDCx5p33_ASAP7_75t_R g6250 ( 
.A(n_5785),
.Y(n_6250)
);

CKINVDCx5p33_ASAP7_75t_R g6251 ( 
.A(n_5787),
.Y(n_6251)
);

INVx1_ASAP7_75t_L g6252 ( 
.A(n_5829),
.Y(n_6252)
);

INVx1_ASAP7_75t_L g6253 ( 
.A(n_5831),
.Y(n_6253)
);

INVx1_ASAP7_75t_L g6254 ( 
.A(n_5832),
.Y(n_6254)
);

INVx1_ASAP7_75t_L g6255 ( 
.A(n_5834),
.Y(n_6255)
);

INVx1_ASAP7_75t_L g6256 ( 
.A(n_5835),
.Y(n_6256)
);

INVx1_ASAP7_75t_L g6257 ( 
.A(n_5837),
.Y(n_6257)
);

INVx1_ASAP7_75t_L g6258 ( 
.A(n_5839),
.Y(n_6258)
);

INVx2_ASAP7_75t_L g6259 ( 
.A(n_5842),
.Y(n_6259)
);

CKINVDCx20_ASAP7_75t_R g6260 ( 
.A(n_5993),
.Y(n_6260)
);

INVx1_ASAP7_75t_L g6261 ( 
.A(n_5845),
.Y(n_6261)
);

CKINVDCx5p33_ASAP7_75t_R g6262 ( 
.A(n_5843),
.Y(n_6262)
);

INVx2_ASAP7_75t_L g6263 ( 
.A(n_5847),
.Y(n_6263)
);

INVx1_ASAP7_75t_L g6264 ( 
.A(n_5850),
.Y(n_6264)
);

INVx1_ASAP7_75t_L g6265 ( 
.A(n_5851),
.Y(n_6265)
);

INVx1_ASAP7_75t_L g6266 ( 
.A(n_5853),
.Y(n_6266)
);

INVx1_ASAP7_75t_L g6267 ( 
.A(n_5857),
.Y(n_6267)
);

INVx1_ASAP7_75t_L g6268 ( 
.A(n_5859),
.Y(n_6268)
);

INVx1_ASAP7_75t_L g6269 ( 
.A(n_5860),
.Y(n_6269)
);

CKINVDCx5p33_ASAP7_75t_R g6270 ( 
.A(n_5844),
.Y(n_6270)
);

INVx1_ASAP7_75t_L g6271 ( 
.A(n_5864),
.Y(n_6271)
);

INVx1_ASAP7_75t_L g6272 ( 
.A(n_5866),
.Y(n_6272)
);

INVx1_ASAP7_75t_L g6273 ( 
.A(n_5868),
.Y(n_6273)
);

INVx1_ASAP7_75t_L g6274 ( 
.A(n_5870),
.Y(n_6274)
);

CKINVDCx20_ASAP7_75t_R g6275 ( 
.A(n_5998),
.Y(n_6275)
);

CKINVDCx5p33_ASAP7_75t_R g6276 ( 
.A(n_5854),
.Y(n_6276)
);

INVx1_ASAP7_75t_L g6277 ( 
.A(n_5872),
.Y(n_6277)
);

CKINVDCx14_ASAP7_75t_R g6278 ( 
.A(n_5809),
.Y(n_6278)
);

INVxp67_ASAP7_75t_L g6279 ( 
.A(n_6051),
.Y(n_6279)
);

INVx1_ASAP7_75t_L g6280 ( 
.A(n_5875),
.Y(n_6280)
);

CKINVDCx5p33_ASAP7_75t_R g6281 ( 
.A(n_5858),
.Y(n_6281)
);

CKINVDCx20_ASAP7_75t_R g6282 ( 
.A(n_6026),
.Y(n_6282)
);

INVx1_ASAP7_75t_L g6283 ( 
.A(n_5876),
.Y(n_6283)
);

INVx1_ASAP7_75t_L g6284 ( 
.A(n_5877),
.Y(n_6284)
);

INVx2_ASAP7_75t_L g6285 ( 
.A(n_5881),
.Y(n_6285)
);

CKINVDCx16_ASAP7_75t_R g6286 ( 
.A(n_5793),
.Y(n_6286)
);

INVx1_ASAP7_75t_L g6287 ( 
.A(n_5886),
.Y(n_6287)
);

INVx1_ASAP7_75t_L g6288 ( 
.A(n_5891),
.Y(n_6288)
);

INVxp33_ASAP7_75t_SL g6289 ( 
.A(n_5771),
.Y(n_6289)
);

INVx2_ASAP7_75t_L g6290 ( 
.A(n_5893),
.Y(n_6290)
);

INVx1_ASAP7_75t_L g6291 ( 
.A(n_5896),
.Y(n_6291)
);

INVx2_ASAP7_75t_L g6292 ( 
.A(n_5899),
.Y(n_6292)
);

CKINVDCx5p33_ASAP7_75t_R g6293 ( 
.A(n_5861),
.Y(n_6293)
);

CKINVDCx5p33_ASAP7_75t_R g6294 ( 
.A(n_5862),
.Y(n_6294)
);

INVx1_ASAP7_75t_L g6295 ( 
.A(n_5903),
.Y(n_6295)
);

CKINVDCx16_ASAP7_75t_R g6296 ( 
.A(n_5830),
.Y(n_6296)
);

CKINVDCx20_ASAP7_75t_R g6297 ( 
.A(n_6027),
.Y(n_6297)
);

CKINVDCx5p33_ASAP7_75t_R g6298 ( 
.A(n_5865),
.Y(n_6298)
);

INVx1_ASAP7_75t_L g6299 ( 
.A(n_5905),
.Y(n_6299)
);

CKINVDCx5p33_ASAP7_75t_R g6300 ( 
.A(n_5869),
.Y(n_6300)
);

INVx1_ASAP7_75t_L g6301 ( 
.A(n_5907),
.Y(n_6301)
);

INVx1_ASAP7_75t_L g6302 ( 
.A(n_5909),
.Y(n_6302)
);

INVx2_ASAP7_75t_L g6303 ( 
.A(n_5910),
.Y(n_6303)
);

INVx1_ASAP7_75t_L g6304 ( 
.A(n_5914),
.Y(n_6304)
);

INVx2_ASAP7_75t_SL g6305 ( 
.A(n_6103),
.Y(n_6305)
);

INVx2_ASAP7_75t_L g6306 ( 
.A(n_5916),
.Y(n_6306)
);

INVxp67_ASAP7_75t_SL g6307 ( 
.A(n_5902),
.Y(n_6307)
);

INVx1_ASAP7_75t_L g6308 ( 
.A(n_5919),
.Y(n_6308)
);

INVx1_ASAP7_75t_L g6309 ( 
.A(n_5920),
.Y(n_6309)
);

INVx1_ASAP7_75t_L g6310 ( 
.A(n_5925),
.Y(n_6310)
);

CKINVDCx16_ASAP7_75t_R g6311 ( 
.A(n_5833),
.Y(n_6311)
);

INVx1_ASAP7_75t_L g6312 ( 
.A(n_5933),
.Y(n_6312)
);

BUFx2_ASAP7_75t_SL g6313 ( 
.A(n_6086),
.Y(n_6313)
);

CKINVDCx5p33_ASAP7_75t_R g6314 ( 
.A(n_5871),
.Y(n_6314)
);

INVxp67_ASAP7_75t_L g6315 ( 
.A(n_6131),
.Y(n_6315)
);

CKINVDCx5p33_ASAP7_75t_R g6316 ( 
.A(n_5878),
.Y(n_6316)
);

INVx1_ASAP7_75t_L g6317 ( 
.A(n_5936),
.Y(n_6317)
);

INVxp67_ASAP7_75t_SL g6318 ( 
.A(n_5931),
.Y(n_6318)
);

INVx1_ASAP7_75t_L g6319 ( 
.A(n_5940),
.Y(n_6319)
);

CKINVDCx16_ASAP7_75t_R g6320 ( 
.A(n_5846),
.Y(n_6320)
);

INVx1_ASAP7_75t_L g6321 ( 
.A(n_5941),
.Y(n_6321)
);

CKINVDCx5p33_ASAP7_75t_R g6322 ( 
.A(n_5879),
.Y(n_6322)
);

INVx1_ASAP7_75t_L g6323 ( 
.A(n_5942),
.Y(n_6323)
);

INVx1_ASAP7_75t_L g6324 ( 
.A(n_5944),
.Y(n_6324)
);

CKINVDCx5p33_ASAP7_75t_R g6325 ( 
.A(n_5880),
.Y(n_6325)
);

INVx2_ASAP7_75t_L g6326 ( 
.A(n_5945),
.Y(n_6326)
);

INVx1_ASAP7_75t_L g6327 ( 
.A(n_5947),
.Y(n_6327)
);

INVx1_ASAP7_75t_L g6328 ( 
.A(n_5952),
.Y(n_6328)
);

INVx1_ASAP7_75t_L g6329 ( 
.A(n_5958),
.Y(n_6329)
);

INVx1_ASAP7_75t_L g6330 ( 
.A(n_5959),
.Y(n_6330)
);

INVx1_ASAP7_75t_L g6331 ( 
.A(n_5962),
.Y(n_6331)
);

CKINVDCx20_ASAP7_75t_R g6332 ( 
.A(n_6028),
.Y(n_6332)
);

CKINVDCx20_ASAP7_75t_R g6333 ( 
.A(n_6056),
.Y(n_6333)
);

INVx1_ASAP7_75t_L g6334 ( 
.A(n_5966),
.Y(n_6334)
);

INVx1_ASAP7_75t_L g6335 ( 
.A(n_5969),
.Y(n_6335)
);

CKINVDCx14_ASAP7_75t_R g6336 ( 
.A(n_5961),
.Y(n_6336)
);

INVxp67_ASAP7_75t_SL g6337 ( 
.A(n_5943),
.Y(n_6337)
);

CKINVDCx20_ASAP7_75t_R g6338 ( 
.A(n_6111),
.Y(n_6338)
);

INVxp67_ASAP7_75t_SL g6339 ( 
.A(n_6013),
.Y(n_6339)
);

CKINVDCx5p33_ASAP7_75t_R g6340 ( 
.A(n_5883),
.Y(n_6340)
);

CKINVDCx5p33_ASAP7_75t_R g6341 ( 
.A(n_5887),
.Y(n_6341)
);

CKINVDCx5p33_ASAP7_75t_R g6342 ( 
.A(n_5889),
.Y(n_6342)
);

INVx1_ASAP7_75t_L g6343 ( 
.A(n_5971),
.Y(n_6343)
);

CKINVDCx5p33_ASAP7_75t_R g6344 ( 
.A(n_5890),
.Y(n_6344)
);

INVx1_ASAP7_75t_L g6345 ( 
.A(n_5973),
.Y(n_6345)
);

INVxp67_ASAP7_75t_SL g6346 ( 
.A(n_6014),
.Y(n_6346)
);

INVx2_ASAP7_75t_L g6347 ( 
.A(n_5974),
.Y(n_6347)
);

BUFx3_ASAP7_75t_L g6348 ( 
.A(n_6049),
.Y(n_6348)
);

CKINVDCx20_ASAP7_75t_R g6349 ( 
.A(n_6135),
.Y(n_6349)
);

INVx1_ASAP7_75t_L g6350 ( 
.A(n_5977),
.Y(n_6350)
);

INVxp67_ASAP7_75t_SL g6351 ( 
.A(n_6059),
.Y(n_6351)
);

CKINVDCx14_ASAP7_75t_R g6352 ( 
.A(n_5982),
.Y(n_6352)
);

INVx1_ASAP7_75t_L g6353 ( 
.A(n_5978),
.Y(n_6353)
);

CKINVDCx20_ASAP7_75t_R g6354 ( 
.A(n_6137),
.Y(n_6354)
);

CKINVDCx5p33_ASAP7_75t_R g6355 ( 
.A(n_5892),
.Y(n_6355)
);

INVx1_ASAP7_75t_L g6356 ( 
.A(n_5979),
.Y(n_6356)
);

CKINVDCx5p33_ASAP7_75t_R g6357 ( 
.A(n_5898),
.Y(n_6357)
);

INVx1_ASAP7_75t_L g6358 ( 
.A(n_5984),
.Y(n_6358)
);

INVx2_ASAP7_75t_L g6359 ( 
.A(n_5986),
.Y(n_6359)
);

INVx1_ASAP7_75t_L g6360 ( 
.A(n_5988),
.Y(n_6360)
);

BUFx2_ASAP7_75t_L g6361 ( 
.A(n_5798),
.Y(n_6361)
);

INVx1_ASAP7_75t_L g6362 ( 
.A(n_5994),
.Y(n_6362)
);

HB1xp67_ASAP7_75t_L g6363 ( 
.A(n_5800),
.Y(n_6363)
);

INVx1_ASAP7_75t_L g6364 ( 
.A(n_6001),
.Y(n_6364)
);

INVx1_ASAP7_75t_L g6365 ( 
.A(n_6007),
.Y(n_6365)
);

INVx1_ASAP7_75t_L g6366 ( 
.A(n_6009),
.Y(n_6366)
);

INVx1_ASAP7_75t_L g6367 ( 
.A(n_6023),
.Y(n_6367)
);

INVx1_ASAP7_75t_L g6368 ( 
.A(n_6025),
.Y(n_6368)
);

INVx1_ASAP7_75t_L g6369 ( 
.A(n_6030),
.Y(n_6369)
);

INVx1_ASAP7_75t_L g6370 ( 
.A(n_6053),
.Y(n_6370)
);

CKINVDCx5p33_ASAP7_75t_R g6371 ( 
.A(n_5906),
.Y(n_6371)
);

CKINVDCx5p33_ASAP7_75t_R g6372 ( 
.A(n_5908),
.Y(n_6372)
);

INVx1_ASAP7_75t_L g6373 ( 
.A(n_6053),
.Y(n_6373)
);

INVx1_ASAP7_75t_L g6374 ( 
.A(n_6053),
.Y(n_6374)
);

INVx1_ASAP7_75t_L g6375 ( 
.A(n_6061),
.Y(n_6375)
);

INVxp67_ASAP7_75t_L g6376 ( 
.A(n_6161),
.Y(n_6376)
);

INVx1_ASAP7_75t_L g6377 ( 
.A(n_6061),
.Y(n_6377)
);

INVx1_ASAP7_75t_L g6378 ( 
.A(n_6061),
.Y(n_6378)
);

HB1xp67_ASAP7_75t_L g6379 ( 
.A(n_5801),
.Y(n_6379)
);

INVx2_ASAP7_75t_L g6380 ( 
.A(n_5776),
.Y(n_6380)
);

INVx1_ASAP7_75t_L g6381 ( 
.A(n_5754),
.Y(n_6381)
);

INVx1_ASAP7_75t_L g6382 ( 
.A(n_5758),
.Y(n_6382)
);

CKINVDCx16_ASAP7_75t_R g6383 ( 
.A(n_5867),
.Y(n_6383)
);

INVx2_ASAP7_75t_L g6384 ( 
.A(n_5777),
.Y(n_6384)
);

CKINVDCx5p33_ASAP7_75t_R g6385 ( 
.A(n_5911),
.Y(n_6385)
);

INVx1_ASAP7_75t_L g6386 ( 
.A(n_5759),
.Y(n_6386)
);

INVxp67_ASAP7_75t_SL g6387 ( 
.A(n_5825),
.Y(n_6387)
);

CKINVDCx5p33_ASAP7_75t_R g6388 ( 
.A(n_5913),
.Y(n_6388)
);

INVx1_ASAP7_75t_L g6389 ( 
.A(n_5760),
.Y(n_6389)
);

INVx1_ASAP7_75t_L g6390 ( 
.A(n_5761),
.Y(n_6390)
);

CKINVDCx5p33_ASAP7_75t_R g6391 ( 
.A(n_5915),
.Y(n_6391)
);

INVx2_ASAP7_75t_L g6392 ( 
.A(n_5779),
.Y(n_6392)
);

HB1xp67_ASAP7_75t_L g6393 ( 
.A(n_5804),
.Y(n_6393)
);

INVx1_ASAP7_75t_L g6394 ( 
.A(n_5762),
.Y(n_6394)
);

CKINVDCx20_ASAP7_75t_R g6395 ( 
.A(n_6177),
.Y(n_6395)
);

BUFx3_ASAP7_75t_L g6396 ( 
.A(n_6035),
.Y(n_6396)
);

INVx1_ASAP7_75t_L g6397 ( 
.A(n_5766),
.Y(n_6397)
);

INVx1_ASAP7_75t_L g6398 ( 
.A(n_5768),
.Y(n_6398)
);

CKINVDCx5p33_ASAP7_75t_R g6399 ( 
.A(n_5918),
.Y(n_6399)
);

CKINVDCx20_ASAP7_75t_R g6400 ( 
.A(n_6184),
.Y(n_6400)
);

INVx1_ASAP7_75t_L g6401 ( 
.A(n_5769),
.Y(n_6401)
);

INVx1_ASAP7_75t_L g6402 ( 
.A(n_5772),
.Y(n_6402)
);

INVx1_ASAP7_75t_L g6403 ( 
.A(n_5778),
.Y(n_6403)
);

INVx1_ASAP7_75t_L g6404 ( 
.A(n_5783),
.Y(n_6404)
);

INVx1_ASAP7_75t_L g6405 ( 
.A(n_5799),
.Y(n_6405)
);

CKINVDCx5p33_ASAP7_75t_R g6406 ( 
.A(n_5921),
.Y(n_6406)
);

INVxp33_ASAP7_75t_SL g6407 ( 
.A(n_5753),
.Y(n_6407)
);

INVx3_ASAP7_75t_L g6408 ( 
.A(n_6173),
.Y(n_6408)
);

CKINVDCx5p33_ASAP7_75t_R g6409 ( 
.A(n_5922),
.Y(n_6409)
);

INVx1_ASAP7_75t_L g6410 ( 
.A(n_5802),
.Y(n_6410)
);

CKINVDCx5p33_ASAP7_75t_R g6411 ( 
.A(n_5923),
.Y(n_6411)
);

CKINVDCx16_ASAP7_75t_R g6412 ( 
.A(n_5885),
.Y(n_6412)
);

CKINVDCx16_ASAP7_75t_R g6413 ( 
.A(n_5956),
.Y(n_6413)
);

CKINVDCx5p33_ASAP7_75t_R g6414 ( 
.A(n_5926),
.Y(n_6414)
);

BUFx3_ASAP7_75t_L g6415 ( 
.A(n_6037),
.Y(n_6415)
);

INVx1_ASAP7_75t_SL g6416 ( 
.A(n_6054),
.Y(n_6416)
);

INVxp67_ASAP7_75t_SL g6417 ( 
.A(n_6000),
.Y(n_6417)
);

INVx1_ASAP7_75t_L g6418 ( 
.A(n_5807),
.Y(n_6418)
);

INVx1_ASAP7_75t_L g6419 ( 
.A(n_5811),
.Y(n_6419)
);

INVx1_ASAP7_75t_L g6420 ( 
.A(n_5812),
.Y(n_6420)
);

INVx1_ASAP7_75t_L g6421 ( 
.A(n_5816),
.Y(n_6421)
);

CKINVDCx5p33_ASAP7_75t_R g6422 ( 
.A(n_5927),
.Y(n_6422)
);

INVx1_ASAP7_75t_L g6423 ( 
.A(n_5820),
.Y(n_6423)
);

INVx1_ASAP7_75t_L g6424 ( 
.A(n_5821),
.Y(n_6424)
);

INVx1_ASAP7_75t_L g6425 ( 
.A(n_5823),
.Y(n_6425)
);

CKINVDCx5p33_ASAP7_75t_R g6426 ( 
.A(n_5929),
.Y(n_6426)
);

INVx1_ASAP7_75t_L g6427 ( 
.A(n_5824),
.Y(n_6427)
);

INVx1_ASAP7_75t_L g6428 ( 
.A(n_6076),
.Y(n_6428)
);

CKINVDCx20_ASAP7_75t_R g6429 ( 
.A(n_5805),
.Y(n_6429)
);

INVx1_ASAP7_75t_L g6430 ( 
.A(n_6079),
.Y(n_6430)
);

INVx1_ASAP7_75t_L g6431 ( 
.A(n_6084),
.Y(n_6431)
);

INVx1_ASAP7_75t_L g6432 ( 
.A(n_6087),
.Y(n_6432)
);

INVxp33_ASAP7_75t_L g6433 ( 
.A(n_5948),
.Y(n_6433)
);

INVx1_ASAP7_75t_L g6434 ( 
.A(n_6088),
.Y(n_6434)
);

CKINVDCx5p33_ASAP7_75t_R g6435 ( 
.A(n_5932),
.Y(n_6435)
);

INVx1_ASAP7_75t_L g6436 ( 
.A(n_6089),
.Y(n_6436)
);

HB1xp67_ASAP7_75t_L g6437 ( 
.A(n_5806),
.Y(n_6437)
);

CKINVDCx20_ASAP7_75t_R g6438 ( 
.A(n_5808),
.Y(n_6438)
);

CKINVDCx20_ASAP7_75t_R g6439 ( 
.A(n_5810),
.Y(n_6439)
);

INVx1_ASAP7_75t_L g6440 ( 
.A(n_6092),
.Y(n_6440)
);

CKINVDCx5p33_ASAP7_75t_R g6441 ( 
.A(n_5934),
.Y(n_6441)
);

CKINVDCx20_ASAP7_75t_R g6442 ( 
.A(n_5813),
.Y(n_6442)
);

CKINVDCx20_ASAP7_75t_R g6443 ( 
.A(n_5815),
.Y(n_6443)
);

INVx1_ASAP7_75t_L g6444 ( 
.A(n_6096),
.Y(n_6444)
);

INVx1_ASAP7_75t_L g6445 ( 
.A(n_6098),
.Y(n_6445)
);

CKINVDCx5p33_ASAP7_75t_R g6446 ( 
.A(n_5935),
.Y(n_6446)
);

INVxp33_ASAP7_75t_SL g6447 ( 
.A(n_5818),
.Y(n_6447)
);

INVx1_ASAP7_75t_L g6448 ( 
.A(n_6104),
.Y(n_6448)
);

INVxp67_ASAP7_75t_L g6449 ( 
.A(n_6125),
.Y(n_6449)
);

INVx1_ASAP7_75t_L g6450 ( 
.A(n_6107),
.Y(n_6450)
);

BUFx6f_ASAP7_75t_L g6451 ( 
.A(n_6173),
.Y(n_6451)
);

XNOR2xp5_ASAP7_75t_L g6452 ( 
.A(n_6136),
.B(n_6183),
.Y(n_6452)
);

INVxp67_ASAP7_75t_SL g6453 ( 
.A(n_6119),
.Y(n_6453)
);

CKINVDCx16_ASAP7_75t_R g6454 ( 
.A(n_6058),
.Y(n_6454)
);

BUFx2_ASAP7_75t_L g6455 ( 
.A(n_5822),
.Y(n_6455)
);

INVx1_ASAP7_75t_SL g6456 ( 
.A(n_6196),
.Y(n_6456)
);

INVx1_ASAP7_75t_L g6457 ( 
.A(n_6110),
.Y(n_6457)
);

INVx1_ASAP7_75t_L g6458 ( 
.A(n_6112),
.Y(n_6458)
);

INVx1_ASAP7_75t_L g6459 ( 
.A(n_6114),
.Y(n_6459)
);

INVx1_ASAP7_75t_L g6460 ( 
.A(n_6116),
.Y(n_6460)
);

INVxp67_ASAP7_75t_SL g6461 ( 
.A(n_6038),
.Y(n_6461)
);

INVx1_ASAP7_75t_L g6462 ( 
.A(n_6117),
.Y(n_6462)
);

INVxp67_ASAP7_75t_SL g6463 ( 
.A(n_6039),
.Y(n_6463)
);

INVx1_ASAP7_75t_L g6464 ( 
.A(n_6124),
.Y(n_6464)
);

INVx1_ASAP7_75t_L g6465 ( 
.A(n_6128),
.Y(n_6465)
);

INVx1_ASAP7_75t_L g6466 ( 
.A(n_6134),
.Y(n_6466)
);

INVx1_ASAP7_75t_L g6467 ( 
.A(n_6138),
.Y(n_6467)
);

INVx1_ASAP7_75t_L g6468 ( 
.A(n_6139),
.Y(n_6468)
);

INVxp33_ASAP7_75t_SL g6469 ( 
.A(n_5827),
.Y(n_6469)
);

BUFx3_ASAP7_75t_L g6470 ( 
.A(n_6041),
.Y(n_6470)
);

INVx1_ASAP7_75t_L g6471 ( 
.A(n_6140),
.Y(n_6471)
);

INVx2_ASAP7_75t_L g6472 ( 
.A(n_5780),
.Y(n_6472)
);

INVxp67_ASAP7_75t_SL g6473 ( 
.A(n_6043),
.Y(n_6473)
);

INVx1_ASAP7_75t_L g6474 ( 
.A(n_6141),
.Y(n_6474)
);

INVx1_ASAP7_75t_L g6475 ( 
.A(n_6143),
.Y(n_6475)
);

CKINVDCx5p33_ASAP7_75t_R g6476 ( 
.A(n_5938),
.Y(n_6476)
);

INVx1_ASAP7_75t_L g6477 ( 
.A(n_6146),
.Y(n_6477)
);

INVxp67_ASAP7_75t_L g6478 ( 
.A(n_6190),
.Y(n_6478)
);

INVxp33_ASAP7_75t_SL g6479 ( 
.A(n_5836),
.Y(n_6479)
);

INVx1_ASAP7_75t_L g6480 ( 
.A(n_6149),
.Y(n_6480)
);

INVx1_ASAP7_75t_L g6481 ( 
.A(n_6151),
.Y(n_6481)
);

INVx1_ASAP7_75t_L g6482 ( 
.A(n_6154),
.Y(n_6482)
);

CKINVDCx20_ASAP7_75t_R g6483 ( 
.A(n_5838),
.Y(n_6483)
);

INVx1_ASAP7_75t_L g6484 ( 
.A(n_6156),
.Y(n_6484)
);

INVx1_ASAP7_75t_L g6485 ( 
.A(n_6158),
.Y(n_6485)
);

INVx1_ASAP7_75t_L g6486 ( 
.A(n_6162),
.Y(n_6486)
);

INVx1_ASAP7_75t_L g6487 ( 
.A(n_6165),
.Y(n_6487)
);

INVx1_ASAP7_75t_L g6488 ( 
.A(n_6169),
.Y(n_6488)
);

INVx1_ASAP7_75t_L g6489 ( 
.A(n_6170),
.Y(n_6489)
);

CKINVDCx5p33_ASAP7_75t_R g6490 ( 
.A(n_5949),
.Y(n_6490)
);

INVx1_ASAP7_75t_L g6491 ( 
.A(n_6172),
.Y(n_6491)
);

CKINVDCx5p33_ASAP7_75t_R g6492 ( 
.A(n_5950),
.Y(n_6492)
);

INVxp67_ASAP7_75t_L g6493 ( 
.A(n_5930),
.Y(n_6493)
);

INVx1_ASAP7_75t_L g6494 ( 
.A(n_6174),
.Y(n_6494)
);

CKINVDCx20_ASAP7_75t_R g6495 ( 
.A(n_5840),
.Y(n_6495)
);

INVx1_ASAP7_75t_L g6496 ( 
.A(n_6175),
.Y(n_6496)
);

INVxp33_ASAP7_75t_SL g6497 ( 
.A(n_5841),
.Y(n_6497)
);

INVx1_ASAP7_75t_L g6498 ( 
.A(n_6179),
.Y(n_6498)
);

INVxp67_ASAP7_75t_SL g6499 ( 
.A(n_6044),
.Y(n_6499)
);

CKINVDCx5p33_ASAP7_75t_R g6500 ( 
.A(n_5953),
.Y(n_6500)
);

INVx1_ASAP7_75t_L g6501 ( 
.A(n_6180),
.Y(n_6501)
);

CKINVDCx5p33_ASAP7_75t_R g6502 ( 
.A(n_5954),
.Y(n_6502)
);

CKINVDCx20_ASAP7_75t_R g6503 ( 
.A(n_5957),
.Y(n_6503)
);

INVx1_ASAP7_75t_L g6504 ( 
.A(n_6186),
.Y(n_6504)
);

INVx1_ASAP7_75t_L g6505 ( 
.A(n_6187),
.Y(n_6505)
);

INVx1_ASAP7_75t_L g6506 ( 
.A(n_6191),
.Y(n_6506)
);

INVx2_ASAP7_75t_L g6507 ( 
.A(n_5794),
.Y(n_6507)
);

INVx1_ASAP7_75t_L g6508 ( 
.A(n_6192),
.Y(n_6508)
);

CKINVDCx20_ASAP7_75t_R g6509 ( 
.A(n_5960),
.Y(n_6509)
);

INVxp33_ASAP7_75t_L g6510 ( 
.A(n_5955),
.Y(n_6510)
);

CKINVDCx20_ASAP7_75t_R g6511 ( 
.A(n_5964),
.Y(n_6511)
);

INVx1_ASAP7_75t_L g6512 ( 
.A(n_6194),
.Y(n_6512)
);

INVxp67_ASAP7_75t_L g6513 ( 
.A(n_6019),
.Y(n_6513)
);

INVxp33_ASAP7_75t_SL g6514 ( 
.A(n_5790),
.Y(n_6514)
);

INVx1_ASAP7_75t_SL g6515 ( 
.A(n_5791),
.Y(n_6515)
);

CKINVDCx5p33_ASAP7_75t_R g6516 ( 
.A(n_5968),
.Y(n_6516)
);

INVx1_ASAP7_75t_L g6517 ( 
.A(n_6195),
.Y(n_6517)
);

INVx1_ASAP7_75t_L g6518 ( 
.A(n_5803),
.Y(n_6518)
);

INVx4_ASAP7_75t_R g6519 ( 
.A(n_5757),
.Y(n_6519)
);

INVx1_ASAP7_75t_L g6520 ( 
.A(n_5817),
.Y(n_6520)
);

INVxp67_ASAP7_75t_SL g6521 ( 
.A(n_6046),
.Y(n_6521)
);

CKINVDCx16_ASAP7_75t_R g6522 ( 
.A(n_6067),
.Y(n_6522)
);

CKINVDCx20_ASAP7_75t_R g6523 ( 
.A(n_5972),
.Y(n_6523)
);

CKINVDCx5p33_ASAP7_75t_R g6524 ( 
.A(n_5980),
.Y(n_6524)
);

INVxp33_ASAP7_75t_L g6525 ( 
.A(n_6152),
.Y(n_6525)
);

BUFx2_ASAP7_75t_L g6526 ( 
.A(n_5981),
.Y(n_6526)
);

INVx1_ASAP7_75t_L g6527 ( 
.A(n_6074),
.Y(n_6527)
);

CKINVDCx5p33_ASAP7_75t_R g6528 ( 
.A(n_5983),
.Y(n_6528)
);

INVx3_ASAP7_75t_L g6529 ( 
.A(n_6173),
.Y(n_6529)
);

INVx1_ASAP7_75t_L g6530 ( 
.A(n_6081),
.Y(n_6530)
);

CKINVDCx20_ASAP7_75t_R g6531 ( 
.A(n_5985),
.Y(n_6531)
);

INVxp33_ASAP7_75t_SL g6532 ( 
.A(n_5792),
.Y(n_6532)
);

CKINVDCx5p33_ASAP7_75t_R g6533 ( 
.A(n_5990),
.Y(n_6533)
);

INVxp67_ASAP7_75t_L g6534 ( 
.A(n_6021),
.Y(n_6534)
);

CKINVDCx5p33_ASAP7_75t_R g6535 ( 
.A(n_5992),
.Y(n_6535)
);

CKINVDCx20_ASAP7_75t_R g6536 ( 
.A(n_5995),
.Y(n_6536)
);

INVx1_ASAP7_75t_L g6537 ( 
.A(n_6085),
.Y(n_6537)
);

BUFx3_ASAP7_75t_L g6538 ( 
.A(n_6052),
.Y(n_6538)
);

CKINVDCx14_ASAP7_75t_R g6539 ( 
.A(n_5773),
.Y(n_6539)
);

INVx1_ASAP7_75t_L g6540 ( 
.A(n_6108),
.Y(n_6540)
);

INVx1_ASAP7_75t_L g6541 ( 
.A(n_6145),
.Y(n_6541)
);

INVx2_ASAP7_75t_L g6542 ( 
.A(n_6193),
.Y(n_6542)
);

CKINVDCx20_ASAP7_75t_R g6543 ( 
.A(n_5997),
.Y(n_6543)
);

INVxp67_ASAP7_75t_L g6544 ( 
.A(n_5939),
.Y(n_6544)
);

CKINVDCx5p33_ASAP7_75t_R g6545 ( 
.A(n_5999),
.Y(n_6545)
);

INVx1_ASAP7_75t_L g6546 ( 
.A(n_6147),
.Y(n_6546)
);

CKINVDCx5p33_ASAP7_75t_R g6547 ( 
.A(n_6003),
.Y(n_6547)
);

INVxp67_ASAP7_75t_SL g6548 ( 
.A(n_6057),
.Y(n_6548)
);

INVx1_ASAP7_75t_L g6549 ( 
.A(n_6168),
.Y(n_6549)
);

CKINVDCx20_ASAP7_75t_R g6550 ( 
.A(n_6004),
.Y(n_6550)
);

INVx1_ASAP7_75t_L g6551 ( 
.A(n_6189),
.Y(n_6551)
);

HB1xp67_ASAP7_75t_L g6552 ( 
.A(n_6005),
.Y(n_6552)
);

CKINVDCx20_ASAP7_75t_R g6553 ( 
.A(n_6006),
.Y(n_6553)
);

CKINVDCx20_ASAP7_75t_R g6554 ( 
.A(n_6010),
.Y(n_6554)
);

INVx1_ASAP7_75t_L g6555 ( 
.A(n_6065),
.Y(n_6555)
);

INVx1_ASAP7_75t_L g6556 ( 
.A(n_6068),
.Y(n_6556)
);

INVx1_ASAP7_75t_L g6557 ( 
.A(n_6071),
.Y(n_6557)
);

INVxp67_ASAP7_75t_SL g6558 ( 
.A(n_6072),
.Y(n_6558)
);

INVx1_ASAP7_75t_L g6559 ( 
.A(n_6073),
.Y(n_6559)
);

INVxp67_ASAP7_75t_SL g6560 ( 
.A(n_5767),
.Y(n_6560)
);

CKINVDCx5p33_ASAP7_75t_R g6561 ( 
.A(n_6015),
.Y(n_6561)
);

INVx1_ASAP7_75t_L g6562 ( 
.A(n_6193),
.Y(n_6562)
);

HB1xp67_ASAP7_75t_L g6563 ( 
.A(n_6016),
.Y(n_6563)
);

CKINVDCx20_ASAP7_75t_R g6564 ( 
.A(n_6017),
.Y(n_6564)
);

INVx1_ASAP7_75t_L g6565 ( 
.A(n_6193),
.Y(n_6565)
);

CKINVDCx5p33_ASAP7_75t_R g6566 ( 
.A(n_6018),
.Y(n_6566)
);

INVxp67_ASAP7_75t_SL g6567 ( 
.A(n_5937),
.Y(n_6567)
);

CKINVDCx5p33_ASAP7_75t_R g6568 ( 
.A(n_6020),
.Y(n_6568)
);

INVx1_ASAP7_75t_L g6569 ( 
.A(n_6002),
.Y(n_6569)
);

INVx1_ASAP7_75t_L g6570 ( 
.A(n_6002),
.Y(n_6570)
);

INVx1_ASAP7_75t_L g6571 ( 
.A(n_6002),
.Y(n_6571)
);

CKINVDCx5p33_ASAP7_75t_R g6572 ( 
.A(n_6022),
.Y(n_6572)
);

BUFx3_ASAP7_75t_L g6573 ( 
.A(n_6002),
.Y(n_6573)
);

INVx1_ASAP7_75t_L g6574 ( 
.A(n_6002),
.Y(n_6574)
);

CKINVDCx16_ASAP7_75t_R g6575 ( 
.A(n_6070),
.Y(n_6575)
);

INVx1_ASAP7_75t_L g6576 ( 
.A(n_6011),
.Y(n_6576)
);

INVx1_ASAP7_75t_L g6577 ( 
.A(n_6011),
.Y(n_6577)
);

INVx1_ASAP7_75t_L g6578 ( 
.A(n_6011),
.Y(n_6578)
);

INVxp67_ASAP7_75t_L g6579 ( 
.A(n_6166),
.Y(n_6579)
);

INVx1_ASAP7_75t_L g6580 ( 
.A(n_6011),
.Y(n_6580)
);

INVx1_ASAP7_75t_L g6581 ( 
.A(n_6011),
.Y(n_6581)
);

CKINVDCx16_ASAP7_75t_R g6582 ( 
.A(n_6121),
.Y(n_6582)
);

INVx1_ASAP7_75t_L g6583 ( 
.A(n_6109),
.Y(n_6583)
);

CKINVDCx20_ASAP7_75t_R g6584 ( 
.A(n_6031),
.Y(n_6584)
);

CKINVDCx5p33_ASAP7_75t_R g6585 ( 
.A(n_6032),
.Y(n_6585)
);

CKINVDCx20_ASAP7_75t_R g6586 ( 
.A(n_6034),
.Y(n_6586)
);

INVx1_ASAP7_75t_L g6587 ( 
.A(n_6109),
.Y(n_6587)
);

CKINVDCx20_ASAP7_75t_R g6588 ( 
.A(n_6036),
.Y(n_6588)
);

INVx1_ASAP7_75t_L g6589 ( 
.A(n_6109),
.Y(n_6589)
);

INVx1_ASAP7_75t_L g6590 ( 
.A(n_6109),
.Y(n_6590)
);

CKINVDCx20_ASAP7_75t_R g6591 ( 
.A(n_6040),
.Y(n_6591)
);

INVx1_ASAP7_75t_L g6592 ( 
.A(n_6109),
.Y(n_6592)
);

CKINVDCx20_ASAP7_75t_R g6593 ( 
.A(n_6042),
.Y(n_6593)
);

INVx1_ASAP7_75t_L g6594 ( 
.A(n_6126),
.Y(n_6594)
);

INVx1_ASAP7_75t_L g6595 ( 
.A(n_6126),
.Y(n_6595)
);

CKINVDCx5p33_ASAP7_75t_R g6596 ( 
.A(n_6045),
.Y(n_6596)
);

CKINVDCx20_ASAP7_75t_R g6597 ( 
.A(n_6047),
.Y(n_6597)
);

INVx1_ASAP7_75t_L g6598 ( 
.A(n_6126),
.Y(n_6598)
);

BUFx3_ASAP7_75t_L g6599 ( 
.A(n_6126),
.Y(n_6599)
);

CKINVDCx5p33_ASAP7_75t_R g6600 ( 
.A(n_6050),
.Y(n_6600)
);

INVx1_ASAP7_75t_L g6601 ( 
.A(n_6126),
.Y(n_6601)
);

BUFx6f_ASAP7_75t_L g6602 ( 
.A(n_6130),
.Y(n_6602)
);

INVxp67_ASAP7_75t_SL g6603 ( 
.A(n_6153),
.Y(n_6603)
);

INVx1_ASAP7_75t_L g6604 ( 
.A(n_5770),
.Y(n_6604)
);

INVxp33_ASAP7_75t_SL g6605 ( 
.A(n_5796),
.Y(n_6605)
);

CKINVDCx16_ASAP7_75t_R g6606 ( 
.A(n_6129),
.Y(n_6606)
);

INVx1_ASAP7_75t_L g6607 ( 
.A(n_5882),
.Y(n_6607)
);

INVx1_ASAP7_75t_L g6608 ( 
.A(n_5882),
.Y(n_6608)
);

INVxp67_ASAP7_75t_L g6609 ( 
.A(n_5764),
.Y(n_6609)
);

CKINVDCx5p33_ASAP7_75t_R g6610 ( 
.A(n_6055),
.Y(n_6610)
);

INVx1_ASAP7_75t_L g6611 ( 
.A(n_5882),
.Y(n_6611)
);

CKINVDCx20_ASAP7_75t_R g6612 ( 
.A(n_6060),
.Y(n_6612)
);

INVx1_ASAP7_75t_L g6613 ( 
.A(n_5882),
.Y(n_6613)
);

INVxp67_ASAP7_75t_SL g6614 ( 
.A(n_6178),
.Y(n_6614)
);

INVx1_ASAP7_75t_L g6615 ( 
.A(n_5882),
.Y(n_6615)
);

INVx1_ASAP7_75t_L g6616 ( 
.A(n_6127),
.Y(n_6616)
);

INVx1_ASAP7_75t_L g6617 ( 
.A(n_6199),
.Y(n_6617)
);

CKINVDCx20_ASAP7_75t_R g6618 ( 
.A(n_6062),
.Y(n_6618)
);

CKINVDCx20_ASAP7_75t_R g6619 ( 
.A(n_6063),
.Y(n_6619)
);

INVx1_ASAP7_75t_L g6620 ( 
.A(n_6064),
.Y(n_6620)
);

INVxp33_ASAP7_75t_SL g6621 ( 
.A(n_6066),
.Y(n_6621)
);

INVx1_ASAP7_75t_L g6622 ( 
.A(n_6075),
.Y(n_6622)
);

INVx2_ASAP7_75t_L g6623 ( 
.A(n_6008),
.Y(n_6623)
);

CKINVDCx16_ASAP7_75t_R g6624 ( 
.A(n_6132),
.Y(n_6624)
);

INVxp67_ASAP7_75t_SL g6625 ( 
.A(n_6185),
.Y(n_6625)
);

CKINVDCx5p33_ASAP7_75t_R g6626 ( 
.A(n_6078),
.Y(n_6626)
);

CKINVDCx5p33_ASAP7_75t_R g6627 ( 
.A(n_6080),
.Y(n_6627)
);

INVx1_ASAP7_75t_SL g6628 ( 
.A(n_5849),
.Y(n_6628)
);

CKINVDCx16_ASAP7_75t_R g6629 ( 
.A(n_6167),
.Y(n_6629)
);

CKINVDCx20_ASAP7_75t_R g6630 ( 
.A(n_6082),
.Y(n_6630)
);

INVx2_ASAP7_75t_SL g6631 ( 
.A(n_5814),
.Y(n_6631)
);

INVxp67_ASAP7_75t_L g6632 ( 
.A(n_5874),
.Y(n_6632)
);

INVxp33_ASAP7_75t_L g6633 ( 
.A(n_6024),
.Y(n_6633)
);

INVx1_ASAP7_75t_L g6634 ( 
.A(n_6198),
.Y(n_6634)
);

CKINVDCx20_ASAP7_75t_R g6635 ( 
.A(n_6083),
.Y(n_6635)
);

INVxp67_ASAP7_75t_L g6636 ( 
.A(n_6090),
.Y(n_6636)
);

INVx1_ASAP7_75t_L g6637 ( 
.A(n_6091),
.Y(n_6637)
);

CKINVDCx5p33_ASAP7_75t_R g6638 ( 
.A(n_6093),
.Y(n_6638)
);

CKINVDCx5p33_ASAP7_75t_R g6639 ( 
.A(n_6094),
.Y(n_6639)
);

CKINVDCx5p33_ASAP7_75t_R g6640 ( 
.A(n_6097),
.Y(n_6640)
);

INVxp67_ASAP7_75t_L g6641 ( 
.A(n_6099),
.Y(n_6641)
);

INVx1_ASAP7_75t_L g6642 ( 
.A(n_6100),
.Y(n_6642)
);

INVx1_ASAP7_75t_L g6643 ( 
.A(n_6101),
.Y(n_6643)
);

INVx2_ASAP7_75t_L g6644 ( 
.A(n_6102),
.Y(n_6644)
);

CKINVDCx5p33_ASAP7_75t_R g6645 ( 
.A(n_6105),
.Y(n_6645)
);

INVx1_ASAP7_75t_L g6646 ( 
.A(n_6106),
.Y(n_6646)
);

INVx2_ASAP7_75t_L g6647 ( 
.A(n_6113),
.Y(n_6647)
);

INVx1_ASAP7_75t_L g6648 ( 
.A(n_6115),
.Y(n_6648)
);

CKINVDCx16_ASAP7_75t_R g6649 ( 
.A(n_5814),
.Y(n_6649)
);

INVxp33_ASAP7_75t_SL g6650 ( 
.A(n_6118),
.Y(n_6650)
);

BUFx2_ASAP7_75t_L g6651 ( 
.A(n_6120),
.Y(n_6651)
);

CKINVDCx5p33_ASAP7_75t_R g6652 ( 
.A(n_6122),
.Y(n_6652)
);

INVxp33_ASAP7_75t_SL g6653 ( 
.A(n_6123),
.Y(n_6653)
);

CKINVDCx5p33_ASAP7_75t_R g6654 ( 
.A(n_6133),
.Y(n_6654)
);

CKINVDCx5p33_ASAP7_75t_R g6655 ( 
.A(n_6142),
.Y(n_6655)
);

INVx1_ASAP7_75t_L g6656 ( 
.A(n_6144),
.Y(n_6656)
);

CKINVDCx5p33_ASAP7_75t_R g6657 ( 
.A(n_6148),
.Y(n_6657)
);

INVx1_ASAP7_75t_L g6658 ( 
.A(n_6150),
.Y(n_6658)
);

CKINVDCx20_ASAP7_75t_R g6659 ( 
.A(n_6155),
.Y(n_6659)
);

CKINVDCx20_ASAP7_75t_R g6660 ( 
.A(n_6157),
.Y(n_6660)
);

BUFx6f_ASAP7_75t_L g6661 ( 
.A(n_6159),
.Y(n_6661)
);

INVx2_ASAP7_75t_L g6662 ( 
.A(n_6160),
.Y(n_6662)
);

CKINVDCx5p33_ASAP7_75t_R g6663 ( 
.A(n_6163),
.Y(n_6663)
);

HB1xp67_ASAP7_75t_L g6664 ( 
.A(n_6164),
.Y(n_6664)
);

INVx1_ASAP7_75t_L g6665 ( 
.A(n_6171),
.Y(n_6665)
);

CKINVDCx5p33_ASAP7_75t_R g6666 ( 
.A(n_6176),
.Y(n_6666)
);

INVx1_ASAP7_75t_L g6667 ( 
.A(n_6181),
.Y(n_6667)
);

INVxp67_ASAP7_75t_L g6668 ( 
.A(n_6182),
.Y(n_6668)
);

INVx2_ASAP7_75t_L g6669 ( 
.A(n_6188),
.Y(n_6669)
);

INVx1_ASAP7_75t_SL g6670 ( 
.A(n_5894),
.Y(n_6670)
);

INVx1_ASAP7_75t_L g6671 ( 
.A(n_5855),
.Y(n_6671)
);

INVx2_ASAP7_75t_L g6672 ( 
.A(n_5755),
.Y(n_6672)
);

INVx2_ASAP7_75t_L g6673 ( 
.A(n_5819),
.Y(n_6673)
);

CKINVDCx5p33_ASAP7_75t_R g6674 ( 
.A(n_6069),
.Y(n_6674)
);

BUFx6f_ASAP7_75t_SL g6675 ( 
.A(n_5894),
.Y(n_6675)
);

CKINVDCx20_ASAP7_75t_R g6676 ( 
.A(n_5928),
.Y(n_6676)
);

CKINVDCx5p33_ASAP7_75t_R g6677 ( 
.A(n_5917),
.Y(n_6677)
);

INVx1_ASAP7_75t_L g6678 ( 
.A(n_5897),
.Y(n_6678)
);

CKINVDCx16_ASAP7_75t_R g6679 ( 
.A(n_5917),
.Y(n_6679)
);

CKINVDCx5p33_ASAP7_75t_R g6680 ( 
.A(n_6077),
.Y(n_6680)
);

INVx1_ASAP7_75t_L g6681 ( 
.A(n_5965),
.Y(n_6681)
);

INVx1_ASAP7_75t_L g6682 ( 
.A(n_5989),
.Y(n_6682)
);

INVxp33_ASAP7_75t_SL g6683 ( 
.A(n_6048),
.Y(n_6683)
);

INVxp67_ASAP7_75t_SL g6684 ( 
.A(n_6197),
.Y(n_6684)
);

INVx1_ASAP7_75t_L g6685 ( 
.A(n_5976),
.Y(n_6685)
);

INVx1_ASAP7_75t_L g6686 ( 
.A(n_6077),
.Y(n_6686)
);

CKINVDCx16_ASAP7_75t_R g6687 ( 
.A(n_6095),
.Y(n_6687)
);

INVxp67_ASAP7_75t_SL g6688 ( 
.A(n_6095),
.Y(n_6688)
);

BUFx2_ASAP7_75t_L g6689 ( 
.A(n_5828),
.Y(n_6689)
);

INVx2_ASAP7_75t_L g6690 ( 
.A(n_5884),
.Y(n_6690)
);

CKINVDCx16_ASAP7_75t_R g6691 ( 
.A(n_5788),
.Y(n_6691)
);

BUFx3_ASAP7_75t_L g6692 ( 
.A(n_5786),
.Y(n_6692)
);

INVx1_ASAP7_75t_L g6693 ( 
.A(n_5774),
.Y(n_6693)
);

INVxp67_ASAP7_75t_SL g6694 ( 
.A(n_5786),
.Y(n_6694)
);

CKINVDCx5p33_ASAP7_75t_R g6695 ( 
.A(n_5775),
.Y(n_6695)
);

CKINVDCx5p33_ASAP7_75t_R g6696 ( 
.A(n_5775),
.Y(n_6696)
);

INVx1_ASAP7_75t_L g6697 ( 
.A(n_5774),
.Y(n_6697)
);

CKINVDCx5p33_ASAP7_75t_R g6698 ( 
.A(n_5775),
.Y(n_6698)
);

INVx1_ASAP7_75t_L g6699 ( 
.A(n_5774),
.Y(n_6699)
);

INVxp67_ASAP7_75t_SL g6700 ( 
.A(n_5786),
.Y(n_6700)
);

INVx1_ASAP7_75t_L g6701 ( 
.A(n_5774),
.Y(n_6701)
);

INVx1_ASAP7_75t_L g6702 ( 
.A(n_5774),
.Y(n_6702)
);

INVx1_ASAP7_75t_L g6703 ( 
.A(n_5774),
.Y(n_6703)
);

INVx1_ASAP7_75t_L g6704 ( 
.A(n_5774),
.Y(n_6704)
);

INVx1_ASAP7_75t_L g6705 ( 
.A(n_5774),
.Y(n_6705)
);

HB1xp67_ASAP7_75t_L g6706 ( 
.A(n_5798),
.Y(n_6706)
);

INVx1_ASAP7_75t_L g6707 ( 
.A(n_5774),
.Y(n_6707)
);

INVx1_ASAP7_75t_L g6708 ( 
.A(n_5774),
.Y(n_6708)
);

INVx1_ASAP7_75t_L g6709 ( 
.A(n_5774),
.Y(n_6709)
);

INVx1_ASAP7_75t_L g6710 ( 
.A(n_5774),
.Y(n_6710)
);

INVxp67_ASAP7_75t_SL g6711 ( 
.A(n_5786),
.Y(n_6711)
);

BUFx2_ASAP7_75t_L g6712 ( 
.A(n_5828),
.Y(n_6712)
);

INVx1_ASAP7_75t_L g6713 ( 
.A(n_5774),
.Y(n_6713)
);

INVxp67_ASAP7_75t_SL g6714 ( 
.A(n_5786),
.Y(n_6714)
);

INVx1_ASAP7_75t_L g6715 ( 
.A(n_5774),
.Y(n_6715)
);

INVxp67_ASAP7_75t_SL g6716 ( 
.A(n_5786),
.Y(n_6716)
);

BUFx6f_ASAP7_75t_L g6717 ( 
.A(n_6451),
.Y(n_6717)
);

INVx3_ASAP7_75t_L g6718 ( 
.A(n_6451),
.Y(n_6718)
);

BUFx6f_ASAP7_75t_L g6719 ( 
.A(n_6451),
.Y(n_6719)
);

OAI22xp5_ASAP7_75t_SL g6720 ( 
.A1(n_6628),
.A2(n_4687),
.B1(n_4691),
.B2(n_4628),
.Y(n_6720)
);

INVx2_ASAP7_75t_L g6721 ( 
.A(n_6542),
.Y(n_6721)
);

INVx1_ASAP7_75t_L g6722 ( 
.A(n_6428),
.Y(n_6722)
);

BUFx6f_ASAP7_75t_L g6723 ( 
.A(n_6348),
.Y(n_6723)
);

OAI22x1_ASAP7_75t_SL g6724 ( 
.A1(n_6674),
.A2(n_4801),
.B1(n_4821),
.B2(n_4790),
.Y(n_6724)
);

BUFx2_ASAP7_75t_L g6725 ( 
.A(n_6609),
.Y(n_6725)
);

INVx2_ASAP7_75t_L g6726 ( 
.A(n_6408),
.Y(n_6726)
);

NAND2xp5_ASAP7_75t_L g6727 ( 
.A(n_6560),
.B(n_4447),
.Y(n_6727)
);

NAND2xp5_ASAP7_75t_L g6728 ( 
.A(n_6604),
.B(n_4455),
.Y(n_6728)
);

INVx2_ASAP7_75t_L g6729 ( 
.A(n_6408),
.Y(n_6729)
);

INVx4_ASAP7_75t_L g6730 ( 
.A(n_6661),
.Y(n_6730)
);

INVx1_ASAP7_75t_L g6731 ( 
.A(n_6430),
.Y(n_6731)
);

INVx3_ASAP7_75t_L g6732 ( 
.A(n_6692),
.Y(n_6732)
);

INVx2_ASAP7_75t_L g6733 ( 
.A(n_6529),
.Y(n_6733)
);

NOR2xp33_ASAP7_75t_L g6734 ( 
.A(n_6567),
.B(n_6387),
.Y(n_6734)
);

OAI22xp5_ASAP7_75t_L g6735 ( 
.A1(n_6417),
.A2(n_4878),
.B1(n_5315),
.B2(n_5195),
.Y(n_6735)
);

INVx3_ASAP7_75t_L g6736 ( 
.A(n_6529),
.Y(n_6736)
);

AOI22xp5_ASAP7_75t_L g6737 ( 
.A1(n_6453),
.A2(n_4525),
.B1(n_4362),
.B2(n_4341),
.Y(n_6737)
);

CKINVDCx16_ASAP7_75t_R g6738 ( 
.A(n_6296),
.Y(n_6738)
);

AND2x2_ASAP7_75t_L g6739 ( 
.A(n_6632),
.B(n_4750),
.Y(n_6739)
);

OAI21x1_ASAP7_75t_L g6740 ( 
.A1(n_6607),
.A2(n_4413),
.B(n_4368),
.Y(n_6740)
);

BUFx6f_ASAP7_75t_L g6741 ( 
.A(n_6396),
.Y(n_6741)
);

NOR2xp33_ASAP7_75t_L g6742 ( 
.A(n_6683),
.B(n_5571),
.Y(n_6742)
);

NAND2xp5_ASAP7_75t_L g6743 ( 
.A(n_6573),
.B(n_4497),
.Y(n_6743)
);

BUFx6f_ASAP7_75t_L g6744 ( 
.A(n_6415),
.Y(n_6744)
);

AND2x4_ASAP7_75t_L g6745 ( 
.A(n_6716),
.B(n_4532),
.Y(n_6745)
);

BUFx12f_ASAP7_75t_L g6746 ( 
.A(n_6262),
.Y(n_6746)
);

NAND2xp5_ASAP7_75t_L g6747 ( 
.A(n_6599),
.B(n_4713),
.Y(n_6747)
);

BUFx12f_ASAP7_75t_L g6748 ( 
.A(n_6270),
.Y(n_6748)
);

INVx5_ASAP7_75t_L g6749 ( 
.A(n_6631),
.Y(n_6749)
);

BUFx6f_ASAP7_75t_L g6750 ( 
.A(n_6470),
.Y(n_6750)
);

BUFx6f_ASAP7_75t_L g6751 ( 
.A(n_6538),
.Y(n_6751)
);

INVx2_ASAP7_75t_L g6752 ( 
.A(n_6562),
.Y(n_6752)
);

AOI22xp5_ASAP7_75t_L g6753 ( 
.A1(n_6617),
.A2(n_4619),
.B1(n_4645),
.B2(n_4612),
.Y(n_6753)
);

BUFx6f_ASAP7_75t_L g6754 ( 
.A(n_6565),
.Y(n_6754)
);

INVx2_ASAP7_75t_L g6755 ( 
.A(n_6235),
.Y(n_6755)
);

INVx2_ASAP7_75t_L g6756 ( 
.A(n_6248),
.Y(n_6756)
);

OA21x2_ASAP7_75t_L g6757 ( 
.A1(n_6569),
.A2(n_4520),
.B(n_4519),
.Y(n_6757)
);

NAND2xp5_ASAP7_75t_L g6758 ( 
.A(n_6381),
.B(n_4728),
.Y(n_6758)
);

BUFx6f_ASAP7_75t_L g6759 ( 
.A(n_6370),
.Y(n_6759)
);

AND2x4_ASAP7_75t_L g6760 ( 
.A(n_6212),
.B(n_4745),
.Y(n_6760)
);

INVx2_ASAP7_75t_SL g6761 ( 
.A(n_6602),
.Y(n_6761)
);

OAI22xp5_ASAP7_75t_L g6762 ( 
.A1(n_6623),
.A2(n_6602),
.B1(n_6622),
.B2(n_6620),
.Y(n_6762)
);

INVx2_ASAP7_75t_L g6763 ( 
.A(n_6690),
.Y(n_6763)
);

INVx5_ASAP7_75t_L g6764 ( 
.A(n_6661),
.Y(n_6764)
);

BUFx6f_ASAP7_75t_L g6765 ( 
.A(n_6373),
.Y(n_6765)
);

AND2x6_ASAP7_75t_L g6766 ( 
.A(n_6661),
.B(n_4698),
.Y(n_6766)
);

NOR2xp33_ASAP7_75t_L g6767 ( 
.A(n_6634),
.B(n_6637),
.Y(n_6767)
);

BUFx12f_ASAP7_75t_L g6768 ( 
.A(n_6276),
.Y(n_6768)
);

INVx3_ASAP7_75t_L g6769 ( 
.A(n_6380),
.Y(n_6769)
);

HB1xp67_ASAP7_75t_L g6770 ( 
.A(n_6416),
.Y(n_6770)
);

AND2x4_ASAP7_75t_L g6771 ( 
.A(n_6220),
.B(n_4772),
.Y(n_6771)
);

NAND2xp5_ASAP7_75t_L g6772 ( 
.A(n_6382),
.B(n_4787),
.Y(n_6772)
);

INVx1_ASAP7_75t_L g6773 ( 
.A(n_6431),
.Y(n_6773)
);

OAI22xp5_ASAP7_75t_L g6774 ( 
.A1(n_6602),
.A2(n_4481),
.B1(n_4483),
.B2(n_4480),
.Y(n_6774)
);

INVx2_ASAP7_75t_L g6775 ( 
.A(n_6384),
.Y(n_6775)
);

CKINVDCx11_ASAP7_75t_R g6776 ( 
.A(n_6214),
.Y(n_6776)
);

INVx2_ASAP7_75t_L g6777 ( 
.A(n_6392),
.Y(n_6777)
);

INVx1_ASAP7_75t_L g6778 ( 
.A(n_6432),
.Y(n_6778)
);

INVx4_ASAP7_75t_L g6779 ( 
.A(n_6207),
.Y(n_6779)
);

INVx2_ASAP7_75t_L g6780 ( 
.A(n_6472),
.Y(n_6780)
);

INVx1_ASAP7_75t_L g6781 ( 
.A(n_6434),
.Y(n_6781)
);

INVx3_ASAP7_75t_L g6782 ( 
.A(n_6507),
.Y(n_6782)
);

CKINVDCx6p67_ASAP7_75t_R g6783 ( 
.A(n_6675),
.Y(n_6783)
);

INVx1_ASAP7_75t_L g6784 ( 
.A(n_6436),
.Y(n_6784)
);

OAI22x1_ASAP7_75t_R g6785 ( 
.A1(n_6311),
.A2(n_4841),
.B1(n_4850),
.B2(n_4834),
.Y(n_6785)
);

CKINVDCx5p33_ASAP7_75t_R g6786 ( 
.A(n_6219),
.Y(n_6786)
);

INVx1_ASAP7_75t_L g6787 ( 
.A(n_6440),
.Y(n_6787)
);

BUFx2_ASAP7_75t_L g6788 ( 
.A(n_6452),
.Y(n_6788)
);

AND2x2_ASAP7_75t_L g6789 ( 
.A(n_6633),
.B(n_4750),
.Y(n_6789)
);

INVx3_ASAP7_75t_L g6790 ( 
.A(n_6374),
.Y(n_6790)
);

INVx1_ASAP7_75t_L g6791 ( 
.A(n_6444),
.Y(n_6791)
);

INVx3_ASAP7_75t_L g6792 ( 
.A(n_6375),
.Y(n_6792)
);

BUFx6f_ASAP7_75t_L g6793 ( 
.A(n_6377),
.Y(n_6793)
);

AOI22xp5_ASAP7_75t_L g6794 ( 
.A1(n_6642),
.A2(n_4792),
.B1(n_4794),
.B2(n_4767),
.Y(n_6794)
);

INVx2_ASAP7_75t_L g6795 ( 
.A(n_6259),
.Y(n_6795)
);

INVx2_ASAP7_75t_L g6796 ( 
.A(n_6263),
.Y(n_6796)
);

AOI22x1_ASAP7_75t_SL g6797 ( 
.A1(n_6206),
.A2(n_4888),
.B1(n_4911),
.B2(n_4859),
.Y(n_6797)
);

OA21x2_ASAP7_75t_L g6798 ( 
.A1(n_6570),
.A2(n_4528),
.B(n_4527),
.Y(n_6798)
);

AND2x6_ASAP7_75t_L g6799 ( 
.A(n_6643),
.B(n_4833),
.Y(n_6799)
);

NAND2xp5_ASAP7_75t_L g6800 ( 
.A(n_6386),
.B(n_6389),
.Y(n_6800)
);

INVx2_ASAP7_75t_L g6801 ( 
.A(n_6285),
.Y(n_6801)
);

INVx1_ASAP7_75t_L g6802 ( 
.A(n_6445),
.Y(n_6802)
);

NOR2xp33_ASAP7_75t_L g6803 ( 
.A(n_6646),
.B(n_4856),
.Y(n_6803)
);

BUFx6f_ASAP7_75t_L g6804 ( 
.A(n_6378),
.Y(n_6804)
);

NAND2xp5_ASAP7_75t_L g6805 ( 
.A(n_6390),
.B(n_4873),
.Y(n_6805)
);

AND2x6_ASAP7_75t_L g6806 ( 
.A(n_6648),
.B(n_4885),
.Y(n_6806)
);

INVx5_ASAP7_75t_L g6807 ( 
.A(n_6320),
.Y(n_6807)
);

INVx2_ASAP7_75t_L g6808 ( 
.A(n_6290),
.Y(n_6808)
);

HB1xp67_ASAP7_75t_L g6809 ( 
.A(n_6456),
.Y(n_6809)
);

INVxp33_ASAP7_75t_SL g6810 ( 
.A(n_6677),
.Y(n_6810)
);

INVx2_ASAP7_75t_L g6811 ( 
.A(n_6292),
.Y(n_6811)
);

INVx2_ASAP7_75t_L g6812 ( 
.A(n_6303),
.Y(n_6812)
);

OAI21x1_ASAP7_75t_L g6813 ( 
.A1(n_6608),
.A2(n_4479),
.B(n_4456),
.Y(n_6813)
);

INVx2_ASAP7_75t_L g6814 ( 
.A(n_6306),
.Y(n_6814)
);

OA21x2_ASAP7_75t_L g6815 ( 
.A1(n_6571),
.A2(n_4536),
.B(n_4533),
.Y(n_6815)
);

BUFx6f_ASAP7_75t_L g6816 ( 
.A(n_6200),
.Y(n_6816)
);

INVx1_ASAP7_75t_L g6817 ( 
.A(n_6448),
.Y(n_6817)
);

AND2x4_ASAP7_75t_L g6818 ( 
.A(n_6242),
.B(n_4919),
.Y(n_6818)
);

AND2x4_ASAP7_75t_L g6819 ( 
.A(n_6307),
.B(n_4920),
.Y(n_6819)
);

BUFx6f_ASAP7_75t_L g6820 ( 
.A(n_6201),
.Y(n_6820)
);

OR2x2_ASAP7_75t_L g6821 ( 
.A(n_6579),
.B(n_4902),
.Y(n_6821)
);

AND2x4_ASAP7_75t_L g6822 ( 
.A(n_6318),
.B(n_4925),
.Y(n_6822)
);

INVx1_ASAP7_75t_L g6823 ( 
.A(n_6450),
.Y(n_6823)
);

AND2x2_ASAP7_75t_L g6824 ( 
.A(n_6313),
.B(n_4756),
.Y(n_6824)
);

INVx2_ASAP7_75t_L g6825 ( 
.A(n_6326),
.Y(n_6825)
);

OAI22xp5_ASAP7_75t_L g6826 ( 
.A1(n_6656),
.A2(n_6665),
.B1(n_6667),
.B2(n_6658),
.Y(n_6826)
);

NAND2xp5_ASAP7_75t_L g6827 ( 
.A(n_6394),
.B(n_4965),
.Y(n_6827)
);

BUFx6f_ASAP7_75t_L g6828 ( 
.A(n_6202),
.Y(n_6828)
);

AND2x2_ASAP7_75t_L g6829 ( 
.A(n_6603),
.B(n_4756),
.Y(n_6829)
);

INVx4_ASAP7_75t_L g6830 ( 
.A(n_6221),
.Y(n_6830)
);

INVx2_ASAP7_75t_L g6831 ( 
.A(n_6347),
.Y(n_6831)
);

AND2x4_ASAP7_75t_L g6832 ( 
.A(n_6337),
.B(n_4978),
.Y(n_6832)
);

AND2x6_ASAP7_75t_L g6833 ( 
.A(n_6644),
.B(n_4907),
.Y(n_6833)
);

BUFx6f_ASAP7_75t_L g6834 ( 
.A(n_6203),
.Y(n_6834)
);

BUFx8_ASAP7_75t_SL g6835 ( 
.A(n_6222),
.Y(n_6835)
);

NOR2x1_ASAP7_75t_L g6836 ( 
.A(n_6647),
.B(n_4946),
.Y(n_6836)
);

INVx2_ASAP7_75t_L g6837 ( 
.A(n_6359),
.Y(n_6837)
);

INVx2_ASAP7_75t_L g6838 ( 
.A(n_6518),
.Y(n_6838)
);

INVx2_ASAP7_75t_SL g6839 ( 
.A(n_6519),
.Y(n_6839)
);

OAI21x1_ASAP7_75t_L g6840 ( 
.A1(n_6611),
.A2(n_4549),
.B(n_4508),
.Y(n_6840)
);

AND2x2_ASAP7_75t_L g6841 ( 
.A(n_6544),
.B(n_4762),
.Y(n_6841)
);

NAND2xp5_ASAP7_75t_L g6842 ( 
.A(n_6397),
.B(n_6398),
.Y(n_6842)
);

INVx1_ASAP7_75t_L g6843 ( 
.A(n_6457),
.Y(n_6843)
);

NOR2x1_ASAP7_75t_L g6844 ( 
.A(n_6662),
.B(n_5140),
.Y(n_6844)
);

INVx1_ASAP7_75t_L g6845 ( 
.A(n_6458),
.Y(n_6845)
);

CKINVDCx16_ASAP7_75t_R g6846 ( 
.A(n_6383),
.Y(n_6846)
);

INVx2_ASAP7_75t_L g6847 ( 
.A(n_6520),
.Y(n_6847)
);

INVx1_ASAP7_75t_L g6848 ( 
.A(n_6459),
.Y(n_6848)
);

AND2x4_ASAP7_75t_L g6849 ( 
.A(n_6339),
.B(n_5010),
.Y(n_6849)
);

BUFx6f_ASAP7_75t_L g6850 ( 
.A(n_6205),
.Y(n_6850)
);

HB1xp67_ASAP7_75t_L g6851 ( 
.A(n_6279),
.Y(n_6851)
);

INVx1_ASAP7_75t_L g6852 ( 
.A(n_6460),
.Y(n_6852)
);

INVx1_ASAP7_75t_L g6853 ( 
.A(n_6462),
.Y(n_6853)
);

BUFx6f_ASAP7_75t_L g6854 ( 
.A(n_6209),
.Y(n_6854)
);

BUFx6f_ASAP7_75t_L g6855 ( 
.A(n_6211),
.Y(n_6855)
);

INVx2_ASAP7_75t_L g6856 ( 
.A(n_6249),
.Y(n_6856)
);

BUFx6f_ASAP7_75t_L g6857 ( 
.A(n_6215),
.Y(n_6857)
);

INVx1_ASAP7_75t_L g6858 ( 
.A(n_6464),
.Y(n_6858)
);

NOR2xp33_ASAP7_75t_L g6859 ( 
.A(n_6669),
.B(n_5061),
.Y(n_6859)
);

INVx1_ASAP7_75t_L g6860 ( 
.A(n_6465),
.Y(n_6860)
);

AND2x6_ASAP7_75t_L g6861 ( 
.A(n_6671),
.B(n_6678),
.Y(n_6861)
);

INVx2_ASAP7_75t_L g6862 ( 
.A(n_6252),
.Y(n_6862)
);

CKINVDCx11_ASAP7_75t_R g6863 ( 
.A(n_6226),
.Y(n_6863)
);

AND2x2_ASAP7_75t_L g6864 ( 
.A(n_6278),
.B(n_4762),
.Y(n_6864)
);

INVx1_ASAP7_75t_L g6865 ( 
.A(n_6466),
.Y(n_6865)
);

BUFx6f_ASAP7_75t_L g6866 ( 
.A(n_6216),
.Y(n_6866)
);

HB1xp67_ASAP7_75t_L g6867 ( 
.A(n_6493),
.Y(n_6867)
);

OAI22xp5_ASAP7_75t_SL g6868 ( 
.A1(n_6676),
.A2(n_4915),
.B1(n_4924),
.B2(n_4912),
.Y(n_6868)
);

INVx1_ASAP7_75t_L g6869 ( 
.A(n_6467),
.Y(n_6869)
);

INVx1_ASAP7_75t_L g6870 ( 
.A(n_6468),
.Y(n_6870)
);

INVx1_ASAP7_75t_L g6871 ( 
.A(n_6471),
.Y(n_6871)
);

OA21x2_ASAP7_75t_L g6872 ( 
.A1(n_6574),
.A2(n_4539),
.B(n_4537),
.Y(n_6872)
);

BUFx8_ASAP7_75t_L g6873 ( 
.A(n_6675),
.Y(n_6873)
);

INVx1_ASAP7_75t_L g6874 ( 
.A(n_6474),
.Y(n_6874)
);

BUFx3_ASAP7_75t_L g6875 ( 
.A(n_6503),
.Y(n_6875)
);

INVx5_ASAP7_75t_L g6876 ( 
.A(n_6412),
.Y(n_6876)
);

INVx3_ASAP7_75t_L g6877 ( 
.A(n_6217),
.Y(n_6877)
);

NAND2xp5_ASAP7_75t_L g6878 ( 
.A(n_6401),
.B(n_5104),
.Y(n_6878)
);

INVx1_ASAP7_75t_L g6879 ( 
.A(n_6475),
.Y(n_6879)
);

CKINVDCx11_ASAP7_75t_R g6880 ( 
.A(n_6232),
.Y(n_6880)
);

BUFx6f_ASAP7_75t_L g6881 ( 
.A(n_6218),
.Y(n_6881)
);

BUFx8_ASAP7_75t_SL g6882 ( 
.A(n_6236),
.Y(n_6882)
);

INVx3_ASAP7_75t_L g6883 ( 
.A(n_6224),
.Y(n_6883)
);

AND2x2_ASAP7_75t_L g6884 ( 
.A(n_6336),
.B(n_4814),
.Y(n_6884)
);

INVx3_ASAP7_75t_L g6885 ( 
.A(n_6227),
.Y(n_6885)
);

BUFx6f_ASAP7_75t_L g6886 ( 
.A(n_6228),
.Y(n_6886)
);

NAND2xp5_ASAP7_75t_L g6887 ( 
.A(n_6402),
.B(n_5127),
.Y(n_6887)
);

BUFx3_ASAP7_75t_L g6888 ( 
.A(n_6509),
.Y(n_6888)
);

INVx2_ASAP7_75t_L g6889 ( 
.A(n_6253),
.Y(n_6889)
);

AOI22xp5_ASAP7_75t_L g6890 ( 
.A1(n_6616),
.A2(n_4949),
.B1(n_4970),
.B2(n_4945),
.Y(n_6890)
);

NAND2xp5_ASAP7_75t_L g6891 ( 
.A(n_6403),
.B(n_5161),
.Y(n_6891)
);

BUFx8_ASAP7_75t_L g6892 ( 
.A(n_6225),
.Y(n_6892)
);

INVx1_ASAP7_75t_L g6893 ( 
.A(n_6477),
.Y(n_6893)
);

OAI21x1_ASAP7_75t_L g6894 ( 
.A1(n_6613),
.A2(n_6615),
.B(n_6577),
.Y(n_6894)
);

INVx2_ASAP7_75t_L g6895 ( 
.A(n_6254),
.Y(n_6895)
);

INVx2_ASAP7_75t_L g6896 ( 
.A(n_6255),
.Y(n_6896)
);

BUFx8_ASAP7_75t_L g6897 ( 
.A(n_6689),
.Y(n_6897)
);

BUFx12f_ASAP7_75t_L g6898 ( 
.A(n_6281),
.Y(n_6898)
);

INVx1_ASAP7_75t_L g6899 ( 
.A(n_6480),
.Y(n_6899)
);

CKINVDCx5p33_ASAP7_75t_R g6900 ( 
.A(n_6234),
.Y(n_6900)
);

INVx2_ASAP7_75t_L g6901 ( 
.A(n_6256),
.Y(n_6901)
);

BUFx3_ASAP7_75t_L g6902 ( 
.A(n_6511),
.Y(n_6902)
);

INVx2_ASAP7_75t_L g6903 ( 
.A(n_6257),
.Y(n_6903)
);

INVx2_ASAP7_75t_L g6904 ( 
.A(n_6258),
.Y(n_6904)
);

INVx3_ASAP7_75t_L g6905 ( 
.A(n_6229),
.Y(n_6905)
);

INVx3_ASAP7_75t_L g6906 ( 
.A(n_6693),
.Y(n_6906)
);

INVx1_ASAP7_75t_L g6907 ( 
.A(n_6481),
.Y(n_6907)
);

BUFx8_ASAP7_75t_L g6908 ( 
.A(n_6712),
.Y(n_6908)
);

INVxp67_ASAP7_75t_L g6909 ( 
.A(n_6614),
.Y(n_6909)
);

BUFx2_ASAP7_75t_L g6910 ( 
.A(n_6429),
.Y(n_6910)
);

INVx5_ASAP7_75t_L g6911 ( 
.A(n_6413),
.Y(n_6911)
);

BUFx6f_ASAP7_75t_L g6912 ( 
.A(n_6697),
.Y(n_6912)
);

INVx1_ASAP7_75t_L g6913 ( 
.A(n_6482),
.Y(n_6913)
);

INVx1_ASAP7_75t_L g6914 ( 
.A(n_6484),
.Y(n_6914)
);

INVxp67_ASAP7_75t_L g6915 ( 
.A(n_6625),
.Y(n_6915)
);

NOR2xp67_ASAP7_75t_L g6916 ( 
.A(n_6636),
.B(n_4279),
.Y(n_6916)
);

AND2x4_ASAP7_75t_L g6917 ( 
.A(n_6346),
.B(n_6351),
.Y(n_6917)
);

BUFx6f_ASAP7_75t_L g6918 ( 
.A(n_6699),
.Y(n_6918)
);

AND2x4_ASAP7_75t_L g6919 ( 
.A(n_6694),
.B(n_5168),
.Y(n_6919)
);

OA21x2_ASAP7_75t_L g6920 ( 
.A1(n_6576),
.A2(n_4546),
.B(n_4543),
.Y(n_6920)
);

INVx2_ASAP7_75t_L g6921 ( 
.A(n_6261),
.Y(n_6921)
);

INVx2_ASAP7_75t_L g6922 ( 
.A(n_6264),
.Y(n_6922)
);

NAND2xp5_ASAP7_75t_L g6923 ( 
.A(n_6404),
.B(n_5245),
.Y(n_6923)
);

INVx3_ASAP7_75t_L g6924 ( 
.A(n_6701),
.Y(n_6924)
);

INVx1_ASAP7_75t_L g6925 ( 
.A(n_6485),
.Y(n_6925)
);

BUFx6f_ASAP7_75t_L g6926 ( 
.A(n_6702),
.Y(n_6926)
);

XNOR2xp5_ASAP7_75t_L g6927 ( 
.A(n_6239),
.B(n_4941),
.Y(n_6927)
);

INVx3_ASAP7_75t_L g6928 ( 
.A(n_6703),
.Y(n_6928)
);

AOI22xp5_ASAP7_75t_L g6929 ( 
.A1(n_6641),
.A2(n_5165),
.B1(n_5173),
.B2(n_5040),
.Y(n_6929)
);

OA21x2_ASAP7_75t_L g6930 ( 
.A1(n_6578),
.A2(n_4555),
.B(n_4553),
.Y(n_6930)
);

BUFx6f_ASAP7_75t_L g6931 ( 
.A(n_6704),
.Y(n_6931)
);

INVx1_ASAP7_75t_L g6932 ( 
.A(n_6486),
.Y(n_6932)
);

INVx2_ASAP7_75t_L g6933 ( 
.A(n_6265),
.Y(n_6933)
);

BUFx8_ASAP7_75t_L g6934 ( 
.A(n_6361),
.Y(n_6934)
);

INVx3_ASAP7_75t_L g6935 ( 
.A(n_6705),
.Y(n_6935)
);

INVx4_ASAP7_75t_L g6936 ( 
.A(n_6250),
.Y(n_6936)
);

BUFx6f_ASAP7_75t_L g6937 ( 
.A(n_6707),
.Y(n_6937)
);

AND2x2_ASAP7_75t_L g6938 ( 
.A(n_6352),
.B(n_4814),
.Y(n_6938)
);

INVx2_ASAP7_75t_L g6939 ( 
.A(n_6266),
.Y(n_6939)
);

BUFx6f_ASAP7_75t_L g6940 ( 
.A(n_6708),
.Y(n_6940)
);

NAND2xp5_ASAP7_75t_L g6941 ( 
.A(n_6405),
.B(n_5438),
.Y(n_6941)
);

INVx1_ASAP7_75t_L g6942 ( 
.A(n_6487),
.Y(n_6942)
);

INVx3_ASAP7_75t_L g6943 ( 
.A(n_6709),
.Y(n_6943)
);

AND2x2_ASAP7_75t_L g6944 ( 
.A(n_6672),
.B(n_4829),
.Y(n_6944)
);

BUFx6f_ASAP7_75t_L g6945 ( 
.A(n_6710),
.Y(n_6945)
);

NAND2xp5_ASAP7_75t_L g6946 ( 
.A(n_6410),
.B(n_5496),
.Y(n_6946)
);

INVx1_ASAP7_75t_L g6947 ( 
.A(n_6488),
.Y(n_6947)
);

AND2x2_ASAP7_75t_L g6948 ( 
.A(n_6673),
.B(n_4829),
.Y(n_6948)
);

NOR2xp33_ASAP7_75t_L g6949 ( 
.A(n_6668),
.B(n_5509),
.Y(n_6949)
);

AOI22xp5_ASAP7_75t_L g6950 ( 
.A1(n_6204),
.A2(n_5265),
.B1(n_5309),
.B2(n_5212),
.Y(n_6950)
);

OAI21x1_ASAP7_75t_L g6951 ( 
.A1(n_6580),
.A2(n_4630),
.B(n_4601),
.Y(n_6951)
);

INVx2_ASAP7_75t_L g6952 ( 
.A(n_6267),
.Y(n_6952)
);

INVx3_ASAP7_75t_L g6953 ( 
.A(n_6713),
.Y(n_6953)
);

CKINVDCx6p67_ASAP7_75t_R g6954 ( 
.A(n_6454),
.Y(n_6954)
);

INVx1_ASAP7_75t_L g6955 ( 
.A(n_6489),
.Y(n_6955)
);

BUFx6f_ASAP7_75t_L g6956 ( 
.A(n_6715),
.Y(n_6956)
);

BUFx6f_ASAP7_75t_L g6957 ( 
.A(n_6491),
.Y(n_6957)
);

AND2x2_ASAP7_75t_L g6958 ( 
.A(n_6433),
.B(n_4917),
.Y(n_6958)
);

OAI22xp5_ASAP7_75t_R g6959 ( 
.A1(n_6680),
.A2(n_4487),
.B1(n_4489),
.B2(n_4485),
.Y(n_6959)
);

INVx2_ASAP7_75t_L g6960 ( 
.A(n_6268),
.Y(n_6960)
);

INVx2_ASAP7_75t_L g6961 ( 
.A(n_6269),
.Y(n_6961)
);

INVx2_ASAP7_75t_L g6962 ( 
.A(n_6271),
.Y(n_6962)
);

NOR2xp33_ASAP7_75t_L g6963 ( 
.A(n_6621),
.B(n_5613),
.Y(n_6963)
);

AOI22xp5_ASAP7_75t_L g6964 ( 
.A1(n_6684),
.A2(n_5329),
.B1(n_5341),
.B2(n_5311),
.Y(n_6964)
);

BUFx6f_ASAP7_75t_L g6965 ( 
.A(n_6494),
.Y(n_6965)
);

BUFx6f_ASAP7_75t_L g6966 ( 
.A(n_6496),
.Y(n_6966)
);

INVx2_ASAP7_75t_L g6967 ( 
.A(n_6272),
.Y(n_6967)
);

AND2x2_ASAP7_75t_L g6968 ( 
.A(n_6510),
.B(n_6525),
.Y(n_6968)
);

NAND2xp5_ASAP7_75t_L g6969 ( 
.A(n_6418),
.B(n_5684),
.Y(n_6969)
);

BUFx6f_ASAP7_75t_L g6970 ( 
.A(n_6498),
.Y(n_6970)
);

INVx1_ASAP7_75t_L g6971 ( 
.A(n_6501),
.Y(n_6971)
);

OA21x2_ASAP7_75t_L g6972 ( 
.A1(n_6581),
.A2(n_4560),
.B(n_4558),
.Y(n_6972)
);

INVx5_ASAP7_75t_L g6973 ( 
.A(n_6522),
.Y(n_6973)
);

OA21x2_ASAP7_75t_L g6974 ( 
.A1(n_6583),
.A2(n_4578),
.B(n_4575),
.Y(n_6974)
);

INVx1_ASAP7_75t_L g6975 ( 
.A(n_6504),
.Y(n_6975)
);

INVx2_ASAP7_75t_L g6976 ( 
.A(n_6273),
.Y(n_6976)
);

BUFx6f_ASAP7_75t_L g6977 ( 
.A(n_6505),
.Y(n_6977)
);

BUFx6f_ASAP7_75t_L g6978 ( 
.A(n_6506),
.Y(n_6978)
);

INVx2_ASAP7_75t_L g6979 ( 
.A(n_6274),
.Y(n_6979)
);

INVx2_ASAP7_75t_L g6980 ( 
.A(n_6277),
.Y(n_6980)
);

INVx2_ASAP7_75t_L g6981 ( 
.A(n_6280),
.Y(n_6981)
);

BUFx6f_ASAP7_75t_L g6982 ( 
.A(n_6508),
.Y(n_6982)
);

INVx1_ASAP7_75t_L g6983 ( 
.A(n_6512),
.Y(n_6983)
);

BUFx6f_ASAP7_75t_L g6984 ( 
.A(n_6517),
.Y(n_6984)
);

OA21x2_ASAP7_75t_L g6985 ( 
.A1(n_6587),
.A2(n_4588),
.B(n_4580),
.Y(n_6985)
);

INVx5_ASAP7_75t_L g6986 ( 
.A(n_6575),
.Y(n_6986)
);

INVx4_ASAP7_75t_L g6987 ( 
.A(n_6251),
.Y(n_6987)
);

AND2x4_ASAP7_75t_L g6988 ( 
.A(n_6700),
.B(n_5722),
.Y(n_6988)
);

INVx2_ASAP7_75t_SL g6989 ( 
.A(n_6685),
.Y(n_6989)
);

OA21x2_ASAP7_75t_L g6990 ( 
.A1(n_6589),
.A2(n_4591),
.B(n_4590),
.Y(n_6990)
);

INVx3_ASAP7_75t_L g6991 ( 
.A(n_6423),
.Y(n_6991)
);

INVx2_ASAP7_75t_L g6992 ( 
.A(n_6283),
.Y(n_6992)
);

INVx2_ASAP7_75t_L g6993 ( 
.A(n_6284),
.Y(n_6993)
);

CKINVDCx20_ASAP7_75t_R g6994 ( 
.A(n_6240),
.Y(n_6994)
);

INVx3_ASAP7_75t_L g6995 ( 
.A(n_6424),
.Y(n_6995)
);

CKINVDCx6p67_ASAP7_75t_R g6996 ( 
.A(n_6582),
.Y(n_6996)
);

CKINVDCx5p33_ASAP7_75t_R g6997 ( 
.A(n_6695),
.Y(n_6997)
);

CKINVDCx5p33_ASAP7_75t_R g6998 ( 
.A(n_6696),
.Y(n_6998)
);

BUFx6f_ASAP7_75t_L g6999 ( 
.A(n_6287),
.Y(n_6999)
);

INVx1_ASAP7_75t_L g7000 ( 
.A(n_6419),
.Y(n_7000)
);

OA21x2_ASAP7_75t_L g7001 ( 
.A1(n_6590),
.A2(n_4609),
.B(n_4598),
.Y(n_7001)
);

HB1xp67_ASAP7_75t_L g7002 ( 
.A(n_6513),
.Y(n_7002)
);

INVx1_ASAP7_75t_L g7003 ( 
.A(n_6420),
.Y(n_7003)
);

NAND2xp5_ASAP7_75t_L g7004 ( 
.A(n_6421),
.B(n_6592),
.Y(n_7004)
);

CKINVDCx11_ASAP7_75t_R g7005 ( 
.A(n_6247),
.Y(n_7005)
);

INVx1_ASAP7_75t_L g7006 ( 
.A(n_6555),
.Y(n_7006)
);

INVx2_ASAP7_75t_L g7007 ( 
.A(n_6288),
.Y(n_7007)
);

HB1xp67_ASAP7_75t_L g7008 ( 
.A(n_6534),
.Y(n_7008)
);

HB1xp67_ASAP7_75t_L g7009 ( 
.A(n_6315),
.Y(n_7009)
);

INVx1_ASAP7_75t_L g7010 ( 
.A(n_6556),
.Y(n_7010)
);

INVx2_ASAP7_75t_L g7011 ( 
.A(n_6291),
.Y(n_7011)
);

OA21x2_ASAP7_75t_L g7012 ( 
.A1(n_6594),
.A2(n_4616),
.B(n_4610),
.Y(n_7012)
);

INVx1_ASAP7_75t_L g7013 ( 
.A(n_6557),
.Y(n_7013)
);

BUFx6f_ASAP7_75t_L g7014 ( 
.A(n_6295),
.Y(n_7014)
);

CKINVDCx20_ASAP7_75t_R g7015 ( 
.A(n_6260),
.Y(n_7015)
);

OAI22xp5_ASAP7_75t_L g7016 ( 
.A1(n_6515),
.A2(n_4492),
.B1(n_4494),
.B2(n_4491),
.Y(n_7016)
);

NAND2xp5_ASAP7_75t_L g7017 ( 
.A(n_6595),
.B(n_5723),
.Y(n_7017)
);

NAND2xp5_ASAP7_75t_L g7018 ( 
.A(n_6598),
.B(n_4634),
.Y(n_7018)
);

INVx1_ASAP7_75t_L g7019 ( 
.A(n_6559),
.Y(n_7019)
);

NAND2xp5_ASAP7_75t_L g7020 ( 
.A(n_6601),
.B(n_4651),
.Y(n_7020)
);

BUFx2_ASAP7_75t_L g7021 ( 
.A(n_6438),
.Y(n_7021)
);

INVx2_ASAP7_75t_L g7022 ( 
.A(n_6299),
.Y(n_7022)
);

AND2x4_ASAP7_75t_L g7023 ( 
.A(n_6711),
.B(n_4617),
.Y(n_7023)
);

BUFx6f_ASAP7_75t_L g7024 ( 
.A(n_6301),
.Y(n_7024)
);

OAI22xp5_ASAP7_75t_SL g7025 ( 
.A1(n_6439),
.A2(n_4957),
.B1(n_4986),
.B2(n_4948),
.Y(n_7025)
);

NAND2xp5_ASAP7_75t_L g7026 ( 
.A(n_6461),
.B(n_4695),
.Y(n_7026)
);

INVx2_ASAP7_75t_L g7027 ( 
.A(n_6302),
.Y(n_7027)
);

OAI22xp5_ASAP7_75t_L g7028 ( 
.A1(n_6681),
.A2(n_6682),
.B1(n_6698),
.B2(n_6653),
.Y(n_7028)
);

INVx1_ASAP7_75t_L g7029 ( 
.A(n_6425),
.Y(n_7029)
);

NAND2xp5_ASAP7_75t_L g7030 ( 
.A(n_6463),
.B(n_4711),
.Y(n_7030)
);

AND2x2_ASAP7_75t_L g7031 ( 
.A(n_6526),
.B(n_4917),
.Y(n_7031)
);

AOI22xp5_ASAP7_75t_L g7032 ( 
.A1(n_6650),
.A2(n_5447),
.B1(n_5467),
.B2(n_5402),
.Y(n_7032)
);

INVx2_ASAP7_75t_SL g7033 ( 
.A(n_6363),
.Y(n_7033)
);

INVx1_ASAP7_75t_L g7034 ( 
.A(n_6427),
.Y(n_7034)
);

BUFx8_ASAP7_75t_SL g7035 ( 
.A(n_6275),
.Y(n_7035)
);

HB1xp67_ASAP7_75t_L g7036 ( 
.A(n_6376),
.Y(n_7036)
);

BUFx6f_ASAP7_75t_L g7037 ( 
.A(n_6304),
.Y(n_7037)
);

INVx2_ASAP7_75t_L g7038 ( 
.A(n_6308),
.Y(n_7038)
);

INVx1_ASAP7_75t_L g7039 ( 
.A(n_6309),
.Y(n_7039)
);

BUFx2_ASAP7_75t_L g7040 ( 
.A(n_6442),
.Y(n_7040)
);

AND2x6_ASAP7_75t_L g7041 ( 
.A(n_6686),
.B(n_5508),
.Y(n_7041)
);

INVx2_ASAP7_75t_L g7042 ( 
.A(n_6310),
.Y(n_7042)
);

INVx1_ASAP7_75t_L g7043 ( 
.A(n_6312),
.Y(n_7043)
);

INVx1_ASAP7_75t_L g7044 ( 
.A(n_6317),
.Y(n_7044)
);

AOI22xp5_ASAP7_75t_L g7045 ( 
.A1(n_6552),
.A2(n_5530),
.B1(n_5567),
.B2(n_5523),
.Y(n_7045)
);

INVx1_ASAP7_75t_L g7046 ( 
.A(n_6319),
.Y(n_7046)
);

BUFx3_ASAP7_75t_L g7047 ( 
.A(n_6523),
.Y(n_7047)
);

OAI21x1_ASAP7_75t_L g7048 ( 
.A1(n_6321),
.A2(n_4764),
.B(n_4724),
.Y(n_7048)
);

INVx3_ASAP7_75t_L g7049 ( 
.A(n_6323),
.Y(n_7049)
);

INVx3_ASAP7_75t_L g7050 ( 
.A(n_6324),
.Y(n_7050)
);

AND2x4_ASAP7_75t_L g7051 ( 
.A(n_6714),
.B(n_4623),
.Y(n_7051)
);

OAI22xp5_ASAP7_75t_L g7052 ( 
.A1(n_6563),
.A2(n_4499),
.B1(n_4500),
.B2(n_4496),
.Y(n_7052)
);

BUFx6f_ASAP7_75t_L g7053 ( 
.A(n_6327),
.Y(n_7053)
);

INVx2_ASAP7_75t_L g7054 ( 
.A(n_6328),
.Y(n_7054)
);

INVx2_ASAP7_75t_L g7055 ( 
.A(n_6329),
.Y(n_7055)
);

INVx2_ASAP7_75t_L g7056 ( 
.A(n_6330),
.Y(n_7056)
);

AND2x2_ASAP7_75t_L g7057 ( 
.A(n_6651),
.B(n_5024),
.Y(n_7057)
);

INVx5_ASAP7_75t_L g7058 ( 
.A(n_6606),
.Y(n_7058)
);

BUFx12f_ASAP7_75t_L g7059 ( 
.A(n_6293),
.Y(n_7059)
);

CKINVDCx11_ASAP7_75t_R g7060 ( 
.A(n_6282),
.Y(n_7060)
);

BUFx3_ASAP7_75t_L g7061 ( 
.A(n_6531),
.Y(n_7061)
);

INVx1_ASAP7_75t_L g7062 ( 
.A(n_6331),
.Y(n_7062)
);

INVx1_ASAP7_75t_L g7063 ( 
.A(n_6334),
.Y(n_7063)
);

INVx1_ASAP7_75t_L g7064 ( 
.A(n_6335),
.Y(n_7064)
);

OA21x2_ASAP7_75t_L g7065 ( 
.A1(n_6473),
.A2(n_4633),
.B(n_4625),
.Y(n_7065)
);

BUFx3_ASAP7_75t_L g7066 ( 
.A(n_6536),
.Y(n_7066)
);

INVx1_ASAP7_75t_L g7067 ( 
.A(n_6343),
.Y(n_7067)
);

INVx3_ASAP7_75t_L g7068 ( 
.A(n_6345),
.Y(n_7068)
);

AOI22xp5_ASAP7_75t_L g7069 ( 
.A1(n_6664),
.A2(n_5636),
.B1(n_5661),
.B2(n_5600),
.Y(n_7069)
);

CKINVDCx8_ASAP7_75t_R g7070 ( 
.A(n_6213),
.Y(n_7070)
);

NOR2xp33_ASAP7_75t_SL g7071 ( 
.A(n_6497),
.B(n_5000),
.Y(n_7071)
);

INVx2_ASAP7_75t_L g7072 ( 
.A(n_6350),
.Y(n_7072)
);

AND2x4_ASAP7_75t_L g7073 ( 
.A(n_6305),
.B(n_4635),
.Y(n_7073)
);

BUFx8_ASAP7_75t_L g7074 ( 
.A(n_6455),
.Y(n_7074)
);

INVx1_ASAP7_75t_L g7075 ( 
.A(n_6353),
.Y(n_7075)
);

BUFx6f_ASAP7_75t_L g7076 ( 
.A(n_6356),
.Y(n_7076)
);

OAI22xp5_ASAP7_75t_L g7077 ( 
.A1(n_6294),
.A2(n_4504),
.B1(n_4505),
.B2(n_4503),
.Y(n_7077)
);

CKINVDCx5p33_ASAP7_75t_R g7078 ( 
.A(n_6298),
.Y(n_7078)
);

INVx2_ASAP7_75t_L g7079 ( 
.A(n_6358),
.Y(n_7079)
);

INVx4_ASAP7_75t_L g7080 ( 
.A(n_6300),
.Y(n_7080)
);

BUFx6f_ASAP7_75t_L g7081 ( 
.A(n_6360),
.Y(n_7081)
);

BUFx3_ASAP7_75t_L g7082 ( 
.A(n_6543),
.Y(n_7082)
);

BUFx6f_ASAP7_75t_L g7083 ( 
.A(n_6362),
.Y(n_7083)
);

BUFx6f_ASAP7_75t_L g7084 ( 
.A(n_6364),
.Y(n_7084)
);

INVx2_ASAP7_75t_L g7085 ( 
.A(n_6365),
.Y(n_7085)
);

INVx2_ASAP7_75t_SL g7086 ( 
.A(n_6379),
.Y(n_7086)
);

BUFx6f_ASAP7_75t_L g7087 ( 
.A(n_6366),
.Y(n_7087)
);

INVx1_ASAP7_75t_L g7088 ( 
.A(n_6367),
.Y(n_7088)
);

BUFx6f_ASAP7_75t_L g7089 ( 
.A(n_6368),
.Y(n_7089)
);

INVxp67_ASAP7_75t_L g7090 ( 
.A(n_6670),
.Y(n_7090)
);

BUFx12f_ASAP7_75t_L g7091 ( 
.A(n_6314),
.Y(n_7091)
);

BUFx2_ASAP7_75t_L g7092 ( 
.A(n_6443),
.Y(n_7092)
);

OAI22xp5_ASAP7_75t_SL g7093 ( 
.A1(n_6483),
.A2(n_5027),
.B1(n_5056),
.B2(n_5016),
.Y(n_7093)
);

BUFx6f_ASAP7_75t_L g7094 ( 
.A(n_6369),
.Y(n_7094)
);

BUFx6f_ASAP7_75t_L g7095 ( 
.A(n_6527),
.Y(n_7095)
);

INVx5_ASAP7_75t_L g7096 ( 
.A(n_6624),
.Y(n_7096)
);

AND2x2_ASAP7_75t_SL g7097 ( 
.A(n_6286),
.B(n_4766),
.Y(n_7097)
);

NOR2x1_ASAP7_75t_L g7098 ( 
.A(n_6530),
.B(n_5254),
.Y(n_7098)
);

BUFx8_ASAP7_75t_SL g7099 ( 
.A(n_6297),
.Y(n_7099)
);

INVx2_ASAP7_75t_L g7100 ( 
.A(n_6230),
.Y(n_7100)
);

CKINVDCx5p33_ASAP7_75t_R g7101 ( 
.A(n_6316),
.Y(n_7101)
);

INVx1_ASAP7_75t_L g7102 ( 
.A(n_6537),
.Y(n_7102)
);

NOR2x1_ASAP7_75t_L g7103 ( 
.A(n_6540),
.B(n_6541),
.Y(n_7103)
);

OAI21x1_ASAP7_75t_L g7104 ( 
.A1(n_6499),
.A2(n_4822),
.B(n_4771),
.Y(n_7104)
);

OA21x2_ASAP7_75t_L g7105 ( 
.A1(n_6521),
.A2(n_4642),
.B(n_4637),
.Y(n_7105)
);

AND2x4_ASAP7_75t_L g7106 ( 
.A(n_6548),
.B(n_4649),
.Y(n_7106)
);

CKINVDCx5p33_ASAP7_75t_R g7107 ( 
.A(n_6322),
.Y(n_7107)
);

BUFx3_ASAP7_75t_L g7108 ( 
.A(n_6550),
.Y(n_7108)
);

BUFx6f_ASAP7_75t_L g7109 ( 
.A(n_6546),
.Y(n_7109)
);

NAND2xp5_ASAP7_75t_L g7110 ( 
.A(n_6558),
.B(n_4852),
.Y(n_7110)
);

INVx1_ASAP7_75t_L g7111 ( 
.A(n_6549),
.Y(n_7111)
);

INVx3_ASAP7_75t_L g7112 ( 
.A(n_6551),
.Y(n_7112)
);

OAI22xp5_ASAP7_75t_L g7113 ( 
.A1(n_6325),
.A2(n_6341),
.B1(n_6342),
.B2(n_6340),
.Y(n_7113)
);

AND2x4_ASAP7_75t_L g7114 ( 
.A(n_6688),
.B(n_4653),
.Y(n_7114)
);

INVx2_ASAP7_75t_L g7115 ( 
.A(n_6231),
.Y(n_7115)
);

BUFx6f_ASAP7_75t_L g7116 ( 
.A(n_6233),
.Y(n_7116)
);

AND2x4_ASAP7_75t_L g7117 ( 
.A(n_6449),
.B(n_4659),
.Y(n_7117)
);

AOI22xp5_ASAP7_75t_L g7118 ( 
.A1(n_6344),
.A2(n_5690),
.B1(n_4513),
.B2(n_4514),
.Y(n_7118)
);

INVx2_ASAP7_75t_L g7119 ( 
.A(n_6238),
.Y(n_7119)
);

BUFx6f_ASAP7_75t_L g7120 ( 
.A(n_6241),
.Y(n_7120)
);

CKINVDCx8_ASAP7_75t_R g7121 ( 
.A(n_6629),
.Y(n_7121)
);

INVx2_ASAP7_75t_L g7122 ( 
.A(n_6243),
.Y(n_7122)
);

BUFx6f_ASAP7_75t_L g7123 ( 
.A(n_6244),
.Y(n_7123)
);

INVx1_ASAP7_75t_L g7124 ( 
.A(n_6245),
.Y(n_7124)
);

BUFx6f_ASAP7_75t_L g7125 ( 
.A(n_6246),
.Y(n_7125)
);

INVx3_ASAP7_75t_L g7126 ( 
.A(n_6355),
.Y(n_7126)
);

BUFx6f_ASAP7_75t_L g7127 ( 
.A(n_6357),
.Y(n_7127)
);

INVx2_ASAP7_75t_L g7128 ( 
.A(n_6478),
.Y(n_7128)
);

AND2x4_ASAP7_75t_L g7129 ( 
.A(n_6393),
.B(n_4661),
.Y(n_7129)
);

AND2x4_ASAP7_75t_L g7130 ( 
.A(n_6437),
.B(n_6706),
.Y(n_7130)
);

INVx3_ASAP7_75t_L g7131 ( 
.A(n_6371),
.Y(n_7131)
);

INVx1_ASAP7_75t_L g7132 ( 
.A(n_6372),
.Y(n_7132)
);

AND2x2_ASAP7_75t_L g7133 ( 
.A(n_6210),
.B(n_5024),
.Y(n_7133)
);

INVx1_ASAP7_75t_L g7134 ( 
.A(n_6385),
.Y(n_7134)
);

BUFx12f_ASAP7_75t_L g7135 ( 
.A(n_6388),
.Y(n_7135)
);

BUFx12f_ASAP7_75t_L g7136 ( 
.A(n_6391),
.Y(n_7136)
);

INVx1_ASAP7_75t_L g7137 ( 
.A(n_6399),
.Y(n_7137)
);

INVx1_ASAP7_75t_L g7138 ( 
.A(n_6406),
.Y(n_7138)
);

BUFx2_ASAP7_75t_L g7139 ( 
.A(n_6495),
.Y(n_7139)
);

INVx2_ASAP7_75t_SL g7140 ( 
.A(n_6409),
.Y(n_7140)
);

INVx2_ASAP7_75t_L g7141 ( 
.A(n_6411),
.Y(n_7141)
);

BUFx12f_ASAP7_75t_L g7142 ( 
.A(n_6414),
.Y(n_7142)
);

OAI22xp5_ASAP7_75t_L g7143 ( 
.A1(n_6422),
.A2(n_4521),
.B1(n_4522),
.B2(n_4512),
.Y(n_7143)
);

INVx1_ASAP7_75t_L g7144 ( 
.A(n_6426),
.Y(n_7144)
);

INVx2_ASAP7_75t_L g7145 ( 
.A(n_6435),
.Y(n_7145)
);

NAND2xp5_ASAP7_75t_L g7146 ( 
.A(n_6441),
.B(n_4863),
.Y(n_7146)
);

NOR2xp33_ASAP7_75t_L g7147 ( 
.A(n_6446),
.B(n_4523),
.Y(n_7147)
);

OAI22xp5_ASAP7_75t_SL g7148 ( 
.A1(n_6553),
.A2(n_5074),
.B1(n_5092),
.B2(n_5062),
.Y(n_7148)
);

OA21x2_ASAP7_75t_L g7149 ( 
.A1(n_6476),
.A2(n_4670),
.B(n_4664),
.Y(n_7149)
);

NAND2xp5_ASAP7_75t_L g7150 ( 
.A(n_6490),
.B(n_4909),
.Y(n_7150)
);

CKINVDCx5p33_ASAP7_75t_R g7151 ( 
.A(n_6492),
.Y(n_7151)
);

BUFx6f_ASAP7_75t_L g7152 ( 
.A(n_6500),
.Y(n_7152)
);

NOR2xp33_ASAP7_75t_L g7153 ( 
.A(n_6502),
.B(n_4524),
.Y(n_7153)
);

BUFx6f_ASAP7_75t_L g7154 ( 
.A(n_6516),
.Y(n_7154)
);

INVx1_ASAP7_75t_L g7155 ( 
.A(n_6524),
.Y(n_7155)
);

INVx3_ASAP7_75t_L g7156 ( 
.A(n_6528),
.Y(n_7156)
);

CKINVDCx5p33_ASAP7_75t_R g7157 ( 
.A(n_6533),
.Y(n_7157)
);

CKINVDCx20_ASAP7_75t_R g7158 ( 
.A(n_6332),
.Y(n_7158)
);

INVx2_ASAP7_75t_L g7159 ( 
.A(n_6535),
.Y(n_7159)
);

BUFx6f_ASAP7_75t_L g7160 ( 
.A(n_6545),
.Y(n_7160)
);

INVx2_ASAP7_75t_L g7161 ( 
.A(n_6547),
.Y(n_7161)
);

OAI21x1_ASAP7_75t_L g7162 ( 
.A1(n_6514),
.A2(n_4960),
.B(n_4950),
.Y(n_7162)
);

INVx2_ASAP7_75t_L g7163 ( 
.A(n_6561),
.Y(n_7163)
);

BUFx6f_ASAP7_75t_L g7164 ( 
.A(n_6566),
.Y(n_7164)
);

INVx1_ASAP7_75t_L g7165 ( 
.A(n_6568),
.Y(n_7165)
);

AOI22xp5_ASAP7_75t_L g7166 ( 
.A1(n_6572),
.A2(n_4531),
.B1(n_4534),
.B2(n_4530),
.Y(n_7166)
);

INVx3_ASAP7_75t_L g7167 ( 
.A(n_6585),
.Y(n_7167)
);

BUFx3_ASAP7_75t_L g7168 ( 
.A(n_6554),
.Y(n_7168)
);

INVx4_ASAP7_75t_L g7169 ( 
.A(n_6596),
.Y(n_7169)
);

NOR2xp33_ASAP7_75t_SL g7170 ( 
.A(n_6447),
.B(n_6469),
.Y(n_7170)
);

INVx1_ASAP7_75t_L g7171 ( 
.A(n_6600),
.Y(n_7171)
);

INVx5_ASAP7_75t_L g7172 ( 
.A(n_6649),
.Y(n_7172)
);

BUFx6f_ASAP7_75t_L g7173 ( 
.A(n_6610),
.Y(n_7173)
);

INVx1_ASAP7_75t_L g7174 ( 
.A(n_6626),
.Y(n_7174)
);

BUFx6f_ASAP7_75t_L g7175 ( 
.A(n_6627),
.Y(n_7175)
);

AND2x2_ASAP7_75t_L g7176 ( 
.A(n_6237),
.B(n_5080),
.Y(n_7176)
);

INVx1_ASAP7_75t_L g7177 ( 
.A(n_6638),
.Y(n_7177)
);

INVx1_ASAP7_75t_L g7178 ( 
.A(n_6639),
.Y(n_7178)
);

HB1xp67_ASAP7_75t_L g7179 ( 
.A(n_6640),
.Y(n_7179)
);

INVx4_ASAP7_75t_L g7180 ( 
.A(n_6645),
.Y(n_7180)
);

INVx2_ASAP7_75t_L g7181 ( 
.A(n_6652),
.Y(n_7181)
);

AND2x2_ASAP7_75t_L g7182 ( 
.A(n_6654),
.B(n_5080),
.Y(n_7182)
);

AND2x6_ASAP7_75t_L g7183 ( 
.A(n_6532),
.B(n_4673),
.Y(n_7183)
);

INVx3_ASAP7_75t_L g7184 ( 
.A(n_6655),
.Y(n_7184)
);

BUFx6f_ASAP7_75t_L g7185 ( 
.A(n_6657),
.Y(n_7185)
);

INVx2_ASAP7_75t_L g7186 ( 
.A(n_6663),
.Y(n_7186)
);

INVx1_ASAP7_75t_L g7187 ( 
.A(n_6666),
.Y(n_7187)
);

INVx2_ASAP7_75t_L g7188 ( 
.A(n_6564),
.Y(n_7188)
);

OAI22xp5_ASAP7_75t_L g7189 ( 
.A1(n_6605),
.A2(n_4538),
.B1(n_4540),
.B2(n_4535),
.Y(n_7189)
);

BUFx6f_ASAP7_75t_L g7190 ( 
.A(n_6479),
.Y(n_7190)
);

OAI21x1_ASAP7_75t_L g7191 ( 
.A1(n_6539),
.A2(n_4985),
.B(n_4967),
.Y(n_7191)
);

NAND2xp5_ASAP7_75t_L g7192 ( 
.A(n_6208),
.B(n_4990),
.Y(n_7192)
);

CKINVDCx5p33_ASAP7_75t_R g7193 ( 
.A(n_6333),
.Y(n_7193)
);

NAND2xp5_ASAP7_75t_L g7194 ( 
.A(n_6223),
.B(n_4999),
.Y(n_7194)
);

BUFx6f_ASAP7_75t_L g7195 ( 
.A(n_6679),
.Y(n_7195)
);

XOR2xp5_ASAP7_75t_L g7196 ( 
.A(n_6338),
.B(n_5115),
.Y(n_7196)
);

INVx1_ASAP7_75t_L g7197 ( 
.A(n_6584),
.Y(n_7197)
);

AND2x2_ASAP7_75t_SL g7198 ( 
.A(n_6691),
.B(n_5053),
.Y(n_7198)
);

BUFx8_ASAP7_75t_L g7199 ( 
.A(n_6407),
.Y(n_7199)
);

BUFx6f_ASAP7_75t_L g7200 ( 
.A(n_6687),
.Y(n_7200)
);

INVx2_ASAP7_75t_SL g7201 ( 
.A(n_6586),
.Y(n_7201)
);

INVx1_ASAP7_75t_L g7202 ( 
.A(n_6588),
.Y(n_7202)
);

INVx1_ASAP7_75t_L g7203 ( 
.A(n_6591),
.Y(n_7203)
);

INVx2_ASAP7_75t_L g7204 ( 
.A(n_6593),
.Y(n_7204)
);

BUFx6f_ASAP7_75t_L g7205 ( 
.A(n_6349),
.Y(n_7205)
);

BUFx6f_ASAP7_75t_L g7206 ( 
.A(n_6354),
.Y(n_7206)
);

BUFx6f_ASAP7_75t_L g7207 ( 
.A(n_6395),
.Y(n_7207)
);

INVx2_ASAP7_75t_L g7208 ( 
.A(n_6597),
.Y(n_7208)
);

INVx2_ASAP7_75t_L g7209 ( 
.A(n_6612),
.Y(n_7209)
);

BUFx6f_ASAP7_75t_L g7210 ( 
.A(n_6400),
.Y(n_7210)
);

BUFx12f_ASAP7_75t_L g7211 ( 
.A(n_6289),
.Y(n_7211)
);

BUFx6f_ASAP7_75t_L g7212 ( 
.A(n_6618),
.Y(n_7212)
);

INVx3_ASAP7_75t_L g7213 ( 
.A(n_6619),
.Y(n_7213)
);

INVx2_ASAP7_75t_L g7214 ( 
.A(n_6630),
.Y(n_7214)
);

BUFx6f_ASAP7_75t_L g7215 ( 
.A(n_6660),
.Y(n_7215)
);

BUFx3_ASAP7_75t_L g7216 ( 
.A(n_6635),
.Y(n_7216)
);

CKINVDCx5p33_ASAP7_75t_R g7217 ( 
.A(n_6659),
.Y(n_7217)
);

INVx3_ASAP7_75t_L g7218 ( 
.A(n_6451),
.Y(n_7218)
);

NAND2xp5_ASAP7_75t_L g7219 ( 
.A(n_6560),
.B(n_5066),
.Y(n_7219)
);

BUFx8_ASAP7_75t_SL g7220 ( 
.A(n_6214),
.Y(n_7220)
);

INVx3_ASAP7_75t_L g7221 ( 
.A(n_6451),
.Y(n_7221)
);

INVx2_ASAP7_75t_L g7222 ( 
.A(n_6542),
.Y(n_7222)
);

BUFx2_ASAP7_75t_L g7223 ( 
.A(n_6609),
.Y(n_7223)
);

AND2x2_ASAP7_75t_L g7224 ( 
.A(n_6609),
.B(n_5139),
.Y(n_7224)
);

BUFx6f_ASAP7_75t_L g7225 ( 
.A(n_6451),
.Y(n_7225)
);

INVx2_ASAP7_75t_L g7226 ( 
.A(n_6542),
.Y(n_7226)
);

BUFx6f_ASAP7_75t_L g7227 ( 
.A(n_6451),
.Y(n_7227)
);

INVx1_ASAP7_75t_L g7228 ( 
.A(n_6428),
.Y(n_7228)
);

NOR2xp33_ASAP7_75t_L g7229 ( 
.A(n_6567),
.B(n_4541),
.Y(n_7229)
);

INVx1_ASAP7_75t_L g7230 ( 
.A(n_6428),
.Y(n_7230)
);

INVx2_ASAP7_75t_L g7231 ( 
.A(n_6542),
.Y(n_7231)
);

INVxp67_ASAP7_75t_L g7232 ( 
.A(n_6628),
.Y(n_7232)
);

BUFx6f_ASAP7_75t_L g7233 ( 
.A(n_6451),
.Y(n_7233)
);

HB1xp67_ASAP7_75t_L g7234 ( 
.A(n_6628),
.Y(n_7234)
);

INVx2_ASAP7_75t_L g7235 ( 
.A(n_6542),
.Y(n_7235)
);

INVx1_ASAP7_75t_L g7236 ( 
.A(n_6428),
.Y(n_7236)
);

INVx2_ASAP7_75t_L g7237 ( 
.A(n_6542),
.Y(n_7237)
);

INVx2_ASAP7_75t_L g7238 ( 
.A(n_6542),
.Y(n_7238)
);

AND2x2_ASAP7_75t_L g7239 ( 
.A(n_6609),
.B(n_5139),
.Y(n_7239)
);

AND2x4_ASAP7_75t_L g7240 ( 
.A(n_6348),
.B(n_4674),
.Y(n_7240)
);

INVx2_ASAP7_75t_L g7241 ( 
.A(n_6542),
.Y(n_7241)
);

AND2x2_ASAP7_75t_L g7242 ( 
.A(n_6609),
.B(n_5166),
.Y(n_7242)
);

BUFx6f_ASAP7_75t_L g7243 ( 
.A(n_6451),
.Y(n_7243)
);

INVx2_ASAP7_75t_L g7244 ( 
.A(n_6542),
.Y(n_7244)
);

AND2x2_ASAP7_75t_L g7245 ( 
.A(n_6609),
.B(n_5166),
.Y(n_7245)
);

BUFx6f_ASAP7_75t_L g7246 ( 
.A(n_6451),
.Y(n_7246)
);

INVx2_ASAP7_75t_L g7247 ( 
.A(n_6542),
.Y(n_7247)
);

INVx2_ASAP7_75t_L g7248 ( 
.A(n_6542),
.Y(n_7248)
);

BUFx12f_ASAP7_75t_L g7249 ( 
.A(n_6262),
.Y(n_7249)
);

AND2x2_ASAP7_75t_L g7250 ( 
.A(n_6609),
.B(n_5206),
.Y(n_7250)
);

INVx1_ASAP7_75t_L g7251 ( 
.A(n_6428),
.Y(n_7251)
);

INVx2_ASAP7_75t_L g7252 ( 
.A(n_6542),
.Y(n_7252)
);

INVx2_ASAP7_75t_L g7253 ( 
.A(n_6542),
.Y(n_7253)
);

BUFx6f_ASAP7_75t_L g7254 ( 
.A(n_6451),
.Y(n_7254)
);

NAND2xp5_ASAP7_75t_L g7255 ( 
.A(n_6560),
.B(n_5107),
.Y(n_7255)
);

CKINVDCx20_ASAP7_75t_R g7256 ( 
.A(n_6206),
.Y(n_7256)
);

INVx4_ASAP7_75t_L g7257 ( 
.A(n_6661),
.Y(n_7257)
);

INVx1_ASAP7_75t_L g7258 ( 
.A(n_6428),
.Y(n_7258)
);

INVx1_ASAP7_75t_L g7259 ( 
.A(n_6428),
.Y(n_7259)
);

NAND2xp5_ASAP7_75t_L g7260 ( 
.A(n_6560),
.B(n_5134),
.Y(n_7260)
);

INVx3_ASAP7_75t_L g7261 ( 
.A(n_6451),
.Y(n_7261)
);

INVx2_ASAP7_75t_L g7262 ( 
.A(n_6542),
.Y(n_7262)
);

HB1xp67_ASAP7_75t_L g7263 ( 
.A(n_6628),
.Y(n_7263)
);

NAND2xp5_ASAP7_75t_L g7264 ( 
.A(n_6560),
.B(n_5151),
.Y(n_7264)
);

NOR2xp33_ASAP7_75t_L g7265 ( 
.A(n_6567),
.B(n_4542),
.Y(n_7265)
);

NOR2xp33_ASAP7_75t_L g7266 ( 
.A(n_6567),
.B(n_4544),
.Y(n_7266)
);

NOR2xp33_ASAP7_75t_L g7267 ( 
.A(n_6567),
.B(n_4545),
.Y(n_7267)
);

INVx5_ASAP7_75t_L g7268 ( 
.A(n_6296),
.Y(n_7268)
);

HB1xp67_ASAP7_75t_L g7269 ( 
.A(n_6628),
.Y(n_7269)
);

INVx1_ASAP7_75t_L g7270 ( 
.A(n_6428),
.Y(n_7270)
);

INVx2_ASAP7_75t_L g7271 ( 
.A(n_6542),
.Y(n_7271)
);

BUFx6f_ASAP7_75t_L g7272 ( 
.A(n_6451),
.Y(n_7272)
);

CKINVDCx14_ASAP7_75t_R g7273 ( 
.A(n_6336),
.Y(n_7273)
);

NOR2xp33_ASAP7_75t_L g7274 ( 
.A(n_6567),
.B(n_4550),
.Y(n_7274)
);

BUFx6f_ASAP7_75t_L g7275 ( 
.A(n_6451),
.Y(n_7275)
);

INVx2_ASAP7_75t_L g7276 ( 
.A(n_6542),
.Y(n_7276)
);

INVx5_ASAP7_75t_L g7277 ( 
.A(n_6296),
.Y(n_7277)
);

BUFx6f_ASAP7_75t_L g7278 ( 
.A(n_6451),
.Y(n_7278)
);

BUFx6f_ASAP7_75t_L g7279 ( 
.A(n_6451),
.Y(n_7279)
);

OAI22x1_ASAP7_75t_R g7280 ( 
.A1(n_6311),
.A2(n_5211),
.B1(n_5257),
.B2(n_5183),
.Y(n_7280)
);

AND2x4_ASAP7_75t_L g7281 ( 
.A(n_6348),
.B(n_4682),
.Y(n_7281)
);

HB1xp67_ASAP7_75t_L g7282 ( 
.A(n_6628),
.Y(n_7282)
);

INVx2_ASAP7_75t_L g7283 ( 
.A(n_6542),
.Y(n_7283)
);

INVx2_ASAP7_75t_L g7284 ( 
.A(n_6542),
.Y(n_7284)
);

INVx1_ASAP7_75t_L g7285 ( 
.A(n_6428),
.Y(n_7285)
);

AND2x6_ASAP7_75t_L g7286 ( 
.A(n_6661),
.B(n_4683),
.Y(n_7286)
);

INVx4_ASAP7_75t_L g7287 ( 
.A(n_6661),
.Y(n_7287)
);

OAI22xp5_ASAP7_75t_L g7288 ( 
.A1(n_6417),
.A2(n_4554),
.B1(n_4557),
.B2(n_4552),
.Y(n_7288)
);

INVx2_ASAP7_75t_L g7289 ( 
.A(n_6542),
.Y(n_7289)
);

INVx2_ASAP7_75t_SL g7290 ( 
.A(n_6628),
.Y(n_7290)
);

BUFx6f_ASAP7_75t_L g7291 ( 
.A(n_6451),
.Y(n_7291)
);

AOI22xp5_ASAP7_75t_L g7292 ( 
.A1(n_6567),
.A2(n_4562),
.B1(n_4563),
.B2(n_4561),
.Y(n_7292)
);

INVx4_ASAP7_75t_L g7293 ( 
.A(n_6661),
.Y(n_7293)
);

BUFx6f_ASAP7_75t_L g7294 ( 
.A(n_6451),
.Y(n_7294)
);

BUFx6f_ASAP7_75t_L g7295 ( 
.A(n_6451),
.Y(n_7295)
);

INVx3_ASAP7_75t_L g7296 ( 
.A(n_6451),
.Y(n_7296)
);

INVx2_ASAP7_75t_L g7297 ( 
.A(n_6542),
.Y(n_7297)
);

NOR2xp33_ASAP7_75t_L g7298 ( 
.A(n_7232),
.B(n_4564),
.Y(n_7298)
);

INVx1_ASAP7_75t_L g7299 ( 
.A(n_6722),
.Y(n_7299)
);

CKINVDCx5p33_ASAP7_75t_R g7300 ( 
.A(n_6835),
.Y(n_7300)
);

CKINVDCx20_ASAP7_75t_R g7301 ( 
.A(n_6882),
.Y(n_7301)
);

CKINVDCx5p33_ASAP7_75t_R g7302 ( 
.A(n_7035),
.Y(n_7302)
);

INVx1_ASAP7_75t_L g7303 ( 
.A(n_6731),
.Y(n_7303)
);

INVx1_ASAP7_75t_L g7304 ( 
.A(n_7285),
.Y(n_7304)
);

INVx3_ASAP7_75t_L g7305 ( 
.A(n_7290),
.Y(n_7305)
);

OAI22xp5_ASAP7_75t_L g7306 ( 
.A1(n_6734),
.A2(n_4569),
.B1(n_4570),
.B2(n_4566),
.Y(n_7306)
);

AND2x2_ASAP7_75t_L g7307 ( 
.A(n_7234),
.B(n_5206),
.Y(n_7307)
);

INVx2_ASAP7_75t_L g7308 ( 
.A(n_6775),
.Y(n_7308)
);

HB1xp67_ASAP7_75t_L g7309 ( 
.A(n_7263),
.Y(n_7309)
);

INVx2_ASAP7_75t_L g7310 ( 
.A(n_6777),
.Y(n_7310)
);

CKINVDCx5p33_ASAP7_75t_R g7311 ( 
.A(n_7099),
.Y(n_7311)
);

INVx2_ASAP7_75t_L g7312 ( 
.A(n_6780),
.Y(n_7312)
);

HB1xp67_ASAP7_75t_L g7313 ( 
.A(n_7282),
.Y(n_7313)
);

CKINVDCx5p33_ASAP7_75t_R g7314 ( 
.A(n_7220),
.Y(n_7314)
);

CKINVDCx5p33_ASAP7_75t_R g7315 ( 
.A(n_6786),
.Y(n_7315)
);

AND2x4_ASAP7_75t_L g7316 ( 
.A(n_6761),
.B(n_4689),
.Y(n_7316)
);

INVx2_ASAP7_75t_L g7317 ( 
.A(n_6755),
.Y(n_7317)
);

BUFx6f_ASAP7_75t_L g7318 ( 
.A(n_6723),
.Y(n_7318)
);

INVx1_ASAP7_75t_L g7319 ( 
.A(n_6773),
.Y(n_7319)
);

INVx2_ASAP7_75t_L g7320 ( 
.A(n_6756),
.Y(n_7320)
);

CKINVDCx8_ASAP7_75t_R g7321 ( 
.A(n_7268),
.Y(n_7321)
);

INVx1_ASAP7_75t_L g7322 ( 
.A(n_6778),
.Y(n_7322)
);

INVx2_ASAP7_75t_L g7323 ( 
.A(n_6763),
.Y(n_7323)
);

INVx1_ASAP7_75t_L g7324 ( 
.A(n_6781),
.Y(n_7324)
);

AND2x2_ASAP7_75t_L g7325 ( 
.A(n_7269),
.B(n_5218),
.Y(n_7325)
);

INVx5_ASAP7_75t_L g7326 ( 
.A(n_6766),
.Y(n_7326)
);

CKINVDCx20_ASAP7_75t_R g7327 ( 
.A(n_6994),
.Y(n_7327)
);

HB1xp67_ASAP7_75t_L g7328 ( 
.A(n_6770),
.Y(n_7328)
);

INVx1_ASAP7_75t_L g7329 ( 
.A(n_6784),
.Y(n_7329)
);

XOR2xp5_ASAP7_75t_L g7330 ( 
.A(n_7015),
.B(n_5266),
.Y(n_7330)
);

BUFx6f_ASAP7_75t_L g7331 ( 
.A(n_6717),
.Y(n_7331)
);

INVx1_ASAP7_75t_L g7332 ( 
.A(n_6787),
.Y(n_7332)
);

INVx1_ASAP7_75t_L g7333 ( 
.A(n_6791),
.Y(n_7333)
);

CKINVDCx20_ASAP7_75t_R g7334 ( 
.A(n_7158),
.Y(n_7334)
);

INVx2_ASAP7_75t_L g7335 ( 
.A(n_6838),
.Y(n_7335)
);

CKINVDCx5p33_ASAP7_75t_R g7336 ( 
.A(n_6900),
.Y(n_7336)
);

CKINVDCx5p33_ASAP7_75t_R g7337 ( 
.A(n_6997),
.Y(n_7337)
);

AND2x4_ASAP7_75t_L g7338 ( 
.A(n_6732),
.B(n_4690),
.Y(n_7338)
);

OR2x2_ASAP7_75t_L g7339 ( 
.A(n_6821),
.B(n_5285),
.Y(n_7339)
);

INVx1_ASAP7_75t_L g7340 ( 
.A(n_6802),
.Y(n_7340)
);

HB1xp67_ASAP7_75t_L g7341 ( 
.A(n_6809),
.Y(n_7341)
);

INVx2_ASAP7_75t_L g7342 ( 
.A(n_6847),
.Y(n_7342)
);

CKINVDCx5p33_ASAP7_75t_R g7343 ( 
.A(n_6998),
.Y(n_7343)
);

CKINVDCx5p33_ASAP7_75t_R g7344 ( 
.A(n_7078),
.Y(n_7344)
);

AND2x2_ASAP7_75t_L g7345 ( 
.A(n_6725),
.B(n_5218),
.Y(n_7345)
);

CKINVDCx5p33_ASAP7_75t_R g7346 ( 
.A(n_7101),
.Y(n_7346)
);

BUFx6f_ASAP7_75t_L g7347 ( 
.A(n_6719),
.Y(n_7347)
);

INVxp67_ASAP7_75t_L g7348 ( 
.A(n_7223),
.Y(n_7348)
);

NAND2xp5_ASAP7_75t_L g7349 ( 
.A(n_7004),
.B(n_7229),
.Y(n_7349)
);

INVx1_ASAP7_75t_L g7350 ( 
.A(n_6817),
.Y(n_7350)
);

AND2x2_ASAP7_75t_L g7351 ( 
.A(n_6824),
.B(n_5220),
.Y(n_7351)
);

BUFx3_ASAP7_75t_L g7352 ( 
.A(n_6741),
.Y(n_7352)
);

INVx3_ASAP7_75t_L g7353 ( 
.A(n_6744),
.Y(n_7353)
);

INVxp67_ASAP7_75t_L g7354 ( 
.A(n_6968),
.Y(n_7354)
);

AND2x4_ASAP7_75t_L g7355 ( 
.A(n_6764),
.B(n_4694),
.Y(n_7355)
);

CKINVDCx5p33_ASAP7_75t_R g7356 ( 
.A(n_7107),
.Y(n_7356)
);

AND2x4_ASAP7_75t_L g7357 ( 
.A(n_6730),
.B(n_4697),
.Y(n_7357)
);

NAND2xp33_ASAP7_75t_R g7358 ( 
.A(n_6788),
.B(n_4571),
.Y(n_7358)
);

CKINVDCx5p33_ASAP7_75t_R g7359 ( 
.A(n_7151),
.Y(n_7359)
);

INVx1_ASAP7_75t_L g7360 ( 
.A(n_6823),
.Y(n_7360)
);

BUFx6f_ASAP7_75t_L g7361 ( 
.A(n_7225),
.Y(n_7361)
);

BUFx3_ASAP7_75t_L g7362 ( 
.A(n_6750),
.Y(n_7362)
);

INVx2_ASAP7_75t_L g7363 ( 
.A(n_6769),
.Y(n_7363)
);

INVx1_ASAP7_75t_L g7364 ( 
.A(n_6843),
.Y(n_7364)
);

INVx6_ASAP7_75t_L g7365 ( 
.A(n_6892),
.Y(n_7365)
);

NOR2xp67_ASAP7_75t_L g7366 ( 
.A(n_7090),
.B(n_4280),
.Y(n_7366)
);

INVx3_ASAP7_75t_L g7367 ( 
.A(n_6751),
.Y(n_7367)
);

NOR2xp33_ASAP7_75t_L g7368 ( 
.A(n_6909),
.B(n_4573),
.Y(n_7368)
);

INVx1_ASAP7_75t_L g7369 ( 
.A(n_6845),
.Y(n_7369)
);

NAND2xp33_ASAP7_75t_R g7370 ( 
.A(n_7149),
.B(n_4574),
.Y(n_7370)
);

INVx1_ASAP7_75t_L g7371 ( 
.A(n_6848),
.Y(n_7371)
);

INVx1_ASAP7_75t_L g7372 ( 
.A(n_6852),
.Y(n_7372)
);

CKINVDCx5p33_ASAP7_75t_R g7373 ( 
.A(n_7157),
.Y(n_7373)
);

INVx1_ASAP7_75t_L g7374 ( 
.A(n_6853),
.Y(n_7374)
);

INVx1_ASAP7_75t_L g7375 ( 
.A(n_6858),
.Y(n_7375)
);

BUFx6f_ASAP7_75t_L g7376 ( 
.A(n_7227),
.Y(n_7376)
);

INVx3_ASAP7_75t_L g7377 ( 
.A(n_7095),
.Y(n_7377)
);

CKINVDCx5p33_ASAP7_75t_R g7378 ( 
.A(n_7193),
.Y(n_7378)
);

INVxp67_ASAP7_75t_SL g7379 ( 
.A(n_6782),
.Y(n_7379)
);

HB1xp67_ASAP7_75t_L g7380 ( 
.A(n_6789),
.Y(n_7380)
);

INVx2_ASAP7_75t_L g7381 ( 
.A(n_6795),
.Y(n_7381)
);

INVx3_ASAP7_75t_L g7382 ( 
.A(n_7109),
.Y(n_7382)
);

HB1xp67_ASAP7_75t_L g7383 ( 
.A(n_6867),
.Y(n_7383)
);

AND2x2_ASAP7_75t_L g7384 ( 
.A(n_6739),
.B(n_5220),
.Y(n_7384)
);

INVx1_ASAP7_75t_L g7385 ( 
.A(n_6860),
.Y(n_7385)
);

CKINVDCx20_ASAP7_75t_R g7386 ( 
.A(n_7256),
.Y(n_7386)
);

HB1xp67_ASAP7_75t_L g7387 ( 
.A(n_7002),
.Y(n_7387)
);

AND2x4_ASAP7_75t_L g7388 ( 
.A(n_7257),
.B(n_4702),
.Y(n_7388)
);

INVx2_ASAP7_75t_L g7389 ( 
.A(n_6796),
.Y(n_7389)
);

CKINVDCx5p33_ASAP7_75t_R g7390 ( 
.A(n_6776),
.Y(n_7390)
);

CKINVDCx20_ASAP7_75t_R g7391 ( 
.A(n_6863),
.Y(n_7391)
);

INVx1_ASAP7_75t_L g7392 ( 
.A(n_6865),
.Y(n_7392)
);

INVx2_ASAP7_75t_L g7393 ( 
.A(n_6801),
.Y(n_7393)
);

OA21x2_ASAP7_75t_L g7394 ( 
.A1(n_6894),
.A2(n_4708),
.B(n_4707),
.Y(n_7394)
);

INVx3_ASAP7_75t_L g7395 ( 
.A(n_6957),
.Y(n_7395)
);

INVxp67_ASAP7_75t_L g7396 ( 
.A(n_7224),
.Y(n_7396)
);

NOR2xp33_ASAP7_75t_L g7397 ( 
.A(n_6915),
.B(n_4577),
.Y(n_7397)
);

NAND3xp33_ASAP7_75t_L g7398 ( 
.A(n_7265),
.B(n_7267),
.C(n_7266),
.Y(n_7398)
);

INVx3_ASAP7_75t_L g7399 ( 
.A(n_6965),
.Y(n_7399)
);

INVx1_ASAP7_75t_L g7400 ( 
.A(n_6869),
.Y(n_7400)
);

INVx1_ASAP7_75t_L g7401 ( 
.A(n_6870),
.Y(n_7401)
);

OAI21x1_ASAP7_75t_L g7402 ( 
.A1(n_7104),
.A2(n_5174),
.B(n_5157),
.Y(n_7402)
);

INVx1_ASAP7_75t_L g7403 ( 
.A(n_6871),
.Y(n_7403)
);

NAND2xp5_ASAP7_75t_SL g7404 ( 
.A(n_7287),
.B(n_4581),
.Y(n_7404)
);

INVx1_ASAP7_75t_L g7405 ( 
.A(n_6874),
.Y(n_7405)
);

CKINVDCx20_ASAP7_75t_R g7406 ( 
.A(n_6880),
.Y(n_7406)
);

INVx2_ASAP7_75t_L g7407 ( 
.A(n_6808),
.Y(n_7407)
);

CKINVDCx20_ASAP7_75t_R g7408 ( 
.A(n_7005),
.Y(n_7408)
);

AND2x2_ASAP7_75t_L g7409 ( 
.A(n_7239),
.B(n_5321),
.Y(n_7409)
);

INVx3_ASAP7_75t_L g7410 ( 
.A(n_6966),
.Y(n_7410)
);

CKINVDCx5p33_ASAP7_75t_R g7411 ( 
.A(n_7060),
.Y(n_7411)
);

CKINVDCx5p33_ASAP7_75t_R g7412 ( 
.A(n_7217),
.Y(n_7412)
);

AOI22xp5_ASAP7_75t_L g7413 ( 
.A1(n_6767),
.A2(n_5348),
.B1(n_5355),
.B2(n_5338),
.Y(n_7413)
);

CKINVDCx20_ASAP7_75t_R g7414 ( 
.A(n_6738),
.Y(n_7414)
);

CKINVDCx5p33_ASAP7_75t_R g7415 ( 
.A(n_6746),
.Y(n_7415)
);

CKINVDCx20_ASAP7_75t_R g7416 ( 
.A(n_6846),
.Y(n_7416)
);

INVx3_ASAP7_75t_L g7417 ( 
.A(n_6970),
.Y(n_7417)
);

INVx2_ASAP7_75t_L g7418 ( 
.A(n_6811),
.Y(n_7418)
);

CKINVDCx20_ASAP7_75t_R g7419 ( 
.A(n_7273),
.Y(n_7419)
);

NAND2xp33_ASAP7_75t_R g7420 ( 
.A(n_7031),
.B(n_4582),
.Y(n_7420)
);

INVx1_ASAP7_75t_L g7421 ( 
.A(n_6879),
.Y(n_7421)
);

BUFx2_ASAP7_75t_L g7422 ( 
.A(n_6833),
.Y(n_7422)
);

BUFx6f_ASAP7_75t_L g7423 ( 
.A(n_7233),
.Y(n_7423)
);

CKINVDCx5p33_ASAP7_75t_R g7424 ( 
.A(n_6748),
.Y(n_7424)
);

INVx1_ASAP7_75t_L g7425 ( 
.A(n_6893),
.Y(n_7425)
);

INVx2_ASAP7_75t_L g7426 ( 
.A(n_6812),
.Y(n_7426)
);

CKINVDCx5p33_ASAP7_75t_R g7427 ( 
.A(n_6768),
.Y(n_7427)
);

AND2x2_ASAP7_75t_L g7428 ( 
.A(n_7242),
.B(n_5321),
.Y(n_7428)
);

OAI21x1_ASAP7_75t_L g7429 ( 
.A1(n_6740),
.A2(n_5272),
.B(n_5240),
.Y(n_7429)
);

BUFx6f_ASAP7_75t_L g7430 ( 
.A(n_7243),
.Y(n_7430)
);

INVx2_ASAP7_75t_L g7431 ( 
.A(n_6814),
.Y(n_7431)
);

INVx1_ASAP7_75t_L g7432 ( 
.A(n_6899),
.Y(n_7432)
);

INVx2_ASAP7_75t_L g7433 ( 
.A(n_6825),
.Y(n_7433)
);

INVx1_ASAP7_75t_L g7434 ( 
.A(n_6907),
.Y(n_7434)
);

CKINVDCx5p33_ASAP7_75t_R g7435 ( 
.A(n_6898),
.Y(n_7435)
);

INVx3_ASAP7_75t_L g7436 ( 
.A(n_6977),
.Y(n_7436)
);

NAND3xp33_ASAP7_75t_L g7437 ( 
.A(n_7274),
.B(n_4586),
.C(n_4585),
.Y(n_7437)
);

INVx3_ASAP7_75t_L g7438 ( 
.A(n_6978),
.Y(n_7438)
);

INVx1_ASAP7_75t_L g7439 ( 
.A(n_6913),
.Y(n_7439)
);

INVxp67_ASAP7_75t_L g7440 ( 
.A(n_7245),
.Y(n_7440)
);

INVx1_ASAP7_75t_L g7441 ( 
.A(n_6914),
.Y(n_7441)
);

INVx2_ASAP7_75t_L g7442 ( 
.A(n_6831),
.Y(n_7442)
);

BUFx2_ASAP7_75t_L g7443 ( 
.A(n_6833),
.Y(n_7443)
);

INVx2_ASAP7_75t_L g7444 ( 
.A(n_6837),
.Y(n_7444)
);

CKINVDCx20_ASAP7_75t_R g7445 ( 
.A(n_6954),
.Y(n_7445)
);

INVx1_ASAP7_75t_L g7446 ( 
.A(n_6925),
.Y(n_7446)
);

INVx1_ASAP7_75t_L g7447 ( 
.A(n_6932),
.Y(n_7447)
);

INVx2_ASAP7_75t_L g7448 ( 
.A(n_7100),
.Y(n_7448)
);

INVx1_ASAP7_75t_L g7449 ( 
.A(n_6942),
.Y(n_7449)
);

OA21x2_ASAP7_75t_L g7450 ( 
.A1(n_6813),
.A2(n_4715),
.B(n_4712),
.Y(n_7450)
);

CKINVDCx5p33_ASAP7_75t_R g7451 ( 
.A(n_7059),
.Y(n_7451)
);

INVx1_ASAP7_75t_L g7452 ( 
.A(n_6947),
.Y(n_7452)
);

AND2x4_ASAP7_75t_L g7453 ( 
.A(n_7293),
.B(n_4731),
.Y(n_7453)
);

BUFx10_ASAP7_75t_L g7454 ( 
.A(n_7195),
.Y(n_7454)
);

CKINVDCx5p33_ASAP7_75t_R g7455 ( 
.A(n_7091),
.Y(n_7455)
);

AND2x6_ASAP7_75t_L g7456 ( 
.A(n_7141),
.B(n_4738),
.Y(n_7456)
);

CKINVDCx6p67_ASAP7_75t_R g7457 ( 
.A(n_7172),
.Y(n_7457)
);

INVx1_ASAP7_75t_L g7458 ( 
.A(n_6955),
.Y(n_7458)
);

AND2x4_ASAP7_75t_L g7459 ( 
.A(n_7240),
.B(n_4739),
.Y(n_7459)
);

CKINVDCx5p33_ASAP7_75t_R g7460 ( 
.A(n_7135),
.Y(n_7460)
);

CKINVDCx5p33_ASAP7_75t_R g7461 ( 
.A(n_7136),
.Y(n_7461)
);

NAND2xp5_ASAP7_75t_L g7462 ( 
.A(n_7000),
.B(n_4587),
.Y(n_7462)
);

INVx1_ASAP7_75t_L g7463 ( 
.A(n_6971),
.Y(n_7463)
);

CKINVDCx5p33_ASAP7_75t_R g7464 ( 
.A(n_7142),
.Y(n_7464)
);

BUFx3_ASAP7_75t_L g7465 ( 
.A(n_7205),
.Y(n_7465)
);

NAND2xp5_ASAP7_75t_L g7466 ( 
.A(n_7003),
.B(n_6800),
.Y(n_7466)
);

BUFx3_ASAP7_75t_L g7467 ( 
.A(n_7206),
.Y(n_7467)
);

CKINVDCx5p33_ASAP7_75t_R g7468 ( 
.A(n_7249),
.Y(n_7468)
);

AND2x2_ASAP7_75t_L g7469 ( 
.A(n_7250),
.B(n_5372),
.Y(n_7469)
);

INVx1_ASAP7_75t_L g7470 ( 
.A(n_6975),
.Y(n_7470)
);

NAND2xp5_ASAP7_75t_L g7471 ( 
.A(n_6842),
.B(n_6983),
.Y(n_7471)
);

INVx1_ASAP7_75t_L g7472 ( 
.A(n_7228),
.Y(n_7472)
);

INVxp67_ASAP7_75t_L g7473 ( 
.A(n_6958),
.Y(n_7473)
);

NAND2xp5_ASAP7_75t_L g7474 ( 
.A(n_7230),
.B(n_4589),
.Y(n_7474)
);

INVx1_ASAP7_75t_L g7475 ( 
.A(n_7236),
.Y(n_7475)
);

INVx1_ASAP7_75t_L g7476 ( 
.A(n_7251),
.Y(n_7476)
);

INVx1_ASAP7_75t_L g7477 ( 
.A(n_7258),
.Y(n_7477)
);

CKINVDCx5p33_ASAP7_75t_R g7478 ( 
.A(n_7211),
.Y(n_7478)
);

NAND2xp5_ASAP7_75t_L g7479 ( 
.A(n_7259),
.B(n_4592),
.Y(n_7479)
);

CKINVDCx5p33_ASAP7_75t_R g7480 ( 
.A(n_7070),
.Y(n_7480)
);

INVx1_ASAP7_75t_L g7481 ( 
.A(n_7270),
.Y(n_7481)
);

CKINVDCx8_ASAP7_75t_R g7482 ( 
.A(n_7277),
.Y(n_7482)
);

INVx3_ASAP7_75t_L g7483 ( 
.A(n_6982),
.Y(n_7483)
);

BUFx2_ASAP7_75t_L g7484 ( 
.A(n_6766),
.Y(n_7484)
);

AND2x6_ASAP7_75t_L g7485 ( 
.A(n_7145),
.B(n_4742),
.Y(n_7485)
);

INVx1_ASAP7_75t_L g7486 ( 
.A(n_7029),
.Y(n_7486)
);

CKINVDCx5p33_ASAP7_75t_R g7487 ( 
.A(n_7127),
.Y(n_7487)
);

INVx2_ASAP7_75t_L g7488 ( 
.A(n_7115),
.Y(n_7488)
);

INVx1_ASAP7_75t_L g7489 ( 
.A(n_7034),
.Y(n_7489)
);

CKINVDCx5p33_ASAP7_75t_R g7490 ( 
.A(n_7152),
.Y(n_7490)
);

INVx2_ASAP7_75t_L g7491 ( 
.A(n_7119),
.Y(n_7491)
);

CKINVDCx5p33_ASAP7_75t_R g7492 ( 
.A(n_7154),
.Y(n_7492)
);

INVx1_ASAP7_75t_L g7493 ( 
.A(n_7039),
.Y(n_7493)
);

NAND2xp5_ASAP7_75t_L g7494 ( 
.A(n_6743),
.B(n_4593),
.Y(n_7494)
);

NAND2xp5_ASAP7_75t_L g7495 ( 
.A(n_6747),
.B(n_6859),
.Y(n_7495)
);

INVx2_ASAP7_75t_L g7496 ( 
.A(n_7122),
.Y(n_7496)
);

INVx1_ASAP7_75t_L g7497 ( 
.A(n_7043),
.Y(n_7497)
);

NAND2xp5_ASAP7_75t_L g7498 ( 
.A(n_6917),
.B(n_4594),
.Y(n_7498)
);

INVx1_ASAP7_75t_L g7499 ( 
.A(n_7044),
.Y(n_7499)
);

INVx2_ASAP7_75t_L g7500 ( 
.A(n_6856),
.Y(n_7500)
);

XOR2xp5_ASAP7_75t_L g7501 ( 
.A(n_6927),
.B(n_5378),
.Y(n_7501)
);

INVx2_ASAP7_75t_L g7502 ( 
.A(n_6862),
.Y(n_7502)
);

INVx1_ASAP7_75t_L g7503 ( 
.A(n_7046),
.Y(n_7503)
);

CKINVDCx5p33_ASAP7_75t_R g7504 ( 
.A(n_7160),
.Y(n_7504)
);

INVx2_ASAP7_75t_L g7505 ( 
.A(n_6889),
.Y(n_7505)
);

NOR2xp33_ASAP7_75t_R g7506 ( 
.A(n_7121),
.B(n_5386),
.Y(n_7506)
);

CKINVDCx5p33_ASAP7_75t_R g7507 ( 
.A(n_7164),
.Y(n_7507)
);

CKINVDCx5p33_ASAP7_75t_R g7508 ( 
.A(n_7173),
.Y(n_7508)
);

CKINVDCx5p33_ASAP7_75t_R g7509 ( 
.A(n_7175),
.Y(n_7509)
);

INVx1_ASAP7_75t_L g7510 ( 
.A(n_7062),
.Y(n_7510)
);

CKINVDCx5p33_ASAP7_75t_R g7511 ( 
.A(n_7185),
.Y(n_7511)
);

INVx1_ASAP7_75t_L g7512 ( 
.A(n_7063),
.Y(n_7512)
);

AND2x4_ASAP7_75t_L g7513 ( 
.A(n_7281),
.B(n_4746),
.Y(n_7513)
);

INVx2_ASAP7_75t_L g7514 ( 
.A(n_6895),
.Y(n_7514)
);

INVx1_ASAP7_75t_L g7515 ( 
.A(n_7064),
.Y(n_7515)
);

INVx1_ASAP7_75t_L g7516 ( 
.A(n_7067),
.Y(n_7516)
);

CKINVDCx5p33_ASAP7_75t_R g7517 ( 
.A(n_7113),
.Y(n_7517)
);

HB1xp67_ASAP7_75t_L g7518 ( 
.A(n_7008),
.Y(n_7518)
);

INVx1_ASAP7_75t_L g7519 ( 
.A(n_7075),
.Y(n_7519)
);

CKINVDCx20_ASAP7_75t_R g7520 ( 
.A(n_6996),
.Y(n_7520)
);

INVx2_ASAP7_75t_L g7521 ( 
.A(n_6896),
.Y(n_7521)
);

CKINVDCx5p33_ASAP7_75t_R g7522 ( 
.A(n_6810),
.Y(n_7522)
);

AND2x2_ASAP7_75t_L g7523 ( 
.A(n_6829),
.B(n_6944),
.Y(n_7523)
);

AND2x2_ASAP7_75t_L g7524 ( 
.A(n_6948),
.B(n_5372),
.Y(n_7524)
);

INVx1_ASAP7_75t_L g7525 ( 
.A(n_7088),
.Y(n_7525)
);

CKINVDCx20_ASAP7_75t_R g7526 ( 
.A(n_6875),
.Y(n_7526)
);

AND2x4_ASAP7_75t_L g7527 ( 
.A(n_6839),
.B(n_4749),
.Y(n_7527)
);

BUFx3_ASAP7_75t_L g7528 ( 
.A(n_7207),
.Y(n_7528)
);

CKINVDCx5p33_ASAP7_75t_R g7529 ( 
.A(n_6888),
.Y(n_7529)
);

CKINVDCx5p33_ASAP7_75t_R g7530 ( 
.A(n_6902),
.Y(n_7530)
);

CKINVDCx5p33_ASAP7_75t_R g7531 ( 
.A(n_7047),
.Y(n_7531)
);

CKINVDCx5p33_ASAP7_75t_R g7532 ( 
.A(n_7061),
.Y(n_7532)
);

CKINVDCx5p33_ASAP7_75t_R g7533 ( 
.A(n_7066),
.Y(n_7533)
);

AND2x2_ASAP7_75t_L g7534 ( 
.A(n_7176),
.B(n_5476),
.Y(n_7534)
);

INVx1_ASAP7_75t_L g7535 ( 
.A(n_7102),
.Y(n_7535)
);

HB1xp67_ASAP7_75t_L g7536 ( 
.A(n_6851),
.Y(n_7536)
);

CKINVDCx5p33_ASAP7_75t_R g7537 ( 
.A(n_7082),
.Y(n_7537)
);

BUFx6f_ASAP7_75t_L g7538 ( 
.A(n_7246),
.Y(n_7538)
);

NAND2xp5_ASAP7_75t_L g7539 ( 
.A(n_6803),
.B(n_4596),
.Y(n_7539)
);

AND2x4_ASAP7_75t_L g7540 ( 
.A(n_7103),
.B(n_4753),
.Y(n_7540)
);

BUFx6f_ASAP7_75t_L g7541 ( 
.A(n_7254),
.Y(n_7541)
);

INVx1_ASAP7_75t_L g7542 ( 
.A(n_7111),
.Y(n_7542)
);

CKINVDCx5p33_ASAP7_75t_R g7543 ( 
.A(n_7108),
.Y(n_7543)
);

INVx1_ASAP7_75t_L g7544 ( 
.A(n_7006),
.Y(n_7544)
);

INVx1_ASAP7_75t_L g7545 ( 
.A(n_7010),
.Y(n_7545)
);

INVx2_ASAP7_75t_L g7546 ( 
.A(n_6901),
.Y(n_7546)
);

CKINVDCx5p33_ASAP7_75t_R g7547 ( 
.A(n_7168),
.Y(n_7547)
);

INVx1_ASAP7_75t_L g7548 ( 
.A(n_7013),
.Y(n_7548)
);

CKINVDCx5p33_ASAP7_75t_R g7549 ( 
.A(n_7216),
.Y(n_7549)
);

INVx1_ASAP7_75t_L g7550 ( 
.A(n_7019),
.Y(n_7550)
);

CKINVDCx5p33_ASAP7_75t_R g7551 ( 
.A(n_7210),
.Y(n_7551)
);

CKINVDCx5p33_ASAP7_75t_R g7552 ( 
.A(n_6779),
.Y(n_7552)
);

INVx1_ASAP7_75t_L g7553 ( 
.A(n_7124),
.Y(n_7553)
);

INVx2_ASAP7_75t_L g7554 ( 
.A(n_6903),
.Y(n_7554)
);

INVx1_ASAP7_75t_L g7555 ( 
.A(n_7112),
.Y(n_7555)
);

CKINVDCx20_ASAP7_75t_R g7556 ( 
.A(n_6897),
.Y(n_7556)
);

INVx1_ASAP7_75t_L g7557 ( 
.A(n_6904),
.Y(n_7557)
);

CKINVDCx5p33_ASAP7_75t_R g7558 ( 
.A(n_6830),
.Y(n_7558)
);

INVx1_ASAP7_75t_L g7559 ( 
.A(n_6921),
.Y(n_7559)
);

INVx1_ASAP7_75t_L g7560 ( 
.A(n_6922),
.Y(n_7560)
);

AND2x4_ASAP7_75t_L g7561 ( 
.A(n_6933),
.B(n_4758),
.Y(n_7561)
);

AND2x2_ASAP7_75t_L g7562 ( 
.A(n_6742),
.B(n_5476),
.Y(n_7562)
);

INVx1_ASAP7_75t_L g7563 ( 
.A(n_6939),
.Y(n_7563)
);

CKINVDCx5p33_ASAP7_75t_R g7564 ( 
.A(n_6936),
.Y(n_7564)
);

INVx2_ASAP7_75t_L g7565 ( 
.A(n_6952),
.Y(n_7565)
);

BUFx2_ASAP7_75t_L g7566 ( 
.A(n_6799),
.Y(n_7566)
);

BUFx6f_ASAP7_75t_L g7567 ( 
.A(n_7272),
.Y(n_7567)
);

INVx1_ASAP7_75t_L g7568 ( 
.A(n_6960),
.Y(n_7568)
);

CKINVDCx5p33_ASAP7_75t_R g7569 ( 
.A(n_6987),
.Y(n_7569)
);

INVx1_ASAP7_75t_L g7570 ( 
.A(n_6961),
.Y(n_7570)
);

CKINVDCx5p33_ASAP7_75t_R g7571 ( 
.A(n_7080),
.Y(n_7571)
);

OA21x2_ASAP7_75t_L g7572 ( 
.A1(n_6840),
.A2(n_4760),
.B(n_4759),
.Y(n_7572)
);

NAND2xp5_ASAP7_75t_L g7573 ( 
.A(n_7017),
.B(n_4597),
.Y(n_7573)
);

CKINVDCx5p33_ASAP7_75t_R g7574 ( 
.A(n_7169),
.Y(n_7574)
);

AND2x2_ASAP7_75t_L g7575 ( 
.A(n_7057),
.B(n_5549),
.Y(n_7575)
);

HB1xp67_ASAP7_75t_L g7576 ( 
.A(n_7009),
.Y(n_7576)
);

INVx1_ASAP7_75t_L g7577 ( 
.A(n_6962),
.Y(n_7577)
);

INVx1_ASAP7_75t_L g7578 ( 
.A(n_6967),
.Y(n_7578)
);

NAND2xp33_ASAP7_75t_R g7579 ( 
.A(n_7130),
.B(n_4599),
.Y(n_7579)
);

CKINVDCx5p33_ASAP7_75t_R g7580 ( 
.A(n_7180),
.Y(n_7580)
);

INVx1_ASAP7_75t_L g7581 ( 
.A(n_6976),
.Y(n_7581)
);

CKINVDCx5p33_ASAP7_75t_R g7582 ( 
.A(n_7199),
.Y(n_7582)
);

NAND2xp5_ASAP7_75t_L g7583 ( 
.A(n_7065),
.B(n_4600),
.Y(n_7583)
);

INVx1_ASAP7_75t_L g7584 ( 
.A(n_6979),
.Y(n_7584)
);

CKINVDCx5p33_ASAP7_75t_R g7585 ( 
.A(n_7190),
.Y(n_7585)
);

NAND2xp5_ASAP7_75t_L g7586 ( 
.A(n_7105),
.B(n_4602),
.Y(n_7586)
);

CKINVDCx5p33_ASAP7_75t_R g7587 ( 
.A(n_7212),
.Y(n_7587)
);

CKINVDCx5p33_ASAP7_75t_R g7588 ( 
.A(n_7215),
.Y(n_7588)
);

INVx2_ASAP7_75t_L g7589 ( 
.A(n_6980),
.Y(n_7589)
);

NAND2xp5_ASAP7_75t_L g7590 ( 
.A(n_7018),
.B(n_4604),
.Y(n_7590)
);

INVx1_ASAP7_75t_L g7591 ( 
.A(n_6981),
.Y(n_7591)
);

INVx1_ASAP7_75t_L g7592 ( 
.A(n_6992),
.Y(n_7592)
);

INVx1_ASAP7_75t_L g7593 ( 
.A(n_6993),
.Y(n_7593)
);

CKINVDCx20_ASAP7_75t_R g7594 ( 
.A(n_6908),
.Y(n_7594)
);

INVx3_ASAP7_75t_L g7595 ( 
.A(n_6984),
.Y(n_7595)
);

INVx2_ASAP7_75t_L g7596 ( 
.A(n_7007),
.Y(n_7596)
);

BUFx8_ASAP7_75t_L g7597 ( 
.A(n_7200),
.Y(n_7597)
);

INVx1_ASAP7_75t_L g7598 ( 
.A(n_7011),
.Y(n_7598)
);

INVx1_ASAP7_75t_SL g7599 ( 
.A(n_6910),
.Y(n_7599)
);

INVx2_ASAP7_75t_L g7600 ( 
.A(n_7022),
.Y(n_7600)
);

INVxp67_ASAP7_75t_L g7601 ( 
.A(n_6963),
.Y(n_7601)
);

INVx3_ASAP7_75t_L g7602 ( 
.A(n_7116),
.Y(n_7602)
);

INVxp67_ASAP7_75t_L g7603 ( 
.A(n_6841),
.Y(n_7603)
);

INVx1_ASAP7_75t_L g7604 ( 
.A(n_7027),
.Y(n_7604)
);

CKINVDCx20_ASAP7_75t_R g7605 ( 
.A(n_7021),
.Y(n_7605)
);

NAND2xp5_ASAP7_75t_L g7606 ( 
.A(n_7020),
.B(n_7146),
.Y(n_7606)
);

INVx1_ASAP7_75t_L g7607 ( 
.A(n_7038),
.Y(n_7607)
);

INVx2_ASAP7_75t_L g7608 ( 
.A(n_7042),
.Y(n_7608)
);

NOR2xp33_ASAP7_75t_L g7609 ( 
.A(n_7150),
.B(n_4605),
.Y(n_7609)
);

CKINVDCx5p33_ASAP7_75t_R g7610 ( 
.A(n_7126),
.Y(n_7610)
);

CKINVDCx5p33_ASAP7_75t_R g7611 ( 
.A(n_7131),
.Y(n_7611)
);

NAND2xp5_ASAP7_75t_SL g7612 ( 
.A(n_6762),
.B(n_4606),
.Y(n_7612)
);

CKINVDCx5p33_ASAP7_75t_R g7613 ( 
.A(n_7156),
.Y(n_7613)
);

INVx2_ASAP7_75t_L g7614 ( 
.A(n_7054),
.Y(n_7614)
);

INVx1_ASAP7_75t_L g7615 ( 
.A(n_7055),
.Y(n_7615)
);

INVx4_ASAP7_75t_L g7616 ( 
.A(n_6807),
.Y(n_7616)
);

INVxp67_ASAP7_75t_L g7617 ( 
.A(n_7196),
.Y(n_7617)
);

INVx1_ASAP7_75t_L g7618 ( 
.A(n_7056),
.Y(n_7618)
);

NAND2xp5_ASAP7_75t_L g7619 ( 
.A(n_6949),
.B(n_4607),
.Y(n_7619)
);

NAND2xp5_ASAP7_75t_L g7620 ( 
.A(n_6991),
.B(n_4608),
.Y(n_7620)
);

CKINVDCx5p33_ASAP7_75t_R g7621 ( 
.A(n_7167),
.Y(n_7621)
);

INVx1_ASAP7_75t_L g7622 ( 
.A(n_7072),
.Y(n_7622)
);

CKINVDCx20_ASAP7_75t_R g7623 ( 
.A(n_7040),
.Y(n_7623)
);

BUFx2_ASAP7_75t_L g7624 ( 
.A(n_6799),
.Y(n_7624)
);

INVx2_ASAP7_75t_L g7625 ( 
.A(n_7079),
.Y(n_7625)
);

CKINVDCx20_ASAP7_75t_R g7626 ( 
.A(n_7092),
.Y(n_7626)
);

NAND2xp5_ASAP7_75t_SL g7627 ( 
.A(n_6989),
.B(n_4611),
.Y(n_7627)
);

INVx2_ASAP7_75t_L g7628 ( 
.A(n_7085),
.Y(n_7628)
);

INVx1_ASAP7_75t_L g7629 ( 
.A(n_6721),
.Y(n_7629)
);

BUFx2_ASAP7_75t_L g7630 ( 
.A(n_6806),
.Y(n_7630)
);

AND2x4_ASAP7_75t_L g7631 ( 
.A(n_6995),
.B(n_6736),
.Y(n_7631)
);

CKINVDCx20_ASAP7_75t_R g7632 ( 
.A(n_7139),
.Y(n_7632)
);

CKINVDCx20_ASAP7_75t_R g7633 ( 
.A(n_6934),
.Y(n_7633)
);

CKINVDCx5p33_ASAP7_75t_R g7634 ( 
.A(n_7184),
.Y(n_7634)
);

HB1xp67_ASAP7_75t_L g7635 ( 
.A(n_7036),
.Y(n_7635)
);

INVx1_ASAP7_75t_L g7636 ( 
.A(n_7222),
.Y(n_7636)
);

BUFx3_ASAP7_75t_L g7637 ( 
.A(n_6876),
.Y(n_7637)
);

INVx1_ASAP7_75t_L g7638 ( 
.A(n_7226),
.Y(n_7638)
);

NOR2xp33_ASAP7_75t_R g7639 ( 
.A(n_7170),
.B(n_5397),
.Y(n_7639)
);

INVx1_ASAP7_75t_L g7640 ( 
.A(n_7231),
.Y(n_7640)
);

INVx1_ASAP7_75t_L g7641 ( 
.A(n_7235),
.Y(n_7641)
);

AND2x4_ASAP7_75t_L g7642 ( 
.A(n_6759),
.B(n_4763),
.Y(n_7642)
);

INVx2_ASAP7_75t_L g7643 ( 
.A(n_6726),
.Y(n_7643)
);

INVx3_ASAP7_75t_L g7644 ( 
.A(n_7120),
.Y(n_7644)
);

CKINVDCx5p33_ASAP7_75t_R g7645 ( 
.A(n_7179),
.Y(n_7645)
);

INVx2_ASAP7_75t_L g7646 ( 
.A(n_6729),
.Y(n_7646)
);

INVx1_ASAP7_75t_L g7647 ( 
.A(n_7237),
.Y(n_7647)
);

INVx1_ASAP7_75t_L g7648 ( 
.A(n_7238),
.Y(n_7648)
);

BUFx3_ASAP7_75t_L g7649 ( 
.A(n_6911),
.Y(n_7649)
);

INVx1_ASAP7_75t_L g7650 ( 
.A(n_7241),
.Y(n_7650)
);

INVx1_ASAP7_75t_L g7651 ( 
.A(n_7244),
.Y(n_7651)
);

CKINVDCx5p33_ASAP7_75t_R g7652 ( 
.A(n_7140),
.Y(n_7652)
);

INVx2_ASAP7_75t_L g7653 ( 
.A(n_6733),
.Y(n_7653)
);

CKINVDCx5p33_ASAP7_75t_R g7654 ( 
.A(n_6973),
.Y(n_7654)
);

AND2x2_ASAP7_75t_L g7655 ( 
.A(n_7128),
.B(n_5549),
.Y(n_7655)
);

AND2x4_ASAP7_75t_L g7656 ( 
.A(n_6765),
.B(n_4765),
.Y(n_7656)
);

XOR2xp5_ASAP7_75t_L g7657 ( 
.A(n_7197),
.B(n_5405),
.Y(n_7657)
);

CKINVDCx5p33_ASAP7_75t_R g7658 ( 
.A(n_6986),
.Y(n_7658)
);

INVxp67_ASAP7_75t_L g7659 ( 
.A(n_7182),
.Y(n_7659)
);

CKINVDCx5p33_ASAP7_75t_R g7660 ( 
.A(n_7058),
.Y(n_7660)
);

INVx1_ASAP7_75t_L g7661 ( 
.A(n_7247),
.Y(n_7661)
);

INVx1_ASAP7_75t_L g7662 ( 
.A(n_7248),
.Y(n_7662)
);

INVx1_ASAP7_75t_L g7663 ( 
.A(n_7252),
.Y(n_7663)
);

INVx3_ASAP7_75t_L g7664 ( 
.A(n_7123),
.Y(n_7664)
);

AND2x2_ASAP7_75t_L g7665 ( 
.A(n_7033),
.B(n_7086),
.Y(n_7665)
);

INVx3_ASAP7_75t_L g7666 ( 
.A(n_7125),
.Y(n_7666)
);

INVx1_ASAP7_75t_L g7667 ( 
.A(n_7253),
.Y(n_7667)
);

CKINVDCx5p33_ASAP7_75t_R g7668 ( 
.A(n_7096),
.Y(n_7668)
);

INVxp67_ASAP7_75t_L g7669 ( 
.A(n_7077),
.Y(n_7669)
);

INVx2_ASAP7_75t_L g7670 ( 
.A(n_7262),
.Y(n_7670)
);

NAND2xp5_ASAP7_75t_L g7671 ( 
.A(n_6861),
.B(n_4613),
.Y(n_7671)
);

HB1xp67_ASAP7_75t_L g7672 ( 
.A(n_7129),
.Y(n_7672)
);

INVx1_ASAP7_75t_L g7673 ( 
.A(n_7271),
.Y(n_7673)
);

NAND2xp5_ASAP7_75t_L g7674 ( 
.A(n_6861),
.B(n_7276),
.Y(n_7674)
);

NOR2xp33_ASAP7_75t_R g7675 ( 
.A(n_7213),
.B(n_5435),
.Y(n_7675)
);

CKINVDCx5p33_ASAP7_75t_R g7676 ( 
.A(n_6783),
.Y(n_7676)
);

CKINVDCx5p33_ASAP7_75t_R g7677 ( 
.A(n_7074),
.Y(n_7677)
);

INVx2_ASAP7_75t_L g7678 ( 
.A(n_7283),
.Y(n_7678)
);

BUFx2_ASAP7_75t_L g7679 ( 
.A(n_6806),
.Y(n_7679)
);

HB1xp67_ASAP7_75t_L g7680 ( 
.A(n_7114),
.Y(n_7680)
);

INVx2_ASAP7_75t_L g7681 ( 
.A(n_7284),
.Y(n_7681)
);

AND2x4_ASAP7_75t_L g7682 ( 
.A(n_6793),
.B(n_4776),
.Y(n_7682)
);

CKINVDCx5p33_ASAP7_75t_R g7683 ( 
.A(n_7159),
.Y(n_7683)
);

BUFx6f_ASAP7_75t_L g7684 ( 
.A(n_7275),
.Y(n_7684)
);

AND2x4_ASAP7_75t_L g7685 ( 
.A(n_6804),
.B(n_6790),
.Y(n_7685)
);

CKINVDCx5p33_ASAP7_75t_R g7686 ( 
.A(n_7161),
.Y(n_7686)
);

CKINVDCx5p33_ASAP7_75t_R g7687 ( 
.A(n_7163),
.Y(n_7687)
);

INVx1_ASAP7_75t_L g7688 ( 
.A(n_7289),
.Y(n_7688)
);

INVx2_ASAP7_75t_L g7689 ( 
.A(n_7297),
.Y(n_7689)
);

INVx1_ASAP7_75t_L g7690 ( 
.A(n_6752),
.Y(n_7690)
);

CKINVDCx20_ASAP7_75t_R g7691 ( 
.A(n_7201),
.Y(n_7691)
);

INVx2_ASAP7_75t_L g7692 ( 
.A(n_6877),
.Y(n_7692)
);

CKINVDCx5p33_ASAP7_75t_R g7693 ( 
.A(n_7181),
.Y(n_7693)
);

NOR2xp67_ASAP7_75t_L g7694 ( 
.A(n_6749),
.B(n_4281),
.Y(n_7694)
);

INVx2_ASAP7_75t_L g7695 ( 
.A(n_6883),
.Y(n_7695)
);

BUFx3_ASAP7_75t_L g7696 ( 
.A(n_7278),
.Y(n_7696)
);

CKINVDCx5p33_ASAP7_75t_R g7697 ( 
.A(n_7186),
.Y(n_7697)
);

OAI22xp5_ASAP7_75t_L g7698 ( 
.A1(n_6826),
.A2(n_4615),
.B1(n_4618),
.B2(n_4614),
.Y(n_7698)
);

CKINVDCx5p33_ASAP7_75t_R g7699 ( 
.A(n_7147),
.Y(n_7699)
);

INVx1_ASAP7_75t_L g7700 ( 
.A(n_7049),
.Y(n_7700)
);

INVx4_ASAP7_75t_L g7701 ( 
.A(n_6999),
.Y(n_7701)
);

CKINVDCx16_ASAP7_75t_R g7702 ( 
.A(n_7071),
.Y(n_7702)
);

INVx1_ASAP7_75t_L g7703 ( 
.A(n_7050),
.Y(n_7703)
);

INVx1_ASAP7_75t_L g7704 ( 
.A(n_7068),
.Y(n_7704)
);

CKINVDCx5p33_ASAP7_75t_R g7705 ( 
.A(n_7153),
.Y(n_7705)
);

NAND2xp5_ASAP7_75t_L g7706 ( 
.A(n_6728),
.B(n_6916),
.Y(n_7706)
);

NAND2xp5_ASAP7_75t_L g7707 ( 
.A(n_7023),
.B(n_4621),
.Y(n_7707)
);

INVx1_ASAP7_75t_L g7708 ( 
.A(n_6757),
.Y(n_7708)
);

INVx2_ASAP7_75t_L g7709 ( 
.A(n_6885),
.Y(n_7709)
);

BUFx2_ASAP7_75t_L g7710 ( 
.A(n_7041),
.Y(n_7710)
);

NAND2xp5_ASAP7_75t_L g7711 ( 
.A(n_7051),
.B(n_4626),
.Y(n_7711)
);

INVx2_ASAP7_75t_L g7712 ( 
.A(n_6905),
.Y(n_7712)
);

INVx4_ASAP7_75t_L g7713 ( 
.A(n_7014),
.Y(n_7713)
);

NOR2xp33_ASAP7_75t_L g7714 ( 
.A(n_7192),
.B(n_4627),
.Y(n_7714)
);

INVx1_ASAP7_75t_L g7715 ( 
.A(n_6798),
.Y(n_7715)
);

INVx3_ASAP7_75t_L g7716 ( 
.A(n_7279),
.Y(n_7716)
);

CKINVDCx5p33_ASAP7_75t_R g7717 ( 
.A(n_7132),
.Y(n_7717)
);

CKINVDCx5p33_ASAP7_75t_R g7718 ( 
.A(n_7134),
.Y(n_7718)
);

CKINVDCx5p33_ASAP7_75t_R g7719 ( 
.A(n_7137),
.Y(n_7719)
);

NAND2xp33_ASAP7_75t_SL g7720 ( 
.A(n_7194),
.B(n_5440),
.Y(n_7720)
);

INVx1_ASAP7_75t_L g7721 ( 
.A(n_6815),
.Y(n_7721)
);

INVx3_ASAP7_75t_L g7722 ( 
.A(n_7291),
.Y(n_7722)
);

INVx3_ASAP7_75t_L g7723 ( 
.A(n_7294),
.Y(n_7723)
);

INVx1_ASAP7_75t_L g7724 ( 
.A(n_6872),
.Y(n_7724)
);

INVx1_ASAP7_75t_L g7725 ( 
.A(n_6920),
.Y(n_7725)
);

INVx1_ASAP7_75t_L g7726 ( 
.A(n_6930),
.Y(n_7726)
);

INVx1_ASAP7_75t_L g7727 ( 
.A(n_6972),
.Y(n_7727)
);

INVx1_ASAP7_75t_L g7728 ( 
.A(n_6974),
.Y(n_7728)
);

NAND2x1_ASAP7_75t_L g7729 ( 
.A(n_6985),
.B(n_4783),
.Y(n_7729)
);

AND2x4_ASAP7_75t_L g7730 ( 
.A(n_6792),
.B(n_7073),
.Y(n_7730)
);

CKINVDCx5p33_ASAP7_75t_R g7731 ( 
.A(n_7138),
.Y(n_7731)
);

AND2x2_ASAP7_75t_L g7732 ( 
.A(n_6727),
.B(n_5588),
.Y(n_7732)
);

CKINVDCx20_ASAP7_75t_R g7733 ( 
.A(n_6873),
.Y(n_7733)
);

CKINVDCx20_ASAP7_75t_R g7734 ( 
.A(n_7025),
.Y(n_7734)
);

AND2x2_ASAP7_75t_L g7735 ( 
.A(n_7117),
.B(n_6745),
.Y(n_7735)
);

INVx1_ASAP7_75t_L g7736 ( 
.A(n_6990),
.Y(n_7736)
);

CKINVDCx5p33_ASAP7_75t_R g7737 ( 
.A(n_7144),
.Y(n_7737)
);

NAND2xp5_ASAP7_75t_L g7738 ( 
.A(n_7106),
.B(n_4629),
.Y(n_7738)
);

BUFx8_ASAP7_75t_L g7739 ( 
.A(n_7188),
.Y(n_7739)
);

INVx2_ASAP7_75t_L g7740 ( 
.A(n_6906),
.Y(n_7740)
);

AND2x6_ASAP7_75t_L g7741 ( 
.A(n_7155),
.B(n_4786),
.Y(n_7741)
);

CKINVDCx5p33_ASAP7_75t_R g7742 ( 
.A(n_7165),
.Y(n_7742)
);

CKINVDCx5p33_ASAP7_75t_R g7743 ( 
.A(n_7171),
.Y(n_7743)
);

INVxp67_ASAP7_75t_L g7744 ( 
.A(n_7143),
.Y(n_7744)
);

BUFx6f_ASAP7_75t_L g7745 ( 
.A(n_7295),
.Y(n_7745)
);

INVx1_ASAP7_75t_L g7746 ( 
.A(n_7001),
.Y(n_7746)
);

INVx2_ASAP7_75t_SL g7747 ( 
.A(n_6760),
.Y(n_7747)
);

INVx1_ASAP7_75t_L g7748 ( 
.A(n_7012),
.Y(n_7748)
);

CKINVDCx5p33_ASAP7_75t_R g7749 ( 
.A(n_7174),
.Y(n_7749)
);

INVx1_ASAP7_75t_L g7750 ( 
.A(n_7219),
.Y(n_7750)
);

INVxp67_ASAP7_75t_L g7751 ( 
.A(n_7189),
.Y(n_7751)
);

INVx1_ASAP7_75t_L g7752 ( 
.A(n_7255),
.Y(n_7752)
);

BUFx2_ASAP7_75t_SL g7753 ( 
.A(n_7204),
.Y(n_7753)
);

INVx2_ASAP7_75t_L g7754 ( 
.A(n_6924),
.Y(n_7754)
);

CKINVDCx20_ASAP7_75t_R g7755 ( 
.A(n_7093),
.Y(n_7755)
);

CKINVDCx20_ASAP7_75t_R g7756 ( 
.A(n_7148),
.Y(n_7756)
);

INVx1_ASAP7_75t_L g7757 ( 
.A(n_7260),
.Y(n_7757)
);

CKINVDCx5p33_ASAP7_75t_R g7758 ( 
.A(n_7177),
.Y(n_7758)
);

AND2x6_ASAP7_75t_L g7759 ( 
.A(n_7178),
.B(n_4795),
.Y(n_7759)
);

INVx2_ASAP7_75t_L g7760 ( 
.A(n_6928),
.Y(n_7760)
);

INVx2_ASAP7_75t_L g7761 ( 
.A(n_6935),
.Y(n_7761)
);

INVx2_ASAP7_75t_L g7762 ( 
.A(n_6943),
.Y(n_7762)
);

INVx2_ASAP7_75t_L g7763 ( 
.A(n_6953),
.Y(n_7763)
);

INVx1_ASAP7_75t_SL g7764 ( 
.A(n_6868),
.Y(n_7764)
);

INVx1_ASAP7_75t_L g7765 ( 
.A(n_7264),
.Y(n_7765)
);

CKINVDCx5p33_ASAP7_75t_R g7766 ( 
.A(n_7187),
.Y(n_7766)
);

INVx1_ASAP7_75t_L g7767 ( 
.A(n_6758),
.Y(n_7767)
);

INVx1_ASAP7_75t_L g7768 ( 
.A(n_6772),
.Y(n_7768)
);

NAND2xp5_ASAP7_75t_SL g7769 ( 
.A(n_6836),
.B(n_4631),
.Y(n_7769)
);

NOR2xp67_ASAP7_75t_L g7770 ( 
.A(n_7166),
.B(n_4282),
.Y(n_7770)
);

INVx2_ASAP7_75t_L g7771 ( 
.A(n_6718),
.Y(n_7771)
);

INVx1_ASAP7_75t_L g7772 ( 
.A(n_6805),
.Y(n_7772)
);

NAND2xp5_ASAP7_75t_L g7773 ( 
.A(n_6771),
.B(n_4632),
.Y(n_7773)
);

CKINVDCx5p33_ASAP7_75t_R g7774 ( 
.A(n_7028),
.Y(n_7774)
);

INVx3_ASAP7_75t_L g7775 ( 
.A(n_6816),
.Y(n_7775)
);

INVx1_ASAP7_75t_L g7776 ( 
.A(n_6827),
.Y(n_7776)
);

INVx1_ASAP7_75t_L g7777 ( 
.A(n_6878),
.Y(n_7777)
);

NOR2xp33_ASAP7_75t_L g7778 ( 
.A(n_7288),
.B(n_4636),
.Y(n_7778)
);

CKINVDCx5p33_ASAP7_75t_R g7779 ( 
.A(n_7208),
.Y(n_7779)
);

INVx1_ASAP7_75t_L g7780 ( 
.A(n_6887),
.Y(n_7780)
);

CKINVDCx5p33_ASAP7_75t_R g7781 ( 
.A(n_7209),
.Y(n_7781)
);

NOR2xp33_ASAP7_75t_L g7782 ( 
.A(n_7292),
.B(n_4638),
.Y(n_7782)
);

INVx1_ASAP7_75t_L g7783 ( 
.A(n_6891),
.Y(n_7783)
);

INVxp67_ASAP7_75t_SL g7784 ( 
.A(n_7218),
.Y(n_7784)
);

INVx2_ASAP7_75t_L g7785 ( 
.A(n_7221),
.Y(n_7785)
);

INVx1_ASAP7_75t_L g7786 ( 
.A(n_6923),
.Y(n_7786)
);

CKINVDCx20_ASAP7_75t_R g7787 ( 
.A(n_7202),
.Y(n_7787)
);

NAND2xp5_ASAP7_75t_L g7788 ( 
.A(n_6818),
.B(n_4639),
.Y(n_7788)
);

BUFx6f_ASAP7_75t_L g7789 ( 
.A(n_6820),
.Y(n_7789)
);

BUFx6f_ASAP7_75t_L g7790 ( 
.A(n_6828),
.Y(n_7790)
);

INVx1_ASAP7_75t_L g7791 ( 
.A(n_6941),
.Y(n_7791)
);

INVx3_ASAP7_75t_L g7792 ( 
.A(n_6834),
.Y(n_7792)
);

CKINVDCx20_ASAP7_75t_R g7793 ( 
.A(n_7203),
.Y(n_7793)
);

INVx2_ASAP7_75t_L g7794 ( 
.A(n_7261),
.Y(n_7794)
);

NAND2xp5_ASAP7_75t_SL g7795 ( 
.A(n_6844),
.B(n_4640),
.Y(n_7795)
);

AOI22xp5_ASAP7_75t_L g7796 ( 
.A1(n_6819),
.A2(n_5465),
.B1(n_5479),
.B2(n_5456),
.Y(n_7796)
);

NAND2xp5_ASAP7_75t_L g7797 ( 
.A(n_6822),
.B(n_4641),
.Y(n_7797)
);

INVx1_ASAP7_75t_L g7798 ( 
.A(n_6946),
.Y(n_7798)
);

NAND2xp33_ASAP7_75t_R g7799 ( 
.A(n_6797),
.B(n_7214),
.Y(n_7799)
);

INVx2_ASAP7_75t_L g7800 ( 
.A(n_7296),
.Y(n_7800)
);

INVx1_ASAP7_75t_L g7801 ( 
.A(n_6969),
.Y(n_7801)
);

CKINVDCx20_ASAP7_75t_R g7802 ( 
.A(n_6785),
.Y(n_7802)
);

INVx2_ASAP7_75t_L g7803 ( 
.A(n_6754),
.Y(n_7803)
);

CKINVDCx5p33_ASAP7_75t_R g7804 ( 
.A(n_7183),
.Y(n_7804)
);

OAI22xp5_ASAP7_75t_SL g7805 ( 
.A1(n_6720),
.A2(n_5494),
.B1(n_5499),
.B2(n_5485),
.Y(n_7805)
);

INVx1_ASAP7_75t_L g7806 ( 
.A(n_7026),
.Y(n_7806)
);

AND2x4_ASAP7_75t_L g7807 ( 
.A(n_6850),
.B(n_4797),
.Y(n_7807)
);

CKINVDCx5p33_ASAP7_75t_R g7808 ( 
.A(n_7183),
.Y(n_7808)
);

BUFx6f_ASAP7_75t_L g7809 ( 
.A(n_6854),
.Y(n_7809)
);

INVx1_ASAP7_75t_L g7810 ( 
.A(n_7030),
.Y(n_7810)
);

AND2x2_ASAP7_75t_L g7811 ( 
.A(n_6832),
.B(n_6849),
.Y(n_7811)
);

CKINVDCx5p33_ASAP7_75t_R g7812 ( 
.A(n_7097),
.Y(n_7812)
);

INVx2_ASAP7_75t_L g7813 ( 
.A(n_7024),
.Y(n_7813)
);

CKINVDCx5p33_ASAP7_75t_R g7814 ( 
.A(n_7198),
.Y(n_7814)
);

INVx1_ASAP7_75t_L g7815 ( 
.A(n_7110),
.Y(n_7815)
);

INVx1_ASAP7_75t_L g7816 ( 
.A(n_7048),
.Y(n_7816)
);

INVx1_ASAP7_75t_L g7817 ( 
.A(n_7037),
.Y(n_7817)
);

INVx1_ASAP7_75t_L g7818 ( 
.A(n_7053),
.Y(n_7818)
);

INVx1_ASAP7_75t_L g7819 ( 
.A(n_7076),
.Y(n_7819)
);

INVx1_ASAP7_75t_L g7820 ( 
.A(n_7081),
.Y(n_7820)
);

HB1xp67_ASAP7_75t_L g7821 ( 
.A(n_6919),
.Y(n_7821)
);

BUFx2_ASAP7_75t_L g7822 ( 
.A(n_7041),
.Y(n_7822)
);

NAND2x1_ASAP7_75t_L g7823 ( 
.A(n_7286),
.B(n_4803),
.Y(n_7823)
);

INVx1_ASAP7_75t_L g7824 ( 
.A(n_7083),
.Y(n_7824)
);

CKINVDCx20_ASAP7_75t_R g7825 ( 
.A(n_7280),
.Y(n_7825)
);

CKINVDCx5p33_ASAP7_75t_R g7826 ( 
.A(n_6959),
.Y(n_7826)
);

AND2x2_ASAP7_75t_SL g7827 ( 
.A(n_6864),
.B(n_5289),
.Y(n_7827)
);

BUFx6f_ASAP7_75t_L g7828 ( 
.A(n_6855),
.Y(n_7828)
);

NAND2x1_ASAP7_75t_L g7829 ( 
.A(n_7286),
.B(n_4805),
.Y(n_7829)
);

INVx1_ASAP7_75t_L g7830 ( 
.A(n_7084),
.Y(n_7830)
);

NAND2xp5_ASAP7_75t_L g7831 ( 
.A(n_6988),
.B(n_4643),
.Y(n_7831)
);

AND2x2_ASAP7_75t_L g7832 ( 
.A(n_6884),
.B(n_5588),
.Y(n_7832)
);

INVx3_ASAP7_75t_L g7833 ( 
.A(n_6857),
.Y(n_7833)
);

CKINVDCx5p33_ASAP7_75t_R g7834 ( 
.A(n_7118),
.Y(n_7834)
);

INVx1_ASAP7_75t_L g7835 ( 
.A(n_7087),
.Y(n_7835)
);

INVx4_ASAP7_75t_L g7836 ( 
.A(n_7089),
.Y(n_7836)
);

CKINVDCx5p33_ASAP7_75t_R g7837 ( 
.A(n_7016),
.Y(n_7837)
);

AND2x4_ASAP7_75t_L g7838 ( 
.A(n_6866),
.B(n_4807),
.Y(n_7838)
);

INVx2_ASAP7_75t_L g7839 ( 
.A(n_7094),
.Y(n_7839)
);

INVx1_ASAP7_75t_L g7840 ( 
.A(n_6951),
.Y(n_7840)
);

INVx1_ASAP7_75t_L g7841 ( 
.A(n_6881),
.Y(n_7841)
);

CKINVDCx5p33_ASAP7_75t_R g7842 ( 
.A(n_7052),
.Y(n_7842)
);

CKINVDCx20_ASAP7_75t_R g7843 ( 
.A(n_7133),
.Y(n_7843)
);

CKINVDCx5p33_ASAP7_75t_R g7844 ( 
.A(n_7032),
.Y(n_7844)
);

INVx2_ASAP7_75t_L g7845 ( 
.A(n_6886),
.Y(n_7845)
);

BUFx8_ASAP7_75t_L g7846 ( 
.A(n_6938),
.Y(n_7846)
);

INVx1_ASAP7_75t_L g7847 ( 
.A(n_6912),
.Y(n_7847)
);

NAND2xp5_ASAP7_75t_L g7848 ( 
.A(n_7162),
.B(n_4644),
.Y(n_7848)
);

CKINVDCx5p33_ASAP7_75t_R g7849 ( 
.A(n_6737),
.Y(n_7849)
);

CKINVDCx5p33_ASAP7_75t_R g7850 ( 
.A(n_6735),
.Y(n_7850)
);

CKINVDCx5p33_ASAP7_75t_R g7851 ( 
.A(n_6724),
.Y(n_7851)
);

NAND2xp5_ASAP7_75t_SL g7852 ( 
.A(n_7098),
.B(n_4646),
.Y(n_7852)
);

OAI21x1_ASAP7_75t_L g7853 ( 
.A1(n_7191),
.A2(n_5394),
.B(n_5318),
.Y(n_7853)
);

CKINVDCx5p33_ASAP7_75t_R g7854 ( 
.A(n_6929),
.Y(n_7854)
);

CKINVDCx5p33_ASAP7_75t_R g7855 ( 
.A(n_7069),
.Y(n_7855)
);

AND2x4_ASAP7_75t_L g7856 ( 
.A(n_6918),
.B(n_4809),
.Y(n_7856)
);

CKINVDCx5p33_ASAP7_75t_R g7857 ( 
.A(n_7045),
.Y(n_7857)
);

NAND2xp5_ASAP7_75t_L g7858 ( 
.A(n_6774),
.B(n_4647),
.Y(n_7858)
);

CKINVDCx5p33_ASAP7_75t_R g7859 ( 
.A(n_6753),
.Y(n_7859)
);

NAND2xp5_ASAP7_75t_L g7860 ( 
.A(n_7349),
.B(n_6794),
.Y(n_7860)
);

INVx2_ASAP7_75t_L g7861 ( 
.A(n_7308),
.Y(n_7861)
);

NOR2xp33_ASAP7_75t_L g7862 ( 
.A(n_7601),
.B(n_6964),
.Y(n_7862)
);

INVx1_ASAP7_75t_L g7863 ( 
.A(n_7299),
.Y(n_7863)
);

INVx3_ASAP7_75t_L g7864 ( 
.A(n_7789),
.Y(n_7864)
);

INVx2_ASAP7_75t_L g7865 ( 
.A(n_7310),
.Y(n_7865)
);

INVx2_ASAP7_75t_L g7866 ( 
.A(n_7312),
.Y(n_7866)
);

INVx4_ASAP7_75t_L g7867 ( 
.A(n_7487),
.Y(n_7867)
);

NAND3xp33_ASAP7_75t_L g7868 ( 
.A(n_7398),
.B(n_6950),
.C(n_6890),
.Y(n_7868)
);

INVx1_ASAP7_75t_L g7869 ( 
.A(n_7303),
.Y(n_7869)
);

INVx5_ASAP7_75t_L g7870 ( 
.A(n_7454),
.Y(n_7870)
);

INVx2_ASAP7_75t_L g7871 ( 
.A(n_7317),
.Y(n_7871)
);

BUFx2_ASAP7_75t_L g7872 ( 
.A(n_7309),
.Y(n_7872)
);

AOI22x1_ASAP7_75t_L g7873 ( 
.A1(n_7708),
.A2(n_6931),
.B1(n_6937),
.B2(n_6926),
.Y(n_7873)
);

INVx1_ASAP7_75t_L g7874 ( 
.A(n_7304),
.Y(n_7874)
);

INVx3_ASAP7_75t_L g7875 ( 
.A(n_7789),
.Y(n_7875)
);

INVx2_ASAP7_75t_L g7876 ( 
.A(n_7320),
.Y(n_7876)
);

INVx2_ASAP7_75t_L g7877 ( 
.A(n_7323),
.Y(n_7877)
);

NOR2xp33_ASAP7_75t_L g7878 ( 
.A(n_7699),
.B(n_5513),
.Y(n_7878)
);

INVx2_ASAP7_75t_L g7879 ( 
.A(n_7381),
.Y(n_7879)
);

INVx2_ASAP7_75t_L g7880 ( 
.A(n_7389),
.Y(n_7880)
);

INVx1_ASAP7_75t_L g7881 ( 
.A(n_7319),
.Y(n_7881)
);

NAND2xp33_ASAP7_75t_L g7882 ( 
.A(n_7552),
.B(n_6940),
.Y(n_7882)
);

INVx1_ASAP7_75t_L g7883 ( 
.A(n_7322),
.Y(n_7883)
);

INVx1_ASAP7_75t_L g7884 ( 
.A(n_7324),
.Y(n_7884)
);

BUFx3_ASAP7_75t_L g7885 ( 
.A(n_7465),
.Y(n_7885)
);

INVx2_ASAP7_75t_SL g7886 ( 
.A(n_7305),
.Y(n_7886)
);

INVx1_ASAP7_75t_L g7887 ( 
.A(n_7329),
.Y(n_7887)
);

CKINVDCx16_ASAP7_75t_R g7888 ( 
.A(n_7506),
.Y(n_7888)
);

INVx2_ASAP7_75t_L g7889 ( 
.A(n_7393),
.Y(n_7889)
);

NAND2xp5_ASAP7_75t_SL g7890 ( 
.A(n_7523),
.B(n_6945),
.Y(n_7890)
);

INVxp33_ASAP7_75t_L g7891 ( 
.A(n_7313),
.Y(n_7891)
);

INVx4_ASAP7_75t_L g7892 ( 
.A(n_7490),
.Y(n_7892)
);

AND2x2_ASAP7_75t_L g7893 ( 
.A(n_7665),
.B(n_6956),
.Y(n_7893)
);

AOI22xp33_ASAP7_75t_L g7894 ( 
.A1(n_7782),
.A2(n_5518),
.B1(n_5540),
.B2(n_5516),
.Y(n_7894)
);

AO21x2_ASAP7_75t_L g7895 ( 
.A1(n_7715),
.A2(n_4813),
.B(n_4810),
.Y(n_7895)
);

INVx2_ASAP7_75t_L g7896 ( 
.A(n_7407),
.Y(n_7896)
);

INVx1_ASAP7_75t_SL g7897 ( 
.A(n_7328),
.Y(n_7897)
);

INVx2_ASAP7_75t_SL g7898 ( 
.A(n_7341),
.Y(n_7898)
);

NAND2xp5_ASAP7_75t_L g7899 ( 
.A(n_7806),
.B(n_4648),
.Y(n_7899)
);

AND2x6_ASAP7_75t_L g7900 ( 
.A(n_7810),
.B(n_4815),
.Y(n_7900)
);

INVx2_ASAP7_75t_L g7901 ( 
.A(n_7418),
.Y(n_7901)
);

INVx4_ASAP7_75t_L g7902 ( 
.A(n_7492),
.Y(n_7902)
);

INVx2_ASAP7_75t_L g7903 ( 
.A(n_7426),
.Y(n_7903)
);

INVx1_ASAP7_75t_L g7904 ( 
.A(n_7332),
.Y(n_7904)
);

HB1xp67_ASAP7_75t_L g7905 ( 
.A(n_7383),
.Y(n_7905)
);

INVx2_ASAP7_75t_L g7906 ( 
.A(n_7431),
.Y(n_7906)
);

INVx2_ASAP7_75t_L g7907 ( 
.A(n_7433),
.Y(n_7907)
);

INVx2_ASAP7_75t_L g7908 ( 
.A(n_7442),
.Y(n_7908)
);

INVx1_ASAP7_75t_L g7909 ( 
.A(n_7333),
.Y(n_7909)
);

AND2x4_ASAP7_75t_L g7910 ( 
.A(n_7467),
.B(n_4819),
.Y(n_7910)
);

NAND2xp5_ASAP7_75t_SL g7911 ( 
.A(n_7827),
.B(n_5575),
.Y(n_7911)
);

AOI22xp5_ASAP7_75t_L g7912 ( 
.A1(n_7815),
.A2(n_5667),
.B1(n_5700),
.B2(n_5607),
.Y(n_7912)
);

INVx2_ASAP7_75t_L g7913 ( 
.A(n_7444),
.Y(n_7913)
);

BUFx6f_ASAP7_75t_L g7914 ( 
.A(n_7331),
.Y(n_7914)
);

AOI21x1_ASAP7_75t_L g7915 ( 
.A1(n_7606),
.A2(n_4840),
.B(n_4838),
.Y(n_7915)
);

INVx2_ASAP7_75t_L g7916 ( 
.A(n_7340),
.Y(n_7916)
);

INVx3_ASAP7_75t_L g7917 ( 
.A(n_7790),
.Y(n_7917)
);

INVxp33_ASAP7_75t_L g7918 ( 
.A(n_7307),
.Y(n_7918)
);

INVx2_ASAP7_75t_L g7919 ( 
.A(n_7350),
.Y(n_7919)
);

INVx2_ASAP7_75t_L g7920 ( 
.A(n_7360),
.Y(n_7920)
);

NOR2x1p5_ASAP7_75t_L g7921 ( 
.A(n_7457),
.B(n_4650),
.Y(n_7921)
);

INVx2_ASAP7_75t_L g7922 ( 
.A(n_7364),
.Y(n_7922)
);

BUFx6f_ASAP7_75t_SL g7923 ( 
.A(n_7637),
.Y(n_7923)
);

INVx2_ASAP7_75t_L g7924 ( 
.A(n_7369),
.Y(n_7924)
);

NAND2xp5_ASAP7_75t_L g7925 ( 
.A(n_7750),
.B(n_4652),
.Y(n_7925)
);

INVx2_ASAP7_75t_L g7926 ( 
.A(n_7371),
.Y(n_7926)
);

INVx1_ASAP7_75t_L g7927 ( 
.A(n_7372),
.Y(n_7927)
);

NAND2xp5_ASAP7_75t_L g7928 ( 
.A(n_7752),
.B(n_7757),
.Y(n_7928)
);

NAND2xp33_ASAP7_75t_L g7929 ( 
.A(n_7558),
.B(n_4654),
.Y(n_7929)
);

INVx2_ASAP7_75t_L g7930 ( 
.A(n_7374),
.Y(n_7930)
);

INVx1_ASAP7_75t_L g7931 ( 
.A(n_7375),
.Y(n_7931)
);

INVx1_ASAP7_75t_L g7932 ( 
.A(n_7385),
.Y(n_7932)
);

INVx1_ASAP7_75t_L g7933 ( 
.A(n_7392),
.Y(n_7933)
);

INVx2_ASAP7_75t_L g7934 ( 
.A(n_7400),
.Y(n_7934)
);

AOI22xp33_ASAP7_75t_L g7935 ( 
.A1(n_7778),
.A2(n_5751),
.B1(n_5718),
.B2(n_5418),
.Y(n_7935)
);

INVx2_ASAP7_75t_L g7936 ( 
.A(n_7401),
.Y(n_7936)
);

BUFx3_ASAP7_75t_L g7937 ( 
.A(n_7528),
.Y(n_7937)
);

INVx2_ASAP7_75t_L g7938 ( 
.A(n_7403),
.Y(n_7938)
);

INVx2_ASAP7_75t_L g7939 ( 
.A(n_7405),
.Y(n_7939)
);

BUFx10_ASAP7_75t_L g7940 ( 
.A(n_7365),
.Y(n_7940)
);

BUFx3_ASAP7_75t_L g7941 ( 
.A(n_7318),
.Y(n_7941)
);

INVx2_ASAP7_75t_L g7942 ( 
.A(n_7421),
.Y(n_7942)
);

NAND2xp5_ASAP7_75t_L g7943 ( 
.A(n_7765),
.B(n_4655),
.Y(n_7943)
);

NAND2xp5_ASAP7_75t_L g7944 ( 
.A(n_7495),
.B(n_7466),
.Y(n_7944)
);

INVx3_ASAP7_75t_L g7945 ( 
.A(n_7790),
.Y(n_7945)
);

NOR2xp33_ASAP7_75t_L g7946 ( 
.A(n_7705),
.B(n_4656),
.Y(n_7946)
);

INVx3_ASAP7_75t_L g7947 ( 
.A(n_7809),
.Y(n_7947)
);

INVx1_ASAP7_75t_L g7948 ( 
.A(n_7425),
.Y(n_7948)
);

AND3x2_ASAP7_75t_L g7949 ( 
.A(n_7484),
.B(n_4844),
.C(n_4843),
.Y(n_7949)
);

INVx5_ASAP7_75t_L g7950 ( 
.A(n_7365),
.Y(n_7950)
);

INVx1_ASAP7_75t_L g7951 ( 
.A(n_7432),
.Y(n_7951)
);

AOI22xp33_ASAP7_75t_L g7952 ( 
.A1(n_7721),
.A2(n_5436),
.B1(n_5453),
.B2(n_5411),
.Y(n_7952)
);

INVx2_ASAP7_75t_L g7953 ( 
.A(n_7434),
.Y(n_7953)
);

INVx2_ASAP7_75t_L g7954 ( 
.A(n_7439),
.Y(n_7954)
);

INVx1_ASAP7_75t_L g7955 ( 
.A(n_7441),
.Y(n_7955)
);

INVx4_ASAP7_75t_L g7956 ( 
.A(n_7504),
.Y(n_7956)
);

INVx2_ASAP7_75t_L g7957 ( 
.A(n_7446),
.Y(n_7957)
);

INVx2_ASAP7_75t_L g7958 ( 
.A(n_7447),
.Y(n_7958)
);

INVx2_ASAP7_75t_L g7959 ( 
.A(n_7449),
.Y(n_7959)
);

INVxp33_ASAP7_75t_SL g7960 ( 
.A(n_7585),
.Y(n_7960)
);

NAND2xp5_ASAP7_75t_SL g7961 ( 
.A(n_7683),
.B(n_7686),
.Y(n_7961)
);

NAND2xp5_ASAP7_75t_SL g7962 ( 
.A(n_7687),
.B(n_4657),
.Y(n_7962)
);

INVx2_ASAP7_75t_L g7963 ( 
.A(n_7452),
.Y(n_7963)
);

INVx1_ASAP7_75t_L g7964 ( 
.A(n_7458),
.Y(n_7964)
);

INVx2_ASAP7_75t_SL g7965 ( 
.A(n_7387),
.Y(n_7965)
);

AND2x2_ASAP7_75t_SL g7966 ( 
.A(n_7702),
.B(n_7413),
.Y(n_7966)
);

CKINVDCx6p67_ASAP7_75t_R g7967 ( 
.A(n_7326),
.Y(n_7967)
);

INVx2_ASAP7_75t_L g7968 ( 
.A(n_7463),
.Y(n_7968)
);

INVx1_ASAP7_75t_L g7969 ( 
.A(n_7470),
.Y(n_7969)
);

INVx2_ASAP7_75t_L g7970 ( 
.A(n_7472),
.Y(n_7970)
);

INVx2_ASAP7_75t_L g7971 ( 
.A(n_7475),
.Y(n_7971)
);

NAND2xp5_ASAP7_75t_SL g7972 ( 
.A(n_7693),
.B(n_4658),
.Y(n_7972)
);

INVx2_ASAP7_75t_SL g7973 ( 
.A(n_7518),
.Y(n_7973)
);

NAND2xp5_ASAP7_75t_L g7974 ( 
.A(n_7471),
.B(n_4660),
.Y(n_7974)
);

NAND2xp5_ASAP7_75t_L g7975 ( 
.A(n_7609),
.B(n_4662),
.Y(n_7975)
);

OR2x2_ASAP7_75t_L g7976 ( 
.A(n_7339),
.B(n_4663),
.Y(n_7976)
);

INVx2_ASAP7_75t_L g7977 ( 
.A(n_7476),
.Y(n_7977)
);

NAND2xp5_ASAP7_75t_L g7978 ( 
.A(n_7767),
.B(n_7768),
.Y(n_7978)
);

INVx2_ASAP7_75t_L g7979 ( 
.A(n_7477),
.Y(n_7979)
);

BUFx3_ASAP7_75t_L g7980 ( 
.A(n_7318),
.Y(n_7980)
);

INVx1_ASAP7_75t_L g7981 ( 
.A(n_7481),
.Y(n_7981)
);

NAND2xp5_ASAP7_75t_SL g7982 ( 
.A(n_7697),
.B(n_4665),
.Y(n_7982)
);

INVx2_ASAP7_75t_L g7983 ( 
.A(n_7486),
.Y(n_7983)
);

NAND2xp5_ASAP7_75t_SL g7984 ( 
.A(n_7326),
.B(n_4666),
.Y(n_7984)
);

NOR2xp33_ASAP7_75t_L g7985 ( 
.A(n_7354),
.B(n_4667),
.Y(n_7985)
);

AND2x2_ASAP7_75t_L g7986 ( 
.A(n_7562),
.B(n_5653),
.Y(n_7986)
);

CKINVDCx5p33_ASAP7_75t_R g7987 ( 
.A(n_7315),
.Y(n_7987)
);

INVx2_ASAP7_75t_L g7988 ( 
.A(n_7489),
.Y(n_7988)
);

INVx2_ASAP7_75t_L g7989 ( 
.A(n_7493),
.Y(n_7989)
);

INVx1_ASAP7_75t_L g7990 ( 
.A(n_7497),
.Y(n_7990)
);

OR2x2_ASAP7_75t_L g7991 ( 
.A(n_7348),
.B(n_4668),
.Y(n_7991)
);

INVx1_ASAP7_75t_L g7992 ( 
.A(n_7499),
.Y(n_7992)
);

INVx1_ASAP7_75t_L g7993 ( 
.A(n_7503),
.Y(n_7993)
);

INVx2_ASAP7_75t_L g7994 ( 
.A(n_7510),
.Y(n_7994)
);

AOI22xp33_ASAP7_75t_L g7995 ( 
.A1(n_7724),
.A2(n_5538),
.B1(n_5547),
.B2(n_5481),
.Y(n_7995)
);

NAND2xp5_ASAP7_75t_L g7996 ( 
.A(n_7772),
.B(n_4671),
.Y(n_7996)
);

INVx1_ASAP7_75t_L g7997 ( 
.A(n_7512),
.Y(n_7997)
);

INVx2_ASAP7_75t_L g7998 ( 
.A(n_7515),
.Y(n_7998)
);

INVx1_ASAP7_75t_L g7999 ( 
.A(n_7516),
.Y(n_7999)
);

INVx3_ASAP7_75t_L g8000 ( 
.A(n_7809),
.Y(n_8000)
);

NAND2xp5_ASAP7_75t_L g8001 ( 
.A(n_7776),
.B(n_4675),
.Y(n_8001)
);

INVx2_ASAP7_75t_L g8002 ( 
.A(n_7519),
.Y(n_8002)
);

INVx1_ASAP7_75t_L g8003 ( 
.A(n_7525),
.Y(n_8003)
);

BUFx6f_ASAP7_75t_L g8004 ( 
.A(n_7331),
.Y(n_8004)
);

INVx1_ASAP7_75t_L g8005 ( 
.A(n_7544),
.Y(n_8005)
);

INVx3_ASAP7_75t_L g8006 ( 
.A(n_7828),
.Y(n_8006)
);

NAND3xp33_ASAP7_75t_L g8007 ( 
.A(n_7298),
.B(n_4678),
.C(n_4676),
.Y(n_8007)
);

INVx3_ASAP7_75t_L g8008 ( 
.A(n_7828),
.Y(n_8008)
);

INVx2_ASAP7_75t_L g8009 ( 
.A(n_7545),
.Y(n_8009)
);

NAND2xp5_ASAP7_75t_SL g8010 ( 
.A(n_7652),
.B(n_4679),
.Y(n_8010)
);

INVx2_ASAP7_75t_L g8011 ( 
.A(n_7548),
.Y(n_8011)
);

NAND2xp5_ASAP7_75t_SL g8012 ( 
.A(n_7396),
.B(n_4680),
.Y(n_8012)
);

INVx2_ASAP7_75t_L g8013 ( 
.A(n_7550),
.Y(n_8013)
);

NAND2xp5_ASAP7_75t_SL g8014 ( 
.A(n_7440),
.B(n_4681),
.Y(n_8014)
);

INVx1_ASAP7_75t_L g8015 ( 
.A(n_7535),
.Y(n_8015)
);

INVx1_ASAP7_75t_L g8016 ( 
.A(n_7542),
.Y(n_8016)
);

AO21x2_ASAP7_75t_L g8017 ( 
.A1(n_7725),
.A2(n_4855),
.B(n_4854),
.Y(n_8017)
);

INVx1_ASAP7_75t_L g8018 ( 
.A(n_7553),
.Y(n_8018)
);

AOI22xp33_ASAP7_75t_L g8019 ( 
.A1(n_7726),
.A2(n_5566),
.B1(n_5585),
.B2(n_5565),
.Y(n_8019)
);

OR2x6_ASAP7_75t_L g8020 ( 
.A(n_7753),
.B(n_7649),
.Y(n_8020)
);

CKINVDCx5p33_ASAP7_75t_R g8021 ( 
.A(n_7336),
.Y(n_8021)
);

INVx2_ASAP7_75t_SL g8022 ( 
.A(n_7536),
.Y(n_8022)
);

INVx2_ASAP7_75t_L g8023 ( 
.A(n_7670),
.Y(n_8023)
);

INVx2_ASAP7_75t_L g8024 ( 
.A(n_7678),
.Y(n_8024)
);

INVx2_ASAP7_75t_L g8025 ( 
.A(n_7681),
.Y(n_8025)
);

BUFx6f_ASAP7_75t_L g8026 ( 
.A(n_7347),
.Y(n_8026)
);

BUFx2_ASAP7_75t_L g8027 ( 
.A(n_7605),
.Y(n_8027)
);

AND2x2_ASAP7_75t_L g8028 ( 
.A(n_7351),
.B(n_5653),
.Y(n_8028)
);

NAND2xp5_ASAP7_75t_SL g8029 ( 
.A(n_7717),
.B(n_4684),
.Y(n_8029)
);

NAND2xp5_ASAP7_75t_SL g8030 ( 
.A(n_7718),
.B(n_4686),
.Y(n_8030)
);

INVx1_ASAP7_75t_L g8031 ( 
.A(n_7557),
.Y(n_8031)
);

NOR2x1p5_ASAP7_75t_L g8032 ( 
.A(n_7616),
.B(n_4688),
.Y(n_8032)
);

INVx2_ASAP7_75t_L g8033 ( 
.A(n_7689),
.Y(n_8033)
);

BUFx6f_ASAP7_75t_SL g8034 ( 
.A(n_7352),
.Y(n_8034)
);

AND2x2_ASAP7_75t_L g8035 ( 
.A(n_7524),
.B(n_4693),
.Y(n_8035)
);

INVx5_ASAP7_75t_L g8036 ( 
.A(n_7456),
.Y(n_8036)
);

INVx1_ASAP7_75t_L g8037 ( 
.A(n_7559),
.Y(n_8037)
);

INVx3_ASAP7_75t_L g8038 ( 
.A(n_7347),
.Y(n_8038)
);

NAND2xp5_ASAP7_75t_L g8039 ( 
.A(n_7777),
.B(n_4696),
.Y(n_8039)
);

OR2x2_ASAP7_75t_L g8040 ( 
.A(n_7380),
.B(n_4699),
.Y(n_8040)
);

NAND2xp5_ASAP7_75t_SL g8041 ( 
.A(n_7719),
.B(n_4700),
.Y(n_8041)
);

INVx1_ASAP7_75t_L g8042 ( 
.A(n_7560),
.Y(n_8042)
);

NAND2xp5_ASAP7_75t_L g8043 ( 
.A(n_7780),
.B(n_4701),
.Y(n_8043)
);

INVx4_ASAP7_75t_L g8044 ( 
.A(n_7507),
.Y(n_8044)
);

NOR2xp33_ASAP7_75t_L g8045 ( 
.A(n_7473),
.B(n_4703),
.Y(n_8045)
);

INVxp67_ASAP7_75t_L g8046 ( 
.A(n_7325),
.Y(n_8046)
);

INVx1_ASAP7_75t_L g8047 ( 
.A(n_7563),
.Y(n_8047)
);

INVx1_ASAP7_75t_L g8048 ( 
.A(n_7568),
.Y(n_8048)
);

BUFx10_ASAP7_75t_L g8049 ( 
.A(n_7337),
.Y(n_8049)
);

INVx2_ASAP7_75t_L g8050 ( 
.A(n_7500),
.Y(n_8050)
);

NOR2xp33_ASAP7_75t_L g8051 ( 
.A(n_7751),
.B(n_4704),
.Y(n_8051)
);

AOI22xp5_ASAP7_75t_L g8052 ( 
.A1(n_7669),
.A2(n_4709),
.B1(n_4714),
.B2(n_4705),
.Y(n_8052)
);

INVx2_ASAP7_75t_L g8053 ( 
.A(n_7502),
.Y(n_8053)
);

INVx2_ASAP7_75t_L g8054 ( 
.A(n_7505),
.Y(n_8054)
);

INVx1_ASAP7_75t_L g8055 ( 
.A(n_7570),
.Y(n_8055)
);

INVx2_ASAP7_75t_L g8056 ( 
.A(n_7514),
.Y(n_8056)
);

AND2x2_ASAP7_75t_L g8057 ( 
.A(n_7534),
.B(n_4716),
.Y(n_8057)
);

INVx2_ASAP7_75t_L g8058 ( 
.A(n_7521),
.Y(n_8058)
);

AND3x2_ASAP7_75t_L g8059 ( 
.A(n_7566),
.B(n_4868),
.C(n_4866),
.Y(n_8059)
);

AOI22xp5_ASAP7_75t_L g8060 ( 
.A1(n_7744),
.A2(n_7783),
.B1(n_7791),
.B2(n_7786),
.Y(n_8060)
);

INVx1_ASAP7_75t_L g8061 ( 
.A(n_7577),
.Y(n_8061)
);

INVx2_ASAP7_75t_L g8062 ( 
.A(n_7546),
.Y(n_8062)
);

INVx2_ASAP7_75t_L g8063 ( 
.A(n_7554),
.Y(n_8063)
);

INVx2_ASAP7_75t_L g8064 ( 
.A(n_7565),
.Y(n_8064)
);

INVx2_ASAP7_75t_L g8065 ( 
.A(n_7589),
.Y(n_8065)
);

INVx2_ASAP7_75t_SL g8066 ( 
.A(n_7576),
.Y(n_8066)
);

INVx8_ASAP7_75t_L g8067 ( 
.A(n_7508),
.Y(n_8067)
);

INVx1_ASAP7_75t_L g8068 ( 
.A(n_7578),
.Y(n_8068)
);

INVxp67_ASAP7_75t_SL g8069 ( 
.A(n_7361),
.Y(n_8069)
);

AND2x6_ASAP7_75t_L g8070 ( 
.A(n_7798),
.B(n_4869),
.Y(n_8070)
);

INVx1_ASAP7_75t_L g8071 ( 
.A(n_7581),
.Y(n_8071)
);

INVx2_ASAP7_75t_L g8072 ( 
.A(n_7596),
.Y(n_8072)
);

NAND2xp5_ASAP7_75t_SL g8073 ( 
.A(n_7731),
.B(n_4717),
.Y(n_8073)
);

NOR2xp33_ASAP7_75t_L g8074 ( 
.A(n_7603),
.B(n_4718),
.Y(n_8074)
);

AND2x2_ASAP7_75t_L g8075 ( 
.A(n_7384),
.B(n_4721),
.Y(n_8075)
);

NAND2xp5_ASAP7_75t_SL g8076 ( 
.A(n_7737),
.B(n_4723),
.Y(n_8076)
);

NAND3xp33_ASAP7_75t_L g8077 ( 
.A(n_7714),
.B(n_7397),
.C(n_7368),
.Y(n_8077)
);

NAND2xp5_ASAP7_75t_L g8078 ( 
.A(n_7801),
.B(n_7706),
.Y(n_8078)
);

NOR3xp33_ASAP7_75t_L g8079 ( 
.A(n_7805),
.B(n_4726),
.C(n_4725),
.Y(n_8079)
);

BUFx10_ASAP7_75t_L g8080 ( 
.A(n_7343),
.Y(n_8080)
);

INVx2_ASAP7_75t_L g8081 ( 
.A(n_7600),
.Y(n_8081)
);

NAND2xp5_ASAP7_75t_L g8082 ( 
.A(n_7590),
.B(n_4730),
.Y(n_8082)
);

INVx2_ASAP7_75t_SL g8083 ( 
.A(n_7635),
.Y(n_8083)
);

NAND2xp5_ASAP7_75t_SL g8084 ( 
.A(n_7742),
.B(n_7743),
.Y(n_8084)
);

NOR2xp33_ASAP7_75t_L g8085 ( 
.A(n_7659),
.B(n_4732),
.Y(n_8085)
);

BUFx6f_ASAP7_75t_L g8086 ( 
.A(n_7361),
.Y(n_8086)
);

INVx1_ASAP7_75t_L g8087 ( 
.A(n_7584),
.Y(n_8087)
);

BUFx2_ASAP7_75t_L g8088 ( 
.A(n_7623),
.Y(n_8088)
);

INVx3_ASAP7_75t_L g8089 ( 
.A(n_7376),
.Y(n_8089)
);

INVxp33_ASAP7_75t_L g8090 ( 
.A(n_7345),
.Y(n_8090)
);

INVx1_ASAP7_75t_L g8091 ( 
.A(n_7591),
.Y(n_8091)
);

INVx2_ASAP7_75t_SL g8092 ( 
.A(n_7338),
.Y(n_8092)
);

INVx4_ASAP7_75t_L g8093 ( 
.A(n_7509),
.Y(n_8093)
);

INVx1_ASAP7_75t_L g8094 ( 
.A(n_7592),
.Y(n_8094)
);

NAND2xp5_ASAP7_75t_L g8095 ( 
.A(n_7539),
.B(n_4733),
.Y(n_8095)
);

INVx1_ASAP7_75t_L g8096 ( 
.A(n_7593),
.Y(n_8096)
);

INVx1_ASAP7_75t_L g8097 ( 
.A(n_7598),
.Y(n_8097)
);

NAND3xp33_ASAP7_75t_L g8098 ( 
.A(n_7437),
.B(n_4735),
.C(n_4734),
.Y(n_8098)
);

BUFx3_ASAP7_75t_L g8099 ( 
.A(n_7597),
.Y(n_8099)
);

INVx2_ASAP7_75t_L g8100 ( 
.A(n_7608),
.Y(n_8100)
);

INVxp33_ASAP7_75t_L g8101 ( 
.A(n_7675),
.Y(n_8101)
);

NOR2xp33_ASAP7_75t_L g8102 ( 
.A(n_7849),
.B(n_4736),
.Y(n_8102)
);

INVx1_ASAP7_75t_L g8103 ( 
.A(n_7604),
.Y(n_8103)
);

INVx2_ASAP7_75t_SL g8104 ( 
.A(n_7357),
.Y(n_8104)
);

NAND2xp5_ASAP7_75t_SL g8105 ( 
.A(n_7749),
.B(n_4737),
.Y(n_8105)
);

INVx2_ASAP7_75t_L g8106 ( 
.A(n_7614),
.Y(n_8106)
);

BUFx2_ASAP7_75t_L g8107 ( 
.A(n_7626),
.Y(n_8107)
);

INVx4_ASAP7_75t_L g8108 ( 
.A(n_7511),
.Y(n_8108)
);

NAND2xp5_ASAP7_75t_L g8109 ( 
.A(n_7619),
.B(n_4740),
.Y(n_8109)
);

NAND2xp5_ASAP7_75t_L g8110 ( 
.A(n_7732),
.B(n_4741),
.Y(n_8110)
);

INVx1_ASAP7_75t_L g8111 ( 
.A(n_7607),
.Y(n_8111)
);

NAND2xp5_ASAP7_75t_SL g8112 ( 
.A(n_7758),
.B(n_4743),
.Y(n_8112)
);

NAND2xp5_ASAP7_75t_SL g8113 ( 
.A(n_7766),
.B(n_4744),
.Y(n_8113)
);

INVx2_ASAP7_75t_L g8114 ( 
.A(n_7625),
.Y(n_8114)
);

INVx3_ASAP7_75t_L g8115 ( 
.A(n_7376),
.Y(n_8115)
);

INVx2_ASAP7_75t_L g8116 ( 
.A(n_7628),
.Y(n_8116)
);

NAND2xp5_ASAP7_75t_L g8117 ( 
.A(n_7494),
.B(n_4747),
.Y(n_8117)
);

NAND2xp5_ASAP7_75t_L g8118 ( 
.A(n_7540),
.B(n_4748),
.Y(n_8118)
);

INVx2_ASAP7_75t_L g8119 ( 
.A(n_7335),
.Y(n_8119)
);

INVx1_ASAP7_75t_L g8120 ( 
.A(n_7615),
.Y(n_8120)
);

INVx3_ASAP7_75t_L g8121 ( 
.A(n_7423),
.Y(n_8121)
);

INVx2_ASAP7_75t_L g8122 ( 
.A(n_7342),
.Y(n_8122)
);

AOI22xp33_ASAP7_75t_L g8123 ( 
.A1(n_7727),
.A2(n_5589),
.B1(n_5616),
.B2(n_5587),
.Y(n_8123)
);

NAND2xp5_ASAP7_75t_L g8124 ( 
.A(n_7573),
.B(n_4751),
.Y(n_8124)
);

OR2x2_ASAP7_75t_L g8125 ( 
.A(n_7599),
.B(n_4754),
.Y(n_8125)
);

NOR2xp33_ASAP7_75t_L g8126 ( 
.A(n_7859),
.B(n_4755),
.Y(n_8126)
);

INVx3_ASAP7_75t_L g8127 ( 
.A(n_7423),
.Y(n_8127)
);

NAND2xp5_ASAP7_75t_SL g8128 ( 
.A(n_7564),
.B(n_4757),
.Y(n_8128)
);

INVx2_ASAP7_75t_L g8129 ( 
.A(n_7448),
.Y(n_8129)
);

INVx4_ASAP7_75t_L g8130 ( 
.A(n_7551),
.Y(n_8130)
);

NAND2xp5_ASAP7_75t_L g8131 ( 
.A(n_7379),
.B(n_4761),
.Y(n_8131)
);

CKINVDCx20_ASAP7_75t_R g8132 ( 
.A(n_7327),
.Y(n_8132)
);

BUFx10_ASAP7_75t_L g8133 ( 
.A(n_7344),
.Y(n_8133)
);

NAND2xp5_ASAP7_75t_SL g8134 ( 
.A(n_7569),
.B(n_4768),
.Y(n_8134)
);

CKINVDCx5p33_ASAP7_75t_R g8135 ( 
.A(n_7346),
.Y(n_8135)
);

CKINVDCx11_ASAP7_75t_R g8136 ( 
.A(n_7556),
.Y(n_8136)
);

AND2x2_ASAP7_75t_L g8137 ( 
.A(n_7409),
.B(n_4769),
.Y(n_8137)
);

INVx2_ASAP7_75t_L g8138 ( 
.A(n_7488),
.Y(n_8138)
);

INVx1_ASAP7_75t_L g8139 ( 
.A(n_7618),
.Y(n_8139)
);

NOR2xp33_ASAP7_75t_L g8140 ( 
.A(n_7850),
.B(n_4770),
.Y(n_8140)
);

BUFx6f_ASAP7_75t_SL g8141 ( 
.A(n_7362),
.Y(n_8141)
);

NAND2xp5_ASAP7_75t_SL g8142 ( 
.A(n_7571),
.B(n_4774),
.Y(n_8142)
);

NAND2xp5_ASAP7_75t_SL g8143 ( 
.A(n_7574),
.B(n_4775),
.Y(n_8143)
);

INVx2_ASAP7_75t_L g8144 ( 
.A(n_7491),
.Y(n_8144)
);

INVx2_ASAP7_75t_L g8145 ( 
.A(n_7496),
.Y(n_8145)
);

NOR2xp33_ASAP7_75t_L g8146 ( 
.A(n_7837),
.B(n_4777),
.Y(n_8146)
);

INVx1_ASAP7_75t_L g8147 ( 
.A(n_7622),
.Y(n_8147)
);

NAND2xp5_ASAP7_75t_L g8148 ( 
.A(n_7700),
.B(n_7703),
.Y(n_8148)
);

INVx1_ASAP7_75t_L g8149 ( 
.A(n_7629),
.Y(n_8149)
);

INVx2_ASAP7_75t_L g8150 ( 
.A(n_7643),
.Y(n_8150)
);

BUFx2_ASAP7_75t_L g8151 ( 
.A(n_7632),
.Y(n_8151)
);

INVx1_ASAP7_75t_L g8152 ( 
.A(n_7636),
.Y(n_8152)
);

INVx2_ASAP7_75t_L g8153 ( 
.A(n_7646),
.Y(n_8153)
);

BUFx3_ASAP7_75t_L g8154 ( 
.A(n_7587),
.Y(n_8154)
);

NAND2xp5_ASAP7_75t_L g8155 ( 
.A(n_7704),
.B(n_4778),
.Y(n_8155)
);

INVx1_ASAP7_75t_L g8156 ( 
.A(n_7638),
.Y(n_8156)
);

INVx2_ASAP7_75t_L g8157 ( 
.A(n_7653),
.Y(n_8157)
);

INVx1_ASAP7_75t_L g8158 ( 
.A(n_7640),
.Y(n_8158)
);

INVx2_ASAP7_75t_L g8159 ( 
.A(n_7641),
.Y(n_8159)
);

BUFx4f_ASAP7_75t_L g8160 ( 
.A(n_7741),
.Y(n_8160)
);

NAND2xp5_ASAP7_75t_SL g8161 ( 
.A(n_7580),
.B(n_4780),
.Y(n_8161)
);

INVx2_ASAP7_75t_L g8162 ( 
.A(n_7647),
.Y(n_8162)
);

INVx2_ASAP7_75t_L g8163 ( 
.A(n_7648),
.Y(n_8163)
);

INVx2_ASAP7_75t_SL g8164 ( 
.A(n_7388),
.Y(n_8164)
);

INVx3_ASAP7_75t_L g8165 ( 
.A(n_7430),
.Y(n_8165)
);

NAND2xp5_ASAP7_75t_L g8166 ( 
.A(n_7428),
.B(n_4781),
.Y(n_8166)
);

INVx2_ASAP7_75t_L g8167 ( 
.A(n_7650),
.Y(n_8167)
);

NAND2xp5_ASAP7_75t_SL g8168 ( 
.A(n_7610),
.B(n_4782),
.Y(n_8168)
);

NAND2xp5_ASAP7_75t_SL g8169 ( 
.A(n_7611),
.B(n_4784),
.Y(n_8169)
);

INVx1_ASAP7_75t_L g8170 ( 
.A(n_7651),
.Y(n_8170)
);

NAND2xp5_ASAP7_75t_L g8171 ( 
.A(n_7469),
.B(n_4785),
.Y(n_8171)
);

INVx2_ASAP7_75t_L g8172 ( 
.A(n_7661),
.Y(n_8172)
);

NAND2xp5_ASAP7_75t_SL g8173 ( 
.A(n_7613),
.B(n_4788),
.Y(n_8173)
);

INVx1_ASAP7_75t_L g8174 ( 
.A(n_7662),
.Y(n_8174)
);

INVx1_ASAP7_75t_L g8175 ( 
.A(n_7663),
.Y(n_8175)
);

NAND2xp5_ASAP7_75t_SL g8176 ( 
.A(n_7621),
.B(n_7634),
.Y(n_8176)
);

BUFx10_ASAP7_75t_L g8177 ( 
.A(n_7356),
.Y(n_8177)
);

BUFx6f_ASAP7_75t_L g8178 ( 
.A(n_7430),
.Y(n_8178)
);

INVx2_ASAP7_75t_SL g8179 ( 
.A(n_7453),
.Y(n_8179)
);

OAI22xp33_ASAP7_75t_L g8180 ( 
.A1(n_7834),
.A2(n_4793),
.B1(n_4796),
.B2(n_4791),
.Y(n_8180)
);

INVx2_ASAP7_75t_L g8181 ( 
.A(n_7667),
.Y(n_8181)
);

BUFx10_ASAP7_75t_L g8182 ( 
.A(n_7359),
.Y(n_8182)
);

INVx1_ASAP7_75t_L g8183 ( 
.A(n_7673),
.Y(n_8183)
);

INVx2_ASAP7_75t_L g8184 ( 
.A(n_7688),
.Y(n_8184)
);

INVx1_ASAP7_75t_L g8185 ( 
.A(n_7690),
.Y(n_8185)
);

CKINVDCx6p67_ASAP7_75t_R g8186 ( 
.A(n_7594),
.Y(n_8186)
);

INVx2_ASAP7_75t_L g8187 ( 
.A(n_7363),
.Y(n_8187)
);

INVx2_ASAP7_75t_L g8188 ( 
.A(n_7692),
.Y(n_8188)
);

BUFx3_ASAP7_75t_L g8189 ( 
.A(n_7588),
.Y(n_8189)
);

INVx1_ASAP7_75t_L g8190 ( 
.A(n_7561),
.Y(n_8190)
);

INVx2_ASAP7_75t_L g8191 ( 
.A(n_7695),
.Y(n_8191)
);

NAND2xp5_ASAP7_75t_SL g8192 ( 
.A(n_7730),
.B(n_4798),
.Y(n_8192)
);

BUFx3_ASAP7_75t_L g8193 ( 
.A(n_7526),
.Y(n_8193)
);

INVx1_ASAP7_75t_L g8194 ( 
.A(n_7555),
.Y(n_8194)
);

INVx2_ASAP7_75t_L g8195 ( 
.A(n_7709),
.Y(n_8195)
);

NOR2xp33_ASAP7_75t_L g8196 ( 
.A(n_7844),
.B(n_4799),
.Y(n_8196)
);

INVx2_ASAP7_75t_L g8197 ( 
.A(n_7712),
.Y(n_8197)
);

NOR2xp33_ASAP7_75t_L g8198 ( 
.A(n_7854),
.B(n_4800),
.Y(n_8198)
);

NOR2x1p5_ASAP7_75t_L g8199 ( 
.A(n_7478),
.B(n_4802),
.Y(n_8199)
);

INVx2_ASAP7_75t_L g8200 ( 
.A(n_7740),
.Y(n_8200)
);

NAND2xp5_ASAP7_75t_L g8201 ( 
.A(n_7498),
.B(n_7575),
.Y(n_8201)
);

INVxp33_ASAP7_75t_L g8202 ( 
.A(n_7330),
.Y(n_8202)
);

INVx1_ASAP7_75t_L g8203 ( 
.A(n_7729),
.Y(n_8203)
);

OR2x2_ASAP7_75t_L g8204 ( 
.A(n_7796),
.B(n_4804),
.Y(n_8204)
);

INVxp67_ASAP7_75t_SL g8205 ( 
.A(n_7538),
.Y(n_8205)
);

INVx2_ASAP7_75t_L g8206 ( 
.A(n_7754),
.Y(n_8206)
);

INVx1_ASAP7_75t_L g8207 ( 
.A(n_7760),
.Y(n_8207)
);

INVx2_ASAP7_75t_L g8208 ( 
.A(n_7761),
.Y(n_8208)
);

BUFx6f_ASAP7_75t_L g8209 ( 
.A(n_7538),
.Y(n_8209)
);

OR2x2_ASAP7_75t_L g8210 ( 
.A(n_7306),
.B(n_4806),
.Y(n_8210)
);

INVx2_ASAP7_75t_L g8211 ( 
.A(n_7762),
.Y(n_8211)
);

NAND2xp33_ASAP7_75t_L g8212 ( 
.A(n_7741),
.B(n_4808),
.Y(n_8212)
);

INVx2_ASAP7_75t_L g8213 ( 
.A(n_7763),
.Y(n_8213)
);

INVx2_ASAP7_75t_L g8214 ( 
.A(n_7771),
.Y(n_8214)
);

NOR2xp33_ASAP7_75t_L g8215 ( 
.A(n_7855),
.B(n_7857),
.Y(n_8215)
);

INVx1_ASAP7_75t_L g8216 ( 
.A(n_7316),
.Y(n_8216)
);

NAND2xp5_ASAP7_75t_SL g8217 ( 
.A(n_7366),
.B(n_4811),
.Y(n_8217)
);

INVx2_ASAP7_75t_L g8218 ( 
.A(n_7785),
.Y(n_8218)
);

NAND2xp5_ASAP7_75t_SL g8219 ( 
.A(n_7631),
.B(n_7517),
.Y(n_8219)
);

NOR2xp33_ASAP7_75t_L g8220 ( 
.A(n_7779),
.B(n_4812),
.Y(n_8220)
);

INVx2_ASAP7_75t_L g8221 ( 
.A(n_7794),
.Y(n_8221)
);

INVxp33_ASAP7_75t_L g8222 ( 
.A(n_7639),
.Y(n_8222)
);

INVx1_ASAP7_75t_L g8223 ( 
.A(n_7800),
.Y(n_8223)
);

NAND2xp5_ASAP7_75t_L g8224 ( 
.A(n_7583),
.B(n_4817),
.Y(n_8224)
);

INVx1_ASAP7_75t_L g8225 ( 
.A(n_7784),
.Y(n_8225)
);

NAND2xp5_ASAP7_75t_SL g8226 ( 
.A(n_7842),
.B(n_7774),
.Y(n_8226)
);

INVx1_ASAP7_75t_L g8227 ( 
.A(n_7685),
.Y(n_8227)
);

AND2x2_ASAP7_75t_L g8228 ( 
.A(n_7655),
.B(n_4820),
.Y(n_8228)
);

INVx4_ASAP7_75t_L g8229 ( 
.A(n_7373),
.Y(n_8229)
);

INVx1_ASAP7_75t_L g8230 ( 
.A(n_7728),
.Y(n_8230)
);

BUFx2_ASAP7_75t_L g8231 ( 
.A(n_7334),
.Y(n_8231)
);

INVx2_ASAP7_75t_L g8232 ( 
.A(n_7736),
.Y(n_8232)
);

INVx1_ASAP7_75t_L g8233 ( 
.A(n_7746),
.Y(n_8233)
);

INVx2_ASAP7_75t_L g8234 ( 
.A(n_7748),
.Y(n_8234)
);

INVx2_ASAP7_75t_SL g8235 ( 
.A(n_7355),
.Y(n_8235)
);

BUFx6f_ASAP7_75t_L g8236 ( 
.A(n_7541),
.Y(n_8236)
);

INVx1_ASAP7_75t_L g8237 ( 
.A(n_7642),
.Y(n_8237)
);

INVx3_ASAP7_75t_L g8238 ( 
.A(n_7541),
.Y(n_8238)
);

INVx3_ASAP7_75t_L g8239 ( 
.A(n_7567),
.Y(n_8239)
);

INVx2_ASAP7_75t_SL g8240 ( 
.A(n_7527),
.Y(n_8240)
);

INVx2_ASAP7_75t_L g8241 ( 
.A(n_7394),
.Y(n_8241)
);

NAND2xp5_ASAP7_75t_SL g8242 ( 
.A(n_7620),
.B(n_7671),
.Y(n_8242)
);

INVx2_ASAP7_75t_L g8243 ( 
.A(n_7816),
.Y(n_8243)
);

INVx1_ASAP7_75t_L g8244 ( 
.A(n_7656),
.Y(n_8244)
);

NAND2xp5_ASAP7_75t_SL g8245 ( 
.A(n_7480),
.B(n_7770),
.Y(n_8245)
);

NAND2xp5_ASAP7_75t_SL g8246 ( 
.A(n_7858),
.B(n_4823),
.Y(n_8246)
);

NAND2xp5_ASAP7_75t_SL g8247 ( 
.A(n_7832),
.B(n_4824),
.Y(n_8247)
);

CKINVDCx5p33_ASAP7_75t_R g8248 ( 
.A(n_7378),
.Y(n_8248)
);

INVxp33_ASAP7_75t_L g8249 ( 
.A(n_7657),
.Y(n_8249)
);

BUFx6f_ASAP7_75t_L g8250 ( 
.A(n_7567),
.Y(n_8250)
);

INVx1_ASAP7_75t_L g8251 ( 
.A(n_7682),
.Y(n_8251)
);

BUFx6f_ASAP7_75t_L g8252 ( 
.A(n_7684),
.Y(n_8252)
);

NAND2xp5_ASAP7_75t_L g8253 ( 
.A(n_7586),
.B(n_4825),
.Y(n_8253)
);

INVx2_ASAP7_75t_SL g8254 ( 
.A(n_7807),
.Y(n_8254)
);

INVx2_ASAP7_75t_L g8255 ( 
.A(n_7838),
.Y(n_8255)
);

NOR2xp33_ASAP7_75t_L g8256 ( 
.A(n_7781),
.B(n_4827),
.Y(n_8256)
);

NAND2xp5_ASAP7_75t_SL g8257 ( 
.A(n_7645),
.B(n_4828),
.Y(n_8257)
);

NAND2xp5_ASAP7_75t_L g8258 ( 
.A(n_7462),
.B(n_4830),
.Y(n_8258)
);

INVx2_ASAP7_75t_L g8259 ( 
.A(n_7856),
.Y(n_8259)
);

BUFx6f_ASAP7_75t_L g8260 ( 
.A(n_7684),
.Y(n_8260)
);

INVx1_ASAP7_75t_L g8261 ( 
.A(n_7674),
.Y(n_8261)
);

NOR2xp33_ASAP7_75t_L g8262 ( 
.A(n_7764),
.B(n_4836),
.Y(n_8262)
);

INVx2_ASAP7_75t_L g8263 ( 
.A(n_7853),
.Y(n_8263)
);

INVx2_ASAP7_75t_SL g8264 ( 
.A(n_7745),
.Y(n_8264)
);

NOR2xp33_ASAP7_75t_L g8265 ( 
.A(n_7812),
.B(n_4837),
.Y(n_8265)
);

INVx1_ASAP7_75t_L g8266 ( 
.A(n_7474),
.Y(n_8266)
);

BUFx2_ASAP7_75t_L g8267 ( 
.A(n_7386),
.Y(n_8267)
);

AND3x2_ASAP7_75t_L g8268 ( 
.A(n_7624),
.B(n_4879),
.C(n_4872),
.Y(n_8268)
);

NAND2xp5_ASAP7_75t_SL g8269 ( 
.A(n_7811),
.B(n_4839),
.Y(n_8269)
);

INVx6_ASAP7_75t_L g8270 ( 
.A(n_7739),
.Y(n_8270)
);

NAND2xp5_ASAP7_75t_L g8271 ( 
.A(n_7479),
.B(n_4842),
.Y(n_8271)
);

BUFx3_ASAP7_75t_L g8272 ( 
.A(n_7745),
.Y(n_8272)
);

INVx2_ASAP7_75t_L g8273 ( 
.A(n_7450),
.Y(n_8273)
);

INVx2_ASAP7_75t_L g8274 ( 
.A(n_7572),
.Y(n_8274)
);

BUFx6f_ASAP7_75t_L g8275 ( 
.A(n_7696),
.Y(n_8275)
);

INVx1_ASAP7_75t_L g8276 ( 
.A(n_7817),
.Y(n_8276)
);

NAND2xp33_ASAP7_75t_L g8277 ( 
.A(n_7741),
.B(n_4845),
.Y(n_8277)
);

INVx1_ASAP7_75t_L g8278 ( 
.A(n_7818),
.Y(n_8278)
);

CKINVDCx20_ASAP7_75t_R g8279 ( 
.A(n_7301),
.Y(n_8279)
);

INVx3_ASAP7_75t_L g8280 ( 
.A(n_7395),
.Y(n_8280)
);

INVx2_ASAP7_75t_L g8281 ( 
.A(n_7840),
.Y(n_8281)
);

INVx2_ASAP7_75t_L g8282 ( 
.A(n_7813),
.Y(n_8282)
);

INVx2_ASAP7_75t_SL g8283 ( 
.A(n_7735),
.Y(n_8283)
);

CKINVDCx6p67_ASAP7_75t_R g8284 ( 
.A(n_7419),
.Y(n_8284)
);

NAND2xp5_ASAP7_75t_SL g8285 ( 
.A(n_7814),
.B(n_4846),
.Y(n_8285)
);

NAND2xp5_ASAP7_75t_SL g8286 ( 
.A(n_7422),
.B(n_4847),
.Y(n_8286)
);

INVx1_ASAP7_75t_L g8287 ( 
.A(n_7819),
.Y(n_8287)
);

BUFx6f_ASAP7_75t_L g8288 ( 
.A(n_7321),
.Y(n_8288)
);

INVx2_ASAP7_75t_SL g8289 ( 
.A(n_7672),
.Y(n_8289)
);

NAND2xp5_ASAP7_75t_SL g8290 ( 
.A(n_7443),
.B(n_4848),
.Y(n_8290)
);

NOR2xp33_ASAP7_75t_L g8291 ( 
.A(n_7630),
.B(n_7679),
.Y(n_8291)
);

INVx2_ASAP7_75t_L g8292 ( 
.A(n_7839),
.Y(n_8292)
);

INVx2_ASAP7_75t_L g8293 ( 
.A(n_7803),
.Y(n_8293)
);

INVx2_ASAP7_75t_L g8294 ( 
.A(n_7845),
.Y(n_8294)
);

INVx1_ASAP7_75t_L g8295 ( 
.A(n_7820),
.Y(n_8295)
);

INVx3_ASAP7_75t_L g8296 ( 
.A(n_7399),
.Y(n_8296)
);

INVx1_ASAP7_75t_L g8297 ( 
.A(n_7824),
.Y(n_8297)
);

INVx1_ASAP7_75t_L g8298 ( 
.A(n_7830),
.Y(n_8298)
);

INVx1_ASAP7_75t_L g8299 ( 
.A(n_7835),
.Y(n_8299)
);

INVx1_ASAP7_75t_L g8300 ( 
.A(n_7841),
.Y(n_8300)
);

INVx3_ASAP7_75t_L g8301 ( 
.A(n_7410),
.Y(n_8301)
);

BUFx10_ASAP7_75t_L g8302 ( 
.A(n_7582),
.Y(n_8302)
);

INVx1_ASAP7_75t_L g8303 ( 
.A(n_7847),
.Y(n_8303)
);

NAND2xp5_ASAP7_75t_SL g8304 ( 
.A(n_7747),
.B(n_4849),
.Y(n_8304)
);

INVx3_ASAP7_75t_L g8305 ( 
.A(n_7417),
.Y(n_8305)
);

INVx1_ASAP7_75t_L g8306 ( 
.A(n_7680),
.Y(n_8306)
);

INVx1_ASAP7_75t_L g8307 ( 
.A(n_7459),
.Y(n_8307)
);

INVx2_ASAP7_75t_L g8308 ( 
.A(n_7429),
.Y(n_8308)
);

INVx2_ASAP7_75t_L g8309 ( 
.A(n_7402),
.Y(n_8309)
);

INVx2_ASAP7_75t_L g8310 ( 
.A(n_7513),
.Y(n_8310)
);

INVx4_ASAP7_75t_L g8311 ( 
.A(n_7701),
.Y(n_8311)
);

OR2x2_ASAP7_75t_SL g8312 ( 
.A(n_7821),
.B(n_5621),
.Y(n_8312)
);

INVx2_ASAP7_75t_L g8313 ( 
.A(n_7377),
.Y(n_8313)
);

INVx2_ASAP7_75t_L g8314 ( 
.A(n_7382),
.Y(n_8314)
);

INVx2_ASAP7_75t_L g8315 ( 
.A(n_7602),
.Y(n_8315)
);

BUFx6f_ASAP7_75t_L g8316 ( 
.A(n_7482),
.Y(n_8316)
);

INVx3_ASAP7_75t_L g8317 ( 
.A(n_7436),
.Y(n_8317)
);

AOI22xp5_ASAP7_75t_L g8318 ( 
.A1(n_7720),
.A2(n_4857),
.B1(n_4858),
.B2(n_4851),
.Y(n_8318)
);

NAND2xp5_ASAP7_75t_SL g8319 ( 
.A(n_7713),
.B(n_4860),
.Y(n_8319)
);

INVx2_ASAP7_75t_L g8320 ( 
.A(n_7644),
.Y(n_8320)
);

INVx6_ASAP7_75t_L g8321 ( 
.A(n_7846),
.Y(n_8321)
);

NAND2xp5_ASAP7_75t_L g8322 ( 
.A(n_7759),
.B(n_7738),
.Y(n_8322)
);

NAND2xp5_ASAP7_75t_L g8323 ( 
.A(n_7759),
.B(n_4861),
.Y(n_8323)
);

INVx1_ASAP7_75t_L g8324 ( 
.A(n_7438),
.Y(n_8324)
);

NOR2xp33_ASAP7_75t_L g8325 ( 
.A(n_7529),
.B(n_4864),
.Y(n_8325)
);

BUFx3_ASAP7_75t_L g8326 ( 
.A(n_7353),
.Y(n_8326)
);

BUFx6f_ASAP7_75t_L g8327 ( 
.A(n_7716),
.Y(n_8327)
);

NAND2xp5_ASAP7_75t_SL g8328 ( 
.A(n_7836),
.B(n_7522),
.Y(n_8328)
);

NAND2xp5_ASAP7_75t_L g8329 ( 
.A(n_7759),
.B(n_4867),
.Y(n_8329)
);

INVx2_ASAP7_75t_L g8330 ( 
.A(n_7664),
.Y(n_8330)
);

INVx2_ASAP7_75t_SL g8331 ( 
.A(n_7722),
.Y(n_8331)
);

INVx2_ASAP7_75t_L g8332 ( 
.A(n_7666),
.Y(n_8332)
);

INVx2_ASAP7_75t_L g8333 ( 
.A(n_7483),
.Y(n_8333)
);

INVx1_ASAP7_75t_L g8334 ( 
.A(n_7595),
.Y(n_8334)
);

INVx1_ASAP7_75t_L g8335 ( 
.A(n_7848),
.Y(n_8335)
);

NAND3xp33_ASAP7_75t_L g8336 ( 
.A(n_7420),
.B(n_4874),
.C(n_4870),
.Y(n_8336)
);

INVx2_ASAP7_75t_L g8337 ( 
.A(n_7775),
.Y(n_8337)
);

INVx1_ASAP7_75t_L g8338 ( 
.A(n_7792),
.Y(n_8338)
);

NAND3xp33_ASAP7_75t_L g8339 ( 
.A(n_7358),
.B(n_4876),
.C(n_4875),
.Y(n_8339)
);

AND2x6_ASAP7_75t_L g8340 ( 
.A(n_7773),
.B(n_4881),
.Y(n_8340)
);

INVx2_ASAP7_75t_L g8341 ( 
.A(n_7833),
.Y(n_8341)
);

INVx1_ASAP7_75t_L g8342 ( 
.A(n_7707),
.Y(n_8342)
);

INVx1_ASAP7_75t_L g8343 ( 
.A(n_7711),
.Y(n_8343)
);

NAND2xp5_ASAP7_75t_SL g8344 ( 
.A(n_7804),
.B(n_4877),
.Y(n_8344)
);

NAND2xp5_ASAP7_75t_L g8345 ( 
.A(n_7788),
.B(n_7797),
.Y(n_8345)
);

BUFx6f_ASAP7_75t_SL g8346 ( 
.A(n_7456),
.Y(n_8346)
);

INVx1_ASAP7_75t_L g8347 ( 
.A(n_7456),
.Y(n_8347)
);

BUFx2_ASAP7_75t_L g8348 ( 
.A(n_7691),
.Y(n_8348)
);

NAND2xp5_ASAP7_75t_L g8349 ( 
.A(n_7831),
.B(n_4880),
.Y(n_8349)
);

INVx2_ASAP7_75t_L g8350 ( 
.A(n_7723),
.Y(n_8350)
);

OR2x2_ASAP7_75t_L g8351 ( 
.A(n_7617),
.B(n_4882),
.Y(n_8351)
);

NAND2xp33_ASAP7_75t_SL g8352 ( 
.A(n_7808),
.B(n_4883),
.Y(n_8352)
);

INVx1_ASAP7_75t_L g8353 ( 
.A(n_7485),
.Y(n_8353)
);

INVx1_ASAP7_75t_L g8354 ( 
.A(n_7485),
.Y(n_8354)
);

NAND2xp5_ASAP7_75t_SL g8355 ( 
.A(n_7710),
.B(n_4884),
.Y(n_8355)
);

INVx6_ASAP7_75t_L g8356 ( 
.A(n_7485),
.Y(n_8356)
);

NAND2xp5_ASAP7_75t_SL g8357 ( 
.A(n_7822),
.B(n_4886),
.Y(n_8357)
);

INVx2_ASAP7_75t_L g8358 ( 
.A(n_7823),
.Y(n_8358)
);

INVx2_ASAP7_75t_L g8359 ( 
.A(n_7829),
.Y(n_8359)
);

INVx2_ASAP7_75t_L g8360 ( 
.A(n_7367),
.Y(n_8360)
);

INVx3_ASAP7_75t_L g8361 ( 
.A(n_7530),
.Y(n_8361)
);

INVx2_ASAP7_75t_L g8362 ( 
.A(n_7627),
.Y(n_8362)
);

INVx2_ASAP7_75t_SL g8363 ( 
.A(n_7531),
.Y(n_8363)
);

INVx2_ASAP7_75t_L g8364 ( 
.A(n_7612),
.Y(n_8364)
);

INVx2_ASAP7_75t_L g8365 ( 
.A(n_7852),
.Y(n_8365)
);

INVx2_ASAP7_75t_L g8366 ( 
.A(n_7769),
.Y(n_8366)
);

NAND2xp5_ASAP7_75t_SL g8367 ( 
.A(n_7694),
.B(n_4887),
.Y(n_8367)
);

AOI22xp33_ASAP7_75t_L g8368 ( 
.A1(n_7698),
.A2(n_5643),
.B1(n_5652),
.B2(n_5629),
.Y(n_8368)
);

CKINVDCx6p67_ASAP7_75t_R g8369 ( 
.A(n_7633),
.Y(n_8369)
);

INVx3_ASAP7_75t_L g8370 ( 
.A(n_7532),
.Y(n_8370)
);

NAND2xp5_ASAP7_75t_L g8371 ( 
.A(n_7795),
.B(n_4891),
.Y(n_8371)
);

OR2x2_ASAP7_75t_L g8372 ( 
.A(n_7501),
.B(n_4892),
.Y(n_8372)
);

INVx1_ASAP7_75t_L g8373 ( 
.A(n_7404),
.Y(n_8373)
);

INVx1_ASAP7_75t_L g8374 ( 
.A(n_7533),
.Y(n_8374)
);

INVx1_ASAP7_75t_L g8375 ( 
.A(n_7537),
.Y(n_8375)
);

NAND2xp5_ASAP7_75t_L g8376 ( 
.A(n_7543),
.B(n_4895),
.Y(n_8376)
);

INVx2_ASAP7_75t_L g8377 ( 
.A(n_7547),
.Y(n_8377)
);

NOR2xp33_ASAP7_75t_L g8378 ( 
.A(n_7549),
.B(n_4897),
.Y(n_8378)
);

OAI22xp5_ASAP7_75t_L g8379 ( 
.A1(n_7843),
.A2(n_4899),
.B1(n_4904),
.B2(n_4898),
.Y(n_8379)
);

INVx1_ASAP7_75t_L g8380 ( 
.A(n_7787),
.Y(n_8380)
);

INVx2_ASAP7_75t_L g8381 ( 
.A(n_7793),
.Y(n_8381)
);

INVx2_ASAP7_75t_L g8382 ( 
.A(n_7654),
.Y(n_8382)
);

INVx1_ASAP7_75t_L g8383 ( 
.A(n_7658),
.Y(n_8383)
);

INVx2_ASAP7_75t_L g8384 ( 
.A(n_7660),
.Y(n_8384)
);

INVx2_ASAP7_75t_L g8385 ( 
.A(n_7668),
.Y(n_8385)
);

NAND2xp5_ASAP7_75t_L g8386 ( 
.A(n_7412),
.B(n_4905),
.Y(n_8386)
);

NAND2xp5_ASAP7_75t_SL g8387 ( 
.A(n_7415),
.B(n_4913),
.Y(n_8387)
);

INVx2_ASAP7_75t_SL g8388 ( 
.A(n_7414),
.Y(n_8388)
);

NOR2xp33_ASAP7_75t_L g8389 ( 
.A(n_7416),
.B(n_4914),
.Y(n_8389)
);

INVx1_ASAP7_75t_L g8390 ( 
.A(n_7734),
.Y(n_8390)
);

INVx1_ASAP7_75t_L g8391 ( 
.A(n_7755),
.Y(n_8391)
);

INVx1_ASAP7_75t_L g8392 ( 
.A(n_7756),
.Y(n_8392)
);

INVx3_ASAP7_75t_L g8393 ( 
.A(n_7390),
.Y(n_8393)
);

CKINVDCx6p67_ASAP7_75t_R g8394 ( 
.A(n_7391),
.Y(n_8394)
);

INVx2_ASAP7_75t_L g8395 ( 
.A(n_7424),
.Y(n_8395)
);

CKINVDCx20_ASAP7_75t_R g8396 ( 
.A(n_7406),
.Y(n_8396)
);

INVx1_ASAP7_75t_L g8397 ( 
.A(n_7427),
.Y(n_8397)
);

INVx1_ASAP7_75t_L g8398 ( 
.A(n_7435),
.Y(n_8398)
);

BUFx10_ASAP7_75t_L g8399 ( 
.A(n_7300),
.Y(n_8399)
);

AO21x2_ASAP7_75t_L g8400 ( 
.A1(n_7370),
.A2(n_4896),
.B(n_4893),
.Y(n_8400)
);

INVx2_ASAP7_75t_L g8401 ( 
.A(n_7451),
.Y(n_8401)
);

INVx1_ASAP7_75t_L g8402 ( 
.A(n_7455),
.Y(n_8402)
);

INVx2_ASAP7_75t_L g8403 ( 
.A(n_7460),
.Y(n_8403)
);

INVx3_ASAP7_75t_L g8404 ( 
.A(n_7411),
.Y(n_8404)
);

INVx2_ASAP7_75t_L g8405 ( 
.A(n_7461),
.Y(n_8405)
);

BUFx2_ASAP7_75t_L g8406 ( 
.A(n_7445),
.Y(n_8406)
);

NAND2xp5_ASAP7_75t_SL g8407 ( 
.A(n_7464),
.B(n_4918),
.Y(n_8407)
);

INVx2_ASAP7_75t_L g8408 ( 
.A(n_7468),
.Y(n_8408)
);

INVx1_ASAP7_75t_L g8409 ( 
.A(n_7802),
.Y(n_8409)
);

NAND2xp5_ASAP7_75t_SL g8410 ( 
.A(n_7676),
.B(n_4921),
.Y(n_8410)
);

INVx1_ASAP7_75t_L g8411 ( 
.A(n_7825),
.Y(n_8411)
);

INVx2_ASAP7_75t_L g8412 ( 
.A(n_7520),
.Y(n_8412)
);

CKINVDCx5p33_ASAP7_75t_R g8413 ( 
.A(n_7302),
.Y(n_8413)
);

INVx1_ASAP7_75t_L g8414 ( 
.A(n_7863),
.Y(n_8414)
);

NAND2xp5_ASAP7_75t_L g8415 ( 
.A(n_7944),
.B(n_4923),
.Y(n_8415)
);

OR2x6_ASAP7_75t_L g8416 ( 
.A(n_8067),
.B(n_7408),
.Y(n_8416)
);

NAND2xp5_ASAP7_75t_L g8417 ( 
.A(n_7928),
.B(n_4926),
.Y(n_8417)
);

INVx1_ASAP7_75t_L g8418 ( 
.A(n_7869),
.Y(n_8418)
);

INVx2_ASAP7_75t_L g8419 ( 
.A(n_7916),
.Y(n_8419)
);

INVx2_ASAP7_75t_L g8420 ( 
.A(n_7919),
.Y(n_8420)
);

NAND2xp5_ASAP7_75t_L g8421 ( 
.A(n_8078),
.B(n_4927),
.Y(n_8421)
);

AND2x4_ASAP7_75t_L g8422 ( 
.A(n_7870),
.B(n_7311),
.Y(n_8422)
);

HB1xp67_ASAP7_75t_L g8423 ( 
.A(n_7872),
.Y(n_8423)
);

INVx1_ASAP7_75t_SL g8424 ( 
.A(n_7897),
.Y(n_8424)
);

AND2x4_ASAP7_75t_L g8425 ( 
.A(n_7870),
.B(n_7314),
.Y(n_8425)
);

NOR2xp33_ASAP7_75t_L g8426 ( 
.A(n_8140),
.B(n_8102),
.Y(n_8426)
);

INVx1_ASAP7_75t_L g8427 ( 
.A(n_7874),
.Y(n_8427)
);

NAND2xp5_ASAP7_75t_SL g8428 ( 
.A(n_8060),
.B(n_7826),
.Y(n_8428)
);

INVxp67_ASAP7_75t_L g8429 ( 
.A(n_7905),
.Y(n_8429)
);

INVx1_ASAP7_75t_L g8430 ( 
.A(n_7881),
.Y(n_8430)
);

INVx1_ASAP7_75t_L g8431 ( 
.A(n_7883),
.Y(n_8431)
);

AND2x4_ASAP7_75t_L g8432 ( 
.A(n_7885),
.B(n_7677),
.Y(n_8432)
);

NAND2xp5_ASAP7_75t_L g8433 ( 
.A(n_7978),
.B(n_4930),
.Y(n_8433)
);

INVx1_ASAP7_75t_L g8434 ( 
.A(n_7884),
.Y(n_8434)
);

AOI22xp5_ASAP7_75t_L g8435 ( 
.A1(n_8077),
.A2(n_7579),
.B1(n_7799),
.B2(n_7851),
.Y(n_8435)
);

INVx1_ASAP7_75t_L g8436 ( 
.A(n_7887),
.Y(n_8436)
);

NAND2xp5_ASAP7_75t_SL g8437 ( 
.A(n_7860),
.B(n_4931),
.Y(n_8437)
);

AND2x2_ASAP7_75t_L g8438 ( 
.A(n_8146),
.B(n_4932),
.Y(n_8438)
);

INVx1_ASAP7_75t_L g8439 ( 
.A(n_7904),
.Y(n_8439)
);

BUFx3_ASAP7_75t_L g8440 ( 
.A(n_8067),
.Y(n_8440)
);

INVx1_ASAP7_75t_L g8441 ( 
.A(n_7909),
.Y(n_8441)
);

INVx1_ASAP7_75t_L g8442 ( 
.A(n_7927),
.Y(n_8442)
);

NAND2xp5_ASAP7_75t_SL g8443 ( 
.A(n_8201),
.B(n_4933),
.Y(n_8443)
);

BUFx10_ASAP7_75t_L g8444 ( 
.A(n_7923),
.Y(n_8444)
);

INVx1_ASAP7_75t_L g8445 ( 
.A(n_7931),
.Y(n_8445)
);

INVx2_ASAP7_75t_L g8446 ( 
.A(n_7920),
.Y(n_8446)
);

INVx1_ASAP7_75t_L g8447 ( 
.A(n_7932),
.Y(n_8447)
);

NOR2xp33_ASAP7_75t_L g8448 ( 
.A(n_8126),
.B(n_4934),
.Y(n_8448)
);

NOR2xp33_ASAP7_75t_L g8449 ( 
.A(n_8198),
.B(n_4936),
.Y(n_8449)
);

BUFx6f_ASAP7_75t_L g8450 ( 
.A(n_7914),
.Y(n_8450)
);

BUFx6f_ASAP7_75t_L g8451 ( 
.A(n_7914),
.Y(n_8451)
);

INVx2_ASAP7_75t_L g8452 ( 
.A(n_7922),
.Y(n_8452)
);

NOR2xp33_ASAP7_75t_L g8453 ( 
.A(n_8196),
.B(n_4937),
.Y(n_8453)
);

BUFx6f_ASAP7_75t_L g8454 ( 
.A(n_8004),
.Y(n_8454)
);

INVx1_ASAP7_75t_L g8455 ( 
.A(n_7933),
.Y(n_8455)
);

AND2x4_ASAP7_75t_L g8456 ( 
.A(n_7937),
.B(n_7733),
.Y(n_8456)
);

CKINVDCx5p33_ASAP7_75t_R g8457 ( 
.A(n_7987),
.Y(n_8457)
);

BUFx6f_ASAP7_75t_L g8458 ( 
.A(n_8004),
.Y(n_8458)
);

OR2x2_ASAP7_75t_L g8459 ( 
.A(n_8381),
.B(n_4942),
.Y(n_8459)
);

INVx1_ASAP7_75t_L g8460 ( 
.A(n_7948),
.Y(n_8460)
);

NAND2xp5_ASAP7_75t_L g8461 ( 
.A(n_8266),
.B(n_4943),
.Y(n_8461)
);

AO22x2_ASAP7_75t_L g8462 ( 
.A1(n_7911),
.A2(n_4906),
.B1(n_4908),
.B2(n_4900),
.Y(n_8462)
);

OR2x2_ASAP7_75t_L g8463 ( 
.A(n_7878),
.B(n_8372),
.Y(n_8463)
);

AND2x2_ASAP7_75t_L g8464 ( 
.A(n_7986),
.B(n_4947),
.Y(n_8464)
);

NAND2xp5_ASAP7_75t_SL g8465 ( 
.A(n_8342),
.B(n_4952),
.Y(n_8465)
);

AND2x4_ASAP7_75t_L g8466 ( 
.A(n_8154),
.B(n_4910),
.Y(n_8466)
);

INVx1_ASAP7_75t_L g8467 ( 
.A(n_7951),
.Y(n_8467)
);

BUFx3_ASAP7_75t_L g8468 ( 
.A(n_8189),
.Y(n_8468)
);

INVx1_ASAP7_75t_L g8469 ( 
.A(n_7955),
.Y(n_8469)
);

BUFx10_ASAP7_75t_L g8470 ( 
.A(n_8325),
.Y(n_8470)
);

INVx1_ASAP7_75t_L g8471 ( 
.A(n_7964),
.Y(n_8471)
);

INVx1_ASAP7_75t_L g8472 ( 
.A(n_7969),
.Y(n_8472)
);

INVx2_ASAP7_75t_L g8473 ( 
.A(n_7924),
.Y(n_8473)
);

CKINVDCx5p33_ASAP7_75t_R g8474 ( 
.A(n_8021),
.Y(n_8474)
);

NAND2xp5_ASAP7_75t_L g8475 ( 
.A(n_8343),
.B(n_4953),
.Y(n_8475)
);

BUFx6f_ASAP7_75t_L g8476 ( 
.A(n_8026),
.Y(n_8476)
);

INVx2_ASAP7_75t_L g8477 ( 
.A(n_7926),
.Y(n_8477)
);

BUFx6f_ASAP7_75t_L g8478 ( 
.A(n_8026),
.Y(n_8478)
);

INVx2_ASAP7_75t_L g8479 ( 
.A(n_7930),
.Y(n_8479)
);

NAND2xp5_ASAP7_75t_L g8480 ( 
.A(n_7974),
.B(n_7975),
.Y(n_8480)
);

INVx1_ASAP7_75t_L g8481 ( 
.A(n_7981),
.Y(n_8481)
);

NOR2xp33_ASAP7_75t_L g8482 ( 
.A(n_8215),
.B(n_4959),
.Y(n_8482)
);

INVx4_ASAP7_75t_L g8483 ( 
.A(n_8086),
.Y(n_8483)
);

INVx5_ASAP7_75t_L g8484 ( 
.A(n_8288),
.Y(n_8484)
);

NAND3x1_ASAP7_75t_L g8485 ( 
.A(n_8079),
.B(n_4928),
.C(n_4916),
.Y(n_8485)
);

NAND2xp5_ASAP7_75t_SL g8486 ( 
.A(n_8160),
.B(n_4961),
.Y(n_8486)
);

INVx2_ASAP7_75t_L g8487 ( 
.A(n_7934),
.Y(n_8487)
);

HB1xp67_ASAP7_75t_L g8488 ( 
.A(n_7965),
.Y(n_8488)
);

INVx2_ASAP7_75t_L g8489 ( 
.A(n_7936),
.Y(n_8489)
);

INVx1_ASAP7_75t_L g8490 ( 
.A(n_7990),
.Y(n_8490)
);

INVx1_ASAP7_75t_L g8491 ( 
.A(n_7992),
.Y(n_8491)
);

BUFx6f_ASAP7_75t_L g8492 ( 
.A(n_8086),
.Y(n_8492)
);

BUFx3_ASAP7_75t_L g8493 ( 
.A(n_7941),
.Y(n_8493)
);

NOR2xp33_ASAP7_75t_L g8494 ( 
.A(n_7862),
.B(n_4963),
.Y(n_8494)
);

INVx1_ASAP7_75t_L g8495 ( 
.A(n_7993),
.Y(n_8495)
);

NAND2xp5_ASAP7_75t_SL g8496 ( 
.A(n_8345),
.B(n_4969),
.Y(n_8496)
);

CKINVDCx5p33_ASAP7_75t_R g8497 ( 
.A(n_8135),
.Y(n_8497)
);

BUFx3_ASAP7_75t_L g8498 ( 
.A(n_7980),
.Y(n_8498)
);

INVx4_ASAP7_75t_L g8499 ( 
.A(n_8178),
.Y(n_8499)
);

AND2x6_ASAP7_75t_L g8500 ( 
.A(n_7893),
.B(n_4935),
.Y(n_8500)
);

BUFx3_ASAP7_75t_L g8501 ( 
.A(n_8178),
.Y(n_8501)
);

INVx1_ASAP7_75t_L g8502 ( 
.A(n_7997),
.Y(n_8502)
);

INVx1_ASAP7_75t_L g8503 ( 
.A(n_7999),
.Y(n_8503)
);

INVx8_ASAP7_75t_L g8504 ( 
.A(n_8034),
.Y(n_8504)
);

INVx6_ASAP7_75t_L g8505 ( 
.A(n_7940),
.Y(n_8505)
);

INVx1_ASAP7_75t_L g8506 ( 
.A(n_8003),
.Y(n_8506)
);

HB1xp67_ASAP7_75t_L g8507 ( 
.A(n_7973),
.Y(n_8507)
);

OR2x6_ASAP7_75t_L g8508 ( 
.A(n_8020),
.B(n_4939),
.Y(n_8508)
);

AND2x4_ASAP7_75t_L g8509 ( 
.A(n_8311),
.B(n_4940),
.Y(n_8509)
);

NAND2xp5_ASAP7_75t_L g8510 ( 
.A(n_8051),
.B(n_4971),
.Y(n_8510)
);

INVx2_ASAP7_75t_L g8511 ( 
.A(n_7938),
.Y(n_8511)
);

NAND2xp5_ASAP7_75t_L g8512 ( 
.A(n_8261),
.B(n_4972),
.Y(n_8512)
);

INVx1_ASAP7_75t_L g8513 ( 
.A(n_8005),
.Y(n_8513)
);

INVx2_ASAP7_75t_L g8514 ( 
.A(n_7939),
.Y(n_8514)
);

AND2x2_ASAP7_75t_L g8515 ( 
.A(n_8228),
.B(n_4973),
.Y(n_8515)
);

INVx1_ASAP7_75t_L g8516 ( 
.A(n_8015),
.Y(n_8516)
);

NOR2xp33_ASAP7_75t_L g8517 ( 
.A(n_7946),
.B(n_4976),
.Y(n_8517)
);

INVx2_ASAP7_75t_SL g8518 ( 
.A(n_7898),
.Y(n_8518)
);

AND2x4_ASAP7_75t_L g8519 ( 
.A(n_8326),
.B(n_8254),
.Y(n_8519)
);

AND2x4_ASAP7_75t_L g8520 ( 
.A(n_8255),
.B(n_4944),
.Y(n_8520)
);

AND2x2_ASAP7_75t_L g8521 ( 
.A(n_8262),
.B(n_8028),
.Y(n_8521)
);

AOI22xp33_ASAP7_75t_L g8522 ( 
.A1(n_7868),
.A2(n_5713),
.B1(n_5735),
.B2(n_5688),
.Y(n_8522)
);

INVx1_ASAP7_75t_L g8523 ( 
.A(n_8016),
.Y(n_8523)
);

CKINVDCx5p33_ASAP7_75t_R g8524 ( 
.A(n_8248),
.Y(n_8524)
);

AND2x4_ASAP7_75t_L g8525 ( 
.A(n_8259),
.B(n_4951),
.Y(n_8525)
);

INVx3_ASAP7_75t_L g8526 ( 
.A(n_8275),
.Y(n_8526)
);

NOR2xp33_ASAP7_75t_L g8527 ( 
.A(n_8265),
.B(n_4977),
.Y(n_8527)
);

INVx1_ASAP7_75t_L g8528 ( 
.A(n_8018),
.Y(n_8528)
);

OA22x2_ASAP7_75t_L g8529 ( 
.A1(n_7912),
.A2(n_4981),
.B1(n_4982),
.B2(n_4979),
.Y(n_8529)
);

INVx2_ASAP7_75t_SL g8530 ( 
.A(n_8022),
.Y(n_8530)
);

INVx4_ASAP7_75t_SL g8531 ( 
.A(n_8270),
.Y(n_8531)
);

NAND2xp5_ASAP7_75t_SL g8532 ( 
.A(n_7966),
.B(n_4983),
.Y(n_8532)
);

NAND3xp33_ASAP7_75t_L g8533 ( 
.A(n_7935),
.B(n_7894),
.C(n_8220),
.Y(n_8533)
);

NOR2xp33_ASAP7_75t_L g8534 ( 
.A(n_8222),
.B(n_4987),
.Y(n_8534)
);

NOR2xp33_ASAP7_75t_L g8535 ( 
.A(n_8226),
.B(n_4988),
.Y(n_8535)
);

INVx2_ASAP7_75t_L g8536 ( 
.A(n_7942),
.Y(n_8536)
);

NAND2xp5_ASAP7_75t_L g8537 ( 
.A(n_8109),
.B(n_4991),
.Y(n_8537)
);

AND2x6_ASAP7_75t_L g8538 ( 
.A(n_8209),
.B(n_4954),
.Y(n_8538)
);

INVx1_ASAP7_75t_L g8539 ( 
.A(n_7953),
.Y(n_8539)
);

INVx2_ASAP7_75t_L g8540 ( 
.A(n_7954),
.Y(n_8540)
);

BUFx2_ASAP7_75t_L g8541 ( 
.A(n_8027),
.Y(n_8541)
);

INVx1_ASAP7_75t_L g8542 ( 
.A(n_7957),
.Y(n_8542)
);

INVx3_ASAP7_75t_L g8543 ( 
.A(n_8275),
.Y(n_8543)
);

INVx1_ASAP7_75t_SL g8544 ( 
.A(n_8088),
.Y(n_8544)
);

BUFx6f_ASAP7_75t_L g8545 ( 
.A(n_8209),
.Y(n_8545)
);

INVx5_ASAP7_75t_L g8546 ( 
.A(n_8288),
.Y(n_8546)
);

AND2x4_ASAP7_75t_L g8547 ( 
.A(n_8104),
.B(n_4955),
.Y(n_8547)
);

INVx2_ASAP7_75t_L g8548 ( 
.A(n_7958),
.Y(n_8548)
);

OAI22xp33_ASAP7_75t_L g8549 ( 
.A1(n_8210),
.A2(n_4994),
.B1(n_4995),
.B2(n_4993),
.Y(n_8549)
);

INVx1_ASAP7_75t_L g8550 ( 
.A(n_7959),
.Y(n_8550)
);

AOI22xp33_ASAP7_75t_L g8551 ( 
.A1(n_7900),
.A2(n_5750),
.B1(n_4962),
.B2(n_4964),
.Y(n_8551)
);

NAND3x1_ASAP7_75t_L g8552 ( 
.A(n_8409),
.B(n_4966),
.C(n_4958),
.Y(n_8552)
);

INVx1_ASAP7_75t_L g8553 ( 
.A(n_7963),
.Y(n_8553)
);

BUFx6f_ASAP7_75t_L g8554 ( 
.A(n_8236),
.Y(n_8554)
);

AND2x2_ASAP7_75t_L g8555 ( 
.A(n_8075),
.B(n_4996),
.Y(n_8555)
);

INVx3_ASAP7_75t_L g8556 ( 
.A(n_7867),
.Y(n_8556)
);

NAND2xp5_ASAP7_75t_L g8557 ( 
.A(n_8095),
.B(n_4997),
.Y(n_8557)
);

NOR2xp33_ASAP7_75t_L g8558 ( 
.A(n_7891),
.B(n_4998),
.Y(n_8558)
);

AND2x2_ASAP7_75t_L g8559 ( 
.A(n_8137),
.B(n_5001),
.Y(n_8559)
);

NAND2xp5_ASAP7_75t_L g8560 ( 
.A(n_8082),
.B(n_7968),
.Y(n_8560)
);

OR2x6_ASAP7_75t_L g8561 ( 
.A(n_8020),
.B(n_4968),
.Y(n_8561)
);

INVx2_ASAP7_75t_L g8562 ( 
.A(n_7970),
.Y(n_8562)
);

AO22x2_ASAP7_75t_L g8563 ( 
.A1(n_8204),
.A2(n_4980),
.B1(n_4989),
.B2(n_4975),
.Y(n_8563)
);

INVx1_ASAP7_75t_L g8564 ( 
.A(n_7971),
.Y(n_8564)
);

INVx1_ASAP7_75t_L g8565 ( 
.A(n_7977),
.Y(n_8565)
);

BUFx3_ASAP7_75t_L g8566 ( 
.A(n_8236),
.Y(n_8566)
);

INVx3_ASAP7_75t_L g8567 ( 
.A(n_7892),
.Y(n_8567)
);

AND2x6_ASAP7_75t_L g8568 ( 
.A(n_8250),
.B(n_4992),
.Y(n_8568)
);

AO22x1_ASAP7_75t_L g8569 ( 
.A1(n_8090),
.A2(n_5004),
.B1(n_5006),
.B2(n_5002),
.Y(n_8569)
);

INVx1_ASAP7_75t_L g8570 ( 
.A(n_7979),
.Y(n_8570)
);

NAND2xp5_ASAP7_75t_SL g8571 ( 
.A(n_8066),
.B(n_5009),
.Y(n_8571)
);

AND2x2_ASAP7_75t_L g8572 ( 
.A(n_8035),
.B(n_5015),
.Y(n_8572)
);

INVx2_ASAP7_75t_SL g8573 ( 
.A(n_8083),
.Y(n_8573)
);

AND2x4_ASAP7_75t_L g8574 ( 
.A(n_8164),
.B(n_5003),
.Y(n_8574)
);

INVx1_ASAP7_75t_L g8575 ( 
.A(n_7983),
.Y(n_8575)
);

NAND2xp5_ASAP7_75t_SL g8576 ( 
.A(n_8046),
.B(n_5017),
.Y(n_8576)
);

INVx1_ASAP7_75t_L g8577 ( 
.A(n_7988),
.Y(n_8577)
);

INVx1_ASAP7_75t_L g8578 ( 
.A(n_7989),
.Y(n_8578)
);

BUFx2_ASAP7_75t_L g8579 ( 
.A(n_8107),
.Y(n_8579)
);

INVx5_ASAP7_75t_L g8580 ( 
.A(n_8316),
.Y(n_8580)
);

NOR2xp33_ASAP7_75t_L g8581 ( 
.A(n_7961),
.B(n_5018),
.Y(n_8581)
);

NAND2x1p5_ASAP7_75t_L g8582 ( 
.A(n_7902),
.B(n_5005),
.Y(n_8582)
);

BUFx3_ASAP7_75t_L g8583 ( 
.A(n_8250),
.Y(n_8583)
);

CKINVDCx5p33_ASAP7_75t_R g8584 ( 
.A(n_8132),
.Y(n_8584)
);

BUFx6f_ASAP7_75t_L g8585 ( 
.A(n_8252),
.Y(n_8585)
);

NAND2xp5_ASAP7_75t_L g8586 ( 
.A(n_7994),
.B(n_5019),
.Y(n_8586)
);

CKINVDCx16_ASAP7_75t_R g8587 ( 
.A(n_7888),
.Y(n_8587)
);

NOR2x1p5_ASAP7_75t_L g8588 ( 
.A(n_7967),
.B(n_5022),
.Y(n_8588)
);

NAND2xp5_ASAP7_75t_L g8589 ( 
.A(n_7998),
.B(n_5025),
.Y(n_8589)
);

INVx1_ASAP7_75t_L g8590 ( 
.A(n_8002),
.Y(n_8590)
);

INVx1_ASAP7_75t_L g8591 ( 
.A(n_8009),
.Y(n_8591)
);

AND2x6_ASAP7_75t_L g8592 ( 
.A(n_8252),
.B(n_5007),
.Y(n_8592)
);

AND2x2_ASAP7_75t_L g8593 ( 
.A(n_8057),
.B(n_5026),
.Y(n_8593)
);

INVx2_ASAP7_75t_SL g8594 ( 
.A(n_8260),
.Y(n_8594)
);

INVx2_ASAP7_75t_L g8595 ( 
.A(n_8011),
.Y(n_8595)
);

INVx2_ASAP7_75t_L g8596 ( 
.A(n_8013),
.Y(n_8596)
);

NOR2xp33_ASAP7_75t_L g8597 ( 
.A(n_7918),
.B(n_8084),
.Y(n_8597)
);

BUFx3_ASAP7_75t_L g8598 ( 
.A(n_8260),
.Y(n_8598)
);

INVx2_ASAP7_75t_SL g8599 ( 
.A(n_8272),
.Y(n_8599)
);

INVx1_ASAP7_75t_L g8600 ( 
.A(n_8149),
.Y(n_8600)
);

AND2x6_ASAP7_75t_L g8601 ( 
.A(n_8374),
.B(n_5011),
.Y(n_8601)
);

BUFx6f_ASAP7_75t_L g8602 ( 
.A(n_8316),
.Y(n_8602)
);

INVx1_ASAP7_75t_L g8603 ( 
.A(n_8152),
.Y(n_8603)
);

BUFx10_ASAP7_75t_L g8604 ( 
.A(n_8378),
.Y(n_8604)
);

INVx4_ASAP7_75t_L g8605 ( 
.A(n_7950),
.Y(n_8605)
);

INVx1_ASAP7_75t_L g8606 ( 
.A(n_8156),
.Y(n_8606)
);

INVx1_ASAP7_75t_L g8607 ( 
.A(n_8158),
.Y(n_8607)
);

NAND2xp5_ASAP7_75t_SL g8608 ( 
.A(n_8363),
.B(n_5030),
.Y(n_8608)
);

INVx1_ASAP7_75t_L g8609 ( 
.A(n_8170),
.Y(n_8609)
);

NAND2xp5_ASAP7_75t_L g8610 ( 
.A(n_7900),
.B(n_5033),
.Y(n_8610)
);

INVxp67_ASAP7_75t_SL g8611 ( 
.A(n_8306),
.Y(n_8611)
);

INVx1_ASAP7_75t_L g8612 ( 
.A(n_8174),
.Y(n_8612)
);

BUFx10_ASAP7_75t_L g8613 ( 
.A(n_8141),
.Y(n_8613)
);

INVx1_ASAP7_75t_L g8614 ( 
.A(n_8175),
.Y(n_8614)
);

NAND2x1p5_ASAP7_75t_L g8615 ( 
.A(n_7956),
.B(n_5013),
.Y(n_8615)
);

BUFx6f_ASAP7_75t_L g8616 ( 
.A(n_7950),
.Y(n_8616)
);

NOR2xp33_ASAP7_75t_L g8617 ( 
.A(n_8386),
.B(n_5036),
.Y(n_8617)
);

AOI22xp33_ASAP7_75t_L g8618 ( 
.A1(n_7900),
.A2(n_5021),
.B1(n_5023),
.B2(n_5014),
.Y(n_8618)
);

NAND3xp33_ASAP7_75t_L g8619 ( 
.A(n_8256),
.B(n_5038),
.C(n_5037),
.Y(n_8619)
);

AND2x4_ASAP7_75t_L g8620 ( 
.A(n_8179),
.B(n_5028),
.Y(n_8620)
);

INVx1_ASAP7_75t_L g8621 ( 
.A(n_8183),
.Y(n_8621)
);

NAND2xp5_ASAP7_75t_L g8622 ( 
.A(n_7899),
.B(n_5039),
.Y(n_8622)
);

INVx2_ASAP7_75t_L g8623 ( 
.A(n_8232),
.Y(n_8623)
);

INVx1_ASAP7_75t_L g8624 ( 
.A(n_8031),
.Y(n_8624)
);

INVx3_ASAP7_75t_L g8625 ( 
.A(n_8044),
.Y(n_8625)
);

INVx1_ASAP7_75t_L g8626 ( 
.A(n_8037),
.Y(n_8626)
);

INVx2_ASAP7_75t_L g8627 ( 
.A(n_8234),
.Y(n_8627)
);

BUFx2_ASAP7_75t_L g8628 ( 
.A(n_8151),
.Y(n_8628)
);

NAND2xp5_ASAP7_75t_SL g8629 ( 
.A(n_8322),
.B(n_5041),
.Y(n_8629)
);

AND2x6_ASAP7_75t_L g8630 ( 
.A(n_8375),
.B(n_5029),
.Y(n_8630)
);

INVx1_ASAP7_75t_L g8631 ( 
.A(n_8042),
.Y(n_8631)
);

INVx2_ASAP7_75t_L g8632 ( 
.A(n_8243),
.Y(n_8632)
);

INVx2_ASAP7_75t_L g8633 ( 
.A(n_8281),
.Y(n_8633)
);

NAND2xp5_ASAP7_75t_SL g8634 ( 
.A(n_8361),
.B(n_5043),
.Y(n_8634)
);

AOI22xp33_ASAP7_75t_L g8635 ( 
.A1(n_8070),
.A2(n_5035),
.B1(n_5042),
.B2(n_5032),
.Y(n_8635)
);

INVx1_ASAP7_75t_L g8636 ( 
.A(n_8047),
.Y(n_8636)
);

NAND2xp5_ASAP7_75t_SL g8637 ( 
.A(n_8370),
.B(n_5044),
.Y(n_8637)
);

AND2x6_ASAP7_75t_L g8638 ( 
.A(n_8373),
.B(n_5054),
.Y(n_8638)
);

NAND2xp5_ASAP7_75t_L g8639 ( 
.A(n_7925),
.B(n_7943),
.Y(n_8639)
);

BUFx8_ASAP7_75t_SL g8640 ( 
.A(n_8396),
.Y(n_8640)
);

INVx1_ASAP7_75t_L g8641 ( 
.A(n_8048),
.Y(n_8641)
);

INVx1_ASAP7_75t_L g8642 ( 
.A(n_8055),
.Y(n_8642)
);

AND2x2_ASAP7_75t_L g8643 ( 
.A(n_7976),
.B(n_5045),
.Y(n_8643)
);

INVx1_ASAP7_75t_L g8644 ( 
.A(n_8061),
.Y(n_8644)
);

AND2x2_ASAP7_75t_L g8645 ( 
.A(n_8377),
.B(n_5047),
.Y(n_8645)
);

AND2x4_ASAP7_75t_L g8646 ( 
.A(n_8235),
.B(n_5059),
.Y(n_8646)
);

OR2x2_ASAP7_75t_L g8647 ( 
.A(n_8351),
.B(n_5048),
.Y(n_8647)
);

CKINVDCx5p33_ASAP7_75t_R g8648 ( 
.A(n_7960),
.Y(n_8648)
);

NAND2xp5_ASAP7_75t_SL g8649 ( 
.A(n_8289),
.B(n_5050),
.Y(n_8649)
);

AND2x2_ASAP7_75t_L g8650 ( 
.A(n_8085),
.B(n_5051),
.Y(n_8650)
);

INVxp33_ASAP7_75t_L g8651 ( 
.A(n_8389),
.Y(n_8651)
);

INVx2_ASAP7_75t_L g8652 ( 
.A(n_7861),
.Y(n_8652)
);

INVx1_ASAP7_75t_L g8653 ( 
.A(n_8068),
.Y(n_8653)
);

INVx2_ASAP7_75t_L g8654 ( 
.A(n_7865),
.Y(n_8654)
);

BUFx6f_ASAP7_75t_L g8655 ( 
.A(n_8327),
.Y(n_8655)
);

INVx4_ASAP7_75t_L g8656 ( 
.A(n_8093),
.Y(n_8656)
);

BUFx6f_ASAP7_75t_L g8657 ( 
.A(n_8327),
.Y(n_8657)
);

INVx1_ASAP7_75t_L g8658 ( 
.A(n_8071),
.Y(n_8658)
);

INVx3_ASAP7_75t_L g8659 ( 
.A(n_8108),
.Y(n_8659)
);

INVx2_ASAP7_75t_L g8660 ( 
.A(n_7866),
.Y(n_8660)
);

NOR2x1p5_ASAP7_75t_L g8661 ( 
.A(n_8099),
.B(n_5052),
.Y(n_8661)
);

BUFx6f_ASAP7_75t_L g8662 ( 
.A(n_8193),
.Y(n_8662)
);

NAND2xp5_ASAP7_75t_L g8663 ( 
.A(n_8124),
.B(n_5055),
.Y(n_8663)
);

BUFx2_ASAP7_75t_L g8664 ( 
.A(n_8348),
.Y(n_8664)
);

INVx2_ASAP7_75t_L g8665 ( 
.A(n_7871),
.Y(n_8665)
);

NAND2xp5_ASAP7_75t_SL g8666 ( 
.A(n_8362),
.B(n_5057),
.Y(n_8666)
);

AND2x2_ASAP7_75t_L g8667 ( 
.A(n_7985),
.B(n_5060),
.Y(n_8667)
);

NAND2xp5_ASAP7_75t_L g8668 ( 
.A(n_8117),
.B(n_5063),
.Y(n_8668)
);

CKINVDCx11_ASAP7_75t_R g8669 ( 
.A(n_8136),
.Y(n_8669)
);

INVx3_ASAP7_75t_L g8670 ( 
.A(n_8130),
.Y(n_8670)
);

INVx2_ASAP7_75t_L g8671 ( 
.A(n_7876),
.Y(n_8671)
);

INVx2_ASAP7_75t_L g8672 ( 
.A(n_7877),
.Y(n_8672)
);

INVx1_ASAP7_75t_L g8673 ( 
.A(n_8087),
.Y(n_8673)
);

INVx2_ASAP7_75t_L g8674 ( 
.A(n_7879),
.Y(n_8674)
);

INVx1_ASAP7_75t_L g8675 ( 
.A(n_8091),
.Y(n_8675)
);

BUFx6f_ASAP7_75t_L g8676 ( 
.A(n_8264),
.Y(n_8676)
);

INVx1_ASAP7_75t_L g8677 ( 
.A(n_8094),
.Y(n_8677)
);

INVx1_ASAP7_75t_L g8678 ( 
.A(n_8096),
.Y(n_8678)
);

NAND2xp5_ASAP7_75t_L g8679 ( 
.A(n_8258),
.B(n_5064),
.Y(n_8679)
);

INVxp33_ASAP7_75t_L g8680 ( 
.A(n_8125),
.Y(n_8680)
);

NAND2xp5_ASAP7_75t_SL g8681 ( 
.A(n_8240),
.B(n_5065),
.Y(n_8681)
);

INVx2_ASAP7_75t_L g8682 ( 
.A(n_7880),
.Y(n_8682)
);

INVx1_ASAP7_75t_L g8683 ( 
.A(n_8097),
.Y(n_8683)
);

NAND2xp5_ASAP7_75t_SL g8684 ( 
.A(n_8271),
.B(n_5068),
.Y(n_8684)
);

INVx2_ASAP7_75t_L g8685 ( 
.A(n_7889),
.Y(n_8685)
);

NAND2xp5_ASAP7_75t_L g8686 ( 
.A(n_8364),
.B(n_5073),
.Y(n_8686)
);

INVx4_ASAP7_75t_L g8687 ( 
.A(n_8038),
.Y(n_8687)
);

INVxp33_ASAP7_75t_L g8688 ( 
.A(n_7991),
.Y(n_8688)
);

INVx1_ASAP7_75t_L g8689 ( 
.A(n_8103),
.Y(n_8689)
);

AND2x4_ASAP7_75t_L g8690 ( 
.A(n_8310),
.B(n_5069),
.Y(n_8690)
);

HB1xp67_ASAP7_75t_L g8691 ( 
.A(n_8380),
.Y(n_8691)
);

INVx2_ASAP7_75t_L g8692 ( 
.A(n_7896),
.Y(n_8692)
);

AND2x2_ASAP7_75t_L g8693 ( 
.A(n_8110),
.B(n_5075),
.Y(n_8693)
);

INVx2_ASAP7_75t_L g8694 ( 
.A(n_7901),
.Y(n_8694)
);

INVx4_ASAP7_75t_L g8695 ( 
.A(n_8089),
.Y(n_8695)
);

INVx1_ASAP7_75t_L g8696 ( 
.A(n_8111),
.Y(n_8696)
);

NAND2xp33_ASAP7_75t_SL g8697 ( 
.A(n_8229),
.B(n_5076),
.Y(n_8697)
);

INVx1_ASAP7_75t_L g8698 ( 
.A(n_8120),
.Y(n_8698)
);

NOR2xp33_ASAP7_75t_L g8699 ( 
.A(n_8101),
.B(n_5077),
.Y(n_8699)
);

NAND2xp5_ASAP7_75t_L g8700 ( 
.A(n_7996),
.B(n_5078),
.Y(n_8700)
);

INVx2_ASAP7_75t_L g8701 ( 
.A(n_7903),
.Y(n_8701)
);

INVx1_ASAP7_75t_L g8702 ( 
.A(n_8139),
.Y(n_8702)
);

AND2x6_ASAP7_75t_L g8703 ( 
.A(n_8216),
.B(n_8307),
.Y(n_8703)
);

NAND2xp5_ASAP7_75t_SL g8704 ( 
.A(n_8283),
.B(n_5079),
.Y(n_8704)
);

CKINVDCx16_ASAP7_75t_R g8705 ( 
.A(n_8279),
.Y(n_8705)
);

INVx3_ASAP7_75t_L g8706 ( 
.A(n_8049),
.Y(n_8706)
);

OR2x6_ASAP7_75t_L g8707 ( 
.A(n_8321),
.B(n_5072),
.Y(n_8707)
);

INVx1_ASAP7_75t_L g8708 ( 
.A(n_8147),
.Y(n_8708)
);

NAND3xp33_ASAP7_75t_L g8709 ( 
.A(n_8339),
.B(n_5082),
.C(n_5081),
.Y(n_8709)
);

INVx1_ASAP7_75t_L g8710 ( 
.A(n_8185),
.Y(n_8710)
);

INVx2_ASAP7_75t_L g8711 ( 
.A(n_7906),
.Y(n_8711)
);

INVx1_ASAP7_75t_L g8712 ( 
.A(n_8159),
.Y(n_8712)
);

INVx1_ASAP7_75t_L g8713 ( 
.A(n_8162),
.Y(n_8713)
);

INVx2_ASAP7_75t_SL g8714 ( 
.A(n_8115),
.Y(n_8714)
);

INVx1_ASAP7_75t_L g8715 ( 
.A(n_8163),
.Y(n_8715)
);

NAND2xp33_ASAP7_75t_L g8716 ( 
.A(n_8070),
.B(n_5083),
.Y(n_8716)
);

CKINVDCx5p33_ASAP7_75t_R g8717 ( 
.A(n_8413),
.Y(n_8717)
);

INVx5_ASAP7_75t_L g8718 ( 
.A(n_8080),
.Y(n_8718)
);

INVx1_ASAP7_75t_L g8719 ( 
.A(n_8167),
.Y(n_8719)
);

OR2x2_ASAP7_75t_L g8720 ( 
.A(n_8388),
.B(n_5084),
.Y(n_8720)
);

NAND2xp5_ASAP7_75t_L g8721 ( 
.A(n_8001),
.B(n_5085),
.Y(n_8721)
);

NAND2xp5_ASAP7_75t_SL g8722 ( 
.A(n_8039),
.B(n_5086),
.Y(n_8722)
);

INVx1_ASAP7_75t_L g8723 ( 
.A(n_8172),
.Y(n_8723)
);

OR2x6_ASAP7_75t_L g8724 ( 
.A(n_8231),
.B(n_5090),
.Y(n_8724)
);

INVx2_ASAP7_75t_SL g8725 ( 
.A(n_8121),
.Y(n_8725)
);

INVx1_ASAP7_75t_L g8726 ( 
.A(n_8181),
.Y(n_8726)
);

AND2x2_ASAP7_75t_SL g8727 ( 
.A(n_8267),
.B(n_5091),
.Y(n_8727)
);

NAND2xp5_ASAP7_75t_SL g8728 ( 
.A(n_8043),
.B(n_5087),
.Y(n_8728)
);

NAND2x1p5_ASAP7_75t_L g8729 ( 
.A(n_7864),
.B(n_5097),
.Y(n_8729)
);

NOR2xp33_ASAP7_75t_L g8730 ( 
.A(n_8376),
.B(n_5089),
.Y(n_8730)
);

INVx3_ASAP7_75t_L g8731 ( 
.A(n_8133),
.Y(n_8731)
);

BUFx3_ASAP7_75t_L g8732 ( 
.A(n_8127),
.Y(n_8732)
);

INVx1_ASAP7_75t_L g8733 ( 
.A(n_8184),
.Y(n_8733)
);

INVx4_ASAP7_75t_SL g8734 ( 
.A(n_8346),
.Y(n_8734)
);

INVx1_ASAP7_75t_L g8735 ( 
.A(n_7907),
.Y(n_8735)
);

INVx1_ASAP7_75t_L g8736 ( 
.A(n_7908),
.Y(n_8736)
);

NAND2x1p5_ASAP7_75t_L g8737 ( 
.A(n_7875),
.B(n_7917),
.Y(n_8737)
);

BUFx2_ASAP7_75t_L g8738 ( 
.A(n_8312),
.Y(n_8738)
);

INVx2_ASAP7_75t_L g8739 ( 
.A(n_7913),
.Y(n_8739)
);

INVxp33_ASAP7_75t_L g8740 ( 
.A(n_8040),
.Y(n_8740)
);

AND2x4_ASAP7_75t_L g8741 ( 
.A(n_8092),
.B(n_5099),
.Y(n_8741)
);

INVx1_ASAP7_75t_L g8742 ( 
.A(n_8023),
.Y(n_8742)
);

NAND2xp5_ASAP7_75t_SL g8743 ( 
.A(n_8036),
.B(n_5093),
.Y(n_8743)
);

AND2x2_ASAP7_75t_L g8744 ( 
.A(n_8074),
.B(n_5094),
.Y(n_8744)
);

INVx2_ASAP7_75t_L g8745 ( 
.A(n_8024),
.Y(n_8745)
);

NOR2xp33_ASAP7_75t_L g8746 ( 
.A(n_8285),
.B(n_5095),
.Y(n_8746)
);

INVx1_ASAP7_75t_L g8747 ( 
.A(n_8025),
.Y(n_8747)
);

INVx1_ASAP7_75t_L g8748 ( 
.A(n_8033),
.Y(n_8748)
);

INVx1_ASAP7_75t_L g8749 ( 
.A(n_8050),
.Y(n_8749)
);

NAND2xp5_ASAP7_75t_SL g8750 ( 
.A(n_8036),
.B(n_5096),
.Y(n_8750)
);

AND2x2_ASAP7_75t_L g8751 ( 
.A(n_8045),
.B(n_5098),
.Y(n_8751)
);

NAND2xp5_ASAP7_75t_SL g8752 ( 
.A(n_8349),
.B(n_5100),
.Y(n_8752)
);

AND2x4_ASAP7_75t_L g8753 ( 
.A(n_8237),
.B(n_5106),
.Y(n_8753)
);

CKINVDCx5p33_ASAP7_75t_R g8754 ( 
.A(n_8394),
.Y(n_8754)
);

INVx2_ASAP7_75t_L g8755 ( 
.A(n_8053),
.Y(n_8755)
);

CKINVDCx5p33_ASAP7_75t_R g8756 ( 
.A(n_8177),
.Y(n_8756)
);

INVx2_ASAP7_75t_L g8757 ( 
.A(n_8054),
.Y(n_8757)
);

CKINVDCx6p67_ASAP7_75t_R g8758 ( 
.A(n_8186),
.Y(n_8758)
);

INVx4_ASAP7_75t_SL g8759 ( 
.A(n_8356),
.Y(n_8759)
);

BUFx2_ASAP7_75t_L g8760 ( 
.A(n_8165),
.Y(n_8760)
);

INVx1_ASAP7_75t_L g8761 ( 
.A(n_8056),
.Y(n_8761)
);

INVx2_ASAP7_75t_L g8762 ( 
.A(n_8058),
.Y(n_8762)
);

INVx1_ASAP7_75t_L g8763 ( 
.A(n_8062),
.Y(n_8763)
);

INVx2_ASAP7_75t_SL g8764 ( 
.A(n_8238),
.Y(n_8764)
);

INVx4_ASAP7_75t_L g8765 ( 
.A(n_8239),
.Y(n_8765)
);

INVx4_ASAP7_75t_L g8766 ( 
.A(n_7945),
.Y(n_8766)
);

INVx1_ASAP7_75t_L g8767 ( 
.A(n_8063),
.Y(n_8767)
);

OR2x2_ASAP7_75t_L g8768 ( 
.A(n_8166),
.B(n_5101),
.Y(n_8768)
);

BUFx10_ASAP7_75t_L g8769 ( 
.A(n_8291),
.Y(n_8769)
);

INVx2_ASAP7_75t_L g8770 ( 
.A(n_8064),
.Y(n_8770)
);

NAND2xp5_ASAP7_75t_SL g8771 ( 
.A(n_8131),
.B(n_5103),
.Y(n_8771)
);

AND2x2_ASAP7_75t_L g8772 ( 
.A(n_8171),
.B(n_5105),
.Y(n_8772)
);

AND2x4_ASAP7_75t_L g8773 ( 
.A(n_8244),
.B(n_5108),
.Y(n_8773)
);

NAND2xp5_ASAP7_75t_L g8774 ( 
.A(n_8224),
.B(n_5110),
.Y(n_8774)
);

NAND2xp5_ASAP7_75t_L g8775 ( 
.A(n_8253),
.B(n_5113),
.Y(n_8775)
);

AND2x2_ASAP7_75t_SL g8776 ( 
.A(n_8406),
.B(n_5111),
.Y(n_8776)
);

INVx2_ASAP7_75t_SL g8777 ( 
.A(n_7947),
.Y(n_8777)
);

INVx2_ASAP7_75t_L g8778 ( 
.A(n_8065),
.Y(n_8778)
);

AND2x4_ASAP7_75t_L g8779 ( 
.A(n_8251),
.B(n_5112),
.Y(n_8779)
);

INVx1_ASAP7_75t_L g8780 ( 
.A(n_8072),
.Y(n_8780)
);

INVxp67_ASAP7_75t_L g8781 ( 
.A(n_7910),
.Y(n_8781)
);

AND2x2_ASAP7_75t_L g8782 ( 
.A(n_8118),
.B(n_8052),
.Y(n_8782)
);

INVx4_ASAP7_75t_L g8783 ( 
.A(n_8000),
.Y(n_8783)
);

BUFx6f_ASAP7_75t_L g8784 ( 
.A(n_8006),
.Y(n_8784)
);

AOI22xp5_ASAP7_75t_L g8785 ( 
.A1(n_8219),
.A2(n_5121),
.B1(n_5123),
.B2(n_5120),
.Y(n_8785)
);

INVx3_ASAP7_75t_L g8786 ( 
.A(n_8182),
.Y(n_8786)
);

INVx3_ASAP7_75t_L g8787 ( 
.A(n_8008),
.Y(n_8787)
);

NAND2xp5_ASAP7_75t_L g8788 ( 
.A(n_8070),
.B(n_8225),
.Y(n_8788)
);

INVx2_ASAP7_75t_L g8789 ( 
.A(n_8081),
.Y(n_8789)
);

INVx1_ASAP7_75t_L g8790 ( 
.A(n_8100),
.Y(n_8790)
);

BUFx8_ASAP7_75t_SL g8791 ( 
.A(n_8393),
.Y(n_8791)
);

INVx1_ASAP7_75t_L g8792 ( 
.A(n_8106),
.Y(n_8792)
);

INVx3_ASAP7_75t_L g8793 ( 
.A(n_8280),
.Y(n_8793)
);

OAI21xp33_ASAP7_75t_L g8794 ( 
.A1(n_8318),
.A2(n_5128),
.B(n_5124),
.Y(n_8794)
);

INVx3_ASAP7_75t_L g8795 ( 
.A(n_8296),
.Y(n_8795)
);

NAND2xp5_ASAP7_75t_SL g8796 ( 
.A(n_8007),
.B(n_5130),
.Y(n_8796)
);

INVx2_ASAP7_75t_L g8797 ( 
.A(n_8114),
.Y(n_8797)
);

BUFx4_ASAP7_75t_L g8798 ( 
.A(n_8397),
.Y(n_8798)
);

INVx1_ASAP7_75t_L g8799 ( 
.A(n_8116),
.Y(n_8799)
);

OR2x2_ASAP7_75t_L g8800 ( 
.A(n_8390),
.B(n_5131),
.Y(n_8800)
);

INVx2_ASAP7_75t_L g8801 ( 
.A(n_8119),
.Y(n_8801)
);

NOR3xp33_ASAP7_75t_L g8802 ( 
.A(n_8336),
.B(n_5133),
.C(n_5132),
.Y(n_8802)
);

NAND2xp5_ASAP7_75t_L g8803 ( 
.A(n_8365),
.B(n_5137),
.Y(n_8803)
);

AND2x4_ASAP7_75t_L g8804 ( 
.A(n_7886),
.B(n_5114),
.Y(n_8804)
);

INVx1_ASAP7_75t_L g8805 ( 
.A(n_8122),
.Y(n_8805)
);

INVx1_ASAP7_75t_L g8806 ( 
.A(n_8129),
.Y(n_8806)
);

BUFx6f_ASAP7_75t_L g8807 ( 
.A(n_8302),
.Y(n_8807)
);

NAND2xp5_ASAP7_75t_L g8808 ( 
.A(n_8366),
.B(n_5138),
.Y(n_8808)
);

NAND2xp5_ASAP7_75t_L g8809 ( 
.A(n_8335),
.B(n_5149),
.Y(n_8809)
);

BUFx6f_ASAP7_75t_L g8810 ( 
.A(n_8284),
.Y(n_8810)
);

BUFx6f_ASAP7_75t_L g8811 ( 
.A(n_8331),
.Y(n_8811)
);

INVx3_ASAP7_75t_L g8812 ( 
.A(n_8301),
.Y(n_8812)
);

AND2x6_ASAP7_75t_L g8813 ( 
.A(n_8227),
.B(n_5116),
.Y(n_8813)
);

NOR2xp33_ASAP7_75t_L g8814 ( 
.A(n_8202),
.B(n_5150),
.Y(n_8814)
);

INVx1_ASAP7_75t_L g8815 ( 
.A(n_8138),
.Y(n_8815)
);

NAND2xp5_ASAP7_75t_SL g8816 ( 
.A(n_8323),
.B(n_5154),
.Y(n_8816)
);

BUFx10_ASAP7_75t_L g8817 ( 
.A(n_8411),
.Y(n_8817)
);

INVx1_ASAP7_75t_L g8818 ( 
.A(n_8144),
.Y(n_8818)
);

INVx1_ASAP7_75t_L g8819 ( 
.A(n_8145),
.Y(n_8819)
);

BUFx6f_ASAP7_75t_L g8820 ( 
.A(n_8360),
.Y(n_8820)
);

AND2x4_ASAP7_75t_L g8821 ( 
.A(n_8069),
.B(n_5119),
.Y(n_8821)
);

AND2x4_ASAP7_75t_L g8822 ( 
.A(n_8205),
.B(n_8305),
.Y(n_8822)
);

BUFx6f_ASAP7_75t_L g8823 ( 
.A(n_8317),
.Y(n_8823)
);

INVx3_ASAP7_75t_L g8824 ( 
.A(n_8350),
.Y(n_8824)
);

AND2x2_ASAP7_75t_L g8825 ( 
.A(n_8391),
.B(n_5156),
.Y(n_8825)
);

AND2x6_ASAP7_75t_L g8826 ( 
.A(n_8190),
.B(n_8347),
.Y(n_8826)
);

BUFx6f_ASAP7_75t_L g8827 ( 
.A(n_8313),
.Y(n_8827)
);

INVx2_ASAP7_75t_L g8828 ( 
.A(n_8150),
.Y(n_8828)
);

INVx1_ASAP7_75t_SL g8829 ( 
.A(n_8176),
.Y(n_8829)
);

INVx2_ASAP7_75t_L g8830 ( 
.A(n_8153),
.Y(n_8830)
);

INVx1_ASAP7_75t_L g8831 ( 
.A(n_8230),
.Y(n_8831)
);

INVx2_ASAP7_75t_L g8832 ( 
.A(n_8157),
.Y(n_8832)
);

BUFx2_ASAP7_75t_L g8833 ( 
.A(n_8392),
.Y(n_8833)
);

OR2x2_ASAP7_75t_L g8834 ( 
.A(n_8412),
.B(n_5158),
.Y(n_8834)
);

INVx1_ASAP7_75t_L g8835 ( 
.A(n_8233),
.Y(n_8835)
);

INVx3_ASAP7_75t_L g8836 ( 
.A(n_8314),
.Y(n_8836)
);

BUFx2_ASAP7_75t_L g8837 ( 
.A(n_8340),
.Y(n_8837)
);

AND2x4_ASAP7_75t_L g8838 ( 
.A(n_8315),
.B(n_5122),
.Y(n_8838)
);

INVx2_ASAP7_75t_L g8839 ( 
.A(n_8187),
.Y(n_8839)
);

INVx2_ASAP7_75t_L g8840 ( 
.A(n_8188),
.Y(n_8840)
);

AND2x2_ASAP7_75t_L g8841 ( 
.A(n_8029),
.B(n_5162),
.Y(n_8841)
);

AND2x6_ASAP7_75t_L g8842 ( 
.A(n_8353),
.B(n_5126),
.Y(n_8842)
);

INVx2_ASAP7_75t_L g8843 ( 
.A(n_8191),
.Y(n_8843)
);

INVx1_ASAP7_75t_L g8844 ( 
.A(n_8194),
.Y(n_8844)
);

INVx5_ASAP7_75t_L g8845 ( 
.A(n_8399),
.Y(n_8845)
);

BUFx3_ASAP7_75t_L g8846 ( 
.A(n_8382),
.Y(n_8846)
);

NOR2xp33_ASAP7_75t_L g8847 ( 
.A(n_8030),
.B(n_5167),
.Y(n_8847)
);

NOR2x1p5_ASAP7_75t_L g8848 ( 
.A(n_8369),
.B(n_8404),
.Y(n_8848)
);

INVx2_ASAP7_75t_L g8849 ( 
.A(n_8195),
.Y(n_8849)
);

NAND2xp5_ASAP7_75t_SL g8850 ( 
.A(n_8329),
.B(n_5170),
.Y(n_8850)
);

INVx1_ASAP7_75t_L g8851 ( 
.A(n_8148),
.Y(n_8851)
);

NAND2xp5_ASAP7_75t_SL g8852 ( 
.A(n_8197),
.B(n_8200),
.Y(n_8852)
);

AND2x2_ASAP7_75t_L g8853 ( 
.A(n_8041),
.B(n_5172),
.Y(n_8853)
);

INVx2_ASAP7_75t_L g8854 ( 
.A(n_8206),
.Y(n_8854)
);

AOI22xp33_ASAP7_75t_L g8855 ( 
.A1(n_8400),
.A2(n_5136),
.B1(n_5142),
.B2(n_5129),
.Y(n_8855)
);

AND2x4_ASAP7_75t_L g8856 ( 
.A(n_8320),
.B(n_5143),
.Y(n_8856)
);

BUFx6f_ASAP7_75t_L g8857 ( 
.A(n_8330),
.Y(n_8857)
);

INVx1_ASAP7_75t_SL g8858 ( 
.A(n_8384),
.Y(n_8858)
);

AND2x4_ASAP7_75t_L g8859 ( 
.A(n_8332),
.B(n_5145),
.Y(n_8859)
);

BUFx3_ASAP7_75t_L g8860 ( 
.A(n_8385),
.Y(n_8860)
);

INVx5_ASAP7_75t_L g8861 ( 
.A(n_8340),
.Y(n_8861)
);

INVx5_ASAP7_75t_L g8862 ( 
.A(n_8340),
.Y(n_8862)
);

BUFx6f_ASAP7_75t_L g8863 ( 
.A(n_8333),
.Y(n_8863)
);

INVx1_ASAP7_75t_L g8864 ( 
.A(n_8207),
.Y(n_8864)
);

NAND2xp5_ASAP7_75t_SL g8865 ( 
.A(n_8208),
.B(n_5175),
.Y(n_8865)
);

INVx1_ASAP7_75t_L g8866 ( 
.A(n_8211),
.Y(n_8866)
);

NAND2x1p5_ASAP7_75t_L g8867 ( 
.A(n_8328),
.B(n_5146),
.Y(n_8867)
);

OR2x2_ASAP7_75t_SL g8868 ( 
.A(n_8395),
.B(n_5147),
.Y(n_8868)
);

HB1xp67_ASAP7_75t_L g8869 ( 
.A(n_8276),
.Y(n_8869)
);

NAND2xp5_ASAP7_75t_L g8870 ( 
.A(n_8242),
.B(n_5176),
.Y(n_8870)
);

AND2x4_ASAP7_75t_L g8871 ( 
.A(n_8337),
.B(n_5148),
.Y(n_8871)
);

NAND2xp5_ASAP7_75t_SL g8872 ( 
.A(n_8213),
.B(n_8245),
.Y(n_8872)
);

AOI22xp5_ASAP7_75t_L g8873 ( 
.A1(n_8246),
.A2(n_5178),
.B1(n_5179),
.B2(n_5177),
.Y(n_8873)
);

INVx1_ASAP7_75t_L g8874 ( 
.A(n_8223),
.Y(n_8874)
);

INVx1_ASAP7_75t_L g8875 ( 
.A(n_8214),
.Y(n_8875)
);

NAND2xp5_ASAP7_75t_SL g8876 ( 
.A(n_8371),
.B(n_8098),
.Y(n_8876)
);

BUFx2_ASAP7_75t_L g8877 ( 
.A(n_8341),
.Y(n_8877)
);

NAND2xp5_ASAP7_75t_L g8878 ( 
.A(n_7952),
.B(n_5180),
.Y(n_8878)
);

INVx1_ASAP7_75t_L g8879 ( 
.A(n_8218),
.Y(n_8879)
);

INVx1_ASAP7_75t_SL g8880 ( 
.A(n_8282),
.Y(n_8880)
);

INVx2_ASAP7_75t_L g8881 ( 
.A(n_8221),
.Y(n_8881)
);

NAND2xp5_ASAP7_75t_L g8882 ( 
.A(n_7995),
.B(n_5181),
.Y(n_8882)
);

INVxp67_ASAP7_75t_L g8883 ( 
.A(n_7962),
.Y(n_8883)
);

OR2x6_ASAP7_75t_L g8884 ( 
.A(n_8401),
.B(n_5152),
.Y(n_8884)
);

INVx1_ASAP7_75t_L g8885 ( 
.A(n_8292),
.Y(n_8885)
);

INVx1_ASAP7_75t_L g8886 ( 
.A(n_8293),
.Y(n_8886)
);

NOR2xp33_ASAP7_75t_L g8887 ( 
.A(n_8073),
.B(n_5184),
.Y(n_8887)
);

INVx5_ASAP7_75t_L g8888 ( 
.A(n_8403),
.Y(n_8888)
);

INVx1_ASAP7_75t_L g8889 ( 
.A(n_8294),
.Y(n_8889)
);

BUFx2_ASAP7_75t_L g8890 ( 
.A(n_8354),
.Y(n_8890)
);

NAND2xp5_ASAP7_75t_L g8891 ( 
.A(n_8019),
.B(n_5185),
.Y(n_8891)
);

INVx1_ASAP7_75t_L g8892 ( 
.A(n_8278),
.Y(n_8892)
);

AOI22xp33_ASAP7_75t_L g8893 ( 
.A1(n_7895),
.A2(n_5155),
.B1(n_5159),
.B2(n_5153),
.Y(n_8893)
);

HB1xp67_ASAP7_75t_L g8894 ( 
.A(n_8287),
.Y(n_8894)
);

AND3x2_ASAP7_75t_L g8895 ( 
.A(n_8398),
.B(n_5171),
.C(n_5160),
.Y(n_8895)
);

NAND2xp5_ASAP7_75t_L g8896 ( 
.A(n_8123),
.B(n_5189),
.Y(n_8896)
);

INVx2_ASAP7_75t_L g8897 ( 
.A(n_8241),
.Y(n_8897)
);

INVx1_ASAP7_75t_L g8898 ( 
.A(n_8295),
.Y(n_8898)
);

AOI22xp33_ASAP7_75t_L g8899 ( 
.A1(n_8017),
.A2(n_8359),
.B1(n_8358),
.B2(n_8212),
.Y(n_8899)
);

INVx1_ASAP7_75t_L g8900 ( 
.A(n_8297),
.Y(n_8900)
);

INVx1_ASAP7_75t_L g8901 ( 
.A(n_8298),
.Y(n_8901)
);

NAND2xp5_ASAP7_75t_L g8902 ( 
.A(n_8155),
.B(n_5190),
.Y(n_8902)
);

AND2x2_ASAP7_75t_L g8903 ( 
.A(n_8076),
.B(n_8105),
.Y(n_8903)
);

CKINVDCx20_ASAP7_75t_R g8904 ( 
.A(n_8352),
.Y(n_8904)
);

NAND2xp5_ASAP7_75t_L g8905 ( 
.A(n_8217),
.B(n_5191),
.Y(n_8905)
);

INVx1_ASAP7_75t_L g8906 ( 
.A(n_8299),
.Y(n_8906)
);

AND2x2_ASAP7_75t_L g8907 ( 
.A(n_8112),
.B(n_5192),
.Y(n_8907)
);

INVx2_ASAP7_75t_L g8908 ( 
.A(n_8273),
.Y(n_8908)
);

AND2x2_ASAP7_75t_L g8909 ( 
.A(n_8113),
.B(n_5194),
.Y(n_8909)
);

INVx2_ASAP7_75t_SL g8910 ( 
.A(n_7949),
.Y(n_8910)
);

NAND2xp5_ASAP7_75t_L g8911 ( 
.A(n_8247),
.B(n_5196),
.Y(n_8911)
);

BUFx3_ASAP7_75t_L g8912 ( 
.A(n_8383),
.Y(n_8912)
);

AND2x2_ASAP7_75t_L g8913 ( 
.A(n_7972),
.B(n_5197),
.Y(n_8913)
);

INVx1_ASAP7_75t_L g8914 ( 
.A(n_8300),
.Y(n_8914)
);

INVx3_ASAP7_75t_L g8915 ( 
.A(n_8324),
.Y(n_8915)
);

INVx1_ASAP7_75t_L g8916 ( 
.A(n_8303),
.Y(n_8916)
);

INVx6_ASAP7_75t_L g8917 ( 
.A(n_7921),
.Y(n_8917)
);

AOI22xp5_ASAP7_75t_L g8918 ( 
.A1(n_7890),
.A2(n_5199),
.B1(n_5200),
.B2(n_5198),
.Y(n_8918)
);

INVx2_ASAP7_75t_L g8919 ( 
.A(n_8274),
.Y(n_8919)
);

NAND2xp5_ASAP7_75t_SL g8920 ( 
.A(n_8180),
.B(n_5201),
.Y(n_8920)
);

CKINVDCx5p33_ASAP7_75t_R g8921 ( 
.A(n_8405),
.Y(n_8921)
);

INVx4_ASAP7_75t_L g8922 ( 
.A(n_8059),
.Y(n_8922)
);

BUFx3_ASAP7_75t_L g8923 ( 
.A(n_8408),
.Y(n_8923)
);

NOR2xp33_ASAP7_75t_L g8924 ( 
.A(n_7982),
.B(n_5202),
.Y(n_8924)
);

O2A1O1Ixp33_ASAP7_75t_L g8925 ( 
.A1(n_8426),
.A2(n_8014),
.B(n_8012),
.C(n_7929),
.Y(n_8925)
);

AND2x2_ASAP7_75t_L g8926 ( 
.A(n_8521),
.B(n_8257),
.Y(n_8926)
);

INVx1_ASAP7_75t_L g8927 ( 
.A(n_8414),
.Y(n_8927)
);

INVxp67_ASAP7_75t_SL g8928 ( 
.A(n_8423),
.Y(n_8928)
);

NOR2xp33_ASAP7_75t_L g8929 ( 
.A(n_8494),
.B(n_8249),
.Y(n_8929)
);

INVx1_ASAP7_75t_L g8930 ( 
.A(n_8418),
.Y(n_8930)
);

NAND2xp5_ASAP7_75t_L g8931 ( 
.A(n_8851),
.B(n_8128),
.Y(n_8931)
);

INVx2_ASAP7_75t_L g8932 ( 
.A(n_8427),
.Y(n_8932)
);

NAND2xp5_ASAP7_75t_L g8933 ( 
.A(n_8480),
.B(n_8134),
.Y(n_8933)
);

INVx2_ASAP7_75t_SL g8934 ( 
.A(n_8484),
.Y(n_8934)
);

INVx2_ASAP7_75t_L g8935 ( 
.A(n_8430),
.Y(n_8935)
);

OAI22xp5_ASAP7_75t_L g8936 ( 
.A1(n_8533),
.A2(n_7873),
.B1(n_8367),
.B2(n_8269),
.Y(n_8936)
);

NAND2xp5_ASAP7_75t_L g8937 ( 
.A(n_8639),
.B(n_8142),
.Y(n_8937)
);

INVx2_ASAP7_75t_SL g8938 ( 
.A(n_8484),
.Y(n_8938)
);

AOI22xp5_ASAP7_75t_L g8939 ( 
.A1(n_8448),
.A2(n_8161),
.B1(n_8143),
.B2(n_8168),
.Y(n_8939)
);

INVx2_ASAP7_75t_L g8940 ( 
.A(n_8431),
.Y(n_8940)
);

NAND2xp5_ASAP7_75t_SL g8941 ( 
.A(n_8470),
.B(n_8402),
.Y(n_8941)
);

INVx2_ASAP7_75t_SL g8942 ( 
.A(n_8546),
.Y(n_8942)
);

NAND2xp5_ASAP7_75t_L g8943 ( 
.A(n_8415),
.B(n_8286),
.Y(n_8943)
);

NAND2xp5_ASAP7_75t_L g8944 ( 
.A(n_8421),
.B(n_8290),
.Y(n_8944)
);

A2O1A1Ixp33_ASAP7_75t_L g8945 ( 
.A1(n_8449),
.A2(n_8277),
.B(n_8304),
.C(n_8355),
.Y(n_8945)
);

INVxp67_ASAP7_75t_SL g8946 ( 
.A(n_8488),
.Y(n_8946)
);

INVx2_ASAP7_75t_L g8947 ( 
.A(n_8434),
.Y(n_8947)
);

NOR2xp33_ASAP7_75t_L g8948 ( 
.A(n_8651),
.B(n_8169),
.Y(n_8948)
);

OAI22xp33_ASAP7_75t_L g8949 ( 
.A1(n_8453),
.A2(n_8379),
.B1(n_8010),
.B2(n_8338),
.Y(n_8949)
);

NAND2xp5_ASAP7_75t_L g8950 ( 
.A(n_8782),
.B(n_8173),
.Y(n_8950)
);

A2O1A1Ixp33_ASAP7_75t_L g8951 ( 
.A1(n_8517),
.A2(n_8357),
.B(n_8203),
.C(n_8192),
.Y(n_8951)
);

NOR2xp33_ASAP7_75t_L g8952 ( 
.A(n_8482),
.B(n_8344),
.Y(n_8952)
);

NAND2xp5_ASAP7_75t_SL g8953 ( 
.A(n_8604),
.B(n_8334),
.Y(n_8953)
);

AND2x2_ASAP7_75t_L g8954 ( 
.A(n_8438),
.B(n_8515),
.Y(n_8954)
);

NAND2xp5_ASAP7_75t_L g8955 ( 
.A(n_8417),
.B(n_8368),
.Y(n_8955)
);

INVx2_ASAP7_75t_L g8956 ( 
.A(n_8436),
.Y(n_8956)
);

AND2x2_ASAP7_75t_L g8957 ( 
.A(n_8555),
.B(n_8199),
.Y(n_8957)
);

NOR3xp33_ASAP7_75t_L g8958 ( 
.A(n_8527),
.B(n_8407),
.C(n_8387),
.Y(n_8958)
);

INVx2_ASAP7_75t_L g8959 ( 
.A(n_8439),
.Y(n_8959)
);

AOI22xp5_ASAP7_75t_L g8960 ( 
.A1(n_8814),
.A2(n_8535),
.B1(n_8597),
.B2(n_8534),
.Y(n_8960)
);

NAND2xp5_ASAP7_75t_L g8961 ( 
.A(n_8433),
.B(n_7882),
.Y(n_8961)
);

CKINVDCx5p33_ASAP7_75t_R g8962 ( 
.A(n_8640),
.Y(n_8962)
);

NAND2xp5_ASAP7_75t_L g8963 ( 
.A(n_8510),
.B(n_7984),
.Y(n_8963)
);

NAND2xp5_ASAP7_75t_SL g8964 ( 
.A(n_8727),
.B(n_8410),
.Y(n_8964)
);

AOI221xp5_ASAP7_75t_L g8965 ( 
.A1(n_8563),
.A2(n_5187),
.B1(n_5188),
.B2(n_5186),
.C(n_5182),
.Y(n_8965)
);

NOR2xp33_ASAP7_75t_L g8966 ( 
.A(n_8463),
.B(n_8319),
.Y(n_8966)
);

OAI22xp33_ASAP7_75t_L g8967 ( 
.A1(n_8435),
.A2(n_7915),
.B1(n_5203),
.B2(n_5208),
.Y(n_8967)
);

NAND2xp5_ASAP7_75t_L g8968 ( 
.A(n_8560),
.B(n_8032),
.Y(n_8968)
);

INVx1_ASAP7_75t_L g8969 ( 
.A(n_8441),
.Y(n_8969)
);

NAND2xp5_ASAP7_75t_L g8970 ( 
.A(n_8730),
.B(n_8268),
.Y(n_8970)
);

OAI22xp5_ASAP7_75t_L g8971 ( 
.A1(n_8442),
.A2(n_8263),
.B1(n_8308),
.B2(n_8309),
.Y(n_8971)
);

BUFx6f_ASAP7_75t_L g8972 ( 
.A(n_8616),
.Y(n_8972)
);

INVxp67_ASAP7_75t_L g8973 ( 
.A(n_8424),
.Y(n_8973)
);

AOI22xp5_ASAP7_75t_L g8974 ( 
.A1(n_8699),
.A2(n_5204),
.B1(n_5210),
.B2(n_5209),
.Y(n_8974)
);

NOR2xp33_ASAP7_75t_L g8975 ( 
.A(n_8680),
.B(n_5213),
.Y(n_8975)
);

NAND2xp5_ASAP7_75t_L g8976 ( 
.A(n_8617),
.B(n_5193),
.Y(n_8976)
);

NAND2xp5_ASAP7_75t_L g8977 ( 
.A(n_8650),
.B(n_8667),
.Y(n_8977)
);

INVx1_ASAP7_75t_L g8978 ( 
.A(n_8445),
.Y(n_8978)
);

INVx3_ASAP7_75t_L g8979 ( 
.A(n_8505),
.Y(n_8979)
);

INVx1_ASAP7_75t_L g8980 ( 
.A(n_8447),
.Y(n_8980)
);

A2O1A1Ixp33_ASAP7_75t_L g8981 ( 
.A1(n_8924),
.A2(n_5217),
.B(n_5228),
.C(n_5207),
.Y(n_8981)
);

INVx2_ASAP7_75t_L g8982 ( 
.A(n_8455),
.Y(n_8982)
);

NOR2xp33_ASAP7_75t_L g8983 ( 
.A(n_8688),
.B(n_5215),
.Y(n_8983)
);

AOI21xp5_ASAP7_75t_L g8984 ( 
.A1(n_8876),
.A2(n_5233),
.B(n_5230),
.Y(n_8984)
);

OAI221xp5_ASAP7_75t_L g8985 ( 
.A1(n_8847),
.A2(n_5242),
.B1(n_5243),
.B2(n_5239),
.C(n_5236),
.Y(n_8985)
);

NAND2xp5_ASAP7_75t_SL g8986 ( 
.A(n_8888),
.B(n_5216),
.Y(n_8986)
);

NAND2xp5_ASAP7_75t_L g8987 ( 
.A(n_8744),
.B(n_5249),
.Y(n_8987)
);

INVx1_ASAP7_75t_L g8988 ( 
.A(n_8460),
.Y(n_8988)
);

NAND2xp5_ASAP7_75t_L g8989 ( 
.A(n_8751),
.B(n_5250),
.Y(n_8989)
);

CKINVDCx5p33_ASAP7_75t_R g8990 ( 
.A(n_8457),
.Y(n_8990)
);

INVxp67_ASAP7_75t_L g8991 ( 
.A(n_8691),
.Y(n_8991)
);

INVx2_ASAP7_75t_L g8992 ( 
.A(n_8467),
.Y(n_8992)
);

AOI21xp5_ASAP7_75t_L g8993 ( 
.A1(n_8629),
.A2(n_5253),
.B(n_5251),
.Y(n_8993)
);

INVx2_ASAP7_75t_L g8994 ( 
.A(n_8469),
.Y(n_8994)
);

NAND2xp5_ASAP7_75t_L g8995 ( 
.A(n_8693),
.B(n_5261),
.Y(n_8995)
);

NAND2xp5_ASAP7_75t_L g8996 ( 
.A(n_8772),
.B(n_5262),
.Y(n_8996)
);

INVx1_ASAP7_75t_L g8997 ( 
.A(n_8471),
.Y(n_8997)
);

INVx4_ASAP7_75t_L g8998 ( 
.A(n_8546),
.Y(n_8998)
);

AOI22xp5_ASAP7_75t_L g8999 ( 
.A1(n_8428),
.A2(n_5221),
.B1(n_5222),
.B2(n_5219),
.Y(n_8999)
);

AOI22xp5_ASAP7_75t_L g9000 ( 
.A1(n_8921),
.A2(n_5224),
.B1(n_5226),
.B2(n_5223),
.Y(n_9000)
);

NAND2xp5_ASAP7_75t_L g9001 ( 
.A(n_8537),
.B(n_5263),
.Y(n_9001)
);

OR2x2_ASAP7_75t_L g9002 ( 
.A(n_8544),
.B(n_5227),
.Y(n_9002)
);

NOR2xp33_ASAP7_75t_L g9003 ( 
.A(n_8740),
.B(n_5229),
.Y(n_9003)
);

INVx2_ASAP7_75t_L g9004 ( 
.A(n_8472),
.Y(n_9004)
);

NAND2xp5_ASAP7_75t_L g9005 ( 
.A(n_8557),
.B(n_5264),
.Y(n_9005)
);

NOR2xp33_ASAP7_75t_SL g9006 ( 
.A(n_8474),
.B(n_5231),
.Y(n_9006)
);

NAND2xp5_ASAP7_75t_L g9007 ( 
.A(n_8663),
.B(n_5267),
.Y(n_9007)
);

NAND2xp5_ASAP7_75t_L g9008 ( 
.A(n_8668),
.B(n_5270),
.Y(n_9008)
);

NAND2xp5_ASAP7_75t_SL g9009 ( 
.A(n_8888),
.B(n_8833),
.Y(n_9009)
);

NAND2xp5_ASAP7_75t_L g9010 ( 
.A(n_8622),
.B(n_5279),
.Y(n_9010)
);

INVx1_ASAP7_75t_L g9011 ( 
.A(n_8481),
.Y(n_9011)
);

NAND2xp5_ASAP7_75t_L g9012 ( 
.A(n_8700),
.B(n_8721),
.Y(n_9012)
);

NAND2xp5_ASAP7_75t_L g9013 ( 
.A(n_8461),
.B(n_5281),
.Y(n_9013)
);

INVx2_ASAP7_75t_L g9014 ( 
.A(n_8490),
.Y(n_9014)
);

INVx2_ASAP7_75t_L g9015 ( 
.A(n_8491),
.Y(n_9015)
);

NAND2xp5_ASAP7_75t_L g9016 ( 
.A(n_8679),
.B(n_5288),
.Y(n_9016)
);

INVx2_ASAP7_75t_L g9017 ( 
.A(n_8495),
.Y(n_9017)
);

NOR2xp33_ASAP7_75t_L g9018 ( 
.A(n_8429),
.B(n_5232),
.Y(n_9018)
);

CKINVDCx5p33_ASAP7_75t_R g9019 ( 
.A(n_8497),
.Y(n_9019)
);

INVx1_ASAP7_75t_L g9020 ( 
.A(n_8502),
.Y(n_9020)
);

OR2x6_ASAP7_75t_L g9021 ( 
.A(n_8504),
.B(n_5290),
.Y(n_9021)
);

INVx8_ASAP7_75t_L g9022 ( 
.A(n_8580),
.Y(n_9022)
);

NAND2xp5_ASAP7_75t_SL g9023 ( 
.A(n_8776),
.B(n_5234),
.Y(n_9023)
);

AND2x4_ASAP7_75t_L g9024 ( 
.A(n_8759),
.B(n_5297),
.Y(n_9024)
);

NOR2xp33_ASAP7_75t_L g9025 ( 
.A(n_8774),
.B(n_5237),
.Y(n_9025)
);

NOR2xp33_ASAP7_75t_L g9026 ( 
.A(n_8775),
.B(n_5238),
.Y(n_9026)
);

NAND2xp5_ASAP7_75t_L g9027 ( 
.A(n_8512),
.B(n_5302),
.Y(n_9027)
);

OAI22xp5_ASAP7_75t_L g9028 ( 
.A1(n_8503),
.A2(n_8513),
.B1(n_8516),
.B2(n_8506),
.Y(n_9028)
);

NAND2xp5_ASAP7_75t_SL g9029 ( 
.A(n_8829),
.B(n_8858),
.Y(n_9029)
);

INVx2_ASAP7_75t_L g9030 ( 
.A(n_8523),
.Y(n_9030)
);

NAND2xp5_ASAP7_75t_SL g9031 ( 
.A(n_8718),
.B(n_5241),
.Y(n_9031)
);

NAND2xp5_ASAP7_75t_L g9032 ( 
.A(n_8475),
.B(n_5303),
.Y(n_9032)
);

BUFx6f_ASAP7_75t_SL g9033 ( 
.A(n_8422),
.Y(n_9033)
);

NAND2xp5_ASAP7_75t_L g9034 ( 
.A(n_8528),
.B(n_5307),
.Y(n_9034)
);

NAND2xp5_ASAP7_75t_L g9035 ( 
.A(n_8809),
.B(n_5312),
.Y(n_9035)
);

NAND2xp5_ASAP7_75t_SL g9036 ( 
.A(n_8718),
.B(n_5246),
.Y(n_9036)
);

NOR2xp33_ASAP7_75t_L g9037 ( 
.A(n_8532),
.B(n_5247),
.Y(n_9037)
);

NOR2xp33_ASAP7_75t_L g9038 ( 
.A(n_8883),
.B(n_5248),
.Y(n_9038)
);

INVx1_ASAP7_75t_L g9039 ( 
.A(n_8831),
.Y(n_9039)
);

INVx1_ASAP7_75t_L g9040 ( 
.A(n_8835),
.Y(n_9040)
);

INVx2_ASAP7_75t_L g9041 ( 
.A(n_8844),
.Y(n_9041)
);

INVx3_ASAP7_75t_L g9042 ( 
.A(n_8616),
.Y(n_9042)
);

AOI22xp5_ASAP7_75t_L g9043 ( 
.A1(n_8581),
.A2(n_5256),
.B1(n_5258),
.B2(n_5252),
.Y(n_9043)
);

OAI22xp5_ASAP7_75t_SL g9044 ( 
.A1(n_8868),
.A2(n_5260),
.B1(n_5268),
.B2(n_5259),
.Y(n_9044)
);

NAND2xp5_ASAP7_75t_L g9045 ( 
.A(n_8539),
.B(n_5313),
.Y(n_9045)
);

NAND2xp5_ASAP7_75t_L g9046 ( 
.A(n_8542),
.B(n_8550),
.Y(n_9046)
);

NAND3xp33_ASAP7_75t_L g9047 ( 
.A(n_8887),
.B(n_5271),
.C(n_5269),
.Y(n_9047)
);

BUFx6f_ASAP7_75t_L g9048 ( 
.A(n_8602),
.Y(n_9048)
);

OR2x6_ASAP7_75t_L g9049 ( 
.A(n_8602),
.B(n_5316),
.Y(n_9049)
);

INVxp67_ASAP7_75t_L g9050 ( 
.A(n_8507),
.Y(n_9050)
);

AND2x2_ASAP7_75t_L g9051 ( 
.A(n_8559),
.B(n_8572),
.Y(n_9051)
);

INVx2_ASAP7_75t_L g9052 ( 
.A(n_8600),
.Y(n_9052)
);

OAI22xp33_ASAP7_75t_SL g9053 ( 
.A1(n_8920),
.A2(n_5275),
.B1(n_5276),
.B2(n_5274),
.Y(n_9053)
);

INVx2_ASAP7_75t_L g9054 ( 
.A(n_8603),
.Y(n_9054)
);

NOR2xp67_ASAP7_75t_L g9055 ( 
.A(n_8556),
.B(n_4283),
.Y(n_9055)
);

INVx2_ASAP7_75t_SL g9056 ( 
.A(n_8580),
.Y(n_9056)
);

AOI22xp33_ASAP7_75t_L g9057 ( 
.A1(n_8462),
.A2(n_5322),
.B1(n_5330),
.B2(n_5319),
.Y(n_9057)
);

AND2x2_ASAP7_75t_L g9058 ( 
.A(n_8593),
.B(n_5277),
.Y(n_9058)
);

NOR2xp33_ASAP7_75t_L g9059 ( 
.A(n_8902),
.B(n_5278),
.Y(n_9059)
);

NAND2xp33_ASAP7_75t_L g9060 ( 
.A(n_8826),
.B(n_5280),
.Y(n_9060)
);

INVx1_ASAP7_75t_L g9061 ( 
.A(n_8606),
.Y(n_9061)
);

NAND2xp5_ASAP7_75t_L g9062 ( 
.A(n_8553),
.B(n_5335),
.Y(n_9062)
);

NAND2xp5_ASAP7_75t_SL g9063 ( 
.A(n_8769),
.B(n_5282),
.Y(n_9063)
);

NAND2xp5_ASAP7_75t_L g9064 ( 
.A(n_8564),
.B(n_5336),
.Y(n_9064)
);

AND2x6_ASAP7_75t_SL g9065 ( 
.A(n_8416),
.B(n_5339),
.Y(n_9065)
);

NAND2xp5_ASAP7_75t_SL g9066 ( 
.A(n_8845),
.B(n_8524),
.Y(n_9066)
);

NOR2xp33_ASAP7_75t_L g9067 ( 
.A(n_8768),
.B(n_5283),
.Y(n_9067)
);

NAND2xp5_ASAP7_75t_L g9068 ( 
.A(n_8565),
.B(n_5344),
.Y(n_9068)
);

NAND2xp5_ASAP7_75t_L g9069 ( 
.A(n_8570),
.B(n_5345),
.Y(n_9069)
);

INVx2_ASAP7_75t_L g9070 ( 
.A(n_8607),
.Y(n_9070)
);

NAND2xp5_ASAP7_75t_SL g9071 ( 
.A(n_8845),
.B(n_5284),
.Y(n_9071)
);

NOR2xp33_ASAP7_75t_L g9072 ( 
.A(n_8496),
.B(n_5286),
.Y(n_9072)
);

INVx2_ASAP7_75t_L g9073 ( 
.A(n_8609),
.Y(n_9073)
);

NAND2xp5_ASAP7_75t_SL g9074 ( 
.A(n_8518),
.B(n_5287),
.Y(n_9074)
);

O2A1O1Ixp33_ASAP7_75t_L g9075 ( 
.A1(n_8437),
.A2(n_5347),
.B(n_5353),
.C(n_5346),
.Y(n_9075)
);

INVx2_ASAP7_75t_L g9076 ( 
.A(n_8612),
.Y(n_9076)
);

NAND2xp5_ASAP7_75t_L g9077 ( 
.A(n_8575),
.B(n_5354),
.Y(n_9077)
);

NOR2xp33_ASAP7_75t_L g9078 ( 
.A(n_8584),
.B(n_5292),
.Y(n_9078)
);

NAND2xp5_ASAP7_75t_L g9079 ( 
.A(n_8577),
.B(n_5360),
.Y(n_9079)
);

INVx1_ASAP7_75t_L g9080 ( 
.A(n_8614),
.Y(n_9080)
);

INVx1_ASAP7_75t_L g9081 ( 
.A(n_8621),
.Y(n_9081)
);

NAND2xp5_ASAP7_75t_SL g9082 ( 
.A(n_8530),
.B(n_5294),
.Y(n_9082)
);

AOI22xp33_ASAP7_75t_L g9083 ( 
.A1(n_8529),
.A2(n_5371),
.B1(n_5373),
.B2(n_5364),
.Y(n_9083)
);

INVx2_ASAP7_75t_L g9084 ( 
.A(n_8624),
.Y(n_9084)
);

BUFx6f_ASAP7_75t_SL g9085 ( 
.A(n_8425),
.Y(n_9085)
);

NAND2xp5_ASAP7_75t_SL g9086 ( 
.A(n_8573),
.B(n_5295),
.Y(n_9086)
);

INVx2_ASAP7_75t_L g9087 ( 
.A(n_8626),
.Y(n_9087)
);

INVx1_ASAP7_75t_L g9088 ( 
.A(n_8631),
.Y(n_9088)
);

BUFx8_ASAP7_75t_L g9089 ( 
.A(n_8810),
.Y(n_9089)
);

INVx2_ASAP7_75t_L g9090 ( 
.A(n_8636),
.Y(n_9090)
);

INVx2_ASAP7_75t_L g9091 ( 
.A(n_8641),
.Y(n_9091)
);

NAND2xp5_ASAP7_75t_SL g9092 ( 
.A(n_8923),
.B(n_5296),
.Y(n_9092)
);

NAND2xp5_ASAP7_75t_L g9093 ( 
.A(n_8578),
.B(n_5374),
.Y(n_9093)
);

OR2x2_ASAP7_75t_L g9094 ( 
.A(n_8541),
.B(n_5298),
.Y(n_9094)
);

NAND3xp33_ASAP7_75t_L g9095 ( 
.A(n_8746),
.B(n_5301),
.C(n_5299),
.Y(n_9095)
);

INVx2_ASAP7_75t_L g9096 ( 
.A(n_8642),
.Y(n_9096)
);

AND2x4_ASAP7_75t_L g9097 ( 
.A(n_8468),
.B(n_5377),
.Y(n_9097)
);

NAND2xp5_ASAP7_75t_L g9098 ( 
.A(n_8590),
.B(n_5381),
.Y(n_9098)
);

NAND2x1_ASAP7_75t_L g9099 ( 
.A(n_8623),
.B(n_5382),
.Y(n_9099)
);

BUFx6f_ASAP7_75t_SL g9100 ( 
.A(n_8613),
.Y(n_9100)
);

NAND2xp5_ASAP7_75t_SL g9101 ( 
.A(n_8662),
.B(n_5304),
.Y(n_9101)
);

INVx1_ASAP7_75t_L g9102 ( 
.A(n_8644),
.Y(n_9102)
);

INVx2_ASAP7_75t_L g9103 ( 
.A(n_8653),
.Y(n_9103)
);

BUFx3_ASAP7_75t_L g9104 ( 
.A(n_8501),
.Y(n_9104)
);

INVx2_ASAP7_75t_L g9105 ( 
.A(n_8658),
.Y(n_9105)
);

INVx1_ASAP7_75t_L g9106 ( 
.A(n_8673),
.Y(n_9106)
);

NAND2xp5_ASAP7_75t_SL g9107 ( 
.A(n_8662),
.B(n_5308),
.Y(n_9107)
);

AND2x4_ASAP7_75t_L g9108 ( 
.A(n_8526),
.B(n_5384),
.Y(n_9108)
);

NAND2xp5_ASAP7_75t_SL g9109 ( 
.A(n_8567),
.B(n_5310),
.Y(n_9109)
);

NAND2xp5_ASAP7_75t_L g9110 ( 
.A(n_8591),
.B(n_5387),
.Y(n_9110)
);

NAND2xp5_ASAP7_75t_L g9111 ( 
.A(n_8675),
.B(n_8677),
.Y(n_9111)
);

NAND2xp5_ASAP7_75t_L g9112 ( 
.A(n_8678),
.B(n_5388),
.Y(n_9112)
);

NAND2xp5_ASAP7_75t_L g9113 ( 
.A(n_8683),
.B(n_5404),
.Y(n_9113)
);

NAND2xp5_ASAP7_75t_SL g9114 ( 
.A(n_8625),
.B(n_5314),
.Y(n_9114)
);

INVx1_ASAP7_75t_L g9115 ( 
.A(n_8689),
.Y(n_9115)
);

NOR2xp33_ASAP7_75t_L g9116 ( 
.A(n_8465),
.B(n_5317),
.Y(n_9116)
);

INVx2_ASAP7_75t_L g9117 ( 
.A(n_8696),
.Y(n_9117)
);

NAND2xp5_ASAP7_75t_L g9118 ( 
.A(n_8698),
.B(n_5410),
.Y(n_9118)
);

INVx3_ASAP7_75t_L g9119 ( 
.A(n_8605),
.Y(n_9119)
);

NAND2xp5_ASAP7_75t_L g9120 ( 
.A(n_8702),
.B(n_5416),
.Y(n_9120)
);

AND2x4_ASAP7_75t_L g9121 ( 
.A(n_8543),
.B(n_5417),
.Y(n_9121)
);

NAND2xp5_ASAP7_75t_SL g9122 ( 
.A(n_8659),
.B(n_5320),
.Y(n_9122)
);

INVx2_ASAP7_75t_L g9123 ( 
.A(n_8708),
.Y(n_9123)
);

A2O1A1Ixp33_ASAP7_75t_L g9124 ( 
.A1(n_8619),
.A2(n_5430),
.B(n_5433),
.C(n_5419),
.Y(n_9124)
);

BUFx6f_ASAP7_75t_L g9125 ( 
.A(n_8450),
.Y(n_9125)
);

NAND2xp5_ASAP7_75t_SL g9126 ( 
.A(n_8670),
.B(n_5325),
.Y(n_9126)
);

INVx2_ASAP7_75t_L g9127 ( 
.A(n_8710),
.Y(n_9127)
);

AND2x2_ASAP7_75t_L g9128 ( 
.A(n_8464),
.B(n_5326),
.Y(n_9128)
);

NAND2xp5_ASAP7_75t_L g9129 ( 
.A(n_8419),
.B(n_5434),
.Y(n_9129)
);

INVx2_ASAP7_75t_L g9130 ( 
.A(n_8897),
.Y(n_9130)
);

AND2x2_ASAP7_75t_L g9131 ( 
.A(n_8643),
.B(n_5327),
.Y(n_9131)
);

NOR2xp33_ASAP7_75t_L g9132 ( 
.A(n_8443),
.B(n_5328),
.Y(n_9132)
);

INVx1_ASAP7_75t_L g9133 ( 
.A(n_8627),
.Y(n_9133)
);

INVx1_ASAP7_75t_L g9134 ( 
.A(n_8892),
.Y(n_9134)
);

INVx1_ASAP7_75t_L g9135 ( 
.A(n_8898),
.Y(n_9135)
);

NAND2xp5_ASAP7_75t_SL g9136 ( 
.A(n_8912),
.B(n_5331),
.Y(n_9136)
);

INVx1_ASAP7_75t_L g9137 ( 
.A(n_8900),
.Y(n_9137)
);

INVx1_ASAP7_75t_L g9138 ( 
.A(n_8901),
.Y(n_9138)
);

AND2x2_ASAP7_75t_L g9139 ( 
.A(n_8825),
.B(n_5332),
.Y(n_9139)
);

INVx1_ASAP7_75t_L g9140 ( 
.A(n_8906),
.Y(n_9140)
);

INVx2_ASAP7_75t_L g9141 ( 
.A(n_8908),
.Y(n_9141)
);

NAND2xp5_ASAP7_75t_L g9142 ( 
.A(n_8420),
.B(n_8446),
.Y(n_9142)
);

AOI22xp33_ASAP7_75t_L g9143 ( 
.A1(n_8794),
.A2(n_5441),
.B1(n_5449),
.B2(n_5437),
.Y(n_9143)
);

NAND2xp33_ASAP7_75t_L g9144 ( 
.A(n_8826),
.B(n_5333),
.Y(n_9144)
);

AOI22xp5_ASAP7_75t_L g9145 ( 
.A1(n_8903),
.A2(n_5340),
.B1(n_5343),
.B2(n_5334),
.Y(n_9145)
);

AOI22xp33_ASAP7_75t_L g9146 ( 
.A1(n_8738),
.A2(n_5452),
.B1(n_5455),
.B2(n_5451),
.Y(n_9146)
);

AOI22xp5_ASAP7_75t_L g9147 ( 
.A1(n_8500),
.A2(n_5350),
.B1(n_5351),
.B2(n_5349),
.Y(n_9147)
);

NAND2xp5_ASAP7_75t_SL g9148 ( 
.A(n_8846),
.B(n_5352),
.Y(n_9148)
);

NAND2xp5_ASAP7_75t_SL g9149 ( 
.A(n_8860),
.B(n_5356),
.Y(n_9149)
);

NAND2xp5_ASAP7_75t_L g9150 ( 
.A(n_8452),
.B(n_5457),
.Y(n_9150)
);

INVx2_ASAP7_75t_L g9151 ( 
.A(n_8919),
.Y(n_9151)
);

CKINVDCx5p33_ASAP7_75t_R g9152 ( 
.A(n_8717),
.Y(n_9152)
);

INVx4_ASAP7_75t_L g9153 ( 
.A(n_8450),
.Y(n_9153)
);

NAND2xp5_ASAP7_75t_L g9154 ( 
.A(n_8473),
.B(n_5461),
.Y(n_9154)
);

NAND2xp5_ASAP7_75t_SL g9155 ( 
.A(n_8587),
.B(n_5357),
.Y(n_9155)
);

NOR2x1p5_ASAP7_75t_L g9156 ( 
.A(n_8758),
.B(n_5358),
.Y(n_9156)
);

CKINVDCx5p33_ASAP7_75t_R g9157 ( 
.A(n_8669),
.Y(n_9157)
);

NAND3xp33_ASAP7_75t_L g9158 ( 
.A(n_8558),
.B(n_5361),
.C(n_5359),
.Y(n_9158)
);

AO22x2_ASAP7_75t_L g9159 ( 
.A1(n_8914),
.A2(n_5475),
.B1(n_5478),
.B2(n_5462),
.Y(n_9159)
);

NAND2xp5_ASAP7_75t_L g9160 ( 
.A(n_8477),
.B(n_5482),
.Y(n_9160)
);

INVx2_ASAP7_75t_L g9161 ( 
.A(n_8479),
.Y(n_9161)
);

INVx1_ASAP7_75t_L g9162 ( 
.A(n_8916),
.Y(n_9162)
);

NAND2xp5_ASAP7_75t_SL g9163 ( 
.A(n_8880),
.B(n_5363),
.Y(n_9163)
);

NAND3xp33_ASAP7_75t_L g9164 ( 
.A(n_8802),
.B(n_5366),
.C(n_5365),
.Y(n_9164)
);

INVx5_ASAP7_75t_L g9165 ( 
.A(n_8451),
.Y(n_9165)
);

NOR2xp33_ASAP7_75t_L g9166 ( 
.A(n_8579),
.B(n_5368),
.Y(n_9166)
);

NAND2xp5_ASAP7_75t_L g9167 ( 
.A(n_8487),
.B(n_5486),
.Y(n_9167)
);

NAND2xp5_ASAP7_75t_L g9168 ( 
.A(n_8489),
.B(n_5487),
.Y(n_9168)
);

NAND2xp5_ASAP7_75t_SL g9169 ( 
.A(n_8822),
.B(n_5369),
.Y(n_9169)
);

NAND2xp5_ASAP7_75t_L g9170 ( 
.A(n_8511),
.B(n_5493),
.Y(n_9170)
);

O2A1O1Ixp5_ASAP7_75t_L g9171 ( 
.A1(n_8816),
.A2(n_8850),
.B(n_8796),
.C(n_8684),
.Y(n_9171)
);

O2A1O1Ixp33_ASAP7_75t_L g9172 ( 
.A1(n_8549),
.A2(n_5500),
.B(n_5502),
.C(n_5498),
.Y(n_9172)
);

NAND2xp5_ASAP7_75t_L g9173 ( 
.A(n_8514),
.B(n_5505),
.Y(n_9173)
);

INVx1_ASAP7_75t_L g9174 ( 
.A(n_8632),
.Y(n_9174)
);

NAND2xp5_ASAP7_75t_L g9175 ( 
.A(n_8536),
.B(n_8540),
.Y(n_9175)
);

NOR2xp67_ASAP7_75t_L g9176 ( 
.A(n_8656),
.B(n_4286),
.Y(n_9176)
);

NAND2xp5_ASAP7_75t_L g9177 ( 
.A(n_8548),
.B(n_5506),
.Y(n_9177)
);

INVx2_ASAP7_75t_L g9178 ( 
.A(n_8562),
.Y(n_9178)
);

NAND2xp5_ASAP7_75t_L g9179 ( 
.A(n_8595),
.B(n_5507),
.Y(n_9179)
);

INVx2_ASAP7_75t_L g9180 ( 
.A(n_8596),
.Y(n_9180)
);

BUFx3_ASAP7_75t_L g9181 ( 
.A(n_8566),
.Y(n_9181)
);

CKINVDCx11_ASAP7_75t_R g9182 ( 
.A(n_8444),
.Y(n_9182)
);

NAND2xp5_ASAP7_75t_L g9183 ( 
.A(n_8712),
.B(n_5515),
.Y(n_9183)
);

INVxp67_ASAP7_75t_L g9184 ( 
.A(n_8628),
.Y(n_9184)
);

INVx5_ASAP7_75t_L g9185 ( 
.A(n_8451),
.Y(n_9185)
);

NAND2xp5_ASAP7_75t_L g9186 ( 
.A(n_8713),
.B(n_5520),
.Y(n_9186)
);

AO221x1_ASAP7_75t_L g9187 ( 
.A1(n_8837),
.A2(n_5535),
.B1(n_5544),
.B2(n_5524),
.C(n_5522),
.Y(n_9187)
);

INVx2_ASAP7_75t_L g9188 ( 
.A(n_8633),
.Y(n_9188)
);

NAND2xp5_ASAP7_75t_L g9189 ( 
.A(n_8715),
.B(n_5552),
.Y(n_9189)
);

NAND2xp5_ASAP7_75t_SL g9190 ( 
.A(n_8788),
.B(n_8648),
.Y(n_9190)
);

INVx1_ASAP7_75t_L g9191 ( 
.A(n_8719),
.Y(n_9191)
);

INVx2_ASAP7_75t_L g9192 ( 
.A(n_8652),
.Y(n_9192)
);

NAND2xp5_ASAP7_75t_L g9193 ( 
.A(n_8723),
.B(n_8726),
.Y(n_9193)
);

INVx1_ASAP7_75t_L g9194 ( 
.A(n_8733),
.Y(n_9194)
);

NOR2xp33_ASAP7_75t_L g9195 ( 
.A(n_8664),
.B(n_5370),
.Y(n_9195)
);

NAND2xp5_ASAP7_75t_L g9196 ( 
.A(n_8686),
.B(n_5555),
.Y(n_9196)
);

INVx2_ASAP7_75t_L g9197 ( 
.A(n_8654),
.Y(n_9197)
);

NAND2xp5_ASAP7_75t_L g9198 ( 
.A(n_8803),
.B(n_5563),
.Y(n_9198)
);

NAND2xp5_ASAP7_75t_L g9199 ( 
.A(n_8808),
.B(n_5568),
.Y(n_9199)
);

INVx1_ASAP7_75t_L g9200 ( 
.A(n_8864),
.Y(n_9200)
);

NAND3xp33_ASAP7_75t_L g9201 ( 
.A(n_8716),
.B(n_5376),
.C(n_5375),
.Y(n_9201)
);

NAND2xp5_ASAP7_75t_L g9202 ( 
.A(n_8870),
.B(n_5570),
.Y(n_9202)
);

NOR2xp33_ASAP7_75t_L g9203 ( 
.A(n_8722),
.B(n_5379),
.Y(n_9203)
);

NAND2xp5_ASAP7_75t_SL g9204 ( 
.A(n_8706),
.B(n_5380),
.Y(n_9204)
);

NAND2xp5_ASAP7_75t_L g9205 ( 
.A(n_8586),
.B(n_5572),
.Y(n_9205)
);

NAND2xp5_ASAP7_75t_L g9206 ( 
.A(n_8589),
.B(n_5591),
.Y(n_9206)
);

NAND2xp5_ASAP7_75t_L g9207 ( 
.A(n_8841),
.B(n_5594),
.Y(n_9207)
);

INVx2_ASAP7_75t_SL g9208 ( 
.A(n_8454),
.Y(n_9208)
);

AND2x2_ASAP7_75t_L g9209 ( 
.A(n_8645),
.B(n_5383),
.Y(n_9209)
);

AND2x4_ASAP7_75t_L g9210 ( 
.A(n_8440),
.B(n_5595),
.Y(n_9210)
);

INVx3_ASAP7_75t_L g9211 ( 
.A(n_8493),
.Y(n_9211)
);

NAND3xp33_ASAP7_75t_L g9212 ( 
.A(n_8522),
.B(n_5391),
.C(n_5385),
.Y(n_9212)
);

INVx1_ASAP7_75t_SL g9213 ( 
.A(n_8498),
.Y(n_9213)
);

INVx2_ASAP7_75t_L g9214 ( 
.A(n_8660),
.Y(n_9214)
);

OR2x2_ASAP7_75t_SL g9215 ( 
.A(n_8705),
.B(n_5596),
.Y(n_9215)
);

NAND2xp5_ASAP7_75t_L g9216 ( 
.A(n_8853),
.B(n_5598),
.Y(n_9216)
);

NAND2xp5_ASAP7_75t_L g9217 ( 
.A(n_8907),
.B(n_5601),
.Y(n_9217)
);

NAND2xp5_ASAP7_75t_L g9218 ( 
.A(n_8909),
.B(n_5614),
.Y(n_9218)
);

NAND2xp5_ASAP7_75t_L g9219 ( 
.A(n_8913),
.B(n_5619),
.Y(n_9219)
);

NOR3xp33_ASAP7_75t_L g9220 ( 
.A(n_8610),
.B(n_5625),
.C(n_5620),
.Y(n_9220)
);

OAI22xp33_ASAP7_75t_L g9221 ( 
.A1(n_8884),
.A2(n_5393),
.B1(n_5395),
.B2(n_5392),
.Y(n_9221)
);

NOR2xp33_ASAP7_75t_L g9222 ( 
.A(n_8728),
.B(n_5396),
.Y(n_9222)
);

NAND2xp5_ASAP7_75t_L g9223 ( 
.A(n_8735),
.B(n_5628),
.Y(n_9223)
);

INVx2_ASAP7_75t_L g9224 ( 
.A(n_8665),
.Y(n_9224)
);

NAND2xp5_ASAP7_75t_L g9225 ( 
.A(n_8736),
.B(n_5633),
.Y(n_9225)
);

INVxp33_ASAP7_75t_L g9226 ( 
.A(n_8720),
.Y(n_9226)
);

NAND2xp5_ASAP7_75t_SL g9227 ( 
.A(n_8731),
.B(n_5398),
.Y(n_9227)
);

INVx1_ASAP7_75t_L g9228 ( 
.A(n_8874),
.Y(n_9228)
);

INVx1_ASAP7_75t_L g9229 ( 
.A(n_8742),
.Y(n_9229)
);

AOI21xp5_ASAP7_75t_L g9230 ( 
.A1(n_8899),
.A2(n_5640),
.B(n_5635),
.Y(n_9230)
);

OAI22xp5_ASAP7_75t_L g9231 ( 
.A1(n_8869),
.A2(n_5400),
.B1(n_5401),
.B2(n_5399),
.Y(n_9231)
);

INVx1_ASAP7_75t_L g9232 ( 
.A(n_8747),
.Y(n_9232)
);

INVx2_ASAP7_75t_L g9233 ( 
.A(n_8671),
.Y(n_9233)
);

NOR2xp33_ASAP7_75t_SL g9234 ( 
.A(n_8756),
.B(n_5403),
.Y(n_9234)
);

NAND2xp5_ASAP7_75t_L g9235 ( 
.A(n_8748),
.B(n_5646),
.Y(n_9235)
);

NAND2xp5_ASAP7_75t_L g9236 ( 
.A(n_8749),
.B(n_5654),
.Y(n_9236)
);

OR2x2_ASAP7_75t_L g9237 ( 
.A(n_8459),
.B(n_5408),
.Y(n_9237)
);

AND2x2_ASAP7_75t_L g9238 ( 
.A(n_8821),
.B(n_5409),
.Y(n_9238)
);

INVx1_ASAP7_75t_SL g9239 ( 
.A(n_8583),
.Y(n_9239)
);

INVx4_ASAP7_75t_L g9240 ( 
.A(n_8454),
.Y(n_9240)
);

INVx1_ASAP7_75t_L g9241 ( 
.A(n_8761),
.Y(n_9241)
);

INVx8_ASAP7_75t_L g9242 ( 
.A(n_8458),
.Y(n_9242)
);

A2O1A1Ixp33_ASAP7_75t_L g9243 ( 
.A1(n_8709),
.A2(n_5660),
.B(n_5668),
.C(n_5656),
.Y(n_9243)
);

INVx1_ASAP7_75t_L g9244 ( 
.A(n_8763),
.Y(n_9244)
);

NOR2xp33_ASAP7_75t_L g9245 ( 
.A(n_8647),
.B(n_5413),
.Y(n_9245)
);

NAND2xp5_ASAP7_75t_SL g9246 ( 
.A(n_8786),
.B(n_5415),
.Y(n_9246)
);

INVx4_ASAP7_75t_L g9247 ( 
.A(n_8458),
.Y(n_9247)
);

NAND2xp5_ASAP7_75t_SL g9248 ( 
.A(n_8877),
.B(n_5420),
.Y(n_9248)
);

AND2x2_ASAP7_75t_L g9249 ( 
.A(n_8804),
.B(n_5421),
.Y(n_9249)
);

NAND2xp5_ASAP7_75t_L g9250 ( 
.A(n_8767),
.B(n_5670),
.Y(n_9250)
);

AND2x2_ASAP7_75t_L g9251 ( 
.A(n_8838),
.B(n_5423),
.Y(n_9251)
);

INVx2_ASAP7_75t_L g9252 ( 
.A(n_8672),
.Y(n_9252)
);

NAND2xp5_ASAP7_75t_L g9253 ( 
.A(n_8780),
.B(n_5672),
.Y(n_9253)
);

NAND3xp33_ASAP7_75t_L g9254 ( 
.A(n_8618),
.B(n_5425),
.C(n_5424),
.Y(n_9254)
);

NAND2xp5_ASAP7_75t_L g9255 ( 
.A(n_8790),
.B(n_5674),
.Y(n_9255)
);

NAND2xp5_ASAP7_75t_SL g9256 ( 
.A(n_8820),
.B(n_5426),
.Y(n_9256)
);

OR2x2_ASAP7_75t_L g9257 ( 
.A(n_8834),
.B(n_5427),
.Y(n_9257)
);

NAND2xp5_ASAP7_75t_L g9258 ( 
.A(n_8792),
.B(n_5675),
.Y(n_9258)
);

NAND2xp5_ASAP7_75t_SL g9259 ( 
.A(n_8820),
.B(n_8827),
.Y(n_9259)
);

AOI22xp33_ASAP7_75t_L g9260 ( 
.A1(n_8638),
.A2(n_5679),
.B1(n_5681),
.B2(n_5677),
.Y(n_9260)
);

NAND2xp5_ASAP7_75t_L g9261 ( 
.A(n_8799),
.B(n_5428),
.Y(n_9261)
);

BUFx2_ASAP7_75t_L g9262 ( 
.A(n_8598),
.Y(n_9262)
);

NAND2xp5_ASAP7_75t_SL g9263 ( 
.A(n_8827),
.B(n_5429),
.Y(n_9263)
);

BUFx6f_ASAP7_75t_L g9264 ( 
.A(n_8476),
.Y(n_9264)
);

AND2x2_ASAP7_75t_L g9265 ( 
.A(n_8856),
.B(n_5431),
.Y(n_9265)
);

CKINVDCx5p33_ASAP7_75t_R g9266 ( 
.A(n_8791),
.Y(n_9266)
);

INVx1_ASAP7_75t_L g9267 ( 
.A(n_8805),
.Y(n_9267)
);

NOR2xp33_ASAP7_75t_L g9268 ( 
.A(n_8800),
.B(n_5432),
.Y(n_9268)
);

BUFx6f_ASAP7_75t_SL g9269 ( 
.A(n_8432),
.Y(n_9269)
);

O2A1O1Ixp5_ASAP7_75t_L g9270 ( 
.A1(n_8752),
.A2(n_9),
.B(n_7),
.C(n_8),
.Y(n_9270)
);

NAND2xp5_ASAP7_75t_L g9271 ( 
.A(n_8806),
.B(n_5439),
.Y(n_9271)
);

NAND2xp5_ASAP7_75t_L g9272 ( 
.A(n_8815),
.B(n_5442),
.Y(n_9272)
);

NAND2xp5_ASAP7_75t_L g9273 ( 
.A(n_8818),
.B(n_5443),
.Y(n_9273)
);

NAND2xp5_ASAP7_75t_L g9274 ( 
.A(n_8819),
.B(n_5444),
.Y(n_9274)
);

INVx4_ASAP7_75t_L g9275 ( 
.A(n_8476),
.Y(n_9275)
);

NOR2xp33_ASAP7_75t_L g9276 ( 
.A(n_8611),
.B(n_5445),
.Y(n_9276)
);

AND2x2_ASAP7_75t_L g9277 ( 
.A(n_8859),
.B(n_8871),
.Y(n_9277)
);

INVx2_ASAP7_75t_L g9278 ( 
.A(n_8674),
.Y(n_9278)
);

INVx2_ASAP7_75t_L g9279 ( 
.A(n_8682),
.Y(n_9279)
);

INVx1_ASAP7_75t_L g9280 ( 
.A(n_8685),
.Y(n_9280)
);

INVx3_ASAP7_75t_L g9281 ( 
.A(n_8655),
.Y(n_9281)
);

NOR2xp33_ASAP7_75t_L g9282 ( 
.A(n_8781),
.B(n_5448),
.Y(n_9282)
);

AND2x2_ASAP7_75t_L g9283 ( 
.A(n_8741),
.B(n_8547),
.Y(n_9283)
);

NAND2xp5_ASAP7_75t_L g9284 ( 
.A(n_8692),
.B(n_5454),
.Y(n_9284)
);

HB1xp67_ASAP7_75t_L g9285 ( 
.A(n_8478),
.Y(n_9285)
);

INVx1_ASAP7_75t_L g9286 ( 
.A(n_8694),
.Y(n_9286)
);

INVx5_ASAP7_75t_L g9287 ( 
.A(n_8478),
.Y(n_9287)
);

INVx1_ASAP7_75t_L g9288 ( 
.A(n_8701),
.Y(n_9288)
);

NAND2xp5_ASAP7_75t_L g9289 ( 
.A(n_8711),
.B(n_5458),
.Y(n_9289)
);

AND2x4_ASAP7_75t_L g9290 ( 
.A(n_8519),
.B(n_4287),
.Y(n_9290)
);

INVx2_ASAP7_75t_L g9291 ( 
.A(n_8739),
.Y(n_9291)
);

INVx2_ASAP7_75t_L g9292 ( 
.A(n_8745),
.Y(n_9292)
);

NAND2xp5_ASAP7_75t_SL g9293 ( 
.A(n_8857),
.B(n_8863),
.Y(n_9293)
);

NAND2xp33_ASAP7_75t_L g9294 ( 
.A(n_8703),
.B(n_5459),
.Y(n_9294)
);

NAND2xp5_ASAP7_75t_SL g9295 ( 
.A(n_8857),
.B(n_5460),
.Y(n_9295)
);

NAND2xp5_ASAP7_75t_L g9296 ( 
.A(n_8755),
.B(n_5463),
.Y(n_9296)
);

AOI22xp5_ASAP7_75t_L g9297 ( 
.A1(n_8500),
.A2(n_5468),
.B1(n_5469),
.B2(n_5464),
.Y(n_9297)
);

NAND2xp5_ASAP7_75t_L g9298 ( 
.A(n_8757),
.B(n_8762),
.Y(n_9298)
);

NAND2xp5_ASAP7_75t_SL g9299 ( 
.A(n_8863),
.B(n_5471),
.Y(n_9299)
);

NAND2xp5_ASAP7_75t_L g9300 ( 
.A(n_8770),
.B(n_5473),
.Y(n_9300)
);

NAND2xp5_ASAP7_75t_L g9301 ( 
.A(n_8778),
.B(n_5474),
.Y(n_9301)
);

AOI22xp33_ASAP7_75t_L g9302 ( 
.A1(n_8638),
.A2(n_5480),
.B1(n_5483),
.B2(n_5477),
.Y(n_9302)
);

NAND3xp33_ASAP7_75t_L g9303 ( 
.A(n_8635),
.B(n_8873),
.C(n_8551),
.Y(n_9303)
);

NOR2xp33_ASAP7_75t_L g9304 ( 
.A(n_8894),
.B(n_5484),
.Y(n_9304)
);

INVx2_ASAP7_75t_SL g9305 ( 
.A(n_8492),
.Y(n_9305)
);

NOR2x1p5_ASAP7_75t_L g9306 ( 
.A(n_8810),
.B(n_5488),
.Y(n_9306)
);

NOR2xp33_ASAP7_75t_L g9307 ( 
.A(n_8666),
.B(n_8771),
.Y(n_9307)
);

INVx2_ASAP7_75t_L g9308 ( 
.A(n_8789),
.Y(n_9308)
);

INVx2_ASAP7_75t_L g9309 ( 
.A(n_8797),
.Y(n_9309)
);

INVx1_ASAP7_75t_L g9310 ( 
.A(n_8801),
.Y(n_9310)
);

OR2x6_ASAP7_75t_L g9311 ( 
.A(n_8807),
.B(n_4288),
.Y(n_9311)
);

INVx8_ASAP7_75t_L g9312 ( 
.A(n_8492),
.Y(n_9312)
);

NAND2xp5_ASAP7_75t_SL g9313 ( 
.A(n_8676),
.B(n_5489),
.Y(n_9313)
);

INVx1_ASAP7_75t_L g9314 ( 
.A(n_8828),
.Y(n_9314)
);

AND2x2_ASAP7_75t_SL g9315 ( 
.A(n_8807),
.B(n_8),
.Y(n_9315)
);

NAND2xp5_ASAP7_75t_L g9316 ( 
.A(n_8830),
.B(n_8832),
.Y(n_9316)
);

NAND2xp5_ASAP7_75t_SL g9317 ( 
.A(n_8676),
.B(n_8861),
.Y(n_9317)
);

INVx2_ASAP7_75t_L g9318 ( 
.A(n_8839),
.Y(n_9318)
);

NAND2xp5_ASAP7_75t_SL g9319 ( 
.A(n_8861),
.B(n_5490),
.Y(n_9319)
);

NAND2xp5_ASAP7_75t_L g9320 ( 
.A(n_8840),
.B(n_5491),
.Y(n_9320)
);

NAND2xp33_ASAP7_75t_L g9321 ( 
.A(n_8703),
.B(n_5492),
.Y(n_9321)
);

INVx1_ASAP7_75t_L g9322 ( 
.A(n_8866),
.Y(n_9322)
);

INVx2_ASAP7_75t_L g9323 ( 
.A(n_8843),
.Y(n_9323)
);

NOR2xp33_ASAP7_75t_L g9324 ( 
.A(n_8911),
.B(n_5495),
.Y(n_9324)
);

NAND2xp5_ASAP7_75t_L g9325 ( 
.A(n_8849),
.B(n_5497),
.Y(n_9325)
);

INVx1_ASAP7_75t_L g9326 ( 
.A(n_8875),
.Y(n_9326)
);

NOR2xp33_ASAP7_75t_L g9327 ( 
.A(n_8576),
.B(n_5504),
.Y(n_9327)
);

NAND2xp5_ASAP7_75t_L g9328 ( 
.A(n_8854),
.B(n_5510),
.Y(n_9328)
);

INVx1_ASAP7_75t_L g9329 ( 
.A(n_8879),
.Y(n_9329)
);

NAND2xp5_ASAP7_75t_L g9330 ( 
.A(n_8881),
.B(n_5511),
.Y(n_9330)
);

AOI22xp5_ASAP7_75t_L g9331 ( 
.A1(n_8904),
.A2(n_5517),
.B1(n_5519),
.B2(n_5512),
.Y(n_9331)
);

AOI22xp5_ASAP7_75t_L g9332 ( 
.A1(n_8571),
.A2(n_8649),
.B1(n_8704),
.B2(n_8697),
.Y(n_9332)
);

INVx2_ASAP7_75t_L g9333 ( 
.A(n_8885),
.Y(n_9333)
);

NAND2xp5_ASAP7_75t_L g9334 ( 
.A(n_8886),
.B(n_5525),
.Y(n_9334)
);

INVx2_ASAP7_75t_L g9335 ( 
.A(n_8889),
.Y(n_9335)
);

NAND2xp33_ASAP7_75t_L g9336 ( 
.A(n_8823),
.B(n_5526),
.Y(n_9336)
);

NAND2xp5_ASAP7_75t_L g9337 ( 
.A(n_8905),
.B(n_8520),
.Y(n_9337)
);

INVx2_ASAP7_75t_SL g9338 ( 
.A(n_8545),
.Y(n_9338)
);

NAND2xp5_ASAP7_75t_L g9339 ( 
.A(n_8525),
.B(n_5529),
.Y(n_9339)
);

NAND2xp5_ASAP7_75t_L g9340 ( 
.A(n_8878),
.B(n_5531),
.Y(n_9340)
);

NOR2xp33_ASAP7_75t_L g9341 ( 
.A(n_8608),
.B(n_5532),
.Y(n_9341)
);

NAND2xp5_ASAP7_75t_SL g9342 ( 
.A(n_8862),
.B(n_5533),
.Y(n_9342)
);

INVx2_ASAP7_75t_L g9343 ( 
.A(n_8852),
.Y(n_9343)
);

NAND2xp5_ASAP7_75t_SL g9344 ( 
.A(n_8862),
.B(n_5534),
.Y(n_9344)
);

INVxp67_ASAP7_75t_L g9345 ( 
.A(n_8760),
.Y(n_9345)
);

INVx1_ASAP7_75t_L g9346 ( 
.A(n_8890),
.Y(n_9346)
);

NAND2xp5_ASAP7_75t_SL g9347 ( 
.A(n_8545),
.B(n_5537),
.Y(n_9347)
);

BUFx6f_ASAP7_75t_L g9348 ( 
.A(n_8554),
.Y(n_9348)
);

INVx3_ASAP7_75t_L g9349 ( 
.A(n_8655),
.Y(n_9349)
);

INVx1_ASAP7_75t_L g9350 ( 
.A(n_8915),
.Y(n_9350)
);

INVx1_ASAP7_75t_L g9351 ( 
.A(n_8824),
.Y(n_9351)
);

AND2x2_ASAP7_75t_L g9352 ( 
.A(n_8574),
.B(n_5539),
.Y(n_9352)
);

INVx2_ASAP7_75t_L g9353 ( 
.A(n_8836),
.Y(n_9353)
);

NOR2xp33_ASAP7_75t_L g9354 ( 
.A(n_8687),
.B(n_5541),
.Y(n_9354)
);

AND2x2_ASAP7_75t_L g9355 ( 
.A(n_8620),
.B(n_5543),
.Y(n_9355)
);

NAND2xp5_ASAP7_75t_SL g9356 ( 
.A(n_8554),
.B(n_5545),
.Y(n_9356)
);

INVx2_ASAP7_75t_SL g9357 ( 
.A(n_8585),
.Y(n_9357)
);

INVx8_ASAP7_75t_L g9358 ( 
.A(n_8585),
.Y(n_9358)
);

NAND2xp5_ASAP7_75t_L g9359 ( 
.A(n_8882),
.B(n_5550),
.Y(n_9359)
);

INVx3_ASAP7_75t_L g9360 ( 
.A(n_8657),
.Y(n_9360)
);

NAND2xp5_ASAP7_75t_L g9361 ( 
.A(n_8891),
.B(n_5551),
.Y(n_9361)
);

NAND2xp5_ASAP7_75t_SL g9362 ( 
.A(n_8657),
.B(n_5554),
.Y(n_9362)
);

NAND2x1p5_ASAP7_75t_L g9363 ( 
.A(n_8483),
.B(n_4289),
.Y(n_9363)
);

OR2x6_ASAP7_75t_L g9364 ( 
.A(n_8499),
.B(n_4290),
.Y(n_9364)
);

NAND2xp5_ASAP7_75t_L g9365 ( 
.A(n_8896),
.B(n_5557),
.Y(n_9365)
);

NAND2x1_ASAP7_75t_L g9366 ( 
.A(n_8695),
.B(n_8765),
.Y(n_9366)
);

NAND2xp33_ASAP7_75t_L g9367 ( 
.A(n_8823),
.B(n_5559),
.Y(n_9367)
);

INVx1_ASAP7_75t_L g9368 ( 
.A(n_8690),
.Y(n_9368)
);

BUFx6f_ASAP7_75t_SL g9369 ( 
.A(n_8456),
.Y(n_9369)
);

BUFx6f_ASAP7_75t_L g9370 ( 
.A(n_8784),
.Y(n_9370)
);

NOR2xp33_ASAP7_75t_L g9371 ( 
.A(n_8766),
.B(n_5560),
.Y(n_9371)
);

NAND2xp5_ASAP7_75t_L g9372 ( 
.A(n_8872),
.B(n_5561),
.Y(n_9372)
);

NAND2xp5_ASAP7_75t_SL g9373 ( 
.A(n_8817),
.B(n_5562),
.Y(n_9373)
);

NOR3xp33_ASAP7_75t_L g9374 ( 
.A(n_8569),
.B(n_5569),
.C(n_5564),
.Y(n_9374)
);

NOR2xp33_ASAP7_75t_L g9375 ( 
.A(n_8783),
.B(n_5573),
.Y(n_9375)
);

INVx1_ASAP7_75t_L g9376 ( 
.A(n_8753),
.Y(n_9376)
);

NAND2xp5_ASAP7_75t_L g9377 ( 
.A(n_8793),
.B(n_5574),
.Y(n_9377)
);

NAND2xp5_ASAP7_75t_L g9378 ( 
.A(n_8795),
.B(n_5576),
.Y(n_9378)
);

HB1xp67_ASAP7_75t_L g9379 ( 
.A(n_8594),
.Y(n_9379)
);

AND2x2_ASAP7_75t_L g9380 ( 
.A(n_8646),
.B(n_5577),
.Y(n_9380)
);

INVx2_ASAP7_75t_L g9381 ( 
.A(n_8812),
.Y(n_9381)
);

INVx1_ASAP7_75t_L g9382 ( 
.A(n_8773),
.Y(n_9382)
);

AND2x4_ASAP7_75t_L g9383 ( 
.A(n_8732),
.B(n_8599),
.Y(n_9383)
);

NAND2xp5_ASAP7_75t_L g9384 ( 
.A(n_8855),
.B(n_5579),
.Y(n_9384)
);

NOR2xp67_ASAP7_75t_L g9385 ( 
.A(n_8787),
.B(n_4291),
.Y(n_9385)
);

INVx2_ASAP7_75t_L g9386 ( 
.A(n_8779),
.Y(n_9386)
);

NAND2xp5_ASAP7_75t_L g9387 ( 
.A(n_8865),
.B(n_5580),
.Y(n_9387)
);

AND2x4_ASAP7_75t_L g9388 ( 
.A(n_8784),
.B(n_8531),
.Y(n_9388)
);

OR2x6_ASAP7_75t_L g9389 ( 
.A(n_8508),
.B(n_4292),
.Y(n_9389)
);

AND2x6_ASAP7_75t_L g9390 ( 
.A(n_8811),
.B(n_4293),
.Y(n_9390)
);

O2A1O1Ixp33_ASAP7_75t_L g9391 ( 
.A1(n_8486),
.A2(n_5582),
.B(n_5583),
.C(n_5581),
.Y(n_9391)
);

NAND2xp5_ASAP7_75t_L g9392 ( 
.A(n_8842),
.B(n_5584),
.Y(n_9392)
);

INVx2_ASAP7_75t_L g9393 ( 
.A(n_8714),
.Y(n_9393)
);

INVx2_ASAP7_75t_L g9394 ( 
.A(n_8725),
.Y(n_9394)
);

INVx2_ASAP7_75t_L g9395 ( 
.A(n_8764),
.Y(n_9395)
);

AOI22xp33_ASAP7_75t_L g9396 ( 
.A1(n_8813),
.A2(n_8681),
.B1(n_8637),
.B2(n_8634),
.Y(n_9396)
);

NAND2xp5_ASAP7_75t_L g9397 ( 
.A(n_8842),
.B(n_5586),
.Y(n_9397)
);

AND2x4_ASAP7_75t_L g9398 ( 
.A(n_8777),
.B(n_4296),
.Y(n_9398)
);

NAND2xp5_ASAP7_75t_SL g9399 ( 
.A(n_8466),
.B(n_5590),
.Y(n_9399)
);

NAND2xp5_ASAP7_75t_L g9400 ( 
.A(n_8893),
.B(n_5592),
.Y(n_9400)
);

NAND2xp5_ASAP7_75t_L g9401 ( 
.A(n_8813),
.B(n_8785),
.Y(n_9401)
);

NAND2xp5_ASAP7_75t_L g9402 ( 
.A(n_8918),
.B(n_5593),
.Y(n_9402)
);

INVx1_ASAP7_75t_L g9403 ( 
.A(n_8737),
.Y(n_9403)
);

INVx2_ASAP7_75t_L g9404 ( 
.A(n_8811),
.Y(n_9404)
);

OR2x2_ASAP7_75t_L g9405 ( 
.A(n_8724),
.B(n_5597),
.Y(n_9405)
);

INVx1_ASAP7_75t_L g9406 ( 
.A(n_8509),
.Y(n_9406)
);

NAND2xp5_ASAP7_75t_L g9407 ( 
.A(n_8601),
.B(n_5602),
.Y(n_9407)
);

AND2x2_ASAP7_75t_L g9408 ( 
.A(n_8867),
.B(n_5603),
.Y(n_9408)
);

NAND2xp5_ASAP7_75t_L g9409 ( 
.A(n_8601),
.B(n_5604),
.Y(n_9409)
);

NOR2xp33_ASAP7_75t_L g9410 ( 
.A(n_8743),
.B(n_5605),
.Y(n_9410)
);

NAND2xp5_ASAP7_75t_L g9411 ( 
.A(n_8630),
.B(n_5606),
.Y(n_9411)
);

NOR2xp67_ASAP7_75t_L g9412 ( 
.A(n_8754),
.B(n_4297),
.Y(n_9412)
);

INVx2_ASAP7_75t_L g9413 ( 
.A(n_8729),
.Y(n_9413)
);

INVx2_ASAP7_75t_SL g9414 ( 
.A(n_8561),
.Y(n_9414)
);

INVx1_ASAP7_75t_L g9415 ( 
.A(n_8750),
.Y(n_9415)
);

INVx2_ASAP7_75t_L g9416 ( 
.A(n_8910),
.Y(n_9416)
);

INVxp67_ASAP7_75t_L g9417 ( 
.A(n_8538),
.Y(n_9417)
);

AND2x4_ASAP7_75t_L g9418 ( 
.A(n_8848),
.B(n_4299),
.Y(n_9418)
);

NAND2xp5_ASAP7_75t_SL g9419 ( 
.A(n_8582),
.B(n_5608),
.Y(n_9419)
);

INVx4_ASAP7_75t_L g9420 ( 
.A(n_8734),
.Y(n_9420)
);

HB1xp67_ASAP7_75t_L g9421 ( 
.A(n_8707),
.Y(n_9421)
);

NAND2xp5_ASAP7_75t_SL g9422 ( 
.A(n_8615),
.B(n_5609),
.Y(n_9422)
);

INVx1_ASAP7_75t_L g9423 ( 
.A(n_8485),
.Y(n_9423)
);

AND2x2_ASAP7_75t_L g9424 ( 
.A(n_8661),
.B(n_5610),
.Y(n_9424)
);

NAND2xp5_ASAP7_75t_L g9425 ( 
.A(n_8630),
.B(n_5611),
.Y(n_9425)
);

HB1xp67_ASAP7_75t_L g9426 ( 
.A(n_8922),
.Y(n_9426)
);

NOR2xp67_ASAP7_75t_L g9427 ( 
.A(n_8798),
.B(n_4300),
.Y(n_9427)
);

NAND2xp5_ASAP7_75t_SL g9428 ( 
.A(n_8552),
.B(n_5612),
.Y(n_9428)
);

O2A1O1Ixp5_ASAP7_75t_L g9429 ( 
.A1(n_8895),
.A2(n_11),
.B(n_9),
.C(n_10),
.Y(n_9429)
);

NAND2xp5_ASAP7_75t_SL g9430 ( 
.A(n_8538),
.B(n_5615),
.Y(n_9430)
);

HB1xp67_ASAP7_75t_L g9431 ( 
.A(n_8568),
.Y(n_9431)
);

OR2x2_ASAP7_75t_L g9432 ( 
.A(n_8588),
.B(n_5617),
.Y(n_9432)
);

INVx1_ASAP7_75t_L g9433 ( 
.A(n_8568),
.Y(n_9433)
);

NAND2xp5_ASAP7_75t_SL g9434 ( 
.A(n_8592),
.B(n_5618),
.Y(n_9434)
);

NAND2xp5_ASAP7_75t_SL g9435 ( 
.A(n_8592),
.B(n_5622),
.Y(n_9435)
);

NOR2xp33_ASAP7_75t_L g9436 ( 
.A(n_8917),
.B(n_5624),
.Y(n_9436)
);

AND2x2_ASAP7_75t_L g9437 ( 
.A(n_8426),
.B(n_5626),
.Y(n_9437)
);

AND2x2_ASAP7_75t_L g9438 ( 
.A(n_8426),
.B(n_5627),
.Y(n_9438)
);

NAND2xp5_ASAP7_75t_L g9439 ( 
.A(n_8426),
.B(n_5630),
.Y(n_9439)
);

NAND2xp5_ASAP7_75t_L g9440 ( 
.A(n_8426),
.B(n_5631),
.Y(n_9440)
);

INVx1_ASAP7_75t_L g9441 ( 
.A(n_8414),
.Y(n_9441)
);

INVx1_ASAP7_75t_L g9442 ( 
.A(n_8414),
.Y(n_9442)
);

NAND2xp5_ASAP7_75t_L g9443 ( 
.A(n_9012),
.B(n_5632),
.Y(n_9443)
);

INVx2_ASAP7_75t_L g9444 ( 
.A(n_8932),
.Y(n_9444)
);

INVx1_ASAP7_75t_SL g9445 ( 
.A(n_9213),
.Y(n_9445)
);

AND2x4_ASAP7_75t_L g9446 ( 
.A(n_8979),
.B(n_4301),
.Y(n_9446)
);

AND2x2_ASAP7_75t_L g9447 ( 
.A(n_9051),
.B(n_5634),
.Y(n_9447)
);

INVx4_ASAP7_75t_L g9448 ( 
.A(n_9022),
.Y(n_9448)
);

INVx2_ASAP7_75t_L g9449 ( 
.A(n_8935),
.Y(n_9449)
);

OAI21xp5_ASAP7_75t_L g9450 ( 
.A1(n_8960),
.A2(n_5638),
.B(n_5637),
.Y(n_9450)
);

NAND2xp5_ASAP7_75t_L g9451 ( 
.A(n_9437),
.B(n_5639),
.Y(n_9451)
);

AND2x2_ASAP7_75t_L g9452 ( 
.A(n_8954),
.B(n_8926),
.Y(n_9452)
);

AND2x2_ASAP7_75t_L g9453 ( 
.A(n_9209),
.B(n_5641),
.Y(n_9453)
);

OAI21x1_ASAP7_75t_L g9454 ( 
.A1(n_8971),
.A2(n_4303),
.B(n_4302),
.Y(n_9454)
);

AOI22xp5_ASAP7_75t_L g9455 ( 
.A1(n_8952),
.A2(n_5645),
.B1(n_5647),
.B2(n_5642),
.Y(n_9455)
);

NAND2xp5_ASAP7_75t_L g9456 ( 
.A(n_9438),
.B(n_5648),
.Y(n_9456)
);

INVx2_ASAP7_75t_L g9457 ( 
.A(n_8940),
.Y(n_9457)
);

BUFx3_ASAP7_75t_L g9458 ( 
.A(n_9022),
.Y(n_9458)
);

INVx2_ASAP7_75t_L g9459 ( 
.A(n_8947),
.Y(n_9459)
);

NAND2xp5_ASAP7_75t_L g9460 ( 
.A(n_8929),
.B(n_5650),
.Y(n_9460)
);

INVx3_ASAP7_75t_L g9461 ( 
.A(n_8998),
.Y(n_9461)
);

NAND2xp5_ASAP7_75t_L g9462 ( 
.A(n_8933),
.B(n_5651),
.Y(n_9462)
);

INVx1_ASAP7_75t_L g9463 ( 
.A(n_9111),
.Y(n_9463)
);

INVx2_ASAP7_75t_L g9464 ( 
.A(n_8956),
.Y(n_9464)
);

NAND2xp5_ASAP7_75t_L g9465 ( 
.A(n_8977),
.B(n_5655),
.Y(n_9465)
);

HB1xp67_ASAP7_75t_L g9466 ( 
.A(n_8973),
.Y(n_9466)
);

BUFx3_ASAP7_75t_L g9467 ( 
.A(n_9242),
.Y(n_9467)
);

INVx2_ASAP7_75t_L g9468 ( 
.A(n_8959),
.Y(n_9468)
);

NAND2xp5_ASAP7_75t_SL g9469 ( 
.A(n_8949),
.B(n_5658),
.Y(n_9469)
);

INVx3_ASAP7_75t_L g9470 ( 
.A(n_9211),
.Y(n_9470)
);

INVx3_ASAP7_75t_L g9471 ( 
.A(n_9370),
.Y(n_9471)
);

NAND2xp5_ASAP7_75t_L g9472 ( 
.A(n_8937),
.B(n_5659),
.Y(n_9472)
);

INVx2_ASAP7_75t_L g9473 ( 
.A(n_8982),
.Y(n_9473)
);

NAND2xp5_ASAP7_75t_SL g9474 ( 
.A(n_8950),
.B(n_5662),
.Y(n_9474)
);

INVx2_ASAP7_75t_L g9475 ( 
.A(n_8992),
.Y(n_9475)
);

AND2x2_ASAP7_75t_L g9476 ( 
.A(n_9139),
.B(n_5663),
.Y(n_9476)
);

INVx2_ASAP7_75t_L g9477 ( 
.A(n_8994),
.Y(n_9477)
);

INVx1_ASAP7_75t_SL g9478 ( 
.A(n_9029),
.Y(n_9478)
);

NAND2xp5_ASAP7_75t_L g9479 ( 
.A(n_9439),
.B(n_5664),
.Y(n_9479)
);

AND2x2_ASAP7_75t_L g9480 ( 
.A(n_9058),
.B(n_5665),
.Y(n_9480)
);

AND2x2_ASAP7_75t_L g9481 ( 
.A(n_9131),
.B(n_5669),
.Y(n_9481)
);

INVx1_ASAP7_75t_L g9482 ( 
.A(n_9004),
.Y(n_9482)
);

INVx2_ASAP7_75t_L g9483 ( 
.A(n_9014),
.Y(n_9483)
);

AND2x4_ASAP7_75t_L g9484 ( 
.A(n_9104),
.B(n_4304),
.Y(n_9484)
);

AND2x2_ASAP7_75t_SL g9485 ( 
.A(n_9315),
.B(n_10),
.Y(n_9485)
);

INVx2_ASAP7_75t_SL g9486 ( 
.A(n_9242),
.Y(n_9486)
);

INVx1_ASAP7_75t_SL g9487 ( 
.A(n_9239),
.Y(n_9487)
);

OR2x2_ASAP7_75t_L g9488 ( 
.A(n_8928),
.B(n_5676),
.Y(n_9488)
);

INVx1_ASAP7_75t_SL g9489 ( 
.A(n_9262),
.Y(n_9489)
);

INVx1_ASAP7_75t_L g9490 ( 
.A(n_9015),
.Y(n_9490)
);

HB1xp67_ASAP7_75t_L g9491 ( 
.A(n_8991),
.Y(n_9491)
);

NAND2xp5_ASAP7_75t_L g9492 ( 
.A(n_9440),
.B(n_5678),
.Y(n_9492)
);

AND2x2_ASAP7_75t_L g9493 ( 
.A(n_9128),
.B(n_5680),
.Y(n_9493)
);

INVxp67_ASAP7_75t_SL g9494 ( 
.A(n_8946),
.Y(n_9494)
);

AND2x4_ASAP7_75t_L g9495 ( 
.A(n_9181),
.B(n_4305),
.Y(n_9495)
);

AND2x2_ASAP7_75t_SL g9496 ( 
.A(n_8958),
.B(n_11),
.Y(n_9496)
);

INVx1_ASAP7_75t_L g9497 ( 
.A(n_9017),
.Y(n_9497)
);

INVx1_ASAP7_75t_L g9498 ( 
.A(n_9030),
.Y(n_9498)
);

INVx2_ASAP7_75t_L g9499 ( 
.A(n_9041),
.Y(n_9499)
);

INVx3_ASAP7_75t_L g9500 ( 
.A(n_9370),
.Y(n_9500)
);

AND2x2_ASAP7_75t_L g9501 ( 
.A(n_9283),
.B(n_9277),
.Y(n_9501)
);

INVx1_ASAP7_75t_L g9502 ( 
.A(n_9052),
.Y(n_9502)
);

NAND2xp5_ASAP7_75t_SL g9503 ( 
.A(n_8961),
.B(n_5682),
.Y(n_9503)
);

BUFx8_ASAP7_75t_L g9504 ( 
.A(n_9100),
.Y(n_9504)
);

NAND2xp5_ASAP7_75t_L g9505 ( 
.A(n_9025),
.B(n_5683),
.Y(n_9505)
);

INVx3_ASAP7_75t_L g9506 ( 
.A(n_9383),
.Y(n_9506)
);

INVx4_ASAP7_75t_L g9507 ( 
.A(n_9165),
.Y(n_9507)
);

INVx2_ASAP7_75t_L g9508 ( 
.A(n_9054),
.Y(n_9508)
);

OAI21xp5_ASAP7_75t_L g9509 ( 
.A1(n_8976),
.A2(n_5692),
.B(n_5687),
.Y(n_9509)
);

INVx2_ASAP7_75t_L g9510 ( 
.A(n_9070),
.Y(n_9510)
);

OR2x2_ASAP7_75t_SL g9511 ( 
.A(n_9431),
.B(n_5698),
.Y(n_9511)
);

NAND2xp5_ASAP7_75t_L g9512 ( 
.A(n_9026),
.B(n_12),
.Y(n_9512)
);

AND2x4_ASAP7_75t_L g9513 ( 
.A(n_9388),
.B(n_4306),
.Y(n_9513)
);

INVx2_ASAP7_75t_L g9514 ( 
.A(n_9073),
.Y(n_9514)
);

BUFx24_ASAP7_75t_L g9515 ( 
.A(n_9215),
.Y(n_9515)
);

INVx2_ASAP7_75t_SL g9516 ( 
.A(n_9312),
.Y(n_9516)
);

HB1xp67_ASAP7_75t_L g9517 ( 
.A(n_9050),
.Y(n_9517)
);

OR2x4_ASAP7_75t_L g9518 ( 
.A(n_9078),
.B(n_12),
.Y(n_9518)
);

AND2x2_ASAP7_75t_L g9519 ( 
.A(n_8957),
.B(n_13),
.Y(n_9519)
);

NOR2xp33_ASAP7_75t_L g9520 ( 
.A(n_8943),
.B(n_4307),
.Y(n_9520)
);

AND2x2_ASAP7_75t_L g9521 ( 
.A(n_9249),
.B(n_14),
.Y(n_9521)
);

AND2x2_ASAP7_75t_L g9522 ( 
.A(n_9352),
.B(n_14),
.Y(n_9522)
);

INVx1_ASAP7_75t_L g9523 ( 
.A(n_9076),
.Y(n_9523)
);

CKINVDCx5p33_ASAP7_75t_R g9524 ( 
.A(n_8990),
.Y(n_9524)
);

AND2x2_ASAP7_75t_L g9525 ( 
.A(n_9355),
.B(n_15),
.Y(n_9525)
);

INVx1_ASAP7_75t_SL g9526 ( 
.A(n_9379),
.Y(n_9526)
);

NAND2xp5_ASAP7_75t_L g9527 ( 
.A(n_9059),
.B(n_15),
.Y(n_9527)
);

NOR2xp33_ASAP7_75t_L g9528 ( 
.A(n_8963),
.B(n_4308),
.Y(n_9528)
);

NOR2xp33_ASAP7_75t_L g9529 ( 
.A(n_8944),
.B(n_4309),
.Y(n_9529)
);

NAND2xp5_ASAP7_75t_L g9530 ( 
.A(n_8931),
.B(n_16),
.Y(n_9530)
);

INVx1_ASAP7_75t_L g9531 ( 
.A(n_9084),
.Y(n_9531)
);

AND2x2_ASAP7_75t_L g9532 ( 
.A(n_9380),
.B(n_17),
.Y(n_9532)
);

AND2x4_ASAP7_75t_L g9533 ( 
.A(n_9042),
.B(n_4310),
.Y(n_9533)
);

CKINVDCx5p33_ASAP7_75t_R g9534 ( 
.A(n_9019),
.Y(n_9534)
);

INVx2_ASAP7_75t_SL g9535 ( 
.A(n_9312),
.Y(n_9535)
);

INVxp67_ASAP7_75t_SL g9536 ( 
.A(n_9346),
.Y(n_9536)
);

AND2x4_ASAP7_75t_L g9537 ( 
.A(n_9404),
.B(n_4312),
.Y(n_9537)
);

NOR2xp33_ASAP7_75t_L g9538 ( 
.A(n_9226),
.B(n_4313),
.Y(n_9538)
);

AND2x2_ASAP7_75t_SL g9539 ( 
.A(n_9423),
.B(n_17),
.Y(n_9539)
);

INVx3_ASAP7_75t_L g9540 ( 
.A(n_9048),
.Y(n_9540)
);

INVx1_ASAP7_75t_L g9541 ( 
.A(n_9087),
.Y(n_9541)
);

INVx4_ASAP7_75t_L g9542 ( 
.A(n_9165),
.Y(n_9542)
);

NAND2xp5_ASAP7_75t_L g9543 ( 
.A(n_8966),
.B(n_19),
.Y(n_9543)
);

INVx1_ASAP7_75t_L g9544 ( 
.A(n_9090),
.Y(n_9544)
);

INVx2_ASAP7_75t_L g9545 ( 
.A(n_9091),
.Y(n_9545)
);

INVx1_ASAP7_75t_L g9546 ( 
.A(n_9096),
.Y(n_9546)
);

AND2x2_ASAP7_75t_L g9547 ( 
.A(n_9304),
.B(n_19),
.Y(n_9547)
);

INVx3_ASAP7_75t_L g9548 ( 
.A(n_9048),
.Y(n_9548)
);

AND2x2_ASAP7_75t_SL g9549 ( 
.A(n_9418),
.B(n_20),
.Y(n_9549)
);

INVx1_ASAP7_75t_L g9550 ( 
.A(n_9103),
.Y(n_9550)
);

HB1xp67_ASAP7_75t_L g9551 ( 
.A(n_9184),
.Y(n_9551)
);

OAI21xp5_ASAP7_75t_L g9552 ( 
.A1(n_9324),
.A2(n_20),
.B(n_21),
.Y(n_9552)
);

HB1xp67_ASAP7_75t_L g9553 ( 
.A(n_9285),
.Y(n_9553)
);

AND2x2_ASAP7_75t_SL g9554 ( 
.A(n_9420),
.B(n_9037),
.Y(n_9554)
);

INVx1_ASAP7_75t_L g9555 ( 
.A(n_9105),
.Y(n_9555)
);

INVx1_ASAP7_75t_SL g9556 ( 
.A(n_9152),
.Y(n_9556)
);

INVxp67_ASAP7_75t_SL g9557 ( 
.A(n_9046),
.Y(n_9557)
);

AND2x2_ASAP7_75t_L g9558 ( 
.A(n_9251),
.B(n_21),
.Y(n_9558)
);

INVx1_ASAP7_75t_L g9559 ( 
.A(n_9117),
.Y(n_9559)
);

INVx1_ASAP7_75t_L g9560 ( 
.A(n_9123),
.Y(n_9560)
);

BUFx6f_ASAP7_75t_L g9561 ( 
.A(n_8972),
.Y(n_9561)
);

INVx2_ASAP7_75t_L g9562 ( 
.A(n_9127),
.Y(n_9562)
);

INVx1_ASAP7_75t_L g9563 ( 
.A(n_8927),
.Y(n_9563)
);

NAND2xp5_ASAP7_75t_L g9564 ( 
.A(n_9067),
.B(n_22),
.Y(n_9564)
);

AND2x2_ASAP7_75t_SL g9565 ( 
.A(n_9396),
.B(n_22),
.Y(n_9565)
);

AND2x2_ASAP7_75t_L g9566 ( 
.A(n_9265),
.B(n_23),
.Y(n_9566)
);

BUFx3_ASAP7_75t_L g9567 ( 
.A(n_9358),
.Y(n_9567)
);

NAND2xp5_ASAP7_75t_L g9568 ( 
.A(n_9337),
.B(n_23),
.Y(n_9568)
);

NAND2xp5_ASAP7_75t_L g9569 ( 
.A(n_8948),
.B(n_24),
.Y(n_9569)
);

INVx1_ASAP7_75t_L g9570 ( 
.A(n_8930),
.Y(n_9570)
);

OR2x2_ASAP7_75t_L g9571 ( 
.A(n_8987),
.B(n_24),
.Y(n_9571)
);

AND2x2_ASAP7_75t_L g9572 ( 
.A(n_9276),
.B(n_25),
.Y(n_9572)
);

BUFx3_ASAP7_75t_L g9573 ( 
.A(n_9358),
.Y(n_9573)
);

INVx1_ASAP7_75t_L g9574 ( 
.A(n_8969),
.Y(n_9574)
);

BUFx6f_ASAP7_75t_L g9575 ( 
.A(n_8972),
.Y(n_9575)
);

NAND2xp5_ASAP7_75t_L g9576 ( 
.A(n_9268),
.B(n_25),
.Y(n_9576)
);

INVx2_ASAP7_75t_L g9577 ( 
.A(n_9161),
.Y(n_9577)
);

BUFx3_ASAP7_75t_L g9578 ( 
.A(n_9125),
.Y(n_9578)
);

INVx1_ASAP7_75t_L g9579 ( 
.A(n_8978),
.Y(n_9579)
);

INVx3_ASAP7_75t_L g9580 ( 
.A(n_9153),
.Y(n_9580)
);

NAND2xp5_ASAP7_75t_L g9581 ( 
.A(n_8995),
.B(n_26),
.Y(n_9581)
);

NAND2xp5_ASAP7_75t_L g9582 ( 
.A(n_8996),
.B(n_26),
.Y(n_9582)
);

NAND2xp5_ASAP7_75t_L g9583 ( 
.A(n_9245),
.B(n_27),
.Y(n_9583)
);

BUFx6f_ASAP7_75t_L g9584 ( 
.A(n_9125),
.Y(n_9584)
);

AND2x2_ASAP7_75t_L g9585 ( 
.A(n_9207),
.B(n_27),
.Y(n_9585)
);

HB1xp67_ASAP7_75t_L g9586 ( 
.A(n_9345),
.Y(n_9586)
);

AND2x2_ASAP7_75t_L g9587 ( 
.A(n_9216),
.B(n_28),
.Y(n_9587)
);

INVx2_ASAP7_75t_L g9588 ( 
.A(n_9178),
.Y(n_9588)
);

BUFx6f_ASAP7_75t_L g9589 ( 
.A(n_9264),
.Y(n_9589)
);

BUFx3_ASAP7_75t_L g9590 ( 
.A(n_9264),
.Y(n_9590)
);

INVx1_ASAP7_75t_L g9591 ( 
.A(n_8980),
.Y(n_9591)
);

AND2x2_ASAP7_75t_L g9592 ( 
.A(n_9217),
.B(n_29),
.Y(n_9592)
);

INVxp67_ASAP7_75t_L g9593 ( 
.A(n_9002),
.Y(n_9593)
);

INVx2_ASAP7_75t_L g9594 ( 
.A(n_9180),
.Y(n_9594)
);

INVx2_ASAP7_75t_L g9595 ( 
.A(n_9188),
.Y(n_9595)
);

NOR2xp33_ASAP7_75t_L g9596 ( 
.A(n_8968),
.B(n_8964),
.Y(n_9596)
);

AND2x2_ASAP7_75t_L g9597 ( 
.A(n_9218),
.B(n_29),
.Y(n_9597)
);

AOI22xp5_ASAP7_75t_L g9598 ( 
.A1(n_9307),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_9598)
);

INVx2_ASAP7_75t_L g9599 ( 
.A(n_9333),
.Y(n_9599)
);

AND2x4_ASAP7_75t_L g9600 ( 
.A(n_9281),
.B(n_4314),
.Y(n_9600)
);

AND2x2_ASAP7_75t_L g9601 ( 
.A(n_9219),
.B(n_31),
.Y(n_9601)
);

NAND2xp5_ASAP7_75t_SL g9602 ( 
.A(n_8925),
.B(n_32),
.Y(n_9602)
);

AND2x2_ASAP7_75t_L g9603 ( 
.A(n_9408),
.B(n_33),
.Y(n_9603)
);

INVx1_ASAP7_75t_SL g9604 ( 
.A(n_9094),
.Y(n_9604)
);

INVx2_ASAP7_75t_L g9605 ( 
.A(n_9335),
.Y(n_9605)
);

AND2x2_ASAP7_75t_L g9606 ( 
.A(n_9238),
.B(n_33),
.Y(n_9606)
);

INVx2_ASAP7_75t_L g9607 ( 
.A(n_9192),
.Y(n_9607)
);

INVx1_ASAP7_75t_L g9608 ( 
.A(n_8988),
.Y(n_9608)
);

BUFx4_ASAP7_75t_SL g9609 ( 
.A(n_9157),
.Y(n_9609)
);

HB1xp67_ASAP7_75t_L g9610 ( 
.A(n_9165),
.Y(n_9610)
);

INVx2_ASAP7_75t_L g9611 ( 
.A(n_9197),
.Y(n_9611)
);

BUFx6f_ASAP7_75t_L g9612 ( 
.A(n_9348),
.Y(n_9612)
);

AND2x4_ASAP7_75t_L g9613 ( 
.A(n_9349),
.B(n_4316),
.Y(n_9613)
);

AND2x2_ASAP7_75t_L g9614 ( 
.A(n_9290),
.B(n_34),
.Y(n_9614)
);

NAND2xp5_ASAP7_75t_L g9615 ( 
.A(n_9038),
.B(n_34),
.Y(n_9615)
);

INVx1_ASAP7_75t_L g9616 ( 
.A(n_8997),
.Y(n_9616)
);

NAND2xp5_ASAP7_75t_L g9617 ( 
.A(n_9001),
.B(n_35),
.Y(n_9617)
);

INVxp67_ASAP7_75t_SL g9618 ( 
.A(n_9193),
.Y(n_9618)
);

CKINVDCx5p33_ASAP7_75t_R g9619 ( 
.A(n_8962),
.Y(n_9619)
);

HB1xp67_ASAP7_75t_L g9620 ( 
.A(n_9185),
.Y(n_9620)
);

INVx2_ASAP7_75t_L g9621 ( 
.A(n_9214),
.Y(n_9621)
);

INVx1_ASAP7_75t_L g9622 ( 
.A(n_9011),
.Y(n_9622)
);

AND2x2_ASAP7_75t_L g9623 ( 
.A(n_9368),
.B(n_35),
.Y(n_9623)
);

NOR2xp33_ASAP7_75t_L g9624 ( 
.A(n_8939),
.B(n_4317),
.Y(n_9624)
);

AND2x4_ASAP7_75t_L g9625 ( 
.A(n_9360),
.B(n_4319),
.Y(n_9625)
);

AND2x2_ASAP7_75t_L g9626 ( 
.A(n_9083),
.B(n_36),
.Y(n_9626)
);

AND2x4_ASAP7_75t_L g9627 ( 
.A(n_9416),
.B(n_9240),
.Y(n_9627)
);

INVx2_ASAP7_75t_L g9628 ( 
.A(n_9224),
.Y(n_9628)
);

INVx1_ASAP7_75t_L g9629 ( 
.A(n_9020),
.Y(n_9629)
);

INVx1_ASAP7_75t_L g9630 ( 
.A(n_9039),
.Y(n_9630)
);

BUFx6f_ASAP7_75t_L g9631 ( 
.A(n_9348),
.Y(n_9631)
);

BUFx6f_ASAP7_75t_L g9632 ( 
.A(n_9185),
.Y(n_9632)
);

BUFx6f_ASAP7_75t_L g9633 ( 
.A(n_9185),
.Y(n_9633)
);

NAND2xp5_ASAP7_75t_L g9634 ( 
.A(n_9005),
.B(n_36),
.Y(n_9634)
);

BUFx6f_ASAP7_75t_L g9635 ( 
.A(n_9287),
.Y(n_9635)
);

INVx2_ASAP7_75t_L g9636 ( 
.A(n_9233),
.Y(n_9636)
);

AND2x2_ASAP7_75t_L g9637 ( 
.A(n_9386),
.B(n_37),
.Y(n_9637)
);

NAND2xp5_ASAP7_75t_L g9638 ( 
.A(n_9007),
.B(n_37),
.Y(n_9638)
);

BUFx2_ASAP7_75t_L g9639 ( 
.A(n_9287),
.Y(n_9639)
);

NAND2xp5_ASAP7_75t_SL g9640 ( 
.A(n_9053),
.B(n_38),
.Y(n_9640)
);

INVx2_ASAP7_75t_L g9641 ( 
.A(n_9252),
.Y(n_9641)
);

NAND2xp5_ASAP7_75t_SL g9642 ( 
.A(n_9332),
.B(n_38),
.Y(n_9642)
);

AND2x2_ASAP7_75t_L g9643 ( 
.A(n_9278),
.B(n_39),
.Y(n_9643)
);

AND2x2_ASAP7_75t_L g9644 ( 
.A(n_9279),
.B(n_39),
.Y(n_9644)
);

INVx3_ASAP7_75t_L g9645 ( 
.A(n_9247),
.Y(n_9645)
);

INVx2_ASAP7_75t_SL g9646 ( 
.A(n_9287),
.Y(n_9646)
);

INVx1_ASAP7_75t_L g9647 ( 
.A(n_9040),
.Y(n_9647)
);

AND2x2_ASAP7_75t_L g9648 ( 
.A(n_9291),
.B(n_40),
.Y(n_9648)
);

INVx2_ASAP7_75t_L g9649 ( 
.A(n_9292),
.Y(n_9649)
);

NAND2xp5_ASAP7_75t_L g9650 ( 
.A(n_9008),
.B(n_40),
.Y(n_9650)
);

INVx2_ASAP7_75t_L g9651 ( 
.A(n_9308),
.Y(n_9651)
);

HB1xp67_ASAP7_75t_L g9652 ( 
.A(n_9208),
.Y(n_9652)
);

AND2x2_ASAP7_75t_L g9653 ( 
.A(n_9309),
.B(n_41),
.Y(n_9653)
);

CKINVDCx5p33_ASAP7_75t_R g9654 ( 
.A(n_9266),
.Y(n_9654)
);

INVx3_ASAP7_75t_L g9655 ( 
.A(n_9275),
.Y(n_9655)
);

INVx1_ASAP7_75t_L g9656 ( 
.A(n_9061),
.Y(n_9656)
);

BUFx6f_ASAP7_75t_L g9657 ( 
.A(n_8934),
.Y(n_9657)
);

AND2x2_ASAP7_75t_L g9658 ( 
.A(n_9318),
.B(n_9323),
.Y(n_9658)
);

HB1xp67_ASAP7_75t_L g9659 ( 
.A(n_9305),
.Y(n_9659)
);

INVx1_ASAP7_75t_L g9660 ( 
.A(n_9080),
.Y(n_9660)
);

AO21x1_ASAP7_75t_L g9661 ( 
.A1(n_8936),
.A2(n_41),
.B(n_42),
.Y(n_9661)
);

INVx1_ASAP7_75t_L g9662 ( 
.A(n_9081),
.Y(n_9662)
);

INVx3_ASAP7_75t_L g9663 ( 
.A(n_9119),
.Y(n_9663)
);

INVx1_ASAP7_75t_L g9664 ( 
.A(n_9088),
.Y(n_9664)
);

NAND2xp5_ASAP7_75t_L g9665 ( 
.A(n_9016),
.B(n_42),
.Y(n_9665)
);

OAI21x1_ASAP7_75t_L g9666 ( 
.A1(n_9230),
.A2(n_4321),
.B(n_4320),
.Y(n_9666)
);

AND2x2_ASAP7_75t_L g9667 ( 
.A(n_8983),
.B(n_43),
.Y(n_9667)
);

NAND2xp5_ASAP7_75t_SL g9668 ( 
.A(n_8955),
.B(n_43),
.Y(n_9668)
);

INVx4_ASAP7_75t_L g9669 ( 
.A(n_9269),
.Y(n_9669)
);

BUFx3_ASAP7_75t_L g9670 ( 
.A(n_9089),
.Y(n_9670)
);

BUFx3_ASAP7_75t_L g9671 ( 
.A(n_9338),
.Y(n_9671)
);

INVx1_ASAP7_75t_L g9672 ( 
.A(n_9102),
.Y(n_9672)
);

NAND2xp5_ASAP7_75t_L g9673 ( 
.A(n_9010),
.B(n_44),
.Y(n_9673)
);

NAND2x1p5_ASAP7_75t_L g9674 ( 
.A(n_9366),
.B(n_44),
.Y(n_9674)
);

NOR2xp67_ASAP7_75t_L g9675 ( 
.A(n_9381),
.B(n_45),
.Y(n_9675)
);

OR2x2_ASAP7_75t_L g9676 ( 
.A(n_8989),
.B(n_46),
.Y(n_9676)
);

NOR2xp33_ASAP7_75t_L g9677 ( 
.A(n_8970),
.B(n_46),
.Y(n_9677)
);

INVxp67_ASAP7_75t_L g9678 ( 
.A(n_9166),
.Y(n_9678)
);

BUFx6f_ASAP7_75t_L g9679 ( 
.A(n_8938),
.Y(n_9679)
);

INVx2_ASAP7_75t_L g9680 ( 
.A(n_9106),
.Y(n_9680)
);

NAND2xp5_ASAP7_75t_L g9681 ( 
.A(n_9013),
.B(n_47),
.Y(n_9681)
);

NAND2xp5_ASAP7_75t_L g9682 ( 
.A(n_9027),
.B(n_47),
.Y(n_9682)
);

AND2x2_ASAP7_75t_L g9683 ( 
.A(n_9018),
.B(n_9003),
.Y(n_9683)
);

INVx1_ASAP7_75t_L g9684 ( 
.A(n_9115),
.Y(n_9684)
);

INVx3_ASAP7_75t_L g9685 ( 
.A(n_9033),
.Y(n_9685)
);

INVx4_ASAP7_75t_L g9686 ( 
.A(n_9085),
.Y(n_9686)
);

INVx2_ASAP7_75t_L g9687 ( 
.A(n_9134),
.Y(n_9687)
);

OAI21xp5_ASAP7_75t_L g9688 ( 
.A1(n_9047),
.A2(n_48),
.B(n_49),
.Y(n_9688)
);

INVx2_ASAP7_75t_L g9689 ( 
.A(n_9135),
.Y(n_9689)
);

NAND2xp5_ASAP7_75t_L g9690 ( 
.A(n_9032),
.B(n_48),
.Y(n_9690)
);

INVx2_ASAP7_75t_L g9691 ( 
.A(n_9137),
.Y(n_9691)
);

INVx1_ASAP7_75t_SL g9692 ( 
.A(n_9009),
.Y(n_9692)
);

INVx1_ASAP7_75t_L g9693 ( 
.A(n_9138),
.Y(n_9693)
);

INVx1_ASAP7_75t_L g9694 ( 
.A(n_9140),
.Y(n_9694)
);

INVx2_ASAP7_75t_L g9695 ( 
.A(n_9162),
.Y(n_9695)
);

BUFx3_ASAP7_75t_L g9696 ( 
.A(n_9357),
.Y(n_9696)
);

INVx3_ASAP7_75t_SL g9697 ( 
.A(n_9049),
.Y(n_9697)
);

NAND2xp5_ASAP7_75t_SL g9698 ( 
.A(n_9401),
.B(n_51),
.Y(n_9698)
);

INVx1_ASAP7_75t_L g9699 ( 
.A(n_9441),
.Y(n_9699)
);

INVx1_ASAP7_75t_L g9700 ( 
.A(n_9442),
.Y(n_9700)
);

AND2x2_ASAP7_75t_L g9701 ( 
.A(n_8975),
.B(n_9195),
.Y(n_9701)
);

INVx2_ASAP7_75t_L g9702 ( 
.A(n_9133),
.Y(n_9702)
);

INVx2_ASAP7_75t_L g9703 ( 
.A(n_9174),
.Y(n_9703)
);

NAND2xp5_ASAP7_75t_SL g9704 ( 
.A(n_8951),
.B(n_51),
.Y(n_9704)
);

AND2x2_ASAP7_75t_L g9705 ( 
.A(n_9376),
.B(n_52),
.Y(n_9705)
);

INVx2_ASAP7_75t_SL g9706 ( 
.A(n_8942),
.Y(n_9706)
);

HB1xp67_ASAP7_75t_L g9707 ( 
.A(n_9382),
.Y(n_9707)
);

INVx1_ASAP7_75t_SL g9708 ( 
.A(n_9393),
.Y(n_9708)
);

INVx1_ASAP7_75t_L g9709 ( 
.A(n_9200),
.Y(n_9709)
);

AND2x2_ASAP7_75t_L g9710 ( 
.A(n_9327),
.B(n_53),
.Y(n_9710)
);

NAND2xp5_ASAP7_75t_L g9711 ( 
.A(n_9035),
.B(n_54),
.Y(n_9711)
);

NAND2xp5_ASAP7_75t_L g9712 ( 
.A(n_9196),
.B(n_55),
.Y(n_9712)
);

INVx2_ASAP7_75t_L g9713 ( 
.A(n_9191),
.Y(n_9713)
);

INVx3_ASAP7_75t_L g9714 ( 
.A(n_9056),
.Y(n_9714)
);

AND2x2_ASAP7_75t_L g9715 ( 
.A(n_9353),
.B(n_55),
.Y(n_9715)
);

NAND2xp5_ASAP7_75t_L g9716 ( 
.A(n_9198),
.B(n_56),
.Y(n_9716)
);

INVx2_ASAP7_75t_L g9717 ( 
.A(n_9194),
.Y(n_9717)
);

INVx1_ASAP7_75t_L g9718 ( 
.A(n_9228),
.Y(n_9718)
);

INVx4_ASAP7_75t_L g9719 ( 
.A(n_9364),
.Y(n_9719)
);

NAND2xp5_ASAP7_75t_L g9720 ( 
.A(n_9199),
.B(n_56),
.Y(n_9720)
);

OAI21xp5_ASAP7_75t_L g9721 ( 
.A1(n_9095),
.A2(n_57),
.B(n_58),
.Y(n_9721)
);

AND2x4_ASAP7_75t_L g9722 ( 
.A(n_9317),
.B(n_57),
.Y(n_9722)
);

OAI21xp5_ASAP7_75t_L g9723 ( 
.A1(n_9303),
.A2(n_58),
.B(n_59),
.Y(n_9723)
);

NAND2xp5_ASAP7_75t_L g9724 ( 
.A(n_9205),
.B(n_9206),
.Y(n_9724)
);

INVx2_ASAP7_75t_L g9725 ( 
.A(n_9280),
.Y(n_9725)
);

INVx1_ASAP7_75t_L g9726 ( 
.A(n_9229),
.Y(n_9726)
);

HB1xp67_ASAP7_75t_L g9727 ( 
.A(n_9394),
.Y(n_9727)
);

AND2x2_ASAP7_75t_L g9728 ( 
.A(n_9146),
.B(n_59),
.Y(n_9728)
);

AND2x4_ASAP7_75t_L g9729 ( 
.A(n_9406),
.B(n_9403),
.Y(n_9729)
);

INVx1_ASAP7_75t_SL g9730 ( 
.A(n_9395),
.Y(n_9730)
);

NAND2xp5_ASAP7_75t_SL g9731 ( 
.A(n_8945),
.B(n_60),
.Y(n_9731)
);

INVx1_ASAP7_75t_L g9732 ( 
.A(n_9232),
.Y(n_9732)
);

INVx2_ASAP7_75t_L g9733 ( 
.A(n_9286),
.Y(n_9733)
);

INVxp67_ASAP7_75t_SL g9734 ( 
.A(n_9142),
.Y(n_9734)
);

BUFx3_ASAP7_75t_L g9735 ( 
.A(n_9414),
.Y(n_9735)
);

INVx1_ASAP7_75t_L g9736 ( 
.A(n_9241),
.Y(n_9736)
);

INVx1_ASAP7_75t_L g9737 ( 
.A(n_9244),
.Y(n_9737)
);

NOR2xp33_ASAP7_75t_L g9738 ( 
.A(n_9158),
.B(n_60),
.Y(n_9738)
);

BUFx3_ASAP7_75t_L g9739 ( 
.A(n_9426),
.Y(n_9739)
);

INVx3_ASAP7_75t_L g9740 ( 
.A(n_9369),
.Y(n_9740)
);

INVxp67_ASAP7_75t_L g9741 ( 
.A(n_9282),
.Y(n_9741)
);

NAND2xp5_ASAP7_75t_L g9742 ( 
.A(n_9202),
.B(n_61),
.Y(n_9742)
);

AND2x4_ASAP7_75t_L g9743 ( 
.A(n_9259),
.B(n_62),
.Y(n_9743)
);

INVx1_ASAP7_75t_L g9744 ( 
.A(n_9267),
.Y(n_9744)
);

AND2x4_ASAP7_75t_L g9745 ( 
.A(n_9293),
.B(n_62),
.Y(n_9745)
);

INVx2_ASAP7_75t_L g9746 ( 
.A(n_9288),
.Y(n_9746)
);

BUFx6f_ASAP7_75t_L g9747 ( 
.A(n_9182),
.Y(n_9747)
);

AND2x2_ASAP7_75t_SL g9748 ( 
.A(n_9220),
.B(n_63),
.Y(n_9748)
);

INVx2_ASAP7_75t_L g9749 ( 
.A(n_9310),
.Y(n_9749)
);

INVx2_ASAP7_75t_SL g9750 ( 
.A(n_9066),
.Y(n_9750)
);

AND2x2_ASAP7_75t_L g9751 ( 
.A(n_9314),
.B(n_63),
.Y(n_9751)
);

INVx2_ASAP7_75t_L g9752 ( 
.A(n_9130),
.Y(n_9752)
);

INVx2_ASAP7_75t_L g9753 ( 
.A(n_9141),
.Y(n_9753)
);

INVx2_ASAP7_75t_L g9754 ( 
.A(n_9151),
.Y(n_9754)
);

NAND2xp5_ASAP7_75t_L g9755 ( 
.A(n_9072),
.B(n_64),
.Y(n_9755)
);

INVx2_ASAP7_75t_L g9756 ( 
.A(n_9322),
.Y(n_9756)
);

NAND2xp5_ASAP7_75t_L g9757 ( 
.A(n_9116),
.B(n_64),
.Y(n_9757)
);

AND2x2_ASAP7_75t_SL g9758 ( 
.A(n_9060),
.B(n_65),
.Y(n_9758)
);

NAND2xp5_ASAP7_75t_L g9759 ( 
.A(n_9132),
.B(n_65),
.Y(n_9759)
);

INVx2_ASAP7_75t_L g9760 ( 
.A(n_9326),
.Y(n_9760)
);

INVx2_ASAP7_75t_L g9761 ( 
.A(n_9329),
.Y(n_9761)
);

AND2x2_ASAP7_75t_L g9762 ( 
.A(n_9108),
.B(n_9121),
.Y(n_9762)
);

AND2x2_ASAP7_75t_L g9763 ( 
.A(n_9143),
.B(n_66),
.Y(n_9763)
);

INVx2_ASAP7_75t_L g9764 ( 
.A(n_9175),
.Y(n_9764)
);

INVx2_ASAP7_75t_L g9765 ( 
.A(n_9298),
.Y(n_9765)
);

AND2x2_ASAP7_75t_L g9766 ( 
.A(n_9237),
.B(n_67),
.Y(n_9766)
);

AND2x2_ASAP7_75t_L g9767 ( 
.A(n_9257),
.B(n_9187),
.Y(n_9767)
);

CKINVDCx5p33_ASAP7_75t_R g9768 ( 
.A(n_9065),
.Y(n_9768)
);

AND2x2_ASAP7_75t_L g9769 ( 
.A(n_9159),
.B(n_67),
.Y(n_9769)
);

AND2x2_ASAP7_75t_L g9770 ( 
.A(n_9159),
.B(n_68),
.Y(n_9770)
);

INVx2_ASAP7_75t_L g9771 ( 
.A(n_9316),
.Y(n_9771)
);

INVx2_ASAP7_75t_L g9772 ( 
.A(n_9343),
.Y(n_9772)
);

NAND2xp5_ASAP7_75t_L g9773 ( 
.A(n_9341),
.B(n_68),
.Y(n_9773)
);

INVx2_ASAP7_75t_L g9774 ( 
.A(n_9350),
.Y(n_9774)
);

AND2x2_ASAP7_75t_L g9775 ( 
.A(n_9311),
.B(n_69),
.Y(n_9775)
);

BUFx6f_ASAP7_75t_L g9776 ( 
.A(n_9049),
.Y(n_9776)
);

INVx1_ASAP7_75t_L g9777 ( 
.A(n_9028),
.Y(n_9777)
);

AND2x2_ASAP7_75t_L g9778 ( 
.A(n_9311),
.B(n_69),
.Y(n_9778)
);

AND2x2_ASAP7_75t_L g9779 ( 
.A(n_9374),
.B(n_70),
.Y(n_9779)
);

INVx1_ASAP7_75t_L g9780 ( 
.A(n_9223),
.Y(n_9780)
);

NAND2xp5_ASAP7_75t_L g9781 ( 
.A(n_9203),
.B(n_70),
.Y(n_9781)
);

NAND2xp5_ASAP7_75t_L g9782 ( 
.A(n_9222),
.B(n_71),
.Y(n_9782)
);

OAI21xp5_ASAP7_75t_L g9783 ( 
.A1(n_9171),
.A2(n_71),
.B(n_72),
.Y(n_9783)
);

HB1xp67_ASAP7_75t_L g9784 ( 
.A(n_9351),
.Y(n_9784)
);

NAND2xp5_ASAP7_75t_SL g9785 ( 
.A(n_9415),
.B(n_72),
.Y(n_9785)
);

AND2x2_ASAP7_75t_L g9786 ( 
.A(n_9145),
.B(n_73),
.Y(n_9786)
);

AND2x4_ASAP7_75t_L g9787 ( 
.A(n_9413),
.B(n_73),
.Y(n_9787)
);

INVx2_ASAP7_75t_L g9788 ( 
.A(n_9129),
.Y(n_9788)
);

INVx2_ASAP7_75t_L g9789 ( 
.A(n_9150),
.Y(n_9789)
);

NOR2xp33_ASAP7_75t_L g9790 ( 
.A(n_9190),
.B(n_9006),
.Y(n_9790)
);

INVx1_ASAP7_75t_L g9791 ( 
.A(n_9225),
.Y(n_9791)
);

INVx3_ASAP7_75t_L g9792 ( 
.A(n_9398),
.Y(n_9792)
);

AND2x2_ASAP7_75t_L g9793 ( 
.A(n_9260),
.B(n_74),
.Y(n_9793)
);

INVx3_ASAP7_75t_L g9794 ( 
.A(n_9210),
.Y(n_9794)
);

INVx2_ASAP7_75t_SL g9795 ( 
.A(n_9421),
.Y(n_9795)
);

AND2x4_ASAP7_75t_L g9796 ( 
.A(n_9169),
.B(n_9364),
.Y(n_9796)
);

INVx1_ASAP7_75t_L g9797 ( 
.A(n_9235),
.Y(n_9797)
);

AND2x2_ASAP7_75t_SL g9798 ( 
.A(n_9144),
.B(n_75),
.Y(n_9798)
);

AND2x2_ASAP7_75t_L g9799 ( 
.A(n_9057),
.B(n_75),
.Y(n_9799)
);

NAND2xp5_ASAP7_75t_L g9800 ( 
.A(n_9354),
.B(n_76),
.Y(n_9800)
);

NAND2xp5_ASAP7_75t_L g9801 ( 
.A(n_9371),
.B(n_76),
.Y(n_9801)
);

AND2x2_ASAP7_75t_L g9802 ( 
.A(n_9410),
.B(n_9424),
.Y(n_9802)
);

INVx3_ASAP7_75t_L g9803 ( 
.A(n_9097),
.Y(n_9803)
);

NOR2xp33_ASAP7_75t_L g9804 ( 
.A(n_9023),
.B(n_77),
.Y(n_9804)
);

NAND2xp5_ASAP7_75t_L g9805 ( 
.A(n_9375),
.B(n_78),
.Y(n_9805)
);

AND2x4_ASAP7_75t_L g9806 ( 
.A(n_8953),
.B(n_78),
.Y(n_9806)
);

INVx2_ASAP7_75t_L g9807 ( 
.A(n_9154),
.Y(n_9807)
);

AND2x2_ASAP7_75t_L g9808 ( 
.A(n_9339),
.B(n_79),
.Y(n_9808)
);

NAND2xp5_ASAP7_75t_SL g9809 ( 
.A(n_8941),
.B(n_79),
.Y(n_9809)
);

AND2x2_ASAP7_75t_L g9810 ( 
.A(n_9340),
.B(n_80),
.Y(n_9810)
);

BUFx5_ASAP7_75t_L g9811 ( 
.A(n_9390),
.Y(n_9811)
);

INVx2_ASAP7_75t_L g9812 ( 
.A(n_9160),
.Y(n_9812)
);

INVx1_ASAP7_75t_SL g9813 ( 
.A(n_9377),
.Y(n_9813)
);

AND2x2_ASAP7_75t_L g9814 ( 
.A(n_9359),
.B(n_9361),
.Y(n_9814)
);

NAND2xp5_ASAP7_75t_L g9815 ( 
.A(n_9365),
.B(n_80),
.Y(n_9815)
);

AND2x2_ASAP7_75t_L g9816 ( 
.A(n_9284),
.B(n_81),
.Y(n_9816)
);

AND2x2_ASAP7_75t_L g9817 ( 
.A(n_9289),
.B(n_81),
.Y(n_9817)
);

OR2x6_ASAP7_75t_L g9818 ( 
.A(n_9389),
.B(n_82),
.Y(n_9818)
);

INVx1_ASAP7_75t_L g9819 ( 
.A(n_9236),
.Y(n_9819)
);

AND2x2_ASAP7_75t_L g9820 ( 
.A(n_9296),
.B(n_82),
.Y(n_9820)
);

INVx4_ASAP7_75t_L g9821 ( 
.A(n_9390),
.Y(n_9821)
);

INVx1_ASAP7_75t_L g9822 ( 
.A(n_9250),
.Y(n_9822)
);

INVx1_ASAP7_75t_L g9823 ( 
.A(n_9253),
.Y(n_9823)
);

INVxp67_ASAP7_75t_L g9824 ( 
.A(n_9378),
.Y(n_9824)
);

INVx2_ASAP7_75t_L g9825 ( 
.A(n_9167),
.Y(n_9825)
);

AND2x2_ASAP7_75t_L g9826 ( 
.A(n_9300),
.B(n_83),
.Y(n_9826)
);

INVx1_ASAP7_75t_L g9827 ( 
.A(n_9255),
.Y(n_9827)
);

AND2x2_ASAP7_75t_L g9828 ( 
.A(n_9301),
.B(n_9320),
.Y(n_9828)
);

INVx2_ASAP7_75t_SL g9829 ( 
.A(n_9433),
.Y(n_9829)
);

NOR2xp67_ASAP7_75t_L g9830 ( 
.A(n_9164),
.B(n_83),
.Y(n_9830)
);

AND2x2_ASAP7_75t_L g9831 ( 
.A(n_9325),
.B(n_84),
.Y(n_9831)
);

OAI21xp5_ASAP7_75t_L g9832 ( 
.A1(n_9402),
.A2(n_84),
.B(n_85),
.Y(n_9832)
);

AND2x2_ASAP7_75t_L g9833 ( 
.A(n_9328),
.B(n_85),
.Y(n_9833)
);

BUFx5_ASAP7_75t_L g9834 ( 
.A(n_9390),
.Y(n_9834)
);

AND2x2_ASAP7_75t_L g9835 ( 
.A(n_9330),
.B(n_86),
.Y(n_9835)
);

INVx1_ASAP7_75t_L g9836 ( 
.A(n_9258),
.Y(n_9836)
);

AND2x4_ASAP7_75t_L g9837 ( 
.A(n_9256),
.B(n_86),
.Y(n_9837)
);

INVx4_ASAP7_75t_L g9838 ( 
.A(n_9389),
.Y(n_9838)
);

NAND2xp5_ASAP7_75t_L g9839 ( 
.A(n_9043),
.B(n_87),
.Y(n_9839)
);

AND2x2_ASAP7_75t_L g9840 ( 
.A(n_9261),
.B(n_88),
.Y(n_9840)
);

AND2x2_ASAP7_75t_L g9841 ( 
.A(n_9271),
.B(n_88),
.Y(n_9841)
);

INVx2_ASAP7_75t_L g9842 ( 
.A(n_9168),
.Y(n_9842)
);

INVx2_ASAP7_75t_L g9843 ( 
.A(n_9170),
.Y(n_9843)
);

NAND2xp5_ASAP7_75t_L g9844 ( 
.A(n_8974),
.B(n_9034),
.Y(n_9844)
);

INVxp67_ASAP7_75t_SL g9845 ( 
.A(n_9173),
.Y(n_9845)
);

NAND2xp5_ASAP7_75t_L g9846 ( 
.A(n_9112),
.B(n_89),
.Y(n_9846)
);

NAND2xp5_ASAP7_75t_SL g9847 ( 
.A(n_9234),
.B(n_89),
.Y(n_9847)
);

AND2x2_ASAP7_75t_L g9848 ( 
.A(n_9272),
.B(n_90),
.Y(n_9848)
);

INVx1_ASAP7_75t_L g9849 ( 
.A(n_9177),
.Y(n_9849)
);

INVx1_ASAP7_75t_L g9850 ( 
.A(n_9179),
.Y(n_9850)
);

INVx1_ASAP7_75t_L g9851 ( 
.A(n_9045),
.Y(n_9851)
);

INVx1_ASAP7_75t_L g9852 ( 
.A(n_9062),
.Y(n_9852)
);

AND2x2_ASAP7_75t_L g9853 ( 
.A(n_9273),
.B(n_90),
.Y(n_9853)
);

INVx2_ASAP7_75t_L g9854 ( 
.A(n_9064),
.Y(n_9854)
);

INVx1_ASAP7_75t_L g9855 ( 
.A(n_9068),
.Y(n_9855)
);

INVx1_ASAP7_75t_L g9856 ( 
.A(n_9069),
.Y(n_9856)
);

NAND2xp5_ASAP7_75t_L g9857 ( 
.A(n_9113),
.B(n_91),
.Y(n_9857)
);

NAND2xp5_ASAP7_75t_L g9858 ( 
.A(n_9118),
.B(n_92),
.Y(n_9858)
);

AND2x2_ASAP7_75t_L g9859 ( 
.A(n_9274),
.B(n_92),
.Y(n_9859)
);

NAND2xp5_ASAP7_75t_L g9860 ( 
.A(n_9120),
.B(n_93),
.Y(n_9860)
);

AND2x2_ASAP7_75t_L g9861 ( 
.A(n_9334),
.B(n_93),
.Y(n_9861)
);

NAND2xp5_ASAP7_75t_SL g9862 ( 
.A(n_9221),
.B(n_94),
.Y(n_9862)
);

NAND2xp5_ASAP7_75t_L g9863 ( 
.A(n_9077),
.B(n_9079),
.Y(n_9863)
);

BUFx3_ASAP7_75t_L g9864 ( 
.A(n_9024),
.Y(n_9864)
);

NAND2xp5_ASAP7_75t_L g9865 ( 
.A(n_9093),
.B(n_94),
.Y(n_9865)
);

AND2x4_ASAP7_75t_L g9866 ( 
.A(n_9263),
.B(n_9295),
.Y(n_9866)
);

NAND2xp5_ASAP7_75t_L g9867 ( 
.A(n_9098),
.B(n_95),
.Y(n_9867)
);

INVx2_ASAP7_75t_L g9868 ( 
.A(n_9110),
.Y(n_9868)
);

INVx1_ASAP7_75t_L g9869 ( 
.A(n_9183),
.Y(n_9869)
);

NAND2xp5_ASAP7_75t_L g9870 ( 
.A(n_9186),
.B(n_95),
.Y(n_9870)
);

INVxp67_ASAP7_75t_SL g9871 ( 
.A(n_9189),
.Y(n_9871)
);

NAND2x1p5_ASAP7_75t_L g9872 ( 
.A(n_9055),
.B(n_96),
.Y(n_9872)
);

HB1xp67_ASAP7_75t_L g9873 ( 
.A(n_9099),
.Y(n_9873)
);

INVx2_ASAP7_75t_L g9874 ( 
.A(n_9270),
.Y(n_9874)
);

NAND2xp5_ASAP7_75t_SL g9875 ( 
.A(n_9419),
.B(n_96),
.Y(n_9875)
);

NAND2xp5_ASAP7_75t_L g9876 ( 
.A(n_9163),
.B(n_8984),
.Y(n_9876)
);

AND2x2_ASAP7_75t_L g9877 ( 
.A(n_9000),
.B(n_8981),
.Y(n_9877)
);

NAND2xp5_ASAP7_75t_L g9878 ( 
.A(n_9372),
.B(n_97),
.Y(n_9878)
);

NOR2xp33_ASAP7_75t_SL g9879 ( 
.A(n_9427),
.B(n_97),
.Y(n_9879)
);

INVx1_ASAP7_75t_L g9880 ( 
.A(n_9075),
.Y(n_9880)
);

INVx1_ASAP7_75t_L g9881 ( 
.A(n_9243),
.Y(n_9881)
);

BUFx5_ASAP7_75t_L g9882 ( 
.A(n_9385),
.Y(n_9882)
);

INVx1_ASAP7_75t_L g9883 ( 
.A(n_9124),
.Y(n_9883)
);

AND2x2_ASAP7_75t_L g9884 ( 
.A(n_9384),
.B(n_98),
.Y(n_9884)
);

INVx2_ASAP7_75t_L g9885 ( 
.A(n_9363),
.Y(n_9885)
);

NOR2xp67_ASAP7_75t_L g9886 ( 
.A(n_9201),
.B(n_98),
.Y(n_9886)
);

NOR2xp33_ASAP7_75t_L g9887 ( 
.A(n_9407),
.B(n_99),
.Y(n_9887)
);

AND2x2_ASAP7_75t_L g9888 ( 
.A(n_9392),
.B(n_99),
.Y(n_9888)
);

AND2x2_ASAP7_75t_L g9889 ( 
.A(n_9397),
.B(n_100),
.Y(n_9889)
);

HB1xp67_ASAP7_75t_L g9890 ( 
.A(n_9248),
.Y(n_9890)
);

INVx1_ASAP7_75t_L g9891 ( 
.A(n_8993),
.Y(n_9891)
);

NAND2xp5_ASAP7_75t_L g9892 ( 
.A(n_8999),
.B(n_100),
.Y(n_9892)
);

INVx1_ASAP7_75t_L g9893 ( 
.A(n_9172),
.Y(n_9893)
);

AND2x2_ASAP7_75t_L g9894 ( 
.A(n_9400),
.B(n_101),
.Y(n_9894)
);

HB1xp67_ASAP7_75t_L g9895 ( 
.A(n_9299),
.Y(n_9895)
);

INVx1_ASAP7_75t_L g9896 ( 
.A(n_8985),
.Y(n_9896)
);

OAI21xp5_ASAP7_75t_L g9897 ( 
.A1(n_8967),
.A2(n_101),
.B(n_102),
.Y(n_9897)
);

AND2x2_ASAP7_75t_L g9898 ( 
.A(n_9331),
.B(n_102),
.Y(n_9898)
);

INVx4_ASAP7_75t_L g9899 ( 
.A(n_9021),
.Y(n_9899)
);

BUFx3_ASAP7_75t_L g9900 ( 
.A(n_9436),
.Y(n_9900)
);

HB1xp67_ASAP7_75t_L g9901 ( 
.A(n_9136),
.Y(n_9901)
);

INVx2_ASAP7_75t_L g9902 ( 
.A(n_9387),
.Y(n_9902)
);

OAI21xp5_ASAP7_75t_L g9903 ( 
.A1(n_9212),
.A2(n_103),
.B(n_104),
.Y(n_9903)
);

NAND2xp5_ASAP7_75t_L g9904 ( 
.A(n_9399),
.B(n_105),
.Y(n_9904)
);

NOR2xp33_ASAP7_75t_L g9905 ( 
.A(n_9409),
.B(n_106),
.Y(n_9905)
);

INVx8_ASAP7_75t_L g9906 ( 
.A(n_9021),
.Y(n_9906)
);

INVxp67_ASAP7_75t_SL g9907 ( 
.A(n_9109),
.Y(n_9907)
);

AND2x2_ASAP7_75t_L g9908 ( 
.A(n_9411),
.B(n_106),
.Y(n_9908)
);

NAND2xp5_ASAP7_75t_L g9909 ( 
.A(n_9231),
.B(n_107),
.Y(n_9909)
);

INVx2_ASAP7_75t_L g9910 ( 
.A(n_9429),
.Y(n_9910)
);

INVx2_ASAP7_75t_L g9911 ( 
.A(n_9092),
.Y(n_9911)
);

BUFx6f_ASAP7_75t_L g9912 ( 
.A(n_9101),
.Y(n_9912)
);

NAND2xp5_ASAP7_75t_SL g9913 ( 
.A(n_9422),
.B(n_107),
.Y(n_9913)
);

AND2x2_ASAP7_75t_L g9914 ( 
.A(n_9425),
.B(n_108),
.Y(n_9914)
);

INVx2_ASAP7_75t_L g9915 ( 
.A(n_9148),
.Y(n_9915)
);

NAND2xp5_ASAP7_75t_L g9916 ( 
.A(n_9302),
.B(n_108),
.Y(n_9916)
);

INVx1_ASAP7_75t_L g9917 ( 
.A(n_9176),
.Y(n_9917)
);

INVx1_ASAP7_75t_SL g9918 ( 
.A(n_9405),
.Y(n_9918)
);

NAND2xp5_ASAP7_75t_SL g9919 ( 
.A(n_9391),
.B(n_109),
.Y(n_9919)
);

INVx2_ASAP7_75t_L g9920 ( 
.A(n_9149),
.Y(n_9920)
);

AND2x6_ASAP7_75t_L g9921 ( 
.A(n_9412),
.B(n_110),
.Y(n_9921)
);

INVx2_ASAP7_75t_L g9922 ( 
.A(n_9313),
.Y(n_9922)
);

AND2x2_ASAP7_75t_SL g9923 ( 
.A(n_9294),
.B(n_110),
.Y(n_9923)
);

INVx1_ASAP7_75t_L g9924 ( 
.A(n_9362),
.Y(n_9924)
);

NOR2xp33_ASAP7_75t_SL g9925 ( 
.A(n_9417),
.B(n_111),
.Y(n_9925)
);

INVx1_ASAP7_75t_L g9926 ( 
.A(n_9347),
.Y(n_9926)
);

INVx1_ASAP7_75t_L g9927 ( 
.A(n_9356),
.Y(n_9927)
);

AND2x2_ASAP7_75t_L g9928 ( 
.A(n_9155),
.B(n_111),
.Y(n_9928)
);

INVx1_ASAP7_75t_L g9929 ( 
.A(n_9321),
.Y(n_9929)
);

INVx2_ASAP7_75t_L g9930 ( 
.A(n_9114),
.Y(n_9930)
);

NOR2xp33_ASAP7_75t_R g9931 ( 
.A(n_9336),
.B(n_112),
.Y(n_9931)
);

NAND2xp5_ASAP7_75t_L g9932 ( 
.A(n_9074),
.B(n_112),
.Y(n_9932)
);

NAND2xp5_ASAP7_75t_L g9933 ( 
.A(n_9082),
.B(n_113),
.Y(n_9933)
);

NOR2xp33_ASAP7_75t_L g9934 ( 
.A(n_9063),
.B(n_113),
.Y(n_9934)
);

INVx1_ASAP7_75t_L g9935 ( 
.A(n_9122),
.Y(n_9935)
);

HB1xp67_ASAP7_75t_L g9936 ( 
.A(n_9086),
.Y(n_9936)
);

BUFx8_ASAP7_75t_SL g9937 ( 
.A(n_9156),
.Y(n_9937)
);

AND2x2_ASAP7_75t_L g9938 ( 
.A(n_9147),
.B(n_114),
.Y(n_9938)
);

NAND2xp5_ASAP7_75t_L g9939 ( 
.A(n_9297),
.B(n_114),
.Y(n_9939)
);

INVx1_ASAP7_75t_L g9940 ( 
.A(n_9126),
.Y(n_9940)
);

INVx3_ASAP7_75t_L g9941 ( 
.A(n_9432),
.Y(n_9941)
);

INVx2_ASAP7_75t_L g9942 ( 
.A(n_9107),
.Y(n_9942)
);

AND2x2_ASAP7_75t_L g9943 ( 
.A(n_8965),
.B(n_115),
.Y(n_9943)
);

AND2x2_ASAP7_75t_SL g9944 ( 
.A(n_9367),
.B(n_115),
.Y(n_9944)
);

INVx2_ASAP7_75t_L g9945 ( 
.A(n_9319),
.Y(n_9945)
);

AND2x2_ASAP7_75t_L g9946 ( 
.A(n_9342),
.B(n_116),
.Y(n_9946)
);

INVx3_ASAP7_75t_L g9947 ( 
.A(n_8986),
.Y(n_9947)
);

INVx3_ASAP7_75t_L g9948 ( 
.A(n_9204),
.Y(n_9948)
);

AND2x2_ASAP7_75t_L g9949 ( 
.A(n_9344),
.B(n_117),
.Y(n_9949)
);

NOR2xp33_ASAP7_75t_L g9950 ( 
.A(n_9373),
.B(n_117),
.Y(n_9950)
);

NOR2xp33_ASAP7_75t_L g9951 ( 
.A(n_9430),
.B(n_118),
.Y(n_9951)
);

INVx2_ASAP7_75t_L g9952 ( 
.A(n_9254),
.Y(n_9952)
);

INVx1_ASAP7_75t_L g9953 ( 
.A(n_9227),
.Y(n_9953)
);

AND2x2_ASAP7_75t_L g9954 ( 
.A(n_9428),
.B(n_118),
.Y(n_9954)
);

NAND2xp5_ASAP7_75t_L g9955 ( 
.A(n_9246),
.B(n_119),
.Y(n_9955)
);

INVx1_ASAP7_75t_SL g9956 ( 
.A(n_9031),
.Y(n_9956)
);

AND2x2_ASAP7_75t_L g9957 ( 
.A(n_9306),
.B(n_119),
.Y(n_9957)
);

INVx2_ASAP7_75t_L g9958 ( 
.A(n_9036),
.Y(n_9958)
);

BUFx6f_ASAP7_75t_L g9959 ( 
.A(n_9071),
.Y(n_9959)
);

INVx4_ASAP7_75t_L g9960 ( 
.A(n_9434),
.Y(n_9960)
);

NOR2xp33_ASAP7_75t_L g9961 ( 
.A(n_9435),
.B(n_120),
.Y(n_9961)
);

HB1xp67_ASAP7_75t_L g9962 ( 
.A(n_9044),
.Y(n_9962)
);

INVx3_ASAP7_75t_L g9963 ( 
.A(n_8998),
.Y(n_9963)
);

AND2x2_ASAP7_75t_L g9964 ( 
.A(n_9051),
.B(n_120),
.Y(n_9964)
);

AND2x2_ASAP7_75t_L g9965 ( 
.A(n_9051),
.B(n_121),
.Y(n_9965)
);

NOR2xp33_ASAP7_75t_L g9966 ( 
.A(n_8929),
.B(n_121),
.Y(n_9966)
);

AND2x2_ASAP7_75t_L g9967 ( 
.A(n_9051),
.B(n_122),
.Y(n_9967)
);

INVx2_ASAP7_75t_L g9968 ( 
.A(n_8932),
.Y(n_9968)
);

CKINVDCx5p33_ASAP7_75t_R g9969 ( 
.A(n_8990),
.Y(n_9969)
);

INVx1_ASAP7_75t_L g9970 ( 
.A(n_9111),
.Y(n_9970)
);

BUFx3_ASAP7_75t_L g9971 ( 
.A(n_9022),
.Y(n_9971)
);

AND2x2_ASAP7_75t_L g9972 ( 
.A(n_9051),
.B(n_122),
.Y(n_9972)
);

INVx2_ASAP7_75t_L g9973 ( 
.A(n_8932),
.Y(n_9973)
);

OAI21xp5_ASAP7_75t_L g9974 ( 
.A1(n_8960),
.A2(n_123),
.B(n_124),
.Y(n_9974)
);

AND2x4_ASAP7_75t_L g9975 ( 
.A(n_8979),
.B(n_123),
.Y(n_9975)
);

CKINVDCx20_ASAP7_75t_R g9976 ( 
.A(n_8962),
.Y(n_9976)
);

AOI22xp5_ASAP7_75t_L g9977 ( 
.A1(n_8960),
.A2(n_126),
.B1(n_124),
.B2(n_125),
.Y(n_9977)
);

INVx2_ASAP7_75t_L g9978 ( 
.A(n_8932),
.Y(n_9978)
);

NAND2xp5_ASAP7_75t_L g9979 ( 
.A(n_9012),
.B(n_126),
.Y(n_9979)
);

INVx1_ASAP7_75t_SL g9980 ( 
.A(n_9213),
.Y(n_9980)
);

INVx3_ASAP7_75t_L g9981 ( 
.A(n_8998),
.Y(n_9981)
);

NAND2xp5_ASAP7_75t_L g9982 ( 
.A(n_9012),
.B(n_127),
.Y(n_9982)
);

BUFx3_ASAP7_75t_L g9983 ( 
.A(n_9022),
.Y(n_9983)
);

AND2x2_ASAP7_75t_L g9984 ( 
.A(n_9051),
.B(n_127),
.Y(n_9984)
);

INVx2_ASAP7_75t_L g9985 ( 
.A(n_8932),
.Y(n_9985)
);

AND2x2_ASAP7_75t_L g9986 ( 
.A(n_9051),
.B(n_128),
.Y(n_9986)
);

NAND2xp5_ASAP7_75t_L g9987 ( 
.A(n_9012),
.B(n_129),
.Y(n_9987)
);

AND2x2_ASAP7_75t_L g9988 ( 
.A(n_9051),
.B(n_130),
.Y(n_9988)
);

AND2x2_ASAP7_75t_L g9989 ( 
.A(n_9051),
.B(n_130),
.Y(n_9989)
);

NAND2xp5_ASAP7_75t_L g9990 ( 
.A(n_9012),
.B(n_131),
.Y(n_9990)
);

BUFx2_ASAP7_75t_L g9991 ( 
.A(n_8973),
.Y(n_9991)
);

AND2x2_ASAP7_75t_SL g9992 ( 
.A(n_9315),
.B(n_131),
.Y(n_9992)
);

INVxp67_ASAP7_75t_L g9993 ( 
.A(n_8928),
.Y(n_9993)
);

INVx2_ASAP7_75t_L g9994 ( 
.A(n_8932),
.Y(n_9994)
);

INVx2_ASAP7_75t_L g9995 ( 
.A(n_8932),
.Y(n_9995)
);

INVx1_ASAP7_75t_L g9996 ( 
.A(n_9111),
.Y(n_9996)
);

HB1xp67_ASAP7_75t_L g9997 ( 
.A(n_8973),
.Y(n_9997)
);

OAI21x1_ASAP7_75t_L g9998 ( 
.A1(n_8971),
.A2(n_132),
.B(n_133),
.Y(n_9998)
);

INVx1_ASAP7_75t_L g9999 ( 
.A(n_9111),
.Y(n_9999)
);

NAND2xp5_ASAP7_75t_L g10000 ( 
.A(n_9012),
.B(n_132),
.Y(n_10000)
);

INVx1_ASAP7_75t_L g10001 ( 
.A(n_9111),
.Y(n_10001)
);

AND2x2_ASAP7_75t_L g10002 ( 
.A(n_9051),
.B(n_133),
.Y(n_10002)
);

NAND2xp5_ASAP7_75t_L g10003 ( 
.A(n_9012),
.B(n_134),
.Y(n_10003)
);

NAND2xp5_ASAP7_75t_L g10004 ( 
.A(n_9012),
.B(n_134),
.Y(n_10004)
);

AND2x2_ASAP7_75t_L g10005 ( 
.A(n_9051),
.B(n_135),
.Y(n_10005)
);

AND2x2_ASAP7_75t_SL g10006 ( 
.A(n_9315),
.B(n_135),
.Y(n_10006)
);

AND2x2_ASAP7_75t_L g10007 ( 
.A(n_9051),
.B(n_136),
.Y(n_10007)
);

NAND2xp5_ASAP7_75t_L g10008 ( 
.A(n_9012),
.B(n_136),
.Y(n_10008)
);

INVx2_ASAP7_75t_L g10009 ( 
.A(n_8932),
.Y(n_10009)
);

AND2x2_ASAP7_75t_L g10010 ( 
.A(n_9051),
.B(n_137),
.Y(n_10010)
);

OR2x2_ASAP7_75t_SL g10011 ( 
.A(n_9431),
.B(n_137),
.Y(n_10011)
);

NAND2xp5_ASAP7_75t_L g10012 ( 
.A(n_9012),
.B(n_138),
.Y(n_10012)
);

AND2x2_ASAP7_75t_L g10013 ( 
.A(n_9051),
.B(n_138),
.Y(n_10013)
);

AND2x2_ASAP7_75t_L g10014 ( 
.A(n_9051),
.B(n_139),
.Y(n_10014)
);

HB1xp67_ASAP7_75t_L g10015 ( 
.A(n_8973),
.Y(n_10015)
);

HB1xp67_ASAP7_75t_L g10016 ( 
.A(n_8973),
.Y(n_10016)
);

INVx3_ASAP7_75t_L g10017 ( 
.A(n_8998),
.Y(n_10017)
);

OAI21xp5_ASAP7_75t_L g10018 ( 
.A1(n_8960),
.A2(n_139),
.B(n_140),
.Y(n_10018)
);

AND2x2_ASAP7_75t_L g10019 ( 
.A(n_9051),
.B(n_140),
.Y(n_10019)
);

AND2x2_ASAP7_75t_L g10020 ( 
.A(n_9051),
.B(n_141),
.Y(n_10020)
);

NAND2xp5_ASAP7_75t_L g10021 ( 
.A(n_9012),
.B(n_141),
.Y(n_10021)
);

NAND2xp5_ASAP7_75t_L g10022 ( 
.A(n_9012),
.B(n_142),
.Y(n_10022)
);

INVx1_ASAP7_75t_L g10023 ( 
.A(n_9111),
.Y(n_10023)
);

OAI21xp5_ASAP7_75t_L g10024 ( 
.A1(n_8960),
.A2(n_142),
.B(n_143),
.Y(n_10024)
);

INVx3_ASAP7_75t_L g10025 ( 
.A(n_8998),
.Y(n_10025)
);

INVx1_ASAP7_75t_L g10026 ( 
.A(n_9111),
.Y(n_10026)
);

INVx1_ASAP7_75t_L g10027 ( 
.A(n_9111),
.Y(n_10027)
);

BUFx6f_ASAP7_75t_L g10028 ( 
.A(n_9022),
.Y(n_10028)
);

INVx3_ASAP7_75t_L g10029 ( 
.A(n_8998),
.Y(n_10029)
);

BUFx3_ASAP7_75t_L g10030 ( 
.A(n_9022),
.Y(n_10030)
);

NAND2xp5_ASAP7_75t_L g10031 ( 
.A(n_9012),
.B(n_144),
.Y(n_10031)
);

INVx2_ASAP7_75t_L g10032 ( 
.A(n_8932),
.Y(n_10032)
);

NAND2xp5_ASAP7_75t_L g10033 ( 
.A(n_9012),
.B(n_144),
.Y(n_10033)
);

NOR2xp33_ASAP7_75t_L g10034 ( 
.A(n_8929),
.B(n_145),
.Y(n_10034)
);

AND2x2_ASAP7_75t_SL g10035 ( 
.A(n_9315),
.B(n_145),
.Y(n_10035)
);

BUFx3_ASAP7_75t_L g10036 ( 
.A(n_9022),
.Y(n_10036)
);

INVx2_ASAP7_75t_L g10037 ( 
.A(n_8932),
.Y(n_10037)
);

AND2x4_ASAP7_75t_L g10038 ( 
.A(n_8979),
.B(n_146),
.Y(n_10038)
);

NAND2xp5_ASAP7_75t_SL g10039 ( 
.A(n_8960),
.B(n_146),
.Y(n_10039)
);

INVx1_ASAP7_75t_L g10040 ( 
.A(n_9111),
.Y(n_10040)
);

AND2x2_ASAP7_75t_L g10041 ( 
.A(n_9051),
.B(n_147),
.Y(n_10041)
);

BUFx6f_ASAP7_75t_L g10042 ( 
.A(n_9022),
.Y(n_10042)
);

AND2x2_ASAP7_75t_L g10043 ( 
.A(n_9051),
.B(n_147),
.Y(n_10043)
);

INVx1_ASAP7_75t_L g10044 ( 
.A(n_9111),
.Y(n_10044)
);

INVx1_ASAP7_75t_L g10045 ( 
.A(n_9111),
.Y(n_10045)
);

AOI21xp5_ASAP7_75t_L g10046 ( 
.A1(n_9731),
.A2(n_148),
.B(n_149),
.Y(n_10046)
);

AOI21xp5_ASAP7_75t_L g10047 ( 
.A1(n_9704),
.A2(n_9624),
.B(n_9783),
.Y(n_10047)
);

AO21x1_ASAP7_75t_L g10048 ( 
.A1(n_9602),
.A2(n_148),
.B(n_149),
.Y(n_10048)
);

NAND2xp5_ASAP7_75t_L g10049 ( 
.A(n_9557),
.B(n_150),
.Y(n_10049)
);

INVx3_ASAP7_75t_L g10050 ( 
.A(n_9470),
.Y(n_10050)
);

NAND2xp5_ASAP7_75t_L g10051 ( 
.A(n_9618),
.B(n_150),
.Y(n_10051)
);

OAI22xp5_ASAP7_75t_L g10052 ( 
.A1(n_9678),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_10052)
);

INVx1_ASAP7_75t_L g10053 ( 
.A(n_9563),
.Y(n_10053)
);

AOI21xp5_ASAP7_75t_L g10054 ( 
.A1(n_9469),
.A2(n_9845),
.B(n_9871),
.Y(n_10054)
);

INVx11_ASAP7_75t_L g10055 ( 
.A(n_9504),
.Y(n_10055)
);

NAND2xp5_ASAP7_75t_SL g10056 ( 
.A(n_9596),
.B(n_151),
.Y(n_10056)
);

NAND2xp5_ASAP7_75t_L g10057 ( 
.A(n_9814),
.B(n_152),
.Y(n_10057)
);

NOR2xp67_ASAP7_75t_SL g10058 ( 
.A(n_9821),
.B(n_153),
.Y(n_10058)
);

A2O1A1Ixp33_ASAP7_75t_L g10059 ( 
.A1(n_9897),
.A2(n_156),
.B(n_154),
.C(n_155),
.Y(n_10059)
);

INVx1_ASAP7_75t_L g10060 ( 
.A(n_9570),
.Y(n_10060)
);

NOR2xp33_ASAP7_75t_L g10061 ( 
.A(n_9701),
.B(n_154),
.Y(n_10061)
);

NAND2xp5_ASAP7_75t_L g10062 ( 
.A(n_9463),
.B(n_155),
.Y(n_10062)
);

INVx1_ASAP7_75t_L g10063 ( 
.A(n_9574),
.Y(n_10063)
);

NAND2xp5_ASAP7_75t_L g10064 ( 
.A(n_9970),
.B(n_156),
.Y(n_10064)
);

OAI22xp5_ASAP7_75t_L g10065 ( 
.A1(n_9565),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.Y(n_10065)
);

NOR2xp33_ASAP7_75t_L g10066 ( 
.A(n_9683),
.B(n_159),
.Y(n_10066)
);

OAI21x1_ASAP7_75t_L g10067 ( 
.A1(n_9454),
.A2(n_160),
.B(n_161),
.Y(n_10067)
);

A2O1A1Ixp33_ASAP7_75t_L g10068 ( 
.A1(n_9552),
.A2(n_162),
.B(n_160),
.C(n_161),
.Y(n_10068)
);

NAND2xp5_ASAP7_75t_SL g10069 ( 
.A(n_9554),
.B(n_162),
.Y(n_10069)
);

OAI21xp33_ASAP7_75t_L g10070 ( 
.A1(n_9974),
.A2(n_163),
.B(n_164),
.Y(n_10070)
);

NAND2xp5_ASAP7_75t_L g10071 ( 
.A(n_9996),
.B(n_165),
.Y(n_10071)
);

NOR2xp33_ASAP7_75t_L g10072 ( 
.A(n_9741),
.B(n_166),
.Y(n_10072)
);

INVx2_ASAP7_75t_L g10073 ( 
.A(n_9444),
.Y(n_10073)
);

AND2x2_ASAP7_75t_L g10074 ( 
.A(n_9452),
.B(n_166),
.Y(n_10074)
);

INVx1_ASAP7_75t_L g10075 ( 
.A(n_9579),
.Y(n_10075)
);

INVx1_ASAP7_75t_L g10076 ( 
.A(n_9591),
.Y(n_10076)
);

AOI21xp5_ASAP7_75t_L g10077 ( 
.A1(n_9863),
.A2(n_167),
.B(n_168),
.Y(n_10077)
);

OAI21xp5_ASAP7_75t_L g10078 ( 
.A1(n_9505),
.A2(n_167),
.B(n_168),
.Y(n_10078)
);

INVx1_ASAP7_75t_L g10079 ( 
.A(n_9608),
.Y(n_10079)
);

NOR2xp33_ASAP7_75t_L g10080 ( 
.A(n_9900),
.B(n_169),
.Y(n_10080)
);

O2A1O1Ixp5_ASAP7_75t_L g10081 ( 
.A1(n_9661),
.A2(n_173),
.B(n_170),
.C(n_171),
.Y(n_10081)
);

AOI21xp5_ASAP7_75t_L g10082 ( 
.A1(n_9724),
.A2(n_9734),
.B(n_9876),
.Y(n_10082)
);

O2A1O1Ixp33_ASAP7_75t_L g10083 ( 
.A1(n_9757),
.A2(n_173),
.B(n_170),
.C(n_171),
.Y(n_10083)
);

HB1xp67_ASAP7_75t_L g10084 ( 
.A(n_9993),
.Y(n_10084)
);

AOI21xp5_ASAP7_75t_L g10085 ( 
.A1(n_9891),
.A2(n_174),
.B(n_175),
.Y(n_10085)
);

AOI21x1_ASAP7_75t_L g10086 ( 
.A1(n_9919),
.A2(n_174),
.B(n_175),
.Y(n_10086)
);

NOR2xp33_ASAP7_75t_SL g10087 ( 
.A(n_9524),
.B(n_176),
.Y(n_10087)
);

AOI21xp5_ASAP7_75t_L g10088 ( 
.A1(n_9844),
.A2(n_176),
.B(n_177),
.Y(n_10088)
);

NOR2xp33_ASAP7_75t_L g10089 ( 
.A(n_9501),
.B(n_9802),
.Y(n_10089)
);

AOI21xp5_ASAP7_75t_L g10090 ( 
.A1(n_10018),
.A2(n_177),
.B(n_178),
.Y(n_10090)
);

NAND3xp33_ASAP7_75t_L g10091 ( 
.A(n_9832),
.B(n_10024),
.C(n_9738),
.Y(n_10091)
);

AO21x1_ASAP7_75t_L g10092 ( 
.A1(n_9723),
.A2(n_178),
.B(n_179),
.Y(n_10092)
);

BUFx2_ASAP7_75t_SL g10093 ( 
.A(n_9632),
.Y(n_10093)
);

OAI21xp5_ASAP7_75t_L g10094 ( 
.A1(n_9450),
.A2(n_179),
.B(n_180),
.Y(n_10094)
);

AOI21xp5_ASAP7_75t_L g10095 ( 
.A1(n_9520),
.A2(n_181),
.B(n_182),
.Y(n_10095)
);

NOR2xp33_ASAP7_75t_L g10096 ( 
.A(n_9445),
.B(n_181),
.Y(n_10096)
);

BUFx6f_ASAP7_75t_L g10097 ( 
.A(n_9632),
.Y(n_10097)
);

OAI21x1_ASAP7_75t_L g10098 ( 
.A1(n_9666),
.A2(n_182),
.B(n_183),
.Y(n_10098)
);

AOI22xp5_ASAP7_75t_L g10099 ( 
.A1(n_9496),
.A2(n_185),
.B1(n_183),
.B2(n_184),
.Y(n_10099)
);

AOI22xp5_ASAP7_75t_L g10100 ( 
.A1(n_9642),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.Y(n_10100)
);

NOR2xp33_ASAP7_75t_L g10101 ( 
.A(n_9980),
.B(n_186),
.Y(n_10101)
);

INVx2_ASAP7_75t_L g10102 ( 
.A(n_9449),
.Y(n_10102)
);

AOI21xp5_ASAP7_75t_L g10103 ( 
.A1(n_9529),
.A2(n_9528),
.B(n_9999),
.Y(n_10103)
);

NOR2xp33_ASAP7_75t_L g10104 ( 
.A(n_9813),
.B(n_187),
.Y(n_10104)
);

OAI321xp33_ASAP7_75t_L g10105 ( 
.A1(n_9688),
.A2(n_189),
.A3(n_191),
.B1(n_187),
.B2(n_188),
.C(n_190),
.Y(n_10105)
);

INVx2_ASAP7_75t_L g10106 ( 
.A(n_9457),
.Y(n_10106)
);

NAND2xp5_ASAP7_75t_L g10107 ( 
.A(n_10001),
.B(n_188),
.Y(n_10107)
);

NOR3xp33_ASAP7_75t_L g10108 ( 
.A(n_9862),
.B(n_190),
.C(n_191),
.Y(n_10108)
);

INVx2_ASAP7_75t_SL g10109 ( 
.A(n_9561),
.Y(n_10109)
);

O2A1O1Ixp5_ASAP7_75t_L g10110 ( 
.A1(n_9721),
.A2(n_194),
.B(n_192),
.C(n_193),
.Y(n_10110)
);

AO21x1_ASAP7_75t_L g10111 ( 
.A1(n_9903),
.A2(n_192),
.B(n_194),
.Y(n_10111)
);

AOI21x1_ASAP7_75t_L g10112 ( 
.A1(n_9910),
.A2(n_196),
.B(n_197),
.Y(n_10112)
);

OAI22xp5_ASAP7_75t_L g10113 ( 
.A1(n_9755),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.Y(n_10113)
);

BUFx8_ASAP7_75t_SL g10114 ( 
.A(n_9976),
.Y(n_10114)
);

INVx4_ASAP7_75t_L g10115 ( 
.A(n_9633),
.Y(n_10115)
);

AOI21xp5_ASAP7_75t_L g10116 ( 
.A1(n_10023),
.A2(n_198),
.B(n_199),
.Y(n_10116)
);

OAI22xp5_ASAP7_75t_L g10117 ( 
.A1(n_9759),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_10117)
);

OAI21xp5_ASAP7_75t_L g10118 ( 
.A1(n_9512),
.A2(n_200),
.B(n_201),
.Y(n_10118)
);

BUFx4f_ASAP7_75t_L g10119 ( 
.A(n_9633),
.Y(n_10119)
);

AOI21x1_ASAP7_75t_L g10120 ( 
.A1(n_9874),
.A2(n_202),
.B(n_204),
.Y(n_10120)
);

AOI21xp5_ASAP7_75t_L g10121 ( 
.A1(n_10026),
.A2(n_202),
.B(n_205),
.Y(n_10121)
);

AOI22xp5_ASAP7_75t_L g10122 ( 
.A1(n_10039),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_10122)
);

O2A1O1Ixp33_ASAP7_75t_L g10123 ( 
.A1(n_9781),
.A2(n_209),
.B(n_207),
.C(n_208),
.Y(n_10123)
);

AOI21xp5_ASAP7_75t_L g10124 ( 
.A1(n_10027),
.A2(n_10044),
.B(n_10040),
.Y(n_10124)
);

NAND2xp5_ASAP7_75t_SL g10125 ( 
.A(n_9854),
.B(n_208),
.Y(n_10125)
);

NOR3xp33_ASAP7_75t_L g10126 ( 
.A(n_9782),
.B(n_209),
.C(n_210),
.Y(n_10126)
);

NAND2xp5_ASAP7_75t_L g10127 ( 
.A(n_10045),
.B(n_210),
.Y(n_10127)
);

NOR2xp33_ASAP7_75t_L g10128 ( 
.A(n_9460),
.B(n_211),
.Y(n_10128)
);

NAND2xp5_ASAP7_75t_L g10129 ( 
.A(n_9780),
.B(n_211),
.Y(n_10129)
);

INVx1_ASAP7_75t_L g10130 ( 
.A(n_9616),
.Y(n_10130)
);

OAI21xp5_ASAP7_75t_L g10131 ( 
.A1(n_9527),
.A2(n_212),
.B(n_213),
.Y(n_10131)
);

INVx3_ASAP7_75t_L g10132 ( 
.A(n_9635),
.Y(n_10132)
);

INVx4_ASAP7_75t_L g10133 ( 
.A(n_9635),
.Y(n_10133)
);

OAI22xp5_ASAP7_75t_L g10134 ( 
.A1(n_9962),
.A2(n_215),
.B1(n_212),
.B2(n_213),
.Y(n_10134)
);

AO22x1_ASAP7_75t_L g10135 ( 
.A1(n_9921),
.A2(n_217),
.B1(n_215),
.B2(n_216),
.Y(n_10135)
);

OAI22xp5_ASAP7_75t_L g10136 ( 
.A1(n_9773),
.A2(n_220),
.B1(n_218),
.B2(n_219),
.Y(n_10136)
);

BUFx4f_ASAP7_75t_L g10137 ( 
.A(n_9747),
.Y(n_10137)
);

INVx2_ASAP7_75t_L g10138 ( 
.A(n_9459),
.Y(n_10138)
);

INVx2_ASAP7_75t_SL g10139 ( 
.A(n_9561),
.Y(n_10139)
);

INVx2_ASAP7_75t_L g10140 ( 
.A(n_9464),
.Y(n_10140)
);

O2A1O1Ixp33_ASAP7_75t_L g10141 ( 
.A1(n_9576),
.A2(n_222),
.B(n_218),
.C(n_221),
.Y(n_10141)
);

OAI21xp5_ASAP7_75t_L g10142 ( 
.A1(n_9564),
.A2(n_9896),
.B(n_9583),
.Y(n_10142)
);

NAND2xp5_ASAP7_75t_L g10143 ( 
.A(n_9791),
.B(n_221),
.Y(n_10143)
);

NAND2xp5_ASAP7_75t_SL g10144 ( 
.A(n_9868),
.B(n_223),
.Y(n_10144)
);

AND2x2_ASAP7_75t_L g10145 ( 
.A(n_9767),
.B(n_223),
.Y(n_10145)
);

INVx1_ASAP7_75t_L g10146 ( 
.A(n_9622),
.Y(n_10146)
);

NAND2xp5_ASAP7_75t_L g10147 ( 
.A(n_9797),
.B(n_224),
.Y(n_10147)
);

NAND2xp5_ASAP7_75t_L g10148 ( 
.A(n_9819),
.B(n_9822),
.Y(n_10148)
);

OAI22xp5_ASAP7_75t_L g10149 ( 
.A1(n_9692),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.Y(n_10149)
);

CKINVDCx8_ASAP7_75t_R g10150 ( 
.A(n_9534),
.Y(n_10150)
);

INVx2_ASAP7_75t_L g10151 ( 
.A(n_9468),
.Y(n_10151)
);

AOI21xp5_ASAP7_75t_L g10152 ( 
.A1(n_9929),
.A2(n_225),
.B(n_226),
.Y(n_10152)
);

INVx1_ASAP7_75t_L g10153 ( 
.A(n_9629),
.Y(n_10153)
);

INVx2_ASAP7_75t_L g10154 ( 
.A(n_9473),
.Y(n_10154)
);

BUFx6f_ASAP7_75t_L g10155 ( 
.A(n_9575),
.Y(n_10155)
);

NAND2xp5_ASAP7_75t_L g10156 ( 
.A(n_9823),
.B(n_227),
.Y(n_10156)
);

OAI21xp5_ASAP7_75t_L g10157 ( 
.A1(n_9509),
.A2(n_228),
.B(n_229),
.Y(n_10157)
);

INVx1_ASAP7_75t_L g10158 ( 
.A(n_9630),
.Y(n_10158)
);

AOI21xp5_ASAP7_75t_L g10159 ( 
.A1(n_9503),
.A2(n_228),
.B(n_229),
.Y(n_10159)
);

AOI21xp5_ASAP7_75t_L g10160 ( 
.A1(n_9788),
.A2(n_230),
.B(n_231),
.Y(n_10160)
);

NAND3xp33_ASAP7_75t_SL g10161 ( 
.A(n_9931),
.B(n_230),
.C(n_231),
.Y(n_10161)
);

NAND2xp5_ASAP7_75t_L g10162 ( 
.A(n_9827),
.B(n_232),
.Y(n_10162)
);

INVx2_ASAP7_75t_L g10163 ( 
.A(n_9475),
.Y(n_10163)
);

INVx2_ASAP7_75t_L g10164 ( 
.A(n_9477),
.Y(n_10164)
);

OAI21xp33_ASAP7_75t_L g10165 ( 
.A1(n_9615),
.A2(n_232),
.B(n_233),
.Y(n_10165)
);

OAI21xp5_ASAP7_75t_L g10166 ( 
.A1(n_9443),
.A2(n_233),
.B(n_234),
.Y(n_10166)
);

NAND2xp5_ASAP7_75t_L g10167 ( 
.A(n_9836),
.B(n_234),
.Y(n_10167)
);

NOR2xp33_ASAP7_75t_L g10168 ( 
.A(n_9487),
.B(n_235),
.Y(n_10168)
);

INVxp33_ASAP7_75t_SL g10169 ( 
.A(n_9609),
.Y(n_10169)
);

OAI21xp5_ASAP7_75t_L g10170 ( 
.A1(n_9479),
.A2(n_235),
.B(n_236),
.Y(n_10170)
);

BUFx6f_ASAP7_75t_L g10171 ( 
.A(n_9575),
.Y(n_10171)
);

NAND2xp33_ASAP7_75t_L g10172 ( 
.A(n_9811),
.B(n_9834),
.Y(n_10172)
);

AOI21xp5_ASAP7_75t_L g10173 ( 
.A1(n_9789),
.A2(n_236),
.B(n_237),
.Y(n_10173)
);

AOI21xp5_ASAP7_75t_L g10174 ( 
.A1(n_9807),
.A2(n_238),
.B(n_239),
.Y(n_10174)
);

BUFx3_ASAP7_75t_L g10175 ( 
.A(n_9578),
.Y(n_10175)
);

OAI22xp5_ASAP7_75t_L g10176 ( 
.A1(n_9604),
.A2(n_241),
.B1(n_238),
.B2(n_240),
.Y(n_10176)
);

NOR2xp33_ASAP7_75t_L g10177 ( 
.A(n_9824),
.B(n_240),
.Y(n_10177)
);

AND2x2_ASAP7_75t_L g10178 ( 
.A(n_9964),
.B(n_242),
.Y(n_10178)
);

AOI21x1_ASAP7_75t_L g10179 ( 
.A1(n_9668),
.A2(n_242),
.B(n_243),
.Y(n_10179)
);

AOI21x1_ASAP7_75t_L g10180 ( 
.A1(n_9893),
.A2(n_243),
.B(n_244),
.Y(n_10180)
);

NAND2xp5_ASAP7_75t_SL g10181 ( 
.A(n_9851),
.B(n_245),
.Y(n_10181)
);

INVx1_ASAP7_75t_L g10182 ( 
.A(n_9647),
.Y(n_10182)
);

NAND2xp5_ASAP7_75t_L g10183 ( 
.A(n_9852),
.B(n_246),
.Y(n_10183)
);

INVx1_ASAP7_75t_L g10184 ( 
.A(n_9656),
.Y(n_10184)
);

NAND2xp5_ASAP7_75t_L g10185 ( 
.A(n_9855),
.B(n_246),
.Y(n_10185)
);

BUFx6f_ASAP7_75t_L g10186 ( 
.A(n_9584),
.Y(n_10186)
);

A2O1A1Ixp33_ASAP7_75t_L g10187 ( 
.A1(n_9877),
.A2(n_249),
.B(n_247),
.C(n_248),
.Y(n_10187)
);

NAND2xp5_ASAP7_75t_L g10188 ( 
.A(n_9856),
.B(n_247),
.Y(n_10188)
);

AOI21xp5_ASAP7_75t_L g10189 ( 
.A1(n_9812),
.A2(n_248),
.B(n_250),
.Y(n_10189)
);

A2O1A1Ixp33_ASAP7_75t_L g10190 ( 
.A1(n_9804),
.A2(n_252),
.B(n_250),
.C(n_251),
.Y(n_10190)
);

NAND2xp5_ASAP7_75t_L g10191 ( 
.A(n_9869),
.B(n_252),
.Y(n_10191)
);

NAND2xp5_ASAP7_75t_L g10192 ( 
.A(n_9849),
.B(n_253),
.Y(n_10192)
);

NAND2xp5_ASAP7_75t_L g10193 ( 
.A(n_9850),
.B(n_253),
.Y(n_10193)
);

AOI21xp5_ASAP7_75t_L g10194 ( 
.A1(n_9825),
.A2(n_254),
.B(n_255),
.Y(n_10194)
);

NAND2xp5_ASAP7_75t_L g10195 ( 
.A(n_9842),
.B(n_254),
.Y(n_10195)
);

OAI22xp5_ASAP7_75t_L g10196 ( 
.A1(n_9593),
.A2(n_258),
.B1(n_256),
.B2(n_257),
.Y(n_10196)
);

AOI21xp5_ASAP7_75t_L g10197 ( 
.A1(n_9843),
.A2(n_257),
.B(n_258),
.Y(n_10197)
);

A2O1A1Ixp33_ASAP7_75t_L g10198 ( 
.A1(n_9887),
.A2(n_261),
.B(n_259),
.C(n_260),
.Y(n_10198)
);

NAND3xp33_ASAP7_75t_SL g10199 ( 
.A(n_9879),
.B(n_259),
.C(n_260),
.Y(n_10199)
);

AOI21xp5_ASAP7_75t_L g10200 ( 
.A1(n_9474),
.A2(n_261),
.B(n_262),
.Y(n_10200)
);

O2A1O1Ixp5_ASAP7_75t_L g10201 ( 
.A1(n_9640),
.A2(n_264),
.B(n_262),
.C(n_263),
.Y(n_10201)
);

NAND2xp5_ASAP7_75t_L g10202 ( 
.A(n_9478),
.B(n_263),
.Y(n_10202)
);

AO21x1_ASAP7_75t_L g10203 ( 
.A1(n_9698),
.A2(n_264),
.B(n_265),
.Y(n_10203)
);

AOI21xp5_ASAP7_75t_L g10204 ( 
.A1(n_9828),
.A2(n_9902),
.B(n_9765),
.Y(n_10204)
);

NAND2xp5_ASAP7_75t_L g10205 ( 
.A(n_9764),
.B(n_266),
.Y(n_10205)
);

AOI21xp5_ASAP7_75t_L g10206 ( 
.A1(n_9771),
.A2(n_267),
.B(n_268),
.Y(n_10206)
);

INVx3_ASAP7_75t_L g10207 ( 
.A(n_9739),
.Y(n_10207)
);

AOI33xp33_ASAP7_75t_L g10208 ( 
.A1(n_9769),
.A2(n_269),
.A3(n_271),
.B1(n_267),
.B2(n_268),
.B3(n_270),
.Y(n_10208)
);

NOR2xp33_ASAP7_75t_L g10209 ( 
.A(n_9556),
.B(n_269),
.Y(n_10209)
);

AND2x6_ASAP7_75t_SL g10210 ( 
.A(n_9966),
.B(n_270),
.Y(n_10210)
);

NAND2xp5_ASAP7_75t_L g10211 ( 
.A(n_9979),
.B(n_271),
.Y(n_10211)
);

INVx1_ASAP7_75t_L g10212 ( 
.A(n_9660),
.Y(n_10212)
);

HB1xp67_ASAP7_75t_L g10213 ( 
.A(n_9494),
.Y(n_10213)
);

O2A1O1Ixp33_ASAP7_75t_L g10214 ( 
.A1(n_9847),
.A2(n_274),
.B(n_272),
.C(n_273),
.Y(n_10214)
);

AOI21xp5_ASAP7_75t_L g10215 ( 
.A1(n_9952),
.A2(n_272),
.B(n_274),
.Y(n_10215)
);

INVx1_ASAP7_75t_L g10216 ( 
.A(n_9662),
.Y(n_10216)
);

OAI21x1_ASAP7_75t_L g10217 ( 
.A1(n_9998),
.A2(n_275),
.B(n_276),
.Y(n_10217)
);

NOR2xp33_ASAP7_75t_L g10218 ( 
.A(n_9991),
.B(n_275),
.Y(n_10218)
);

OAI21xp33_ASAP7_75t_L g10219 ( 
.A1(n_9839),
.A2(n_276),
.B(n_277),
.Y(n_10219)
);

AO32x1_ASAP7_75t_L g10220 ( 
.A1(n_9777),
.A2(n_279),
.A3(n_277),
.B1(n_278),
.B2(n_280),
.Y(n_10220)
);

A2O1A1Ixp33_ASAP7_75t_L g10221 ( 
.A1(n_9905),
.A2(n_281),
.B(n_278),
.C(n_279),
.Y(n_10221)
);

INVx4_ASAP7_75t_L g10222 ( 
.A(n_9584),
.Y(n_10222)
);

AOI21x1_ASAP7_75t_L g10223 ( 
.A1(n_9880),
.A2(n_281),
.B(n_282),
.Y(n_10223)
);

NAND2xp5_ASAP7_75t_SL g10224 ( 
.A(n_9790),
.B(n_282),
.Y(n_10224)
);

NOR2xp67_ASAP7_75t_L g10225 ( 
.A(n_9663),
.B(n_283),
.Y(n_10225)
);

INVx3_ASAP7_75t_L g10226 ( 
.A(n_9471),
.Y(n_10226)
);

BUFx6f_ASAP7_75t_L g10227 ( 
.A(n_9589),
.Y(n_10227)
);

OAI321xp33_ASAP7_75t_L g10228 ( 
.A1(n_9977),
.A2(n_286),
.A3(n_288),
.B1(n_283),
.B2(n_284),
.C(n_287),
.Y(n_10228)
);

INVx1_ASAP7_75t_L g10229 ( 
.A(n_9664),
.Y(n_10229)
);

INVx2_ASAP7_75t_L g10230 ( 
.A(n_9483),
.Y(n_10230)
);

INVx2_ASAP7_75t_L g10231 ( 
.A(n_9499),
.Y(n_10231)
);

BUFx8_ASAP7_75t_L g10232 ( 
.A(n_9747),
.Y(n_10232)
);

NAND2xp5_ASAP7_75t_L g10233 ( 
.A(n_9982),
.B(n_284),
.Y(n_10233)
);

AOI21xp5_ASAP7_75t_L g10234 ( 
.A1(n_9885),
.A2(n_286),
.B(n_287),
.Y(n_10234)
);

NAND2xp5_ASAP7_75t_L g10235 ( 
.A(n_9987),
.B(n_288),
.Y(n_10235)
);

AOI21xp5_ASAP7_75t_L g10236 ( 
.A1(n_9990),
.A2(n_289),
.B(n_290),
.Y(n_10236)
);

AOI22xp33_ASAP7_75t_L g10237 ( 
.A1(n_9748),
.A2(n_291),
.B1(n_289),
.B2(n_290),
.Y(n_10237)
);

INVx2_ASAP7_75t_L g10238 ( 
.A(n_9508),
.Y(n_10238)
);

AOI21xp5_ASAP7_75t_L g10239 ( 
.A1(n_10000),
.A2(n_291),
.B(n_292),
.Y(n_10239)
);

NAND2xp5_ASAP7_75t_L g10240 ( 
.A(n_10003),
.B(n_292),
.Y(n_10240)
);

NAND2xp5_ASAP7_75t_L g10241 ( 
.A(n_10004),
.B(n_293),
.Y(n_10241)
);

NOR2xp33_ASAP7_75t_L g10242 ( 
.A(n_9918),
.B(n_293),
.Y(n_10242)
);

NOR2xp33_ASAP7_75t_L g10243 ( 
.A(n_9549),
.B(n_295),
.Y(n_10243)
);

NAND2xp5_ASAP7_75t_L g10244 ( 
.A(n_10008),
.B(n_295),
.Y(n_10244)
);

NOR2x1_ASAP7_75t_L g10245 ( 
.A(n_9719),
.B(n_296),
.Y(n_10245)
);

INVx2_ASAP7_75t_L g10246 ( 
.A(n_9510),
.Y(n_10246)
);

BUFx6f_ASAP7_75t_L g10247 ( 
.A(n_9589),
.Y(n_10247)
);

A2O1A1Ixp33_ASAP7_75t_L g10248 ( 
.A1(n_9800),
.A2(n_298),
.B(n_296),
.C(n_297),
.Y(n_10248)
);

NAND2xp5_ASAP7_75t_SL g10249 ( 
.A(n_9811),
.B(n_297),
.Y(n_10249)
);

AOI22xp33_ASAP7_75t_L g10250 ( 
.A1(n_9710),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.Y(n_10250)
);

AOI21xp5_ASAP7_75t_L g10251 ( 
.A1(n_10012),
.A2(n_299),
.B(n_300),
.Y(n_10251)
);

OAI21xp5_ASAP7_75t_L g10252 ( 
.A1(n_9492),
.A2(n_301),
.B(n_302),
.Y(n_10252)
);

AOI21xp5_ASAP7_75t_L g10253 ( 
.A1(n_10021),
.A2(n_303),
.B(n_304),
.Y(n_10253)
);

OAI21xp5_ASAP7_75t_L g10254 ( 
.A1(n_9455),
.A2(n_304),
.B(n_305),
.Y(n_10254)
);

NAND2xp5_ASAP7_75t_L g10255 ( 
.A(n_10022),
.B(n_306),
.Y(n_10255)
);

NAND2xp5_ASAP7_75t_L g10256 ( 
.A(n_10031),
.B(n_306),
.Y(n_10256)
);

AOI21xp5_ASAP7_75t_L g10257 ( 
.A1(n_10033),
.A2(n_307),
.B(n_308),
.Y(n_10257)
);

INVx1_ASAP7_75t_L g10258 ( 
.A(n_9672),
.Y(n_10258)
);

AOI21xp5_ASAP7_75t_L g10259 ( 
.A1(n_9881),
.A2(n_307),
.B(n_308),
.Y(n_10259)
);

OAI22xp5_ASAP7_75t_L g10260 ( 
.A1(n_9543),
.A2(n_311),
.B1(n_309),
.B2(n_310),
.Y(n_10260)
);

AOI21xp5_ASAP7_75t_L g10261 ( 
.A1(n_9883),
.A2(n_9917),
.B(n_9798),
.Y(n_10261)
);

OAI21xp5_ASAP7_75t_L g10262 ( 
.A1(n_9801),
.A2(n_309),
.B(n_310),
.Y(n_10262)
);

AOI21xp5_ASAP7_75t_L g10263 ( 
.A1(n_9758),
.A2(n_311),
.B(n_312),
.Y(n_10263)
);

INVx3_ASAP7_75t_L g10264 ( 
.A(n_9500),
.Y(n_10264)
);

INVx3_ASAP7_75t_L g10265 ( 
.A(n_9467),
.Y(n_10265)
);

AOI21xp5_ASAP7_75t_L g10266 ( 
.A1(n_9923),
.A2(n_312),
.B(n_313),
.Y(n_10266)
);

AOI21xp5_ASAP7_75t_L g10267 ( 
.A1(n_9907),
.A2(n_313),
.B(n_314),
.Y(n_10267)
);

O2A1O1Ixp33_ASAP7_75t_L g10268 ( 
.A1(n_9805),
.A2(n_317),
.B(n_315),
.C(n_316),
.Y(n_10268)
);

NAND2xp5_ASAP7_75t_L g10269 ( 
.A(n_9466),
.B(n_9997),
.Y(n_10269)
);

NOR2xp67_ASAP7_75t_L g10270 ( 
.A(n_9941),
.B(n_315),
.Y(n_10270)
);

AOI21xp5_ASAP7_75t_L g10271 ( 
.A1(n_9462),
.A2(n_316),
.B(n_317),
.Y(n_10271)
);

OAI22xp5_ASAP7_75t_L g10272 ( 
.A1(n_9485),
.A2(n_320),
.B1(n_318),
.B2(n_319),
.Y(n_10272)
);

O2A1O1Ixp33_ASAP7_75t_L g10273 ( 
.A1(n_9909),
.A2(n_320),
.B(n_318),
.C(n_319),
.Y(n_10273)
);

AOI21xp5_ASAP7_75t_L g10274 ( 
.A1(n_9472),
.A2(n_322),
.B(n_323),
.Y(n_10274)
);

OAI21xp5_ASAP7_75t_L g10275 ( 
.A1(n_9892),
.A2(n_322),
.B(n_324),
.Y(n_10275)
);

NOR2xp33_ASAP7_75t_L g10276 ( 
.A(n_10015),
.B(n_324),
.Y(n_10276)
);

OA21x2_ASAP7_75t_L g10277 ( 
.A1(n_9684),
.A2(n_325),
.B(n_326),
.Y(n_10277)
);

NAND2xp5_ASAP7_75t_SL g10278 ( 
.A(n_9811),
.B(n_326),
.Y(n_10278)
);

INVx1_ASAP7_75t_L g10279 ( 
.A(n_9693),
.Y(n_10279)
);

INVx1_ASAP7_75t_L g10280 ( 
.A(n_9694),
.Y(n_10280)
);

INVx2_ASAP7_75t_SL g10281 ( 
.A(n_9612),
.Y(n_10281)
);

INVx2_ASAP7_75t_L g10282 ( 
.A(n_9514),
.Y(n_10282)
);

O2A1O1Ixp5_ASAP7_75t_L g10283 ( 
.A1(n_9785),
.A2(n_329),
.B(n_327),
.C(n_328),
.Y(n_10283)
);

NAND2xp5_ASAP7_75t_L g10284 ( 
.A(n_10016),
.B(n_9491),
.Y(n_10284)
);

AOI21xp5_ASAP7_75t_L g10285 ( 
.A1(n_9815),
.A2(n_327),
.B(n_328),
.Y(n_10285)
);

AOI21xp5_ASAP7_75t_L g10286 ( 
.A1(n_9772),
.A2(n_329),
.B(n_330),
.Y(n_10286)
);

AND2x2_ASAP7_75t_SL g10287 ( 
.A(n_9992),
.B(n_330),
.Y(n_10287)
);

INVx1_ASAP7_75t_SL g10288 ( 
.A(n_9489),
.Y(n_10288)
);

INVx2_ASAP7_75t_L g10289 ( 
.A(n_9545),
.Y(n_10289)
);

NAND2xp5_ASAP7_75t_L g10290 ( 
.A(n_9658),
.B(n_331),
.Y(n_10290)
);

AND2x2_ASAP7_75t_L g10291 ( 
.A(n_9965),
.B(n_331),
.Y(n_10291)
);

NAND2xp33_ASAP7_75t_L g10292 ( 
.A(n_9834),
.B(n_332),
.Y(n_10292)
);

AOI21xp5_ASAP7_75t_L g10293 ( 
.A1(n_9599),
.A2(n_333),
.B(n_335),
.Y(n_10293)
);

A2O1A1Ixp33_ASAP7_75t_L g10294 ( 
.A1(n_9951),
.A2(n_336),
.B(n_333),
.C(n_335),
.Y(n_10294)
);

NAND2xp5_ASAP7_75t_L g10295 ( 
.A(n_9562),
.B(n_336),
.Y(n_10295)
);

AOI21xp5_ASAP7_75t_L g10296 ( 
.A1(n_9605),
.A2(n_337),
.B(n_338),
.Y(n_10296)
);

NAND2xp5_ASAP7_75t_L g10297 ( 
.A(n_9968),
.B(n_337),
.Y(n_10297)
);

NAND2xp5_ASAP7_75t_SL g10298 ( 
.A(n_9834),
.B(n_338),
.Y(n_10298)
);

AOI22xp5_ASAP7_75t_L g10299 ( 
.A1(n_10034),
.A2(n_341),
.B1(n_339),
.B2(n_340),
.Y(n_10299)
);

NOR2xp33_ASAP7_75t_L g10300 ( 
.A(n_9960),
.B(n_339),
.Y(n_10300)
);

INVx2_ASAP7_75t_SL g10301 ( 
.A(n_9612),
.Y(n_10301)
);

NAND2x1p5_ASAP7_75t_L g10302 ( 
.A(n_9507),
.B(n_340),
.Y(n_10302)
);

NAND2xp5_ASAP7_75t_SL g10303 ( 
.A(n_9750),
.B(n_341),
.Y(n_10303)
);

NAND2xp5_ASAP7_75t_L g10304 ( 
.A(n_9973),
.B(n_342),
.Y(n_10304)
);

NOR2xp33_ASAP7_75t_L g10305 ( 
.A(n_9956),
.B(n_342),
.Y(n_10305)
);

AND2x2_ASAP7_75t_L g10306 ( 
.A(n_9967),
.B(n_343),
.Y(n_10306)
);

AND2x2_ASAP7_75t_L g10307 ( 
.A(n_9972),
.B(n_344),
.Y(n_10307)
);

AOI21xp5_ASAP7_75t_L g10308 ( 
.A1(n_9978),
.A2(n_344),
.B(n_345),
.Y(n_10308)
);

A2O1A1Ixp33_ASAP7_75t_L g10309 ( 
.A1(n_9961),
.A2(n_347),
.B(n_345),
.C(n_346),
.Y(n_10309)
);

OAI21xp5_ASAP7_75t_L g10310 ( 
.A1(n_9742),
.A2(n_347),
.B(n_348),
.Y(n_10310)
);

AOI21x1_ASAP7_75t_L g10311 ( 
.A1(n_9873),
.A2(n_9530),
.B(n_9886),
.Y(n_10311)
);

AO32x2_ASAP7_75t_L g10312 ( 
.A1(n_9829),
.A2(n_351),
.A3(n_349),
.B1(n_350),
.B2(n_352),
.Y(n_10312)
);

OAI21xp5_ASAP7_75t_L g10313 ( 
.A1(n_9617),
.A2(n_350),
.B(n_351),
.Y(n_10313)
);

NOR2xp67_ASAP7_75t_L g10314 ( 
.A(n_9461),
.B(n_353),
.Y(n_10314)
);

O2A1O1Ixp33_ASAP7_75t_L g10315 ( 
.A1(n_9939),
.A2(n_355),
.B(n_353),
.C(n_354),
.Y(n_10315)
);

NAND2xp5_ASAP7_75t_SL g10316 ( 
.A(n_9882),
.B(n_9796),
.Y(n_10316)
);

OAI21xp5_ASAP7_75t_L g10317 ( 
.A1(n_9634),
.A2(n_355),
.B(n_356),
.Y(n_10317)
);

O2A1O1Ixp5_ASAP7_75t_L g10318 ( 
.A1(n_9809),
.A2(n_358),
.B(n_356),
.C(n_357),
.Y(n_10318)
);

AO22x1_ASAP7_75t_L g10319 ( 
.A1(n_9921),
.A2(n_360),
.B1(n_358),
.B2(n_359),
.Y(n_10319)
);

NOR2xp33_ASAP7_75t_R g10320 ( 
.A(n_9969),
.B(n_359),
.Y(n_10320)
);

NAND2xp5_ASAP7_75t_L g10321 ( 
.A(n_9985),
.B(n_360),
.Y(n_10321)
);

INVx1_ASAP7_75t_L g10322 ( 
.A(n_9699),
.Y(n_10322)
);

OAI22xp5_ASAP7_75t_L g10323 ( 
.A1(n_10006),
.A2(n_363),
.B1(n_361),
.B2(n_362),
.Y(n_10323)
);

INVxp67_ASAP7_75t_L g10324 ( 
.A(n_9551),
.Y(n_10324)
);

NAND2xp5_ASAP7_75t_L g10325 ( 
.A(n_9994),
.B(n_9995),
.Y(n_10325)
);

NOR2xp67_ASAP7_75t_SL g10326 ( 
.A(n_9670),
.B(n_361),
.Y(n_10326)
);

NAND2xp5_ASAP7_75t_SL g10327 ( 
.A(n_9882),
.B(n_362),
.Y(n_10327)
);

AO21x1_ASAP7_75t_L g10328 ( 
.A1(n_9950),
.A2(n_363),
.B(n_364),
.Y(n_10328)
);

NAND2xp5_ASAP7_75t_L g10329 ( 
.A(n_10009),
.B(n_364),
.Y(n_10329)
);

INVx1_ASAP7_75t_L g10330 ( 
.A(n_9700),
.Y(n_10330)
);

NOR2xp33_ASAP7_75t_L g10331 ( 
.A(n_9901),
.B(n_366),
.Y(n_10331)
);

AOI21xp5_ASAP7_75t_L g10332 ( 
.A1(n_10032),
.A2(n_366),
.B(n_367),
.Y(n_10332)
);

NAND2xp5_ASAP7_75t_L g10333 ( 
.A(n_10037),
.B(n_367),
.Y(n_10333)
);

HB1xp67_ASAP7_75t_L g10334 ( 
.A(n_9536),
.Y(n_10334)
);

AOI21xp5_ASAP7_75t_L g10335 ( 
.A1(n_9935),
.A2(n_368),
.B(n_369),
.Y(n_10335)
);

INVx2_ASAP7_75t_L g10336 ( 
.A(n_9680),
.Y(n_10336)
);

NAND2xp5_ASAP7_75t_L g10337 ( 
.A(n_9517),
.B(n_368),
.Y(n_10337)
);

A2O1A1Ixp33_ASAP7_75t_L g10338 ( 
.A1(n_9934),
.A2(n_371),
.B(n_369),
.C(n_370),
.Y(n_10338)
);

AOI21xp5_ASAP7_75t_L g10339 ( 
.A1(n_9940),
.A2(n_371),
.B(n_372),
.Y(n_10339)
);

AOI21xp5_ASAP7_75t_L g10340 ( 
.A1(n_9713),
.A2(n_373),
.B(n_374),
.Y(n_10340)
);

BUFx12f_ASAP7_75t_L g10341 ( 
.A(n_9654),
.Y(n_10341)
);

AOI21xp5_ASAP7_75t_L g10342 ( 
.A1(n_9717),
.A2(n_374),
.B(n_375),
.Y(n_10342)
);

AOI211xp5_ASAP7_75t_L g10343 ( 
.A1(n_9943),
.A2(n_377),
.B(n_375),
.C(n_376),
.Y(n_10343)
);

INVx2_ASAP7_75t_L g10344 ( 
.A(n_9687),
.Y(n_10344)
);

O2A1O1Ixp33_ASAP7_75t_L g10345 ( 
.A1(n_9875),
.A2(n_9913),
.B(n_9569),
.C(n_9916),
.Y(n_10345)
);

NOR2xp33_ASAP7_75t_L g10346 ( 
.A(n_9506),
.B(n_377),
.Y(n_10346)
);

AOI21xp5_ASAP7_75t_L g10347 ( 
.A1(n_9756),
.A2(n_378),
.B(n_379),
.Y(n_10347)
);

NOR2xp33_ASAP7_75t_L g10348 ( 
.A(n_9762),
.B(n_378),
.Y(n_10348)
);

AND2x4_ASAP7_75t_L g10349 ( 
.A(n_9685),
.B(n_380),
.Y(n_10349)
);

AOI21xp5_ASAP7_75t_L g10350 ( 
.A1(n_9760),
.A2(n_380),
.B(n_381),
.Y(n_10350)
);

NAND2xp5_ASAP7_75t_L g10351 ( 
.A(n_9482),
.B(n_381),
.Y(n_10351)
);

AOI21xp5_ASAP7_75t_L g10352 ( 
.A1(n_9761),
.A2(n_382),
.B(n_383),
.Y(n_10352)
);

AOI21x1_ASAP7_75t_L g10353 ( 
.A1(n_9726),
.A2(n_383),
.B(n_384),
.Y(n_10353)
);

OAI21xp5_ASAP7_75t_L g10354 ( 
.A1(n_9638),
.A2(n_384),
.B(n_385),
.Y(n_10354)
);

AND2x2_ASAP7_75t_L g10355 ( 
.A(n_9984),
.B(n_385),
.Y(n_10355)
);

AND2x2_ASAP7_75t_L g10356 ( 
.A(n_9986),
.B(n_386),
.Y(n_10356)
);

INVx1_ASAP7_75t_L g10357 ( 
.A(n_9709),
.Y(n_10357)
);

AOI21xp5_ASAP7_75t_L g10358 ( 
.A1(n_9878),
.A2(n_387),
.B(n_388),
.Y(n_10358)
);

AOI21xp5_ASAP7_75t_L g10359 ( 
.A1(n_9930),
.A2(n_387),
.B(n_388),
.Y(n_10359)
);

AO21x1_ASAP7_75t_L g10360 ( 
.A1(n_9598),
.A2(n_9665),
.B(n_9650),
.Y(n_10360)
);

AO21x1_ASAP7_75t_L g10361 ( 
.A1(n_9673),
.A2(n_389),
.B(n_390),
.Y(n_10361)
);

BUFx12f_ASAP7_75t_L g10362 ( 
.A(n_9619),
.Y(n_10362)
);

INVx1_ASAP7_75t_L g10363 ( 
.A(n_9718),
.Y(n_10363)
);

NOR2x1_ASAP7_75t_L g10364 ( 
.A(n_9838),
.B(n_389),
.Y(n_10364)
);

OAI21xp5_ASAP7_75t_L g10365 ( 
.A1(n_9465),
.A2(n_9682),
.B(n_9681),
.Y(n_10365)
);

NAND2xp5_ASAP7_75t_SL g10366 ( 
.A(n_9882),
.B(n_391),
.Y(n_10366)
);

AOI21xp5_ASAP7_75t_L g10367 ( 
.A1(n_9689),
.A2(n_391),
.B(n_392),
.Y(n_10367)
);

AOI21xp5_ASAP7_75t_L g10368 ( 
.A1(n_9691),
.A2(n_392),
.B(n_393),
.Y(n_10368)
);

NAND2xp5_ASAP7_75t_L g10369 ( 
.A(n_9490),
.B(n_393),
.Y(n_10369)
);

AOI21xp5_ASAP7_75t_L g10370 ( 
.A1(n_9695),
.A2(n_394),
.B(n_395),
.Y(n_10370)
);

AOI22xp33_ASAP7_75t_L g10371 ( 
.A1(n_9786),
.A2(n_397),
.B1(n_394),
.B2(n_396),
.Y(n_10371)
);

INVx1_ASAP7_75t_L g10372 ( 
.A(n_9732),
.Y(n_10372)
);

OAI21xp33_ASAP7_75t_L g10373 ( 
.A1(n_9690),
.A2(n_397),
.B(n_398),
.Y(n_10373)
);

OAI21x1_ASAP7_75t_L g10374 ( 
.A1(n_9736),
.A2(n_398),
.B(n_399),
.Y(n_10374)
);

AOI21xp5_ASAP7_75t_L g10375 ( 
.A1(n_9702),
.A2(n_400),
.B(n_401),
.Y(n_10375)
);

AOI21xp5_ASAP7_75t_L g10376 ( 
.A1(n_9703),
.A2(n_402),
.B(n_403),
.Y(n_10376)
);

AOI21xp5_ASAP7_75t_L g10377 ( 
.A1(n_9725),
.A2(n_402),
.B(n_403),
.Y(n_10377)
);

AND2x4_ASAP7_75t_L g10378 ( 
.A(n_9795),
.B(n_9740),
.Y(n_10378)
);

AND2x2_ASAP7_75t_L g10379 ( 
.A(n_9988),
.B(n_404),
.Y(n_10379)
);

NOR2xp33_ASAP7_75t_SL g10380 ( 
.A(n_9669),
.B(n_404),
.Y(n_10380)
);

NAND2xp5_ASAP7_75t_L g10381 ( 
.A(n_9497),
.B(n_405),
.Y(n_10381)
);

AOI33xp33_ASAP7_75t_L g10382 ( 
.A1(n_9770),
.A2(n_9572),
.A3(n_9547),
.B1(n_9898),
.B2(n_9938),
.B3(n_9592),
.Y(n_10382)
);

OAI22xp5_ASAP7_75t_L g10383 ( 
.A1(n_10035),
.A2(n_407),
.B1(n_405),
.B2(n_406),
.Y(n_10383)
);

A2O1A1Ixp33_ASAP7_75t_L g10384 ( 
.A1(n_9711),
.A2(n_409),
.B(n_407),
.C(n_408),
.Y(n_10384)
);

BUFx2_ASAP7_75t_L g10385 ( 
.A(n_9553),
.Y(n_10385)
);

OAI21xp5_ASAP7_75t_L g10386 ( 
.A1(n_9712),
.A2(n_408),
.B(n_410),
.Y(n_10386)
);

NAND2xp5_ASAP7_75t_L g10387 ( 
.A(n_9498),
.B(n_410),
.Y(n_10387)
);

BUFx8_ASAP7_75t_L g10388 ( 
.A(n_10028),
.Y(n_10388)
);

AOI21xp5_ASAP7_75t_L g10389 ( 
.A1(n_9733),
.A2(n_411),
.B(n_412),
.Y(n_10389)
);

AND2x2_ASAP7_75t_L g10390 ( 
.A(n_9989),
.B(n_412),
.Y(n_10390)
);

BUFx6f_ASAP7_75t_L g10391 ( 
.A(n_9631),
.Y(n_10391)
);

A2O1A1Ixp33_ASAP7_75t_L g10392 ( 
.A1(n_9716),
.A2(n_415),
.B(n_413),
.C(n_414),
.Y(n_10392)
);

AOI21xp5_ASAP7_75t_L g10393 ( 
.A1(n_9746),
.A2(n_413),
.B(n_414),
.Y(n_10393)
);

INVx1_ASAP7_75t_L g10394 ( 
.A(n_9737),
.Y(n_10394)
);

A2O1A1Ixp33_ASAP7_75t_L g10395 ( 
.A1(n_9720),
.A2(n_418),
.B(n_416),
.C(n_417),
.Y(n_10395)
);

INVx1_ASAP7_75t_L g10396 ( 
.A(n_9744),
.Y(n_10396)
);

INVx2_ASAP7_75t_L g10397 ( 
.A(n_9577),
.Y(n_10397)
);

INVx1_ASAP7_75t_L g10398 ( 
.A(n_9502),
.Y(n_10398)
);

AOI21x1_ASAP7_75t_L g10399 ( 
.A1(n_9830),
.A2(n_416),
.B(n_417),
.Y(n_10399)
);

OAI22xp5_ASAP7_75t_L g10400 ( 
.A1(n_9944),
.A2(n_421),
.B1(n_419),
.B2(n_420),
.Y(n_10400)
);

AOI21xp5_ASAP7_75t_L g10401 ( 
.A1(n_9749),
.A2(n_419),
.B(n_421),
.Y(n_10401)
);

NAND2xp5_ASAP7_75t_SL g10402 ( 
.A(n_9866),
.B(n_422),
.Y(n_10402)
);

OAI21xp5_ASAP7_75t_L g10403 ( 
.A1(n_9451),
.A2(n_422),
.B(n_423),
.Y(n_10403)
);

OAI21xp5_ASAP7_75t_L g10404 ( 
.A1(n_9456),
.A2(n_423),
.B(n_424),
.Y(n_10404)
);

AOI21xp5_ASAP7_75t_L g10405 ( 
.A1(n_9523),
.A2(n_424),
.B(n_425),
.Y(n_10405)
);

INVx11_ASAP7_75t_L g10406 ( 
.A(n_9921),
.Y(n_10406)
);

NOR2xp33_ASAP7_75t_L g10407 ( 
.A(n_9936),
.B(n_425),
.Y(n_10407)
);

OAI21xp5_ASAP7_75t_L g10408 ( 
.A1(n_9581),
.A2(n_426),
.B(n_427),
.Y(n_10408)
);

BUFx8_ASAP7_75t_SL g10409 ( 
.A(n_9937),
.Y(n_10409)
);

AOI21xp5_ASAP7_75t_L g10410 ( 
.A1(n_9531),
.A2(n_9544),
.B(n_9541),
.Y(n_10410)
);

NAND2xp5_ASAP7_75t_SL g10411 ( 
.A(n_9948),
.B(n_426),
.Y(n_10411)
);

OR2x2_ASAP7_75t_L g10412 ( 
.A(n_9546),
.B(n_427),
.Y(n_10412)
);

NAND2xp5_ASAP7_75t_SL g10413 ( 
.A(n_9953),
.B(n_428),
.Y(n_10413)
);

AOI21xp5_ASAP7_75t_L g10414 ( 
.A1(n_9550),
.A2(n_429),
.B(n_430),
.Y(n_10414)
);

A2O1A1Ixp33_ASAP7_75t_L g10415 ( 
.A1(n_9582),
.A2(n_431),
.B(n_429),
.C(n_430),
.Y(n_10415)
);

O2A1O1Ixp5_ASAP7_75t_L g10416 ( 
.A1(n_9865),
.A2(n_9870),
.B(n_9867),
.C(n_9857),
.Y(n_10416)
);

AOI21xp5_ASAP7_75t_L g10417 ( 
.A1(n_9555),
.A2(n_431),
.B(n_432),
.Y(n_10417)
);

AOI21xp5_ASAP7_75t_L g10418 ( 
.A1(n_9559),
.A2(n_9560),
.B(n_9911),
.Y(n_10418)
);

NOR2xp33_ASAP7_75t_L g10419 ( 
.A(n_9890),
.B(n_9895),
.Y(n_10419)
);

AOI21xp5_ASAP7_75t_L g10420 ( 
.A1(n_9915),
.A2(n_432),
.B(n_433),
.Y(n_10420)
);

OAI22xp5_ASAP7_75t_L g10421 ( 
.A1(n_9818),
.A2(n_435),
.B1(n_433),
.B2(n_434),
.Y(n_10421)
);

AOI22xp5_ASAP7_75t_L g10422 ( 
.A1(n_9779),
.A2(n_437),
.B1(n_434),
.B2(n_436),
.Y(n_10422)
);

CKINVDCx10_ASAP7_75t_R g10423 ( 
.A(n_9818),
.Y(n_10423)
);

NOR3xp33_ASAP7_75t_L g10424 ( 
.A(n_9947),
.B(n_436),
.C(n_437),
.Y(n_10424)
);

CKINVDCx5p33_ASAP7_75t_R g10425 ( 
.A(n_9515),
.Y(n_10425)
);

AOI21xp5_ASAP7_75t_L g10426 ( 
.A1(n_9920),
.A2(n_438),
.B(n_439),
.Y(n_10426)
);

INVx2_ASAP7_75t_L g10427 ( 
.A(n_9588),
.Y(n_10427)
);

AOI22xp5_ASAP7_75t_L g10428 ( 
.A1(n_9837),
.A2(n_441),
.B1(n_439),
.B2(n_440),
.Y(n_10428)
);

INVx3_ASAP7_75t_L g10429 ( 
.A(n_9567),
.Y(n_10429)
);

OAI22xp5_ASAP7_75t_L g10430 ( 
.A1(n_9942),
.A2(n_442),
.B1(n_440),
.B2(n_441),
.Y(n_10430)
);

NAND2xp5_ASAP7_75t_L g10431 ( 
.A(n_9586),
.B(n_442),
.Y(n_10431)
);

AOI21xp5_ASAP7_75t_L g10432 ( 
.A1(n_9872),
.A2(n_443),
.B(n_444),
.Y(n_10432)
);

INVx5_ASAP7_75t_L g10433 ( 
.A(n_9542),
.Y(n_10433)
);

BUFx2_ASAP7_75t_L g10434 ( 
.A(n_9639),
.Y(n_10434)
);

AOI21xp5_ASAP7_75t_L g10435 ( 
.A1(n_9846),
.A2(n_443),
.B(n_444),
.Y(n_10435)
);

AOI21x1_ASAP7_75t_L g10436 ( 
.A1(n_9784),
.A2(n_445),
.B(n_446),
.Y(n_10436)
);

BUFx6f_ASAP7_75t_L g10437 ( 
.A(n_9631),
.Y(n_10437)
);

NOR2xp33_ASAP7_75t_L g10438 ( 
.A(n_9792),
.B(n_446),
.Y(n_10438)
);

INVx1_ASAP7_75t_L g10439 ( 
.A(n_9594),
.Y(n_10439)
);

AOI21xp5_ASAP7_75t_L g10440 ( 
.A1(n_9858),
.A2(n_447),
.B(n_448),
.Y(n_10440)
);

INVx2_ASAP7_75t_SL g10441 ( 
.A(n_9590),
.Y(n_10441)
);

AOI21xp5_ASAP7_75t_L g10442 ( 
.A1(n_9860),
.A2(n_447),
.B(n_448),
.Y(n_10442)
);

NAND2xp5_ASAP7_75t_L g10443 ( 
.A(n_9595),
.B(n_449),
.Y(n_10443)
);

NOR2xp33_ASAP7_75t_L g10444 ( 
.A(n_9958),
.B(n_449),
.Y(n_10444)
);

NOR2xp33_ASAP7_75t_L g10445 ( 
.A(n_9538),
.B(n_450),
.Y(n_10445)
);

AOI21xp5_ASAP7_75t_L g10446 ( 
.A1(n_9607),
.A2(n_451),
.B(n_452),
.Y(n_10446)
);

NOR2xp33_ASAP7_75t_L g10447 ( 
.A(n_9945),
.B(n_451),
.Y(n_10447)
);

O2A1O1Ixp33_ASAP7_75t_L g10448 ( 
.A1(n_9925),
.A2(n_454),
.B(n_452),
.C(n_453),
.Y(n_10448)
);

NAND2xp5_ASAP7_75t_L g10449 ( 
.A(n_9611),
.B(n_453),
.Y(n_10449)
);

NAND2xp5_ASAP7_75t_L g10450 ( 
.A(n_9621),
.B(n_9628),
.Y(n_10450)
);

NOR2xp33_ASAP7_75t_L g10451 ( 
.A(n_9697),
.B(n_454),
.Y(n_10451)
);

AOI21xp5_ASAP7_75t_L g10452 ( 
.A1(n_9636),
.A2(n_456),
.B(n_457),
.Y(n_10452)
);

BUFx6f_ASAP7_75t_L g10453 ( 
.A(n_10028),
.Y(n_10453)
);

CKINVDCx14_ASAP7_75t_R g10454 ( 
.A(n_9768),
.Y(n_10454)
);

NAND3xp33_ASAP7_75t_L g10455 ( 
.A(n_9677),
.B(n_456),
.C(n_457),
.Y(n_10455)
);

NAND2xp5_ASAP7_75t_L g10456 ( 
.A(n_9641),
.B(n_458),
.Y(n_10456)
);

NAND2xp5_ASAP7_75t_L g10457 ( 
.A(n_9649),
.B(n_458),
.Y(n_10457)
);

NAND2xp5_ASAP7_75t_L g10458 ( 
.A(n_9651),
.B(n_459),
.Y(n_10458)
);

NAND3xp33_ASAP7_75t_L g10459 ( 
.A(n_9763),
.B(n_459),
.C(n_460),
.Y(n_10459)
);

INVx1_ASAP7_75t_L g10460 ( 
.A(n_9752),
.Y(n_10460)
);

BUFx3_ASAP7_75t_L g10461 ( 
.A(n_9573),
.Y(n_10461)
);

NAND2xp33_ASAP7_75t_L g10462 ( 
.A(n_10042),
.B(n_460),
.Y(n_10462)
);

INVx2_ASAP7_75t_L g10463 ( 
.A(n_9753),
.Y(n_10463)
);

NAND2xp5_ASAP7_75t_SL g10464 ( 
.A(n_9912),
.B(n_9922),
.Y(n_10464)
);

NAND2xp5_ASAP7_75t_L g10465 ( 
.A(n_9754),
.B(n_461),
.Y(n_10465)
);

INVx1_ASAP7_75t_L g10466 ( 
.A(n_9774),
.Y(n_10466)
);

AOI21xp5_ASAP7_75t_L g10467 ( 
.A1(n_9924),
.A2(n_462),
.B(n_463),
.Y(n_10467)
);

NAND2xp5_ASAP7_75t_L g10468 ( 
.A(n_9568),
.B(n_462),
.Y(n_10468)
);

AOI21xp5_ASAP7_75t_L g10469 ( 
.A1(n_9926),
.A2(n_463),
.B(n_464),
.Y(n_10469)
);

NAND2xp5_ASAP7_75t_L g10470 ( 
.A(n_9626),
.B(n_464),
.Y(n_10470)
);

OAI21xp5_ASAP7_75t_L g10471 ( 
.A1(n_9927),
.A2(n_465),
.B(n_466),
.Y(n_10471)
);

AOI21xp5_ASAP7_75t_L g10472 ( 
.A1(n_9884),
.A2(n_465),
.B(n_466),
.Y(n_10472)
);

HB1xp67_ASAP7_75t_L g10473 ( 
.A(n_9707),
.Y(n_10473)
);

HB1xp67_ASAP7_75t_L g10474 ( 
.A(n_9727),
.Y(n_10474)
);

INVx2_ASAP7_75t_L g10475 ( 
.A(n_9729),
.Y(n_10475)
);

AOI21xp5_ASAP7_75t_L g10476 ( 
.A1(n_9894),
.A2(n_467),
.B(n_468),
.Y(n_10476)
);

AOI21xp5_ASAP7_75t_L g10477 ( 
.A1(n_9810),
.A2(n_467),
.B(n_469),
.Y(n_10477)
);

INVx2_ASAP7_75t_L g10478 ( 
.A(n_9643),
.Y(n_10478)
);

OAI21x1_ASAP7_75t_L g10479 ( 
.A1(n_9674),
.A2(n_469),
.B(n_470),
.Y(n_10479)
);

NAND2xp5_ASAP7_75t_L g10480 ( 
.A(n_9799),
.B(n_471),
.Y(n_10480)
);

AOI21xp5_ASAP7_75t_L g10481 ( 
.A1(n_9955),
.A2(n_9904),
.B(n_9932),
.Y(n_10481)
);

AOI21xp5_ASAP7_75t_L g10482 ( 
.A1(n_9933),
.A2(n_472),
.B(n_473),
.Y(n_10482)
);

INVx2_ASAP7_75t_L g10483 ( 
.A(n_9644),
.Y(n_10483)
);

NAND2xp5_ASAP7_75t_L g10484 ( 
.A(n_9585),
.B(n_472),
.Y(n_10484)
);

HB1xp67_ASAP7_75t_L g10485 ( 
.A(n_9526),
.Y(n_10485)
);

AOI21xp5_ASAP7_75t_L g10486 ( 
.A1(n_9675),
.A2(n_473),
.B(n_474),
.Y(n_10486)
);

NOR2xp67_ASAP7_75t_L g10487 ( 
.A(n_9963),
.B(n_474),
.Y(n_10487)
);

NAND2xp5_ASAP7_75t_L g10488 ( 
.A(n_9587),
.B(n_9597),
.Y(n_10488)
);

OAI21xp5_ASAP7_75t_L g10489 ( 
.A1(n_9453),
.A2(n_475),
.B(n_476),
.Y(n_10489)
);

A2O1A1Ixp33_ASAP7_75t_L g10490 ( 
.A1(n_9601),
.A2(n_478),
.B(n_475),
.C(n_476),
.Y(n_10490)
);

AOI21xp5_ASAP7_75t_L g10491 ( 
.A1(n_9816),
.A2(n_478),
.B(n_479),
.Y(n_10491)
);

BUFx2_ASAP7_75t_L g10492 ( 
.A(n_9610),
.Y(n_10492)
);

OAI21xp33_ASAP7_75t_L g10493 ( 
.A1(n_9793),
.A2(n_479),
.B(n_480),
.Y(n_10493)
);

OAI21xp5_ASAP7_75t_L g10494 ( 
.A1(n_9476),
.A2(n_480),
.B(n_481),
.Y(n_10494)
);

AND2x2_ASAP7_75t_L g10495 ( 
.A(n_10002),
.B(n_482),
.Y(n_10495)
);

NOR2xp33_ASAP7_75t_L g10496 ( 
.A(n_9803),
.B(n_482),
.Y(n_10496)
);

OAI21xp5_ASAP7_75t_L g10497 ( 
.A1(n_9481),
.A2(n_483),
.B(n_484),
.Y(n_10497)
);

NAND2xp5_ASAP7_75t_L g10498 ( 
.A(n_9728),
.B(n_483),
.Y(n_10498)
);

HB1xp67_ASAP7_75t_L g10499 ( 
.A(n_9620),
.Y(n_10499)
);

NOR2x1p5_ASAP7_75t_SL g10500 ( 
.A(n_9571),
.B(n_484),
.Y(n_10500)
);

NAND2xp5_ASAP7_75t_L g10501 ( 
.A(n_9676),
.B(n_9708),
.Y(n_10501)
);

AOI21xp33_ASAP7_75t_L g10502 ( 
.A1(n_9480),
.A2(n_485),
.B(n_486),
.Y(n_10502)
);

AOI21xp5_ASAP7_75t_L g10503 ( 
.A1(n_9817),
.A2(n_485),
.B(n_486),
.Y(n_10503)
);

NAND2xp5_ASAP7_75t_L g10504 ( 
.A(n_9730),
.B(n_487),
.Y(n_10504)
);

HB1xp67_ASAP7_75t_L g10505 ( 
.A(n_9652),
.Y(n_10505)
);

AOI21xp5_ASAP7_75t_L g10506 ( 
.A1(n_9820),
.A2(n_487),
.B(n_488),
.Y(n_10506)
);

AND2x2_ASAP7_75t_L g10507 ( 
.A(n_10005),
.B(n_488),
.Y(n_10507)
);

O2A1O1Ixp33_ASAP7_75t_L g10508 ( 
.A1(n_9667),
.A2(n_9954),
.B(n_9888),
.C(n_9908),
.Y(n_10508)
);

NAND2x1p5_ASAP7_75t_L g10509 ( 
.A(n_9448),
.B(n_9686),
.Y(n_10509)
);

AOI21xp5_ASAP7_75t_L g10510 ( 
.A1(n_9826),
.A2(n_489),
.B(n_490),
.Y(n_10510)
);

AOI21xp5_ASAP7_75t_L g10511 ( 
.A1(n_9831),
.A2(n_489),
.B(n_490),
.Y(n_10511)
);

NOR2xp33_ASAP7_75t_L g10512 ( 
.A(n_9912),
.B(n_491),
.Y(n_10512)
);

INVx1_ASAP7_75t_L g10513 ( 
.A(n_9648),
.Y(n_10513)
);

NOR2x1_ASAP7_75t_R g10514 ( 
.A(n_9864),
.B(n_491),
.Y(n_10514)
);

AOI21xp5_ASAP7_75t_L g10515 ( 
.A1(n_9833),
.A2(n_492),
.B(n_493),
.Y(n_10515)
);

INVx2_ASAP7_75t_SL g10516 ( 
.A(n_10042),
.Y(n_10516)
);

OAI21xp5_ASAP7_75t_L g10517 ( 
.A1(n_9493),
.A2(n_494),
.B(n_495),
.Y(n_10517)
);

AO22x1_ASAP7_75t_L g10518 ( 
.A1(n_9775),
.A2(n_497),
.B1(n_494),
.B2(n_496),
.Y(n_10518)
);

NAND2xp5_ASAP7_75t_L g10519 ( 
.A(n_9835),
.B(n_497),
.Y(n_10519)
);

AOI21x1_ASAP7_75t_L g10520 ( 
.A1(n_9840),
.A2(n_498),
.B(n_499),
.Y(n_10520)
);

AOI22xp5_ASAP7_75t_L g10521 ( 
.A1(n_9889),
.A2(n_500),
.B1(n_498),
.B2(n_499),
.Y(n_10521)
);

CKINVDCx5p33_ASAP7_75t_R g10522 ( 
.A(n_9906),
.Y(n_10522)
);

AOI21xp5_ASAP7_75t_L g10523 ( 
.A1(n_9841),
.A2(n_9853),
.B(n_9848),
.Y(n_10523)
);

OAI21xp33_ASAP7_75t_L g10524 ( 
.A1(n_9859),
.A2(n_500),
.B(n_501),
.Y(n_10524)
);

NAND2xp33_ASAP7_75t_L g10525 ( 
.A(n_9959),
.B(n_502),
.Y(n_10525)
);

AND2x2_ASAP7_75t_L g10526 ( 
.A(n_10007),
.B(n_502),
.Y(n_10526)
);

OAI22xp5_ASAP7_75t_L g10527 ( 
.A1(n_9539),
.A2(n_505),
.B1(n_503),
.B2(n_504),
.Y(n_10527)
);

NAND3xp33_ASAP7_75t_L g10528 ( 
.A(n_9914),
.B(n_503),
.C(n_504),
.Y(n_10528)
);

NAND2xp5_ASAP7_75t_L g10529 ( 
.A(n_9861),
.B(n_505),
.Y(n_10529)
);

AOI21xp5_ASAP7_75t_L g10530 ( 
.A1(n_9484),
.A2(n_506),
.B(n_507),
.Y(n_10530)
);

NAND2xp5_ASAP7_75t_L g10531 ( 
.A(n_9806),
.B(n_9743),
.Y(n_10531)
);

INVx11_ASAP7_75t_L g10532 ( 
.A(n_9540),
.Y(n_10532)
);

BUFx12f_ASAP7_75t_L g10533 ( 
.A(n_9776),
.Y(n_10533)
);

AND2x2_ASAP7_75t_L g10534 ( 
.A(n_10010),
.B(n_506),
.Y(n_10534)
);

INVx1_ASAP7_75t_L g10535 ( 
.A(n_9653),
.Y(n_10535)
);

AOI221xp5_ASAP7_75t_L g10536 ( 
.A1(n_9766),
.A2(n_510),
.B1(n_508),
.B2(n_509),
.C(n_511),
.Y(n_10536)
);

AOI21xp5_ASAP7_75t_L g10537 ( 
.A1(n_9495),
.A2(n_510),
.B(n_511),
.Y(n_10537)
);

INVx1_ASAP7_75t_L g10538 ( 
.A(n_9751),
.Y(n_10538)
);

OAI21xp5_ASAP7_75t_L g10539 ( 
.A1(n_9447),
.A2(n_512),
.B(n_513),
.Y(n_10539)
);

INVx3_ASAP7_75t_L g10540 ( 
.A(n_9671),
.Y(n_10540)
);

INVx1_ASAP7_75t_L g10541 ( 
.A(n_9715),
.Y(n_10541)
);

AOI21x1_ASAP7_75t_L g10542 ( 
.A1(n_9488),
.A2(n_513),
.B(n_514),
.Y(n_10542)
);

AOI21xp5_ASAP7_75t_L g10543 ( 
.A1(n_9600),
.A2(n_515),
.B(n_516),
.Y(n_10543)
);

AOI21xp5_ASAP7_75t_L g10544 ( 
.A1(n_9613),
.A2(n_9625),
.B(n_9537),
.Y(n_10544)
);

NAND2xp5_ASAP7_75t_L g10545 ( 
.A(n_9745),
.B(n_515),
.Y(n_10545)
);

AOI21xp5_ASAP7_75t_L g10546 ( 
.A1(n_9533),
.A2(n_517),
.B(n_518),
.Y(n_10546)
);

O2A1O1Ixp33_ASAP7_75t_L g10547 ( 
.A1(n_9946),
.A2(n_522),
.B(n_519),
.C(n_520),
.Y(n_10547)
);

AOI21xp5_ASAP7_75t_L g10548 ( 
.A1(n_9808),
.A2(n_519),
.B(n_523),
.Y(n_10548)
);

INVx2_ASAP7_75t_L g10549 ( 
.A(n_9659),
.Y(n_10549)
);

NAND2xp5_ASAP7_75t_L g10550 ( 
.A(n_10013),
.B(n_523),
.Y(n_10550)
);

NOR2xp33_ASAP7_75t_L g10551 ( 
.A(n_9794),
.B(n_524),
.Y(n_10551)
);

INVx2_ASAP7_75t_L g10552 ( 
.A(n_9637),
.Y(n_10552)
);

NAND2xp5_ASAP7_75t_L g10553 ( 
.A(n_10014),
.B(n_524),
.Y(n_10553)
);

AOI22xp5_ASAP7_75t_L g10554 ( 
.A1(n_9959),
.A2(n_528),
.B1(n_525),
.B2(n_526),
.Y(n_10554)
);

AND2x2_ASAP7_75t_L g10555 ( 
.A(n_10019),
.B(n_525),
.Y(n_10555)
);

NAND2xp5_ASAP7_75t_L g10556 ( 
.A(n_10020),
.B(n_526),
.Y(n_10556)
);

AOI21xp5_ASAP7_75t_L g10557 ( 
.A1(n_9603),
.A2(n_528),
.B(n_529),
.Y(n_10557)
);

NAND2xp5_ASAP7_75t_L g10558 ( 
.A(n_10041),
.B(n_529),
.Y(n_10558)
);

NAND3xp33_ASAP7_75t_L g10559 ( 
.A(n_9949),
.B(n_9928),
.C(n_9606),
.Y(n_10559)
);

AOI21xp5_ASAP7_75t_L g10560 ( 
.A1(n_9518),
.A2(n_530),
.B(n_531),
.Y(n_10560)
);

INVx2_ASAP7_75t_L g10561 ( 
.A(n_9646),
.Y(n_10561)
);

NAND2xp5_ASAP7_75t_L g10562 ( 
.A(n_10043),
.B(n_530),
.Y(n_10562)
);

AOI21xp5_ASAP7_75t_L g10563 ( 
.A1(n_9614),
.A2(n_531),
.B(n_532),
.Y(n_10563)
);

INVxp67_ASAP7_75t_L g10564 ( 
.A(n_9696),
.Y(n_10564)
);

AOI21xp5_ASAP7_75t_L g10565 ( 
.A1(n_9778),
.A2(n_532),
.B(n_533),
.Y(n_10565)
);

INVx11_ASAP7_75t_L g10566 ( 
.A(n_9548),
.Y(n_10566)
);

INVx3_ASAP7_75t_L g10567 ( 
.A(n_9580),
.Y(n_10567)
);

AND2x2_ASAP7_75t_L g10568 ( 
.A(n_9519),
.B(n_534),
.Y(n_10568)
);

NAND2xp5_ASAP7_75t_L g10569 ( 
.A(n_9722),
.B(n_534),
.Y(n_10569)
);

OR2x2_ASAP7_75t_L g10570 ( 
.A(n_9511),
.B(n_535),
.Y(n_10570)
);

AOI21xp5_ASAP7_75t_L g10571 ( 
.A1(n_9513),
.A2(n_535),
.B(n_536),
.Y(n_10571)
);

AND2x4_ASAP7_75t_L g10572 ( 
.A(n_9735),
.B(n_536),
.Y(n_10572)
);

AOI21xp5_ASAP7_75t_L g10573 ( 
.A1(n_9787),
.A2(n_537),
.B(n_539),
.Y(n_10573)
);

AOI21xp5_ASAP7_75t_L g10574 ( 
.A1(n_9446),
.A2(n_537),
.B(n_540),
.Y(n_10574)
);

AOI21xp33_ASAP7_75t_L g10575 ( 
.A1(n_9558),
.A2(n_541),
.B(n_542),
.Y(n_10575)
);

AOI21x1_ASAP7_75t_L g10576 ( 
.A1(n_9627),
.A2(n_543),
.B(n_544),
.Y(n_10576)
);

NOR2xp33_ASAP7_75t_SL g10577 ( 
.A(n_9899),
.B(n_544),
.Y(n_10577)
);

NAND2xp5_ASAP7_75t_L g10578 ( 
.A(n_9623),
.B(n_545),
.Y(n_10578)
);

INVx1_ASAP7_75t_SL g10579 ( 
.A(n_9714),
.Y(n_10579)
);

AOI21xp5_ASAP7_75t_L g10580 ( 
.A1(n_9566),
.A2(n_545),
.B(n_546),
.Y(n_10580)
);

AOI21x1_ASAP7_75t_L g10581 ( 
.A1(n_9705),
.A2(n_546),
.B(n_547),
.Y(n_10581)
);

BUFx8_ASAP7_75t_L g10582 ( 
.A(n_9776),
.Y(n_10582)
);

NAND2xp5_ASAP7_75t_L g10583 ( 
.A(n_9521),
.B(n_547),
.Y(n_10583)
);

AOI21xp5_ASAP7_75t_L g10584 ( 
.A1(n_9522),
.A2(n_548),
.B(n_549),
.Y(n_10584)
);

INVx3_ASAP7_75t_L g10585 ( 
.A(n_9645),
.Y(n_10585)
);

AOI21xp5_ASAP7_75t_L g10586 ( 
.A1(n_9525),
.A2(n_548),
.B(n_549),
.Y(n_10586)
);

OAI21xp5_ASAP7_75t_L g10587 ( 
.A1(n_9532),
.A2(n_550),
.B(n_551),
.Y(n_10587)
);

AOI21xp5_ASAP7_75t_L g10588 ( 
.A1(n_9957),
.A2(n_10017),
.B(n_9981),
.Y(n_10588)
);

NAND2xp33_ASAP7_75t_L g10589 ( 
.A(n_9906),
.B(n_550),
.Y(n_10589)
);

NAND2xp5_ASAP7_75t_SL g10590 ( 
.A(n_10025),
.B(n_551),
.Y(n_10590)
);

NOR2xp33_ASAP7_75t_L g10591 ( 
.A(n_9975),
.B(n_552),
.Y(n_10591)
);

AOI21xp5_ASAP7_75t_L g10592 ( 
.A1(n_10029),
.A2(n_552),
.B(n_553),
.Y(n_10592)
);

NOR2xp33_ASAP7_75t_SL g10593 ( 
.A(n_9458),
.B(n_553),
.Y(n_10593)
);

INVx1_ASAP7_75t_L g10594 ( 
.A(n_9706),
.Y(n_10594)
);

INVx1_ASAP7_75t_L g10595 ( 
.A(n_9657),
.Y(n_10595)
);

AOI21xp5_ASAP7_75t_L g10596 ( 
.A1(n_9486),
.A2(n_9535),
.B(n_9516),
.Y(n_10596)
);

NOR2xp33_ASAP7_75t_L g10597 ( 
.A(n_10038),
.B(n_555),
.Y(n_10597)
);

NAND2xp5_ASAP7_75t_SL g10598 ( 
.A(n_9657),
.B(n_555),
.Y(n_10598)
);

AOI21xp5_ASAP7_75t_L g10599 ( 
.A1(n_9655),
.A2(n_556),
.B(n_558),
.Y(n_10599)
);

HB1xp67_ASAP7_75t_L g10600 ( 
.A(n_9679),
.Y(n_10600)
);

AOI21xp5_ASAP7_75t_L g10601 ( 
.A1(n_9971),
.A2(n_556),
.B(n_558),
.Y(n_10601)
);

OAI21xp5_ASAP7_75t_L g10602 ( 
.A1(n_9983),
.A2(n_559),
.B(n_560),
.Y(n_10602)
);

O2A1O1Ixp5_ASAP7_75t_L g10603 ( 
.A1(n_10011),
.A2(n_561),
.B(n_559),
.C(n_560),
.Y(n_10603)
);

AOI21xp5_ASAP7_75t_L g10604 ( 
.A1(n_10030),
.A2(n_561),
.B(n_562),
.Y(n_10604)
);

NOR3xp33_ASAP7_75t_L g10605 ( 
.A(n_10036),
.B(n_562),
.C(n_563),
.Y(n_10605)
);

CKINVDCx10_ASAP7_75t_R g10606 ( 
.A(n_9679),
.Y(n_10606)
);

INVx1_ASAP7_75t_L g10607 ( 
.A(n_9563),
.Y(n_10607)
);

INVx2_ASAP7_75t_SL g10608 ( 
.A(n_9561),
.Y(n_10608)
);

AOI22xp33_ASAP7_75t_L g10609 ( 
.A1(n_9565),
.A2(n_565),
.B1(n_563),
.B2(n_564),
.Y(n_10609)
);

OAI21xp5_ASAP7_75t_L g10610 ( 
.A1(n_9469),
.A2(n_565),
.B(n_566),
.Y(n_10610)
);

INVx1_ASAP7_75t_L g10611 ( 
.A(n_9563),
.Y(n_10611)
);

OAI22xp5_ASAP7_75t_L g10612 ( 
.A1(n_9678),
.A2(n_569),
.B1(n_567),
.B2(n_568),
.Y(n_10612)
);

AOI21xp5_ASAP7_75t_L g10613 ( 
.A1(n_9731),
.A2(n_567),
.B(n_568),
.Y(n_10613)
);

NAND2xp5_ASAP7_75t_L g10614 ( 
.A(n_9557),
.B(n_569),
.Y(n_10614)
);

AOI21xp5_ASAP7_75t_L g10615 ( 
.A1(n_9731),
.A2(n_570),
.B(n_571),
.Y(n_10615)
);

INVx2_ASAP7_75t_L g10616 ( 
.A(n_9444),
.Y(n_10616)
);

INVx1_ASAP7_75t_L g10617 ( 
.A(n_9563),
.Y(n_10617)
);

NAND2xp5_ASAP7_75t_L g10618 ( 
.A(n_9557),
.B(n_570),
.Y(n_10618)
);

OAI22xp5_ASAP7_75t_L g10619 ( 
.A1(n_9678),
.A2(n_574),
.B1(n_572),
.B2(n_573),
.Y(n_10619)
);

AOI21xp5_ASAP7_75t_L g10620 ( 
.A1(n_9731),
.A2(n_573),
.B(n_574),
.Y(n_10620)
);

NAND2xp5_ASAP7_75t_L g10621 ( 
.A(n_9557),
.B(n_575),
.Y(n_10621)
);

A2O1A1Ixp33_ASAP7_75t_L g10622 ( 
.A1(n_9624),
.A2(n_577),
.B(n_575),
.C(n_576),
.Y(n_10622)
);

NAND2xp5_ASAP7_75t_L g10623 ( 
.A(n_9557),
.B(n_577),
.Y(n_10623)
);

OAI21xp5_ASAP7_75t_L g10624 ( 
.A1(n_9469),
.A2(n_578),
.B(n_579),
.Y(n_10624)
);

INVx2_ASAP7_75t_L g10625 ( 
.A(n_9444),
.Y(n_10625)
);

NAND2xp5_ASAP7_75t_L g10626 ( 
.A(n_9557),
.B(n_578),
.Y(n_10626)
);

NAND2xp5_ASAP7_75t_SL g10627 ( 
.A(n_9596),
.B(n_580),
.Y(n_10627)
);

AOI21xp5_ASAP7_75t_L g10628 ( 
.A1(n_9731),
.A2(n_580),
.B(n_581),
.Y(n_10628)
);

AOI21xp5_ASAP7_75t_L g10629 ( 
.A1(n_9731),
.A2(n_581),
.B(n_582),
.Y(n_10629)
);

NOR2xp33_ASAP7_75t_L g10630 ( 
.A(n_9678),
.B(n_582),
.Y(n_10630)
);

NAND2xp5_ASAP7_75t_L g10631 ( 
.A(n_9557),
.B(n_583),
.Y(n_10631)
);

AOI21xp33_ASAP7_75t_L g10632 ( 
.A1(n_9469),
.A2(n_583),
.B(n_584),
.Y(n_10632)
);

NAND2xp5_ASAP7_75t_L g10633 ( 
.A(n_9557),
.B(n_584),
.Y(n_10633)
);

INVx2_ASAP7_75t_L g10634 ( 
.A(n_9444),
.Y(n_10634)
);

NAND2xp5_ASAP7_75t_L g10635 ( 
.A(n_9557),
.B(n_585),
.Y(n_10635)
);

AND2x4_ASAP7_75t_L g10636 ( 
.A(n_9739),
.B(n_585),
.Y(n_10636)
);

AOI21xp5_ASAP7_75t_L g10637 ( 
.A1(n_9731),
.A2(n_586),
.B(n_587),
.Y(n_10637)
);

AND2x4_ASAP7_75t_L g10638 ( 
.A(n_9739),
.B(n_586),
.Y(n_10638)
);

NAND2x1_ASAP7_75t_L g10639 ( 
.A(n_9821),
.B(n_587),
.Y(n_10639)
);

INVx2_ASAP7_75t_L g10640 ( 
.A(n_9444),
.Y(n_10640)
);

NAND2xp5_ASAP7_75t_SL g10641 ( 
.A(n_9596),
.B(n_588),
.Y(n_10641)
);

OAI21xp5_ASAP7_75t_L g10642 ( 
.A1(n_9469),
.A2(n_588),
.B(n_589),
.Y(n_10642)
);

AND2x4_ASAP7_75t_L g10643 ( 
.A(n_9739),
.B(n_589),
.Y(n_10643)
);

NAND2xp5_ASAP7_75t_SL g10644 ( 
.A(n_9596),
.B(n_590),
.Y(n_10644)
);

NOR2xp33_ASAP7_75t_L g10645 ( 
.A(n_9678),
.B(n_590),
.Y(n_10645)
);

NAND2xp5_ASAP7_75t_L g10646 ( 
.A(n_9557),
.B(n_591),
.Y(n_10646)
);

INVx1_ASAP7_75t_L g10647 ( 
.A(n_9563),
.Y(n_10647)
);

NAND2xp5_ASAP7_75t_L g10648 ( 
.A(n_9557),
.B(n_591),
.Y(n_10648)
);

NAND2xp5_ASAP7_75t_SL g10649 ( 
.A(n_9596),
.B(n_592),
.Y(n_10649)
);

A2O1A1Ixp33_ASAP7_75t_L g10650 ( 
.A1(n_9624),
.A2(n_594),
.B(n_592),
.C(n_593),
.Y(n_10650)
);

AOI21xp5_ASAP7_75t_L g10651 ( 
.A1(n_9731),
.A2(n_593),
.B(n_594),
.Y(n_10651)
);

AOI21xp5_ASAP7_75t_L g10652 ( 
.A1(n_9731),
.A2(n_595),
.B(n_596),
.Y(n_10652)
);

OR2x6_ASAP7_75t_L g10653 ( 
.A(n_9821),
.B(n_595),
.Y(n_10653)
);

AOI21xp33_ASAP7_75t_L g10654 ( 
.A1(n_9469),
.A2(n_596),
.B(n_597),
.Y(n_10654)
);

AOI21xp5_ASAP7_75t_L g10655 ( 
.A1(n_9731),
.A2(n_598),
.B(n_599),
.Y(n_10655)
);

INVx1_ASAP7_75t_L g10656 ( 
.A(n_9563),
.Y(n_10656)
);

NAND2xp33_ASAP7_75t_L g10657 ( 
.A(n_9811),
.B(n_599),
.Y(n_10657)
);

NAND2xp5_ASAP7_75t_SL g10658 ( 
.A(n_9596),
.B(n_600),
.Y(n_10658)
);

INVx1_ASAP7_75t_L g10659 ( 
.A(n_9563),
.Y(n_10659)
);

AOI21xp5_ASAP7_75t_L g10660 ( 
.A1(n_9731),
.A2(n_601),
.B(n_602),
.Y(n_10660)
);

AOI21xp5_ASAP7_75t_L g10661 ( 
.A1(n_9731),
.A2(n_601),
.B(n_602),
.Y(n_10661)
);

BUFx6f_ASAP7_75t_L g10662 ( 
.A(n_9632),
.Y(n_10662)
);

AOI22x1_ASAP7_75t_L g10663 ( 
.A1(n_9783),
.A2(n_605),
.B1(n_603),
.B2(n_604),
.Y(n_10663)
);

NAND2xp5_ASAP7_75t_SL g10664 ( 
.A(n_9596),
.B(n_604),
.Y(n_10664)
);

AOI21xp5_ASAP7_75t_L g10665 ( 
.A1(n_9731),
.A2(n_605),
.B(n_606),
.Y(n_10665)
);

NAND2xp5_ASAP7_75t_L g10666 ( 
.A(n_9557),
.B(n_606),
.Y(n_10666)
);

O2A1O1Ixp33_ASAP7_75t_L g10667 ( 
.A1(n_9552),
.A2(n_609),
.B(n_607),
.C(n_608),
.Y(n_10667)
);

INVx3_ASAP7_75t_L g10668 ( 
.A(n_9470),
.Y(n_10668)
);

AOI21xp5_ASAP7_75t_L g10669 ( 
.A1(n_9731),
.A2(n_607),
.B(n_608),
.Y(n_10669)
);

INVx1_ASAP7_75t_L g10670 ( 
.A(n_9563),
.Y(n_10670)
);

AOI21xp5_ASAP7_75t_L g10671 ( 
.A1(n_9731),
.A2(n_610),
.B(n_611),
.Y(n_10671)
);

NAND2xp5_ASAP7_75t_SL g10672 ( 
.A(n_9596),
.B(n_611),
.Y(n_10672)
);

OAI21xp5_ASAP7_75t_L g10673 ( 
.A1(n_9469),
.A2(n_612),
.B(n_613),
.Y(n_10673)
);

OAI21xp5_ASAP7_75t_L g10674 ( 
.A1(n_9469),
.A2(n_612),
.B(n_613),
.Y(n_10674)
);

OAI21xp5_ASAP7_75t_L g10675 ( 
.A1(n_9469),
.A2(n_614),
.B(n_616),
.Y(n_10675)
);

INVx2_ASAP7_75t_L g10676 ( 
.A(n_9444),
.Y(n_10676)
);

NAND2xp5_ASAP7_75t_L g10677 ( 
.A(n_9557),
.B(n_614),
.Y(n_10677)
);

AOI21xp5_ASAP7_75t_L g10678 ( 
.A1(n_9731),
.A2(n_616),
.B(n_617),
.Y(n_10678)
);

NAND2xp5_ASAP7_75t_L g10679 ( 
.A(n_9557),
.B(n_617),
.Y(n_10679)
);

NAND2xp5_ASAP7_75t_L g10680 ( 
.A(n_9557),
.B(n_618),
.Y(n_10680)
);

AOI21xp5_ASAP7_75t_L g10681 ( 
.A1(n_9731),
.A2(n_618),
.B(n_620),
.Y(n_10681)
);

BUFx6f_ASAP7_75t_L g10682 ( 
.A(n_9632),
.Y(n_10682)
);

AO21x1_ASAP7_75t_L g10683 ( 
.A1(n_9704),
.A2(n_620),
.B(n_621),
.Y(n_10683)
);

BUFx6f_ASAP7_75t_L g10684 ( 
.A(n_9632),
.Y(n_10684)
);

OAI21xp5_ASAP7_75t_L g10685 ( 
.A1(n_9469),
.A2(n_621),
.B(n_622),
.Y(n_10685)
);

O2A1O1Ixp33_ASAP7_75t_L g10686 ( 
.A1(n_9552),
.A2(n_624),
.B(n_622),
.C(n_623),
.Y(n_10686)
);

AOI22xp33_ASAP7_75t_L g10687 ( 
.A1(n_9565),
.A2(n_625),
.B1(n_623),
.B2(n_624),
.Y(n_10687)
);

O2A1O1Ixp33_ASAP7_75t_L g10688 ( 
.A1(n_9552),
.A2(n_628),
.B(n_626),
.C(n_627),
.Y(n_10688)
);

AO21x1_ASAP7_75t_L g10689 ( 
.A1(n_9704),
.A2(n_626),
.B(n_628),
.Y(n_10689)
);

NAND2xp5_ASAP7_75t_L g10690 ( 
.A(n_9557),
.B(n_629),
.Y(n_10690)
);

INVx3_ASAP7_75t_L g10691 ( 
.A(n_9470),
.Y(n_10691)
);

NAND2xp5_ASAP7_75t_SL g10692 ( 
.A(n_9596),
.B(n_630),
.Y(n_10692)
);

INVx2_ASAP7_75t_L g10693 ( 
.A(n_9444),
.Y(n_10693)
);

AOI21xp5_ASAP7_75t_L g10694 ( 
.A1(n_9731),
.A2(n_630),
.B(n_631),
.Y(n_10694)
);

O2A1O1Ixp33_ASAP7_75t_L g10695 ( 
.A1(n_9552),
.A2(n_633),
.B(n_631),
.C(n_632),
.Y(n_10695)
);

OAI21x1_ASAP7_75t_L g10696 ( 
.A1(n_9454),
.A2(n_632),
.B(n_633),
.Y(n_10696)
);

AO21x1_ASAP7_75t_L g10697 ( 
.A1(n_9704),
.A2(n_635),
.B(n_636),
.Y(n_10697)
);

INVx1_ASAP7_75t_L g10698 ( 
.A(n_9563),
.Y(n_10698)
);

O2A1O1Ixp33_ASAP7_75t_L g10699 ( 
.A1(n_9552),
.A2(n_637),
.B(n_635),
.C(n_636),
.Y(n_10699)
);

AOI21xp5_ASAP7_75t_L g10700 ( 
.A1(n_9731),
.A2(n_637),
.B(n_639),
.Y(n_10700)
);

A2O1A1Ixp33_ASAP7_75t_L g10701 ( 
.A1(n_9624),
.A2(n_642),
.B(n_640),
.C(n_641),
.Y(n_10701)
);

INVx1_ASAP7_75t_L g10702 ( 
.A(n_9563),
.Y(n_10702)
);

AOI21xp5_ASAP7_75t_L g10703 ( 
.A1(n_9731),
.A2(n_640),
.B(n_641),
.Y(n_10703)
);

OAI21xp5_ASAP7_75t_L g10704 ( 
.A1(n_9469),
.A2(n_642),
.B(n_643),
.Y(n_10704)
);

AOI21xp5_ASAP7_75t_L g10705 ( 
.A1(n_9731),
.A2(n_643),
.B(n_644),
.Y(n_10705)
);

BUFx12f_ASAP7_75t_L g10706 ( 
.A(n_9504),
.Y(n_10706)
);

NAND2xp5_ASAP7_75t_L g10707 ( 
.A(n_9557),
.B(n_644),
.Y(n_10707)
);

INVx2_ASAP7_75t_SL g10708 ( 
.A(n_9561),
.Y(n_10708)
);

INVxp67_ASAP7_75t_L g10709 ( 
.A(n_9466),
.Y(n_10709)
);

NAND2xp5_ASAP7_75t_SL g10710 ( 
.A(n_9596),
.B(n_645),
.Y(n_10710)
);

NAND2xp5_ASAP7_75t_L g10711 ( 
.A(n_9557),
.B(n_646),
.Y(n_10711)
);

OAI21xp5_ASAP7_75t_L g10712 ( 
.A1(n_9469),
.A2(n_646),
.B(n_647),
.Y(n_10712)
);

AOI21xp5_ASAP7_75t_L g10713 ( 
.A1(n_9731),
.A2(n_647),
.B(n_648),
.Y(n_10713)
);

NOR2xp33_ASAP7_75t_L g10714 ( 
.A(n_9678),
.B(n_648),
.Y(n_10714)
);

INVxp67_ASAP7_75t_L g10715 ( 
.A(n_9466),
.Y(n_10715)
);

NAND2xp5_ASAP7_75t_L g10716 ( 
.A(n_9557),
.B(n_649),
.Y(n_10716)
);

INVx2_ASAP7_75t_L g10717 ( 
.A(n_9444),
.Y(n_10717)
);

OAI22xp5_ASAP7_75t_L g10718 ( 
.A1(n_9678),
.A2(n_652),
.B1(n_650),
.B2(n_651),
.Y(n_10718)
);

NAND2xp5_ASAP7_75t_SL g10719 ( 
.A(n_9596),
.B(n_650),
.Y(n_10719)
);

AOI21xp5_ASAP7_75t_L g10720 ( 
.A1(n_9731),
.A2(n_651),
.B(n_653),
.Y(n_10720)
);

O2A1O1Ixp33_ASAP7_75t_L g10721 ( 
.A1(n_9552),
.A2(n_655),
.B(n_653),
.C(n_654),
.Y(n_10721)
);

INVx1_ASAP7_75t_L g10722 ( 
.A(n_9563),
.Y(n_10722)
);

NAND2xp5_ASAP7_75t_L g10723 ( 
.A(n_9557),
.B(n_655),
.Y(n_10723)
);

INVx1_ASAP7_75t_SL g10724 ( 
.A(n_9487),
.Y(n_10724)
);

AOI21xp5_ASAP7_75t_L g10725 ( 
.A1(n_9731),
.A2(n_656),
.B(n_657),
.Y(n_10725)
);

NAND3xp33_ASAP7_75t_L g10726 ( 
.A(n_9552),
.B(n_656),
.C(n_657),
.Y(n_10726)
);

AND2x2_ASAP7_75t_L g10727 ( 
.A(n_9452),
.B(n_658),
.Y(n_10727)
);

OAI22xp5_ASAP7_75t_L g10728 ( 
.A1(n_9678),
.A2(n_660),
.B1(n_658),
.B2(n_659),
.Y(n_10728)
);

BUFx3_ASAP7_75t_L g10729 ( 
.A(n_9578),
.Y(n_10729)
);

AOI21xp5_ASAP7_75t_L g10730 ( 
.A1(n_9731),
.A2(n_659),
.B(n_661),
.Y(n_10730)
);

O2A1O1Ixp5_ASAP7_75t_L g10731 ( 
.A1(n_9783),
.A2(n_663),
.B(n_661),
.C(n_662),
.Y(n_10731)
);

AOI21xp33_ASAP7_75t_L g10732 ( 
.A1(n_9469),
.A2(n_662),
.B(n_663),
.Y(n_10732)
);

INVx1_ASAP7_75t_L g10733 ( 
.A(n_9563),
.Y(n_10733)
);

NOR3xp33_ASAP7_75t_L g10734 ( 
.A(n_9552),
.B(n_664),
.C(n_665),
.Y(n_10734)
);

NAND2xp5_ASAP7_75t_SL g10735 ( 
.A(n_9596),
.B(n_666),
.Y(n_10735)
);

INVx1_ASAP7_75t_L g10736 ( 
.A(n_9563),
.Y(n_10736)
);

INVx1_ASAP7_75t_L g10737 ( 
.A(n_9563),
.Y(n_10737)
);

NOR2xp33_ASAP7_75t_L g10738 ( 
.A(n_9678),
.B(n_666),
.Y(n_10738)
);

NOR2xp33_ASAP7_75t_L g10739 ( 
.A(n_9678),
.B(n_667),
.Y(n_10739)
);

NAND2xp5_ASAP7_75t_SL g10740 ( 
.A(n_9596),
.B(n_667),
.Y(n_10740)
);

OAI22xp5_ASAP7_75t_L g10741 ( 
.A1(n_9678),
.A2(n_670),
.B1(n_668),
.B2(n_669),
.Y(n_10741)
);

CKINVDCx20_ASAP7_75t_R g10742 ( 
.A(n_9976),
.Y(n_10742)
);

OAI21xp33_ASAP7_75t_L g10743 ( 
.A1(n_9552),
.A2(n_668),
.B(n_669),
.Y(n_10743)
);

AOI21xp5_ASAP7_75t_L g10744 ( 
.A1(n_9731),
.A2(n_670),
.B(n_671),
.Y(n_10744)
);

AND2x4_ASAP7_75t_L g10745 ( 
.A(n_9739),
.B(n_671),
.Y(n_10745)
);

INVx1_ASAP7_75t_L g10746 ( 
.A(n_9563),
.Y(n_10746)
);

NAND3xp33_ASAP7_75t_L g10747 ( 
.A(n_9552),
.B(n_672),
.C(n_673),
.Y(n_10747)
);

NAND2xp5_ASAP7_75t_SL g10748 ( 
.A(n_9596),
.B(n_672),
.Y(n_10748)
);

OAI321xp33_ASAP7_75t_L g10749 ( 
.A1(n_9974),
.A2(n_675),
.A3(n_677),
.B1(n_673),
.B2(n_674),
.C(n_676),
.Y(n_10749)
);

NAND2xp5_ASAP7_75t_L g10750 ( 
.A(n_9557),
.B(n_674),
.Y(n_10750)
);

AO21x1_ASAP7_75t_L g10751 ( 
.A1(n_9704),
.A2(n_675),
.B(n_676),
.Y(n_10751)
);

BUFx4f_ASAP7_75t_L g10752 ( 
.A(n_9632),
.Y(n_10752)
);

NOR2xp67_ASAP7_75t_L g10753 ( 
.A(n_9678),
.B(n_677),
.Y(n_10753)
);

NAND2xp5_ASAP7_75t_SL g10754 ( 
.A(n_9596),
.B(n_678),
.Y(n_10754)
);

INVx2_ASAP7_75t_L g10755 ( 
.A(n_9444),
.Y(n_10755)
);

INVxp67_ASAP7_75t_L g10756 ( 
.A(n_9466),
.Y(n_10756)
);

NOR2xp33_ASAP7_75t_L g10757 ( 
.A(n_9678),
.B(n_678),
.Y(n_10757)
);

NAND2xp5_ASAP7_75t_L g10758 ( 
.A(n_9557),
.B(n_679),
.Y(n_10758)
);

OAI21xp5_ASAP7_75t_L g10759 ( 
.A1(n_9469),
.A2(n_679),
.B(n_680),
.Y(n_10759)
);

NAND2xp5_ASAP7_75t_L g10760 ( 
.A(n_9557),
.B(n_680),
.Y(n_10760)
);

AOI21x1_ASAP7_75t_L g10761 ( 
.A1(n_9602),
.A2(n_681),
.B(n_682),
.Y(n_10761)
);

AND2x2_ASAP7_75t_L g10762 ( 
.A(n_9452),
.B(n_681),
.Y(n_10762)
);

NAND2xp5_ASAP7_75t_L g10763 ( 
.A(n_9557),
.B(n_682),
.Y(n_10763)
);

AOI21xp5_ASAP7_75t_L g10764 ( 
.A1(n_9731),
.A2(n_683),
.B(n_684),
.Y(n_10764)
);

O2A1O1Ixp33_ASAP7_75t_L g10765 ( 
.A1(n_9552),
.A2(n_685),
.B(n_683),
.C(n_684),
.Y(n_10765)
);

NAND2xp5_ASAP7_75t_L g10766 ( 
.A(n_9557),
.B(n_685),
.Y(n_10766)
);

A2O1A1Ixp33_ASAP7_75t_L g10767 ( 
.A1(n_9624),
.A2(n_688),
.B(n_686),
.C(n_687),
.Y(n_10767)
);

AOI21xp5_ASAP7_75t_L g10768 ( 
.A1(n_9731),
.A2(n_687),
.B(n_688),
.Y(n_10768)
);

AO21x1_ASAP7_75t_L g10769 ( 
.A1(n_9704),
.A2(n_689),
.B(n_690),
.Y(n_10769)
);

AND2x4_ASAP7_75t_L g10770 ( 
.A(n_9739),
.B(n_691),
.Y(n_10770)
);

NAND2xp5_ASAP7_75t_L g10771 ( 
.A(n_9557),
.B(n_691),
.Y(n_10771)
);

AND2x2_ASAP7_75t_L g10772 ( 
.A(n_9452),
.B(n_692),
.Y(n_10772)
);

O2A1O1Ixp5_ASAP7_75t_L g10773 ( 
.A1(n_9783),
.A2(n_694),
.B(n_692),
.C(n_693),
.Y(n_10773)
);

NOR2xp67_ASAP7_75t_L g10774 ( 
.A(n_9678),
.B(n_694),
.Y(n_10774)
);

NOR2xp33_ASAP7_75t_L g10775 ( 
.A(n_9678),
.B(n_695),
.Y(n_10775)
);

AOI21xp33_ASAP7_75t_L g10776 ( 
.A1(n_9469),
.A2(n_695),
.B(n_696),
.Y(n_10776)
);

CKINVDCx10_ASAP7_75t_R g10777 ( 
.A(n_9818),
.Y(n_10777)
);

NAND2xp5_ASAP7_75t_L g10778 ( 
.A(n_9557),
.B(n_696),
.Y(n_10778)
);

NOR2xp33_ASAP7_75t_L g10779 ( 
.A(n_9678),
.B(n_697),
.Y(n_10779)
);

NOR2xp33_ASAP7_75t_L g10780 ( 
.A(n_9678),
.B(n_698),
.Y(n_10780)
);

BUFx5_ASAP7_75t_L g10781 ( 
.A(n_9891),
.Y(n_10781)
);

AOI21xp5_ASAP7_75t_L g10782 ( 
.A1(n_9731),
.A2(n_698),
.B(n_699),
.Y(n_10782)
);

AOI21xp5_ASAP7_75t_L g10783 ( 
.A1(n_9731),
.A2(n_699),
.B(n_700),
.Y(n_10783)
);

NAND2xp5_ASAP7_75t_L g10784 ( 
.A(n_9557),
.B(n_700),
.Y(n_10784)
);

AOI21xp5_ASAP7_75t_L g10785 ( 
.A1(n_9731),
.A2(n_701),
.B(n_702),
.Y(n_10785)
);

INVx2_ASAP7_75t_L g10786 ( 
.A(n_9444),
.Y(n_10786)
);

OAI21x1_ASAP7_75t_L g10787 ( 
.A1(n_9454),
.A2(n_702),
.B(n_703),
.Y(n_10787)
);

OAI22xp5_ASAP7_75t_L g10788 ( 
.A1(n_9678),
.A2(n_705),
.B1(n_703),
.B2(n_704),
.Y(n_10788)
);

INVx1_ASAP7_75t_L g10789 ( 
.A(n_9563),
.Y(n_10789)
);

OR2x2_ASAP7_75t_L g10790 ( 
.A(n_10334),
.B(n_704),
.Y(n_10790)
);

INVx1_ASAP7_75t_L g10791 ( 
.A(n_10053),
.Y(n_10791)
);

BUFx3_ASAP7_75t_L g10792 ( 
.A(n_10175),
.Y(n_10792)
);

NOR2xp33_ASAP7_75t_L g10793 ( 
.A(n_10724),
.B(n_705),
.Y(n_10793)
);

AOI21xp5_ASAP7_75t_L g10794 ( 
.A1(n_10103),
.A2(n_706),
.B(n_707),
.Y(n_10794)
);

AOI21xp5_ASAP7_75t_L g10795 ( 
.A1(n_10047),
.A2(n_10657),
.B(n_10292),
.Y(n_10795)
);

INVx1_ASAP7_75t_L g10796 ( 
.A(n_10060),
.Y(n_10796)
);

AOI21xp5_ASAP7_75t_L g10797 ( 
.A1(n_10082),
.A2(n_706),
.B(n_707),
.Y(n_10797)
);

OAI22xp5_ASAP7_75t_SL g10798 ( 
.A1(n_10287),
.A2(n_710),
.B1(n_708),
.B2(n_709),
.Y(n_10798)
);

NAND2xp5_ASAP7_75t_L g10799 ( 
.A(n_10204),
.B(n_708),
.Y(n_10799)
);

AND2x4_ASAP7_75t_L g10800 ( 
.A(n_10385),
.B(n_709),
.Y(n_10800)
);

INVx1_ASAP7_75t_SL g10801 ( 
.A(n_10288),
.Y(n_10801)
);

OAI22xp5_ASAP7_75t_L g10802 ( 
.A1(n_10091),
.A2(n_712),
.B1(n_710),
.B2(n_711),
.Y(n_10802)
);

NOR2xp33_ASAP7_75t_SL g10803 ( 
.A(n_10169),
.B(n_711),
.Y(n_10803)
);

CKINVDCx5p33_ASAP7_75t_R g10804 ( 
.A(n_10114),
.Y(n_10804)
);

NOR3xp33_ASAP7_75t_L g10805 ( 
.A(n_10726),
.B(n_712),
.C(n_713),
.Y(n_10805)
);

CKINVDCx5p33_ASAP7_75t_R g10806 ( 
.A(n_10409),
.Y(n_10806)
);

NOR2xp33_ASAP7_75t_SL g10807 ( 
.A(n_10150),
.B(n_713),
.Y(n_10807)
);

INVx3_ASAP7_75t_L g10808 ( 
.A(n_10532),
.Y(n_10808)
);

INVx1_ASAP7_75t_L g10809 ( 
.A(n_10063),
.Y(n_10809)
);

BUFx4f_ASAP7_75t_L g10810 ( 
.A(n_10706),
.Y(n_10810)
);

AOI21xp5_ASAP7_75t_L g10811 ( 
.A1(n_10124),
.A2(n_714),
.B(n_715),
.Y(n_10811)
);

BUFx3_ASAP7_75t_L g10812 ( 
.A(n_10729),
.Y(n_10812)
);

AND2x2_ASAP7_75t_L g10813 ( 
.A(n_10089),
.B(n_714),
.Y(n_10813)
);

AOI21xp5_ASAP7_75t_L g10814 ( 
.A1(n_10172),
.A2(n_715),
.B(n_716),
.Y(n_10814)
);

NAND2xp5_ASAP7_75t_L g10815 ( 
.A(n_10213),
.B(n_716),
.Y(n_10815)
);

BUFx2_ASAP7_75t_L g10816 ( 
.A(n_10492),
.Y(n_10816)
);

BUFx6f_ASAP7_75t_L g10817 ( 
.A(n_10155),
.Y(n_10817)
);

INVx1_ASAP7_75t_L g10818 ( 
.A(n_10075),
.Y(n_10818)
);

NOR2xp33_ASAP7_75t_L g10819 ( 
.A(n_10269),
.B(n_717),
.Y(n_10819)
);

A2O1A1Ixp33_ASAP7_75t_L g10820 ( 
.A1(n_10090),
.A2(n_10070),
.B(n_10743),
.C(n_10686),
.Y(n_10820)
);

NAND2xp5_ASAP7_75t_L g10821 ( 
.A(n_10474),
.B(n_717),
.Y(n_10821)
);

OAI22xp5_ASAP7_75t_L g10822 ( 
.A1(n_10609),
.A2(n_720),
.B1(n_718),
.B2(n_719),
.Y(n_10822)
);

OAI22xp5_ASAP7_75t_L g10823 ( 
.A1(n_10687),
.A2(n_10099),
.B1(n_10237),
.B2(n_10343),
.Y(n_10823)
);

AOI22xp33_ASAP7_75t_L g10824 ( 
.A1(n_10734),
.A2(n_721),
.B1(n_718),
.B2(n_719),
.Y(n_10824)
);

AND2x2_ASAP7_75t_L g10825 ( 
.A(n_10478),
.B(n_10483),
.Y(n_10825)
);

BUFx8_ASAP7_75t_SL g10826 ( 
.A(n_10742),
.Y(n_10826)
);

OR2x2_ASAP7_75t_L g10827 ( 
.A(n_10473),
.B(n_721),
.Y(n_10827)
);

INVx1_ASAP7_75t_L g10828 ( 
.A(n_10076),
.Y(n_10828)
);

NOR2xp33_ASAP7_75t_L g10829 ( 
.A(n_10284),
.B(n_722),
.Y(n_10829)
);

OAI21x1_ASAP7_75t_L g10830 ( 
.A1(n_10787),
.A2(n_722),
.B(n_723),
.Y(n_10830)
);

OAI321xp33_ASAP7_75t_L g10831 ( 
.A1(n_10094),
.A2(n_726),
.A3(n_728),
.B1(n_723),
.B2(n_725),
.C(n_727),
.Y(n_10831)
);

INVx5_ASAP7_75t_L g10832 ( 
.A(n_10653),
.Y(n_10832)
);

INVx5_ASAP7_75t_L g10833 ( 
.A(n_10653),
.Y(n_10833)
);

INVx2_ASAP7_75t_L g10834 ( 
.A(n_10336),
.Y(n_10834)
);

NAND2xp5_ASAP7_75t_L g10835 ( 
.A(n_10084),
.B(n_727),
.Y(n_10835)
);

INVx1_ASAP7_75t_L g10836 ( 
.A(n_10079),
.Y(n_10836)
);

A2O1A1Ixp33_ASAP7_75t_L g10837 ( 
.A1(n_10667),
.A2(n_732),
.B(n_730),
.C(n_731),
.Y(n_10837)
);

A2O1A1Ixp33_ASAP7_75t_L g10838 ( 
.A1(n_10688),
.A2(n_733),
.B(n_730),
.C(n_732),
.Y(n_10838)
);

AOI21xp5_ASAP7_75t_L g10839 ( 
.A1(n_10157),
.A2(n_10699),
.B(n_10695),
.Y(n_10839)
);

OAI22xp5_ASAP7_75t_L g10840 ( 
.A1(n_10747),
.A2(n_10059),
.B1(n_10122),
.B2(n_10068),
.Y(n_10840)
);

INVx1_ASAP7_75t_L g10841 ( 
.A(n_10130),
.Y(n_10841)
);

AOI21xp5_ASAP7_75t_L g10842 ( 
.A1(n_10721),
.A2(n_733),
.B(n_735),
.Y(n_10842)
);

INVx1_ASAP7_75t_L g10843 ( 
.A(n_10146),
.Y(n_10843)
);

O2A1O1Ixp33_ASAP7_75t_L g10844 ( 
.A1(n_10622),
.A2(n_738),
.B(n_736),
.C(n_737),
.Y(n_10844)
);

A2O1A1Ixp33_ASAP7_75t_SL g10845 ( 
.A1(n_10078),
.A2(n_10058),
.B(n_10252),
.C(n_10170),
.Y(n_10845)
);

AOI21xp5_ASAP7_75t_L g10846 ( 
.A1(n_10765),
.A2(n_736),
.B(n_738),
.Y(n_10846)
);

O2A1O1Ixp33_ASAP7_75t_L g10847 ( 
.A1(n_10650),
.A2(n_741),
.B(n_739),
.C(n_740),
.Y(n_10847)
);

NAND2xp5_ASAP7_75t_L g10848 ( 
.A(n_10485),
.B(n_739),
.Y(n_10848)
);

OAI22xp5_ASAP7_75t_L g10849 ( 
.A1(n_10100),
.A2(n_744),
.B1(n_742),
.B2(n_743),
.Y(n_10849)
);

AOI21xp5_ASAP7_75t_L g10850 ( 
.A1(n_10054),
.A2(n_742),
.B(n_744),
.Y(n_10850)
);

NAND2xp5_ASAP7_75t_L g10851 ( 
.A(n_10709),
.B(n_745),
.Y(n_10851)
);

AOI21xp5_ASAP7_75t_L g10852 ( 
.A1(n_10663),
.A2(n_745),
.B(n_746),
.Y(n_10852)
);

INVx1_ASAP7_75t_L g10853 ( 
.A(n_10153),
.Y(n_10853)
);

NAND2xp5_ASAP7_75t_L g10854 ( 
.A(n_10715),
.B(n_746),
.Y(n_10854)
);

OAI22xp5_ASAP7_75t_L g10855 ( 
.A1(n_10299),
.A2(n_750),
.B1(n_748),
.B2(n_749),
.Y(n_10855)
);

NAND2xp5_ASAP7_75t_L g10856 ( 
.A(n_10756),
.B(n_748),
.Y(n_10856)
);

NOR2xp33_ASAP7_75t_SL g10857 ( 
.A(n_10137),
.B(n_749),
.Y(n_10857)
);

BUFx2_ASAP7_75t_L g10858 ( 
.A(n_10434),
.Y(n_10858)
);

INVx1_ASAP7_75t_L g10859 ( 
.A(n_10158),
.Y(n_10859)
);

AOI21x1_ASAP7_75t_L g10860 ( 
.A1(n_10120),
.A2(n_10112),
.B(n_10311),
.Y(n_10860)
);

OA22x2_ASAP7_75t_L g10861 ( 
.A1(n_10602),
.A2(n_752),
.B1(n_750),
.B2(n_751),
.Y(n_10861)
);

OR2x2_ASAP7_75t_L g10862 ( 
.A(n_10182),
.B(n_751),
.Y(n_10862)
);

INVxp67_ASAP7_75t_L g10863 ( 
.A(n_10505),
.Y(n_10863)
);

AOI21xp5_ASAP7_75t_L g10864 ( 
.A1(n_10731),
.A2(n_752),
.B(n_753),
.Y(n_10864)
);

INVx1_ASAP7_75t_SL g10865 ( 
.A(n_10579),
.Y(n_10865)
);

NAND2xp5_ASAP7_75t_L g10866 ( 
.A(n_10324),
.B(n_753),
.Y(n_10866)
);

O2A1O1Ixp33_ASAP7_75t_L g10867 ( 
.A1(n_10701),
.A2(n_756),
.B(n_754),
.C(n_755),
.Y(n_10867)
);

INVx2_ASAP7_75t_L g10868 ( 
.A(n_10344),
.Y(n_10868)
);

BUFx3_ASAP7_75t_L g10869 ( 
.A(n_10155),
.Y(n_10869)
);

A2O1A1Ixp33_ASAP7_75t_L g10870 ( 
.A1(n_10254),
.A2(n_757),
.B(n_755),
.C(n_756),
.Y(n_10870)
);

BUFx6f_ASAP7_75t_L g10871 ( 
.A(n_10171),
.Y(n_10871)
);

INVx1_ASAP7_75t_SL g10872 ( 
.A(n_10207),
.Y(n_10872)
);

AOI22xp33_ASAP7_75t_L g10873 ( 
.A1(n_10126),
.A2(n_759),
.B1(n_757),
.B2(n_758),
.Y(n_10873)
);

INVx2_ASAP7_75t_L g10874 ( 
.A(n_10466),
.Y(n_10874)
);

INVx2_ASAP7_75t_L g10875 ( 
.A(n_10398),
.Y(n_10875)
);

INVx1_ASAP7_75t_L g10876 ( 
.A(n_10184),
.Y(n_10876)
);

AOI21xp5_ASAP7_75t_L g10877 ( 
.A1(n_10773),
.A2(n_758),
.B(n_759),
.Y(n_10877)
);

AOI22x1_ASAP7_75t_L g10878 ( 
.A1(n_10095),
.A2(n_763),
.B1(n_760),
.B2(n_761),
.Y(n_10878)
);

BUFx3_ASAP7_75t_L g10879 ( 
.A(n_10171),
.Y(n_10879)
);

BUFx8_ASAP7_75t_SL g10880 ( 
.A(n_10341),
.Y(n_10880)
);

NOR2xp33_ASAP7_75t_L g10881 ( 
.A(n_10464),
.B(n_760),
.Y(n_10881)
);

NAND2xp5_ASAP7_75t_SL g10882 ( 
.A(n_10142),
.B(n_761),
.Y(n_10882)
);

AOI21xp5_ASAP7_75t_L g10883 ( 
.A1(n_10481),
.A2(n_763),
.B(n_764),
.Y(n_10883)
);

A2O1A1Ixp33_ASAP7_75t_L g10884 ( 
.A1(n_10345),
.A2(n_766),
.B(n_764),
.C(n_765),
.Y(n_10884)
);

NOR2xp33_ASAP7_75t_L g10885 ( 
.A(n_10419),
.B(n_765),
.Y(n_10885)
);

AOI22xp5_ASAP7_75t_L g10886 ( 
.A1(n_10108),
.A2(n_769),
.B1(n_767),
.B2(n_768),
.Y(n_10886)
);

O2A1O1Ixp5_ASAP7_75t_L g10887 ( 
.A1(n_10092),
.A2(n_770),
.B(n_767),
.C(n_768),
.Y(n_10887)
);

AOI21xp5_ASAP7_75t_L g10888 ( 
.A1(n_10365),
.A2(n_770),
.B(n_771),
.Y(n_10888)
);

INVx1_ASAP7_75t_L g10889 ( 
.A(n_10212),
.Y(n_10889)
);

INVx1_ASAP7_75t_L g10890 ( 
.A(n_10216),
.Y(n_10890)
);

BUFx2_ASAP7_75t_L g10891 ( 
.A(n_10499),
.Y(n_10891)
);

AO21x1_ASAP7_75t_L g10892 ( 
.A1(n_10261),
.A2(n_771),
.B(n_772),
.Y(n_10892)
);

NAND2xp5_ASAP7_75t_L g10893 ( 
.A(n_10148),
.B(n_10501),
.Y(n_10893)
);

NAND2xp5_ASAP7_75t_L g10894 ( 
.A(n_10439),
.B(n_772),
.Y(n_10894)
);

NAND2xp5_ASAP7_75t_SL g10895 ( 
.A(n_10588),
.B(n_773),
.Y(n_10895)
);

OAI21xp33_ASAP7_75t_L g10896 ( 
.A1(n_10767),
.A2(n_10166),
.B(n_10165),
.Y(n_10896)
);

AOI22xp33_ASAP7_75t_L g10897 ( 
.A1(n_10243),
.A2(n_10111),
.B1(n_10445),
.B2(n_10455),
.Y(n_10897)
);

NAND2xp5_ASAP7_75t_SL g10898 ( 
.A(n_10360),
.B(n_773),
.Y(n_10898)
);

OAI21xp33_ASAP7_75t_L g10899 ( 
.A1(n_10471),
.A2(n_774),
.B(n_775),
.Y(n_10899)
);

AOI21xp5_ASAP7_75t_L g10900 ( 
.A1(n_10749),
.A2(n_774),
.B(n_775),
.Y(n_10900)
);

OAI22xp5_ASAP7_75t_SL g10901 ( 
.A1(n_10425),
.A2(n_778),
.B1(n_776),
.B2(n_777),
.Y(n_10901)
);

A2O1A1Ixp33_ASAP7_75t_L g10902 ( 
.A1(n_10403),
.A2(n_778),
.B(n_776),
.C(n_777),
.Y(n_10902)
);

AND2x4_ASAP7_75t_L g10903 ( 
.A(n_10549),
.B(n_779),
.Y(n_10903)
);

INVx1_ASAP7_75t_L g10904 ( 
.A(n_10229),
.Y(n_10904)
);

A2O1A1Ixp33_ASAP7_75t_L g10905 ( 
.A1(n_10404),
.A2(n_781),
.B(n_779),
.C(n_780),
.Y(n_10905)
);

HB1xp67_ASAP7_75t_L g10906 ( 
.A(n_10258),
.Y(n_10906)
);

AND2x4_ASAP7_75t_L g10907 ( 
.A(n_10475),
.B(n_780),
.Y(n_10907)
);

NAND2xp5_ASAP7_75t_SL g10908 ( 
.A(n_10416),
.B(n_781),
.Y(n_10908)
);

INVxp67_ASAP7_75t_L g10909 ( 
.A(n_10594),
.Y(n_10909)
);

INVx2_ASAP7_75t_L g10910 ( 
.A(n_10279),
.Y(n_10910)
);

NAND2xp5_ASAP7_75t_L g10911 ( 
.A(n_10460),
.B(n_782),
.Y(n_10911)
);

INVx2_ASAP7_75t_L g10912 ( 
.A(n_10280),
.Y(n_10912)
);

OR2x2_ASAP7_75t_L g10913 ( 
.A(n_10322),
.B(n_782),
.Y(n_10913)
);

INVx1_ASAP7_75t_L g10914 ( 
.A(n_10330),
.Y(n_10914)
);

OAI22xp5_ASAP7_75t_L g10915 ( 
.A1(n_10559),
.A2(n_785),
.B1(n_783),
.B2(n_784),
.Y(n_10915)
);

CKINVDCx20_ASAP7_75t_R g10916 ( 
.A(n_10232),
.Y(n_10916)
);

OAI22xp5_ASAP7_75t_L g10917 ( 
.A1(n_10065),
.A2(n_785),
.B1(n_783),
.B2(n_784),
.Y(n_10917)
);

NAND2xp5_ASAP7_75t_L g10918 ( 
.A(n_10073),
.B(n_786),
.Y(n_10918)
);

NAND2xp5_ASAP7_75t_SL g10919 ( 
.A(n_10382),
.B(n_786),
.Y(n_10919)
);

HB1xp67_ASAP7_75t_L g10920 ( 
.A(n_10357),
.Y(n_10920)
);

OAI21x1_ASAP7_75t_L g10921 ( 
.A1(n_10067),
.A2(n_787),
.B(n_788),
.Y(n_10921)
);

O2A1O1Ixp33_ASAP7_75t_L g10922 ( 
.A1(n_10198),
.A2(n_790),
.B(n_788),
.C(n_789),
.Y(n_10922)
);

NOR2xp33_ASAP7_75t_L g10923 ( 
.A(n_10061),
.B(n_789),
.Y(n_10923)
);

INVx8_ASAP7_75t_L g10924 ( 
.A(n_10362),
.Y(n_10924)
);

NAND2xp5_ASAP7_75t_SL g10925 ( 
.A(n_10523),
.B(n_790),
.Y(n_10925)
);

O2A1O1Ixp5_ASAP7_75t_L g10926 ( 
.A1(n_10328),
.A2(n_793),
.B(n_791),
.C(n_792),
.Y(n_10926)
);

AOI21xp5_ASAP7_75t_L g10927 ( 
.A1(n_10220),
.A2(n_791),
.B(n_792),
.Y(n_10927)
);

BUFx2_ASAP7_75t_R g10928 ( 
.A(n_10522),
.Y(n_10928)
);

NAND2xp5_ASAP7_75t_L g10929 ( 
.A(n_10102),
.B(n_793),
.Y(n_10929)
);

INVx2_ASAP7_75t_L g10930 ( 
.A(n_10363),
.Y(n_10930)
);

NAND2xp5_ASAP7_75t_L g10931 ( 
.A(n_10106),
.B(n_794),
.Y(n_10931)
);

AOI21xp5_ASAP7_75t_L g10932 ( 
.A1(n_10220),
.A2(n_795),
.B(n_796),
.Y(n_10932)
);

INVx2_ASAP7_75t_L g10933 ( 
.A(n_10372),
.Y(n_10933)
);

INVx3_ASAP7_75t_L g10934 ( 
.A(n_10566),
.Y(n_10934)
);

NAND2xp5_ASAP7_75t_L g10935 ( 
.A(n_10138),
.B(n_796),
.Y(n_10935)
);

OAI21xp33_ASAP7_75t_SL g10936 ( 
.A1(n_10208),
.A2(n_797),
.B(n_798),
.Y(n_10936)
);

BUFx6f_ASAP7_75t_L g10937 ( 
.A(n_10391),
.Y(n_10937)
);

O2A1O1Ixp33_ASAP7_75t_L g10938 ( 
.A1(n_10221),
.A2(n_801),
.B(n_799),
.C(n_800),
.Y(n_10938)
);

NAND2xp5_ASAP7_75t_SL g10939 ( 
.A(n_10508),
.B(n_799),
.Y(n_10939)
);

BUFx6f_ASAP7_75t_L g10940 ( 
.A(n_10391),
.Y(n_10940)
);

INVx11_ASAP7_75t_L g10941 ( 
.A(n_10388),
.Y(n_10941)
);

INVx1_ASAP7_75t_L g10942 ( 
.A(n_10394),
.Y(n_10942)
);

AOI21xp5_ASAP7_75t_L g10943 ( 
.A1(n_10544),
.A2(n_800),
.B(n_801),
.Y(n_10943)
);

HB1xp67_ASAP7_75t_L g10944 ( 
.A(n_10396),
.Y(n_10944)
);

NAND3xp33_ASAP7_75t_L g10945 ( 
.A(n_10088),
.B(n_802),
.C(n_803),
.Y(n_10945)
);

NAND2xp5_ASAP7_75t_SL g10946 ( 
.A(n_10262),
.B(n_802),
.Y(n_10946)
);

AOI21xp5_ASAP7_75t_L g10947 ( 
.A1(n_10418),
.A2(n_803),
.B(n_804),
.Y(n_10947)
);

AOI21xp5_ASAP7_75t_L g10948 ( 
.A1(n_10105),
.A2(n_805),
.B(n_806),
.Y(n_10948)
);

INVxp33_ASAP7_75t_SL g10949 ( 
.A(n_10600),
.Y(n_10949)
);

OAI21x1_ASAP7_75t_L g10950 ( 
.A1(n_10696),
.A2(n_805),
.B(n_806),
.Y(n_10950)
);

AOI22xp5_ASAP7_75t_L g10951 ( 
.A1(n_10589),
.A2(n_809),
.B1(n_807),
.B2(n_808),
.Y(n_10951)
);

O2A1O1Ixp33_ASAP7_75t_L g10952 ( 
.A1(n_10338),
.A2(n_810),
.B(n_807),
.C(n_809),
.Y(n_10952)
);

HB1xp67_ASAP7_75t_L g10953 ( 
.A(n_10607),
.Y(n_10953)
);

INVx1_ASAP7_75t_L g10954 ( 
.A(n_10611),
.Y(n_10954)
);

AOI21xp5_ASAP7_75t_L g10955 ( 
.A1(n_10110),
.A2(n_810),
.B(n_811),
.Y(n_10955)
);

AND2x2_ASAP7_75t_L g10956 ( 
.A(n_10552),
.B(n_811),
.Y(n_10956)
);

NAND2xp5_ASAP7_75t_L g10957 ( 
.A(n_10140),
.B(n_812),
.Y(n_10957)
);

A2O1A1Ixp33_ASAP7_75t_L g10958 ( 
.A1(n_10083),
.A2(n_814),
.B(n_812),
.C(n_813),
.Y(n_10958)
);

NOR2xp33_ASAP7_75t_SL g10959 ( 
.A(n_10514),
.B(n_813),
.Y(n_10959)
);

OR2x6_ASAP7_75t_L g10960 ( 
.A(n_10316),
.B(n_814),
.Y(n_10960)
);

OAI21xp5_ASAP7_75t_L g10961 ( 
.A1(n_10271),
.A2(n_815),
.B(n_816),
.Y(n_10961)
);

NAND2xp5_ASAP7_75t_L g10962 ( 
.A(n_10151),
.B(n_815),
.Y(n_10962)
);

AO31x2_ASAP7_75t_L g10963 ( 
.A1(n_10048),
.A2(n_819),
.A3(n_817),
.B(n_818),
.Y(n_10963)
);

NAND2xp5_ASAP7_75t_SL g10964 ( 
.A(n_10118),
.B(n_817),
.Y(n_10964)
);

AOI21x1_ASAP7_75t_L g10965 ( 
.A1(n_10086),
.A2(n_818),
.B(n_819),
.Y(n_10965)
);

INVx2_ASAP7_75t_L g10966 ( 
.A(n_10617),
.Y(n_10966)
);

NOR2xp67_ASAP7_75t_L g10967 ( 
.A(n_10567),
.B(n_820),
.Y(n_10967)
);

AND2x2_ASAP7_75t_L g10968 ( 
.A(n_10513),
.B(n_820),
.Y(n_10968)
);

INVx6_ASAP7_75t_SL g10969 ( 
.A(n_10378),
.Y(n_10969)
);

INVx1_ASAP7_75t_L g10970 ( 
.A(n_10647),
.Y(n_10970)
);

BUFx6f_ASAP7_75t_L g10971 ( 
.A(n_10186),
.Y(n_10971)
);

OAI22xp5_ASAP7_75t_L g10972 ( 
.A1(n_10371),
.A2(n_824),
.B1(n_822),
.B2(n_823),
.Y(n_10972)
);

NOR2xp33_ASAP7_75t_R g10973 ( 
.A(n_10454),
.B(n_823),
.Y(n_10973)
);

A2O1A1Ixp33_ASAP7_75t_L g10974 ( 
.A1(n_10123),
.A2(n_826),
.B(n_824),
.C(n_825),
.Y(n_10974)
);

INVx2_ASAP7_75t_L g10975 ( 
.A(n_10656),
.Y(n_10975)
);

BUFx12f_ASAP7_75t_L g10976 ( 
.A(n_10582),
.Y(n_10976)
);

NAND2xp5_ASAP7_75t_SL g10977 ( 
.A(n_10131),
.B(n_825),
.Y(n_10977)
);

NOR2xp33_ASAP7_75t_L g10978 ( 
.A(n_10066),
.B(n_826),
.Y(n_10978)
);

INVx1_ASAP7_75t_L g10979 ( 
.A(n_10659),
.Y(n_10979)
);

OAI22xp5_ASAP7_75t_SL g10980 ( 
.A1(n_10527),
.A2(n_829),
.B1(n_827),
.B2(n_828),
.Y(n_10980)
);

OAI21xp5_ASAP7_75t_L g10981 ( 
.A1(n_10274),
.A2(n_827),
.B(n_829),
.Y(n_10981)
);

OAI22xp5_ASAP7_75t_L g10982 ( 
.A1(n_10428),
.A2(n_832),
.B1(n_830),
.B2(n_831),
.Y(n_10982)
);

INVxp67_ASAP7_75t_SL g10983 ( 
.A(n_10410),
.Y(n_10983)
);

A2O1A1Ixp33_ASAP7_75t_SL g10984 ( 
.A1(n_10310),
.A2(n_832),
.B(n_830),
.C(n_831),
.Y(n_10984)
);

AOI21xp5_ASAP7_75t_L g10985 ( 
.A1(n_10610),
.A2(n_833),
.B(n_834),
.Y(n_10985)
);

AOI21xp5_ASAP7_75t_L g10986 ( 
.A1(n_10624),
.A2(n_10673),
.B(n_10642),
.Y(n_10986)
);

INVx1_ASAP7_75t_L g10987 ( 
.A(n_10670),
.Y(n_10987)
);

INVx1_ASAP7_75t_SL g10988 ( 
.A(n_10540),
.Y(n_10988)
);

NOR2xp33_ASAP7_75t_L g10989 ( 
.A(n_10488),
.B(n_834),
.Y(n_10989)
);

AOI21xp33_ASAP7_75t_L g10990 ( 
.A1(n_10315),
.A2(n_835),
.B(n_836),
.Y(n_10990)
);

INVx2_ASAP7_75t_L g10991 ( 
.A(n_10698),
.Y(n_10991)
);

AOI21xp5_ASAP7_75t_L g10992 ( 
.A1(n_10674),
.A2(n_835),
.B(n_836),
.Y(n_10992)
);

AND2x2_ASAP7_75t_L g10993 ( 
.A(n_10535),
.B(n_837),
.Y(n_10993)
);

NOR3xp33_ASAP7_75t_SL g10994 ( 
.A(n_10161),
.B(n_837),
.C(n_838),
.Y(n_10994)
);

NOR2xp33_ASAP7_75t_SL g10995 ( 
.A(n_10087),
.B(n_838),
.Y(n_10995)
);

INVx2_ASAP7_75t_L g10996 ( 
.A(n_10702),
.Y(n_10996)
);

OAI22xp5_ASAP7_75t_L g10997 ( 
.A1(n_10069),
.A2(n_841),
.B1(n_839),
.B2(n_840),
.Y(n_10997)
);

OAI22xp5_ASAP7_75t_L g10998 ( 
.A1(n_10190),
.A2(n_843),
.B1(n_840),
.B2(n_842),
.Y(n_10998)
);

CKINVDCx6p67_ASAP7_75t_R g10999 ( 
.A(n_10606),
.Y(n_10999)
);

INVx1_ASAP7_75t_L g11000 ( 
.A(n_10722),
.Y(n_11000)
);

AND2x2_ASAP7_75t_L g11001 ( 
.A(n_10538),
.B(n_842),
.Y(n_11001)
);

O2A1O1Ixp5_ASAP7_75t_L g11002 ( 
.A1(n_10135),
.A2(n_846),
.B(n_844),
.C(n_845),
.Y(n_11002)
);

NAND2xp5_ASAP7_75t_SL g11003 ( 
.A(n_10049),
.B(n_10051),
.Y(n_11003)
);

NAND2xp5_ASAP7_75t_SL g11004 ( 
.A(n_10614),
.B(n_10618),
.Y(n_11004)
);

OAI22xp5_ASAP7_75t_L g11005 ( 
.A1(n_10422),
.A2(n_847),
.B1(n_845),
.B2(n_846),
.Y(n_11005)
);

NAND2xp5_ASAP7_75t_L g11006 ( 
.A(n_10154),
.B(n_847),
.Y(n_11006)
);

INVx2_ASAP7_75t_L g11007 ( 
.A(n_10733),
.Y(n_11007)
);

AOI21xp5_ASAP7_75t_L g11008 ( 
.A1(n_10675),
.A2(n_848),
.B(n_849),
.Y(n_11008)
);

AND2x4_ASAP7_75t_L g11009 ( 
.A(n_10441),
.B(n_848),
.Y(n_11009)
);

AOI21xp5_ASAP7_75t_L g11010 ( 
.A1(n_10685),
.A2(n_10712),
.B(n_10704),
.Y(n_11010)
);

AOI21xp5_ASAP7_75t_L g11011 ( 
.A1(n_10759),
.A2(n_849),
.B(n_850),
.Y(n_11011)
);

INVx2_ASAP7_75t_L g11012 ( 
.A(n_10736),
.Y(n_11012)
);

AOI21xp5_ASAP7_75t_L g11013 ( 
.A1(n_10085),
.A2(n_850),
.B(n_851),
.Y(n_11013)
);

BUFx3_ASAP7_75t_L g11014 ( 
.A(n_10461),
.Y(n_11014)
);

INVx2_ASAP7_75t_L g11015 ( 
.A(n_10737),
.Y(n_11015)
);

NAND2xp5_ASAP7_75t_L g11016 ( 
.A(n_10163),
.B(n_851),
.Y(n_11016)
);

AOI21xp5_ASAP7_75t_L g11017 ( 
.A1(n_10275),
.A2(n_852),
.B(n_853),
.Y(n_11017)
);

O2A1O1Ixp5_ASAP7_75t_L g11018 ( 
.A1(n_10319),
.A2(n_855),
.B(n_853),
.C(n_854),
.Y(n_11018)
);

NOR2xp33_ASAP7_75t_L g11019 ( 
.A(n_10050),
.B(n_854),
.Y(n_11019)
);

BUFx2_ASAP7_75t_L g11020 ( 
.A(n_10533),
.Y(n_11020)
);

INVx2_ASAP7_75t_L g11021 ( 
.A(n_10746),
.Y(n_11021)
);

INVx1_ASAP7_75t_L g11022 ( 
.A(n_10789),
.Y(n_11022)
);

AND2x4_ASAP7_75t_L g11023 ( 
.A(n_10164),
.B(n_855),
.Y(n_11023)
);

AOI22xp33_ASAP7_75t_SL g11024 ( 
.A1(n_10313),
.A2(n_858),
.B1(n_856),
.B2(n_857),
.Y(n_11024)
);

AOI21xp5_ASAP7_75t_L g11025 ( 
.A1(n_10259),
.A2(n_856),
.B(n_858),
.Y(n_11025)
);

AND2x2_ASAP7_75t_SL g11026 ( 
.A(n_10525),
.B(n_859),
.Y(n_11026)
);

BUFx6f_ASAP7_75t_L g11027 ( 
.A(n_10186),
.Y(n_11027)
);

CKINVDCx5p33_ASAP7_75t_R g11028 ( 
.A(n_10055),
.Y(n_11028)
);

OAI22xp5_ASAP7_75t_L g11029 ( 
.A1(n_10294),
.A2(n_861),
.B1(n_859),
.B2(n_860),
.Y(n_11029)
);

AOI21xp5_ASAP7_75t_L g11030 ( 
.A1(n_10317),
.A2(n_860),
.B(n_861),
.Y(n_11030)
);

AND2x4_ASAP7_75t_L g11031 ( 
.A(n_10230),
.B(n_862),
.Y(n_11031)
);

NAND3xp33_ASAP7_75t_SL g11032 ( 
.A(n_10489),
.B(n_863),
.C(n_865),
.Y(n_11032)
);

NAND2xp5_ASAP7_75t_L g11033 ( 
.A(n_10231),
.B(n_863),
.Y(n_11033)
);

NAND2xp5_ASAP7_75t_SL g11034 ( 
.A(n_10621),
.B(n_865),
.Y(n_11034)
);

AND2x4_ASAP7_75t_L g11035 ( 
.A(n_10238),
.B(n_866),
.Y(n_11035)
);

BUFx6f_ASAP7_75t_L g11036 ( 
.A(n_10186),
.Y(n_11036)
);

INVx2_ASAP7_75t_L g11037 ( 
.A(n_10246),
.Y(n_11037)
);

NOR2xp33_ASAP7_75t_R g11038 ( 
.A(n_10423),
.B(n_10777),
.Y(n_11038)
);

NAND2xp5_ASAP7_75t_L g11039 ( 
.A(n_10282),
.B(n_866),
.Y(n_11039)
);

AND2x2_ASAP7_75t_L g11040 ( 
.A(n_10145),
.B(n_10541),
.Y(n_11040)
);

AND3x1_ASAP7_75t_SL g11041 ( 
.A(n_10536),
.B(n_867),
.C(n_868),
.Y(n_11041)
);

NOR2xp33_ASAP7_75t_R g11042 ( 
.A(n_10119),
.B(n_867),
.Y(n_11042)
);

INVx1_ASAP7_75t_L g11043 ( 
.A(n_10289),
.Y(n_11043)
);

OAI21xp5_ASAP7_75t_L g11044 ( 
.A1(n_10215),
.A2(n_869),
.B(n_870),
.Y(n_11044)
);

NOR2xp33_ASAP7_75t_L g11045 ( 
.A(n_10668),
.B(n_10691),
.Y(n_11045)
);

NOR2xp33_ASAP7_75t_SL g11046 ( 
.A(n_10115),
.B(n_869),
.Y(n_11046)
);

BUFx6f_ASAP7_75t_L g11047 ( 
.A(n_10227),
.Y(n_11047)
);

AND2x2_ASAP7_75t_SL g11048 ( 
.A(n_10462),
.B(n_870),
.Y(n_11048)
);

INVx3_ASAP7_75t_L g11049 ( 
.A(n_10227),
.Y(n_11049)
);

BUFx2_ASAP7_75t_L g11050 ( 
.A(n_10133),
.Y(n_11050)
);

INVx2_ASAP7_75t_L g11051 ( 
.A(n_10616),
.Y(n_11051)
);

INVxp67_ASAP7_75t_L g11052 ( 
.A(n_10109),
.Y(n_11052)
);

NOR2xp33_ASAP7_75t_L g11053 ( 
.A(n_10531),
.B(n_871),
.Y(n_11053)
);

NAND2xp5_ASAP7_75t_L g11054 ( 
.A(n_10625),
.B(n_871),
.Y(n_11054)
);

AND2x6_ASAP7_75t_L g11055 ( 
.A(n_10245),
.B(n_872),
.Y(n_11055)
);

HB1xp67_ASAP7_75t_L g11056 ( 
.A(n_10634),
.Y(n_11056)
);

INVx1_ASAP7_75t_L g11057 ( 
.A(n_10640),
.Y(n_11057)
);

AOI22xp5_ASAP7_75t_L g11058 ( 
.A1(n_10219),
.A2(n_874),
.B1(n_872),
.B2(n_873),
.Y(n_11058)
);

AOI21xp5_ASAP7_75t_L g11059 ( 
.A1(n_10354),
.A2(n_873),
.B(n_874),
.Y(n_11059)
);

OAI21x1_ASAP7_75t_L g11060 ( 
.A1(n_10098),
.A2(n_875),
.B(n_876),
.Y(n_11060)
);

INVx2_ASAP7_75t_L g11061 ( 
.A(n_10676),
.Y(n_11061)
);

OAI22xp5_ASAP7_75t_L g11062 ( 
.A1(n_10309),
.A2(n_10406),
.B1(n_10187),
.B2(n_10521),
.Y(n_11062)
);

INVx1_ASAP7_75t_L g11063 ( 
.A(n_10693),
.Y(n_11063)
);

BUFx6f_ASAP7_75t_L g11064 ( 
.A(n_10227),
.Y(n_11064)
);

NOR2xp33_ASAP7_75t_L g11065 ( 
.A(n_10128),
.B(n_875),
.Y(n_11065)
);

AOI21xp5_ASAP7_75t_L g11066 ( 
.A1(n_10386),
.A2(n_876),
.B(n_877),
.Y(n_11066)
);

BUFx2_ASAP7_75t_L g11067 ( 
.A(n_10561),
.Y(n_11067)
);

INVx2_ASAP7_75t_L g11068 ( 
.A(n_10717),
.Y(n_11068)
);

NAND2xp5_ASAP7_75t_SL g11069 ( 
.A(n_10623),
.B(n_877),
.Y(n_11069)
);

BUFx6f_ASAP7_75t_L g11070 ( 
.A(n_10247),
.Y(n_11070)
);

AND2x2_ASAP7_75t_L g11071 ( 
.A(n_10074),
.B(n_878),
.Y(n_11071)
);

BUFx6f_ASAP7_75t_L g11072 ( 
.A(n_10247),
.Y(n_11072)
);

INVxp33_ASAP7_75t_L g11073 ( 
.A(n_10247),
.Y(n_11073)
);

A2O1A1Ixp33_ASAP7_75t_L g11074 ( 
.A1(n_10141),
.A2(n_881),
.B(n_879),
.C(n_880),
.Y(n_11074)
);

OA22x2_ASAP7_75t_L g11075 ( 
.A1(n_10494),
.A2(n_883),
.B1(n_879),
.B2(n_882),
.Y(n_11075)
);

OR2x6_ASAP7_75t_L g11076 ( 
.A(n_10093),
.B(n_882),
.Y(n_11076)
);

BUFx6f_ASAP7_75t_L g11077 ( 
.A(n_10437),
.Y(n_11077)
);

AOI21xp5_ASAP7_75t_L g11078 ( 
.A1(n_10408),
.A2(n_884),
.B(n_885),
.Y(n_11078)
);

NOR2xp33_ASAP7_75t_SL g11079 ( 
.A(n_10752),
.B(n_884),
.Y(n_11079)
);

NOR2xp33_ASAP7_75t_SL g11080 ( 
.A(n_10593),
.B(n_885),
.Y(n_11080)
);

CKINVDCx5p33_ASAP7_75t_R g11081 ( 
.A(n_10320),
.Y(n_11081)
);

BUFx12f_ASAP7_75t_L g11082 ( 
.A(n_10453),
.Y(n_11082)
);

AOI21xp5_ASAP7_75t_L g11083 ( 
.A1(n_10046),
.A2(n_886),
.B(n_887),
.Y(n_11083)
);

NOR3xp33_ASAP7_75t_SL g11084 ( 
.A(n_10199),
.B(n_888),
.C(n_889),
.Y(n_11084)
);

INVx1_ASAP7_75t_L g11085 ( 
.A(n_10755),
.Y(n_11085)
);

NAND2xp5_ASAP7_75t_SL g11086 ( 
.A(n_10626),
.B(n_888),
.Y(n_11086)
);

AOI21xp5_ASAP7_75t_L g11087 ( 
.A1(n_10613),
.A2(n_890),
.B(n_891),
.Y(n_11087)
);

BUFx6f_ASAP7_75t_L g11088 ( 
.A(n_10437),
.Y(n_11088)
);

AND2x2_ASAP7_75t_L g11089 ( 
.A(n_10727),
.B(n_891),
.Y(n_11089)
);

NAND2xp5_ASAP7_75t_SL g11090 ( 
.A(n_10631),
.B(n_892),
.Y(n_11090)
);

O2A1O1Ixp5_ASAP7_75t_L g11091 ( 
.A1(n_10081),
.A2(n_10361),
.B(n_10517),
.C(n_10497),
.Y(n_11091)
);

OR2x2_ASAP7_75t_L g11092 ( 
.A(n_10633),
.B(n_892),
.Y(n_11092)
);

O2A1O1Ixp33_ASAP7_75t_L g11093 ( 
.A1(n_10248),
.A2(n_895),
.B(n_893),
.C(n_894),
.Y(n_11093)
);

BUFx6f_ASAP7_75t_L g11094 ( 
.A(n_10437),
.Y(n_11094)
);

NAND2xp5_ASAP7_75t_L g11095 ( 
.A(n_10786),
.B(n_893),
.Y(n_11095)
);

INVx1_ASAP7_75t_L g11096 ( 
.A(n_10397),
.Y(n_11096)
);

INVx1_ASAP7_75t_L g11097 ( 
.A(n_10427),
.Y(n_11097)
);

NAND2xp5_ASAP7_75t_SL g11098 ( 
.A(n_10635),
.B(n_894),
.Y(n_11098)
);

NAND2xp5_ASAP7_75t_L g11099 ( 
.A(n_10463),
.B(n_895),
.Y(n_11099)
);

BUFx12f_ASAP7_75t_L g11100 ( 
.A(n_10453),
.Y(n_11100)
);

NOR2xp33_ASAP7_75t_L g11101 ( 
.A(n_10564),
.B(n_896),
.Y(n_11101)
);

OAI22xp5_ASAP7_75t_L g11102 ( 
.A1(n_10528),
.A2(n_898),
.B1(n_896),
.B2(n_897),
.Y(n_11102)
);

AOI22xp5_ASAP7_75t_L g11103 ( 
.A1(n_10424),
.A2(n_899),
.B1(n_897),
.B2(n_898),
.Y(n_11103)
);

NAND2xp5_ASAP7_75t_SL g11104 ( 
.A(n_10646),
.B(n_900),
.Y(n_11104)
);

OAI22x1_ASAP7_75t_L g11105 ( 
.A1(n_10224),
.A2(n_902),
.B1(n_900),
.B2(n_901),
.Y(n_11105)
);

A2O1A1Ixp33_ASAP7_75t_L g11106 ( 
.A1(n_10268),
.A2(n_903),
.B(n_901),
.C(n_902),
.Y(n_11106)
);

BUFx6f_ASAP7_75t_L g11107 ( 
.A(n_10097),
.Y(n_11107)
);

OAI22xp5_ASAP7_75t_L g11108 ( 
.A1(n_10250),
.A2(n_905),
.B1(n_903),
.B2(n_904),
.Y(n_11108)
);

INVx1_ASAP7_75t_L g11109 ( 
.A(n_10325),
.Y(n_11109)
);

INVx2_ASAP7_75t_L g11110 ( 
.A(n_10450),
.Y(n_11110)
);

AOI22xp5_ASAP7_75t_L g11111 ( 
.A1(n_10373),
.A2(n_906),
.B1(n_904),
.B2(n_905),
.Y(n_11111)
);

AND2x2_ASAP7_75t_L g11112 ( 
.A(n_10762),
.B(n_906),
.Y(n_11112)
);

NOR2xp33_ASAP7_75t_L g11113 ( 
.A(n_10057),
.B(n_907),
.Y(n_11113)
);

A2O1A1Ixp33_ASAP7_75t_L g11114 ( 
.A1(n_10448),
.A2(n_911),
.B(n_908),
.C(n_910),
.Y(n_11114)
);

AND2x2_ASAP7_75t_L g11115 ( 
.A(n_10772),
.B(n_910),
.Y(n_11115)
);

NAND2xp5_ASAP7_75t_SL g11116 ( 
.A(n_10648),
.B(n_911),
.Y(n_11116)
);

OAI22xp5_ASAP7_75t_L g11117 ( 
.A1(n_10459),
.A2(n_914),
.B1(n_912),
.B2(n_913),
.Y(n_11117)
);

OAI22xp5_ASAP7_75t_L g11118 ( 
.A1(n_10554),
.A2(n_914),
.B1(n_912),
.B2(n_913),
.Y(n_11118)
);

OAI21xp33_ASAP7_75t_L g11119 ( 
.A1(n_10493),
.A2(n_915),
.B(n_916),
.Y(n_11119)
);

NOR2xp33_ASAP7_75t_L g11120 ( 
.A(n_10348),
.B(n_915),
.Y(n_11120)
);

NAND2xp5_ASAP7_75t_SL g11121 ( 
.A(n_10666),
.B(n_917),
.Y(n_11121)
);

INVx2_ASAP7_75t_L g11122 ( 
.A(n_10781),
.Y(n_11122)
);

AOI21xp5_ASAP7_75t_L g11123 ( 
.A1(n_10615),
.A2(n_10628),
.B(n_10620),
.Y(n_11123)
);

O2A1O1Ixp5_ASAP7_75t_L g11124 ( 
.A1(n_10077),
.A2(n_920),
.B(n_918),
.C(n_919),
.Y(n_11124)
);

AND2x4_ASAP7_75t_L g11125 ( 
.A(n_10595),
.B(n_918),
.Y(n_11125)
);

A2O1A1Ixp33_ASAP7_75t_L g11126 ( 
.A1(n_10273),
.A2(n_922),
.B(n_920),
.C(n_921),
.Y(n_11126)
);

AND2x2_ASAP7_75t_SL g11127 ( 
.A(n_10577),
.B(n_921),
.Y(n_11127)
);

AND2x2_ASAP7_75t_L g11128 ( 
.A(n_10178),
.B(n_923),
.Y(n_11128)
);

O2A1O1Ixp33_ASAP7_75t_L g11129 ( 
.A1(n_10384),
.A2(n_925),
.B(n_923),
.C(n_924),
.Y(n_11129)
);

NOR3xp33_ASAP7_75t_L g11130 ( 
.A(n_10228),
.B(n_924),
.C(n_926),
.Y(n_11130)
);

NAND2xp5_ASAP7_75t_SL g11131 ( 
.A(n_10677),
.B(n_926),
.Y(n_11131)
);

HB1xp67_ASAP7_75t_L g11132 ( 
.A(n_10679),
.Y(n_11132)
);

AOI21x1_ASAP7_75t_L g11133 ( 
.A1(n_10761),
.A2(n_927),
.B(n_928),
.Y(n_11133)
);

O2A1O1Ixp33_ASAP7_75t_L g11134 ( 
.A1(n_10392),
.A2(n_929),
.B(n_927),
.C(n_928),
.Y(n_11134)
);

AOI21xp5_ASAP7_75t_L g11135 ( 
.A1(n_10629),
.A2(n_929),
.B(n_930),
.Y(n_11135)
);

INVx1_ASAP7_75t_L g11136 ( 
.A(n_10277),
.Y(n_11136)
);

NAND2xp5_ASAP7_75t_L g11137 ( 
.A(n_10680),
.B(n_931),
.Y(n_11137)
);

AOI21xp5_ASAP7_75t_L g11138 ( 
.A1(n_10637),
.A2(n_931),
.B(n_932),
.Y(n_11138)
);

AOI22xp5_ASAP7_75t_L g11139 ( 
.A1(n_10402),
.A2(n_10380),
.B1(n_10524),
.B2(n_10056),
.Y(n_11139)
);

NAND2xp5_ASAP7_75t_SL g11140 ( 
.A(n_10690),
.B(n_933),
.Y(n_11140)
);

O2A1O1Ixp33_ASAP7_75t_L g11141 ( 
.A1(n_10395),
.A2(n_10415),
.B(n_10490),
.C(n_10547),
.Y(n_11141)
);

A2O1A1Ixp33_ASAP7_75t_L g11142 ( 
.A1(n_10539),
.A2(n_935),
.B(n_933),
.C(n_934),
.Y(n_11142)
);

OAI22xp5_ASAP7_75t_L g11143 ( 
.A1(n_10263),
.A2(n_10266),
.B1(n_10400),
.B2(n_10323),
.Y(n_11143)
);

OAI22xp5_ASAP7_75t_SL g11144 ( 
.A1(n_10272),
.A2(n_937),
.B1(n_935),
.B2(n_936),
.Y(n_11144)
);

CKINVDCx5p33_ASAP7_75t_R g11145 ( 
.A(n_10097),
.Y(n_11145)
);

NAND2xp5_ASAP7_75t_L g11146 ( 
.A(n_10707),
.B(n_10711),
.Y(n_11146)
);

BUFx6f_ASAP7_75t_L g11147 ( 
.A(n_10662),
.Y(n_11147)
);

NAND3xp33_ASAP7_75t_L g11148 ( 
.A(n_10267),
.B(n_938),
.C(n_939),
.Y(n_11148)
);

INVx3_ASAP7_75t_L g11149 ( 
.A(n_10222),
.Y(n_11149)
);

NAND2xp5_ASAP7_75t_L g11150 ( 
.A(n_10716),
.B(n_939),
.Y(n_11150)
);

NAND2xp5_ASAP7_75t_L g11151 ( 
.A(n_10723),
.B(n_940),
.Y(n_11151)
);

HB1xp67_ASAP7_75t_L g11152 ( 
.A(n_10750),
.Y(n_11152)
);

AOI21xp5_ASAP7_75t_L g11153 ( 
.A1(n_10651),
.A2(n_940),
.B(n_941),
.Y(n_11153)
);

A2O1A1Ixp33_ASAP7_75t_L g11154 ( 
.A1(n_10652),
.A2(n_943),
.B(n_941),
.C(n_942),
.Y(n_11154)
);

NAND2xp5_ASAP7_75t_L g11155 ( 
.A(n_10758),
.B(n_942),
.Y(n_11155)
);

A2O1A1Ixp33_ASAP7_75t_L g11156 ( 
.A1(n_10655),
.A2(n_945),
.B(n_943),
.C(n_944),
.Y(n_11156)
);

O2A1O1Ixp33_ASAP7_75t_L g11157 ( 
.A1(n_10627),
.A2(n_947),
.B(n_945),
.C(n_946),
.Y(n_11157)
);

BUFx6f_ASAP7_75t_SL g11158 ( 
.A(n_10349),
.Y(n_11158)
);

NAND2xp5_ASAP7_75t_L g11159 ( 
.A(n_10760),
.B(n_946),
.Y(n_11159)
);

NAND2xp5_ASAP7_75t_L g11160 ( 
.A(n_10763),
.B(n_948),
.Y(n_11160)
);

INVx2_ASAP7_75t_L g11161 ( 
.A(n_10781),
.Y(n_11161)
);

O2A1O1Ixp33_ASAP7_75t_L g11162 ( 
.A1(n_10641),
.A2(n_950),
.B(n_948),
.C(n_949),
.Y(n_11162)
);

AOI21xp5_ASAP7_75t_L g11163 ( 
.A1(n_10660),
.A2(n_950),
.B(n_951),
.Y(n_11163)
);

OAI22xp5_ASAP7_75t_L g11164 ( 
.A1(n_10383),
.A2(n_954),
.B1(n_952),
.B2(n_953),
.Y(n_11164)
);

O2A1O1Ixp33_ASAP7_75t_SL g11165 ( 
.A1(n_10632),
.A2(n_955),
.B(n_952),
.C(n_953),
.Y(n_11165)
);

AOI21xp5_ASAP7_75t_L g11166 ( 
.A1(n_10661),
.A2(n_955),
.B(n_956),
.Y(n_11166)
);

NAND2xp5_ASAP7_75t_L g11167 ( 
.A(n_10766),
.B(n_956),
.Y(n_11167)
);

AND2x6_ASAP7_75t_L g11168 ( 
.A(n_10364),
.B(n_957),
.Y(n_11168)
);

NOR2xp33_ASAP7_75t_L g11169 ( 
.A(n_10210),
.B(n_957),
.Y(n_11169)
);

A2O1A1Ixp33_ASAP7_75t_L g11170 ( 
.A1(n_10665),
.A2(n_960),
.B(n_958),
.C(n_959),
.Y(n_11170)
);

AOI22xp5_ASAP7_75t_L g11171 ( 
.A1(n_10644),
.A2(n_960),
.B1(n_958),
.B2(n_959),
.Y(n_11171)
);

INVx6_ASAP7_75t_L g11172 ( 
.A(n_10662),
.Y(n_11172)
);

NAND2xp5_ASAP7_75t_L g11173 ( 
.A(n_10771),
.B(n_961),
.Y(n_11173)
);

NAND2xp5_ASAP7_75t_L g11174 ( 
.A(n_10778),
.B(n_961),
.Y(n_11174)
);

INVx1_ASAP7_75t_L g11175 ( 
.A(n_10277),
.Y(n_11175)
);

AOI21xp5_ASAP7_75t_L g11176 ( 
.A1(n_10669),
.A2(n_962),
.B(n_963),
.Y(n_11176)
);

BUFx2_ASAP7_75t_SL g11177 ( 
.A(n_10585),
.Y(n_11177)
);

INVx2_ASAP7_75t_L g11178 ( 
.A(n_10781),
.Y(n_11178)
);

INVx1_ASAP7_75t_L g11179 ( 
.A(n_10781),
.Y(n_11179)
);

AOI21xp5_ASAP7_75t_L g11180 ( 
.A1(n_10671),
.A2(n_962),
.B(n_964),
.Y(n_11180)
);

AND2x2_ASAP7_75t_L g11181 ( 
.A(n_10291),
.B(n_965),
.Y(n_11181)
);

CKINVDCx5p33_ASAP7_75t_R g11182 ( 
.A(n_10682),
.Y(n_11182)
);

NAND2xp5_ASAP7_75t_L g11183 ( 
.A(n_10784),
.B(n_965),
.Y(n_11183)
);

INVx1_ASAP7_75t_L g11184 ( 
.A(n_10353),
.Y(n_11184)
);

BUFx6f_ASAP7_75t_L g11185 ( 
.A(n_10682),
.Y(n_11185)
);

NOR2xp33_ASAP7_75t_L g11186 ( 
.A(n_10570),
.B(n_966),
.Y(n_11186)
);

AOI21xp5_ASAP7_75t_L g11187 ( 
.A1(n_10678),
.A2(n_967),
.B(n_968),
.Y(n_11187)
);

INVx2_ASAP7_75t_L g11188 ( 
.A(n_10351),
.Y(n_11188)
);

NAND2x1_ASAP7_75t_L g11189 ( 
.A(n_10265),
.B(n_967),
.Y(n_11189)
);

AOI21xp5_ASAP7_75t_L g11190 ( 
.A1(n_10681),
.A2(n_968),
.B(n_969),
.Y(n_11190)
);

O2A1O1Ixp33_ASAP7_75t_L g11191 ( 
.A1(n_10649),
.A2(n_971),
.B(n_969),
.C(n_970),
.Y(n_11191)
);

CKINVDCx10_ASAP7_75t_R g11192 ( 
.A(n_10326),
.Y(n_11192)
);

HB1xp67_ASAP7_75t_L g11193 ( 
.A(n_10217),
.Y(n_11193)
);

BUFx3_ASAP7_75t_L g11194 ( 
.A(n_10429),
.Y(n_11194)
);

INVx1_ASAP7_75t_L g11195 ( 
.A(n_10312),
.Y(n_11195)
);

NAND2xp5_ASAP7_75t_L g11196 ( 
.A(n_10498),
.B(n_970),
.Y(n_11196)
);

AO22x1_ASAP7_75t_L g11197 ( 
.A1(n_10587),
.A2(n_974),
.B1(n_972),
.B2(n_973),
.Y(n_11197)
);

O2A1O1Ixp5_ASAP7_75t_L g11198 ( 
.A1(n_10603),
.A2(n_974),
.B(n_972),
.C(n_973),
.Y(n_11198)
);

NAND2x1p5_ASAP7_75t_L g11199 ( 
.A(n_10433),
.B(n_975),
.Y(n_11199)
);

OR2x2_ASAP7_75t_L g11200 ( 
.A(n_10290),
.B(n_10412),
.Y(n_11200)
);

NAND2xp5_ASAP7_75t_L g11201 ( 
.A(n_10470),
.B(n_10205),
.Y(n_11201)
);

NAND2xp5_ASAP7_75t_L g11202 ( 
.A(n_10480),
.B(n_975),
.Y(n_11202)
);

INVx2_ASAP7_75t_L g11203 ( 
.A(n_10369),
.Y(n_11203)
);

INVx3_ASAP7_75t_L g11204 ( 
.A(n_10684),
.Y(n_11204)
);

AND2x4_ASAP7_75t_L g11205 ( 
.A(n_10132),
.B(n_976),
.Y(n_11205)
);

CKINVDCx8_ASAP7_75t_R g11206 ( 
.A(n_10684),
.Y(n_11206)
);

BUFx6f_ASAP7_75t_L g11207 ( 
.A(n_10139),
.Y(n_11207)
);

NAND2xp5_ASAP7_75t_L g11208 ( 
.A(n_10062),
.B(n_977),
.Y(n_11208)
);

NAND2xp5_ASAP7_75t_SL g11209 ( 
.A(n_10203),
.B(n_978),
.Y(n_11209)
);

NAND2xp5_ASAP7_75t_L g11210 ( 
.A(n_10064),
.B(n_978),
.Y(n_11210)
);

BUFx2_ASAP7_75t_L g11211 ( 
.A(n_10509),
.Y(n_11211)
);

INVx1_ASAP7_75t_L g11212 ( 
.A(n_10312),
.Y(n_11212)
);

INVx1_ASAP7_75t_L g11213 ( 
.A(n_10312),
.Y(n_11213)
);

AOI21xp5_ASAP7_75t_L g11214 ( 
.A1(n_10694),
.A2(n_980),
.B(n_981),
.Y(n_11214)
);

AOI21xp5_ASAP7_75t_L g11215 ( 
.A1(n_10700),
.A2(n_980),
.B(n_981),
.Y(n_11215)
);

AOI21xp5_ASAP7_75t_L g11216 ( 
.A1(n_10703),
.A2(n_982),
.B(n_983),
.Y(n_11216)
);

AOI21xp5_ASAP7_75t_L g11217 ( 
.A1(n_10705),
.A2(n_10720),
.B(n_10713),
.Y(n_11217)
);

BUFx6f_ASAP7_75t_L g11218 ( 
.A(n_10281),
.Y(n_11218)
);

AND2x2_ASAP7_75t_L g11219 ( 
.A(n_10306),
.B(n_983),
.Y(n_11219)
);

BUFx3_ASAP7_75t_L g11220 ( 
.A(n_10301),
.Y(n_11220)
);

INVx1_ASAP7_75t_SL g11221 ( 
.A(n_10226),
.Y(n_11221)
);

CKINVDCx16_ASAP7_75t_R g11222 ( 
.A(n_10568),
.Y(n_11222)
);

HB1xp67_ASAP7_75t_L g11223 ( 
.A(n_10295),
.Y(n_11223)
);

AOI21xp5_ASAP7_75t_L g11224 ( 
.A1(n_10725),
.A2(n_984),
.B(n_985),
.Y(n_11224)
);

NAND2xp5_ASAP7_75t_L g11225 ( 
.A(n_10071),
.B(n_984),
.Y(n_11225)
);

INVx2_ASAP7_75t_SL g11226 ( 
.A(n_10608),
.Y(n_11226)
);

AOI21xp5_ASAP7_75t_L g11227 ( 
.A1(n_10730),
.A2(n_985),
.B(n_986),
.Y(n_11227)
);

INVx1_ASAP7_75t_L g11228 ( 
.A(n_10381),
.Y(n_11228)
);

AOI21xp5_ASAP7_75t_L g11229 ( 
.A1(n_10744),
.A2(n_986),
.B(n_987),
.Y(n_11229)
);

OAI22x1_ASAP7_75t_L g11230 ( 
.A1(n_10300),
.A2(n_989),
.B1(n_987),
.B2(n_988),
.Y(n_11230)
);

NAND2xp5_ASAP7_75t_SL g11231 ( 
.A(n_10683),
.B(n_10689),
.Y(n_11231)
);

NAND2xp5_ASAP7_75t_L g11232 ( 
.A(n_10107),
.B(n_988),
.Y(n_11232)
);

A2O1A1Ixp33_ASAP7_75t_L g11233 ( 
.A1(n_10764),
.A2(n_991),
.B(n_989),
.C(n_990),
.Y(n_11233)
);

AOI21xp5_ASAP7_75t_L g11234 ( 
.A1(n_10768),
.A2(n_990),
.B(n_991),
.Y(n_11234)
);

AND2x2_ASAP7_75t_L g11235 ( 
.A(n_10307),
.B(n_992),
.Y(n_11235)
);

AOI221xp5_ASAP7_75t_L g11236 ( 
.A1(n_10113),
.A2(n_995),
.B1(n_993),
.B2(n_994),
.C(n_996),
.Y(n_11236)
);

INVx3_ASAP7_75t_L g11237 ( 
.A(n_10264),
.Y(n_11237)
);

NAND2xp5_ASAP7_75t_SL g11238 ( 
.A(n_10697),
.B(n_993),
.Y(n_11238)
);

OAI22xp5_ASAP7_75t_SL g11239 ( 
.A1(n_10407),
.A2(n_997),
.B1(n_995),
.B2(n_996),
.Y(n_11239)
);

NAND2xp5_ASAP7_75t_L g11240 ( 
.A(n_10127),
.B(n_997),
.Y(n_11240)
);

NOR2xp33_ASAP7_75t_SL g11241 ( 
.A(n_10080),
.B(n_998),
.Y(n_11241)
);

INVx2_ASAP7_75t_L g11242 ( 
.A(n_10387),
.Y(n_11242)
);

INVx2_ASAP7_75t_L g11243 ( 
.A(n_10297),
.Y(n_11243)
);

INVx6_ASAP7_75t_L g11244 ( 
.A(n_10636),
.Y(n_11244)
);

NAND2xp5_ASAP7_75t_L g11245 ( 
.A(n_10192),
.B(n_998),
.Y(n_11245)
);

INVx1_ASAP7_75t_L g11246 ( 
.A(n_10436),
.Y(n_11246)
);

BUFx3_ASAP7_75t_L g11247 ( 
.A(n_10708),
.Y(n_11247)
);

INVx2_ASAP7_75t_L g11248 ( 
.A(n_10304),
.Y(n_11248)
);

INVx1_ASAP7_75t_L g11249 ( 
.A(n_10500),
.Y(n_11249)
);

O2A1O1Ixp33_ASAP7_75t_L g11250 ( 
.A1(n_10658),
.A2(n_1001),
.B(n_999),
.C(n_1000),
.Y(n_11250)
);

NOR2xp33_ASAP7_75t_L g11251 ( 
.A(n_10591),
.B(n_999),
.Y(n_11251)
);

NOR2xp33_ASAP7_75t_SL g11252 ( 
.A(n_10516),
.B(n_1000),
.Y(n_11252)
);

INVx2_ASAP7_75t_L g11253 ( 
.A(n_10321),
.Y(n_11253)
);

INVx1_ASAP7_75t_L g11254 ( 
.A(n_10374),
.Y(n_11254)
);

A2O1A1Ixp33_ASAP7_75t_L g11255 ( 
.A1(n_10782),
.A2(n_1003),
.B(n_1001),
.C(n_1002),
.Y(n_11255)
);

NAND2xp5_ASAP7_75t_L g11256 ( 
.A(n_10193),
.B(n_1002),
.Y(n_11256)
);

NOR2xp33_ASAP7_75t_L g11257 ( 
.A(n_10597),
.B(n_1004),
.Y(n_11257)
);

NOR2xp33_ASAP7_75t_R g11258 ( 
.A(n_10399),
.B(n_1004),
.Y(n_11258)
);

INVx1_ASAP7_75t_L g11259 ( 
.A(n_10329),
.Y(n_11259)
);

AOI22xp5_ASAP7_75t_L g11260 ( 
.A1(n_10664),
.A2(n_10692),
.B1(n_10710),
.B2(n_10672),
.Y(n_11260)
);

OAI22xp5_ASAP7_75t_L g11261 ( 
.A1(n_10783),
.A2(n_1007),
.B1(n_1005),
.B2(n_1006),
.Y(n_11261)
);

HB1xp67_ASAP7_75t_L g11262 ( 
.A(n_10333),
.Y(n_11262)
);

O2A1O1Ixp33_ASAP7_75t_L g11263 ( 
.A1(n_10719),
.A2(n_1008),
.B(n_1005),
.C(n_1007),
.Y(n_11263)
);

INVx2_ASAP7_75t_L g11264 ( 
.A(n_10443),
.Y(n_11264)
);

AND2x2_ASAP7_75t_L g11265 ( 
.A(n_10355),
.B(n_1009),
.Y(n_11265)
);

NOR2xp33_ASAP7_75t_SL g11266 ( 
.A(n_10630),
.B(n_10645),
.Y(n_11266)
);

BUFx3_ASAP7_75t_L g11267 ( 
.A(n_10638),
.Y(n_11267)
);

AOI21xp5_ASAP7_75t_L g11268 ( 
.A1(n_10785),
.A2(n_1009),
.B(n_1010),
.Y(n_11268)
);

AOI22xp5_ASAP7_75t_L g11269 ( 
.A1(n_10735),
.A2(n_1012),
.B1(n_1010),
.B2(n_1011),
.Y(n_11269)
);

AND2x2_ASAP7_75t_L g11270 ( 
.A(n_10356),
.B(n_1011),
.Y(n_11270)
);

NAND2xp5_ASAP7_75t_L g11271 ( 
.A(n_10195),
.B(n_1012),
.Y(n_11271)
);

INVx2_ASAP7_75t_L g11272 ( 
.A(n_10449),
.Y(n_11272)
);

AOI21xp5_ASAP7_75t_L g11273 ( 
.A1(n_10206),
.A2(n_1013),
.B(n_1014),
.Y(n_11273)
);

NAND2xp5_ASAP7_75t_SL g11274 ( 
.A(n_10751),
.B(n_1013),
.Y(n_11274)
);

INVx2_ASAP7_75t_SL g11275 ( 
.A(n_10643),
.Y(n_11275)
);

O2A1O1Ixp33_ASAP7_75t_L g11276 ( 
.A1(n_10740),
.A2(n_1016),
.B(n_1014),
.C(n_1015),
.Y(n_11276)
);

NAND2xp5_ASAP7_75t_L g11277 ( 
.A(n_10129),
.B(n_1015),
.Y(n_11277)
);

OAI22x1_ASAP7_75t_L g11278 ( 
.A1(n_10748),
.A2(n_1018),
.B1(n_1016),
.B2(n_1017),
.Y(n_11278)
);

OAI22xp5_ASAP7_75t_L g11279 ( 
.A1(n_10754),
.A2(n_1019),
.B1(n_1017),
.B2(n_1018),
.Y(n_11279)
);

NAND2xp5_ASAP7_75t_L g11280 ( 
.A(n_10143),
.B(n_10147),
.Y(n_11280)
);

NAND2xp5_ASAP7_75t_SL g11281 ( 
.A(n_10769),
.B(n_1019),
.Y(n_11281)
);

NAND2xp5_ASAP7_75t_L g11282 ( 
.A(n_10156),
.B(n_1020),
.Y(n_11282)
);

OAI22xp5_ASAP7_75t_L g11283 ( 
.A1(n_10211),
.A2(n_1022),
.B1(n_1020),
.B2(n_1021),
.Y(n_11283)
);

AND2x2_ASAP7_75t_L g11284 ( 
.A(n_10379),
.B(n_1021),
.Y(n_11284)
);

BUFx2_ASAP7_75t_L g11285 ( 
.A(n_10433),
.Y(n_11285)
);

NAND2xp5_ASAP7_75t_L g11286 ( 
.A(n_10162),
.B(n_1022),
.Y(n_11286)
);

INVx2_ASAP7_75t_SL g11287 ( 
.A(n_10745),
.Y(n_11287)
);

AND2x2_ASAP7_75t_L g11288 ( 
.A(n_10390),
.B(n_1023),
.Y(n_11288)
);

O2A1O1Ixp33_ASAP7_75t_L g11289 ( 
.A1(n_10117),
.A2(n_1025),
.B(n_1023),
.C(n_1024),
.Y(n_11289)
);

AND2x2_ASAP7_75t_L g11290 ( 
.A(n_10495),
.B(n_10507),
.Y(n_11290)
);

NOR2xp33_ASAP7_75t_L g11291 ( 
.A(n_10512),
.B(n_1025),
.Y(n_11291)
);

OAI21xp5_ASAP7_75t_L g11292 ( 
.A1(n_10358),
.A2(n_1026),
.B(n_1027),
.Y(n_11292)
);

INVx3_ASAP7_75t_L g11293 ( 
.A(n_10770),
.Y(n_11293)
);

INVx1_ASAP7_75t_L g11294 ( 
.A(n_10223),
.Y(n_11294)
);

AOI21xp5_ASAP7_75t_L g11295 ( 
.A1(n_10340),
.A2(n_1026),
.B(n_1027),
.Y(n_11295)
);

BUFx6f_ASAP7_75t_L g11296 ( 
.A(n_10572),
.Y(n_11296)
);

O2A1O1Ixp5_ASAP7_75t_L g11297 ( 
.A1(n_10335),
.A2(n_1030),
.B(n_1028),
.C(n_1029),
.Y(n_11297)
);

INVx4_ASAP7_75t_L g11298 ( 
.A(n_10433),
.Y(n_11298)
);

INVx2_ASAP7_75t_L g11299 ( 
.A(n_10456),
.Y(n_11299)
);

BUFx2_ASAP7_75t_L g11300 ( 
.A(n_10457),
.Y(n_11300)
);

NAND2xp5_ASAP7_75t_L g11301 ( 
.A(n_10167),
.B(n_1028),
.Y(n_11301)
);

NAND2xp5_ASAP7_75t_L g11302 ( 
.A(n_10183),
.B(n_10185),
.Y(n_11302)
);

INVx1_ASAP7_75t_SL g11303 ( 
.A(n_10504),
.Y(n_11303)
);

NAND2xp5_ASAP7_75t_SL g11304 ( 
.A(n_10270),
.B(n_1029),
.Y(n_11304)
);

AOI21xp5_ASAP7_75t_L g11305 ( 
.A1(n_10342),
.A2(n_10350),
.B(n_10347),
.Y(n_11305)
);

INVx2_ASAP7_75t_SL g11306 ( 
.A(n_10337),
.Y(n_11306)
);

INVx1_ASAP7_75t_L g11307 ( 
.A(n_10458),
.Y(n_11307)
);

INVx3_ASAP7_75t_L g11308 ( 
.A(n_10639),
.Y(n_11308)
);

INVx1_ASAP7_75t_L g11309 ( 
.A(n_10465),
.Y(n_11309)
);

BUFx5_ASAP7_75t_L g11310 ( 
.A(n_10180),
.Y(n_11310)
);

AOI21xp5_ASAP7_75t_L g11311 ( 
.A1(n_10352),
.A2(n_10368),
.B(n_10367),
.Y(n_11311)
);

BUFx3_ASAP7_75t_L g11312 ( 
.A(n_10431),
.Y(n_11312)
);

NAND2xp5_ASAP7_75t_L g11313 ( 
.A(n_10188),
.B(n_1030),
.Y(n_11313)
);

INVx2_ASAP7_75t_L g11314 ( 
.A(n_10191),
.Y(n_11314)
);

AOI21xp5_ASAP7_75t_L g11315 ( 
.A1(n_10370),
.A2(n_1031),
.B(n_1032),
.Y(n_11315)
);

NAND3xp33_ASAP7_75t_SL g11316 ( 
.A(n_10285),
.B(n_1032),
.C(n_1033),
.Y(n_11316)
);

INVx3_ASAP7_75t_L g11317 ( 
.A(n_10302),
.Y(n_11317)
);

NAND2xp5_ASAP7_75t_SL g11318 ( 
.A(n_10201),
.B(n_1033),
.Y(n_11318)
);

BUFx12f_ASAP7_75t_L g11319 ( 
.A(n_10526),
.Y(n_11319)
);

AOI22xp5_ASAP7_75t_L g11320 ( 
.A1(n_10136),
.A2(n_1036),
.B1(n_1034),
.B2(n_1035),
.Y(n_11320)
);

O2A1O1Ixp33_ASAP7_75t_L g11321 ( 
.A1(n_10214),
.A2(n_1037),
.B(n_1034),
.C(n_1036),
.Y(n_11321)
);

OAI21x1_ASAP7_75t_SL g11322 ( 
.A1(n_10179),
.A2(n_1037),
.B(n_1038),
.Y(n_11322)
);

O2A1O1Ixp33_ASAP7_75t_SL g11323 ( 
.A1(n_10654),
.A2(n_1040),
.B(n_1038),
.C(n_1039),
.Y(n_11323)
);

INVxp33_ASAP7_75t_SL g11324 ( 
.A(n_10242),
.Y(n_11324)
);

NOR2xp33_ASAP7_75t_L g11325 ( 
.A(n_10529),
.B(n_1039),
.Y(n_11325)
);

AND2x2_ASAP7_75t_L g11326 ( 
.A(n_10534),
.B(n_1040),
.Y(n_11326)
);

A2O1A1Ixp33_ASAP7_75t_SL g11327 ( 
.A1(n_10605),
.A2(n_1043),
.B(n_1041),
.C(n_1042),
.Y(n_11327)
);

NAND3xp33_ASAP7_75t_SL g11328 ( 
.A(n_10236),
.B(n_1041),
.C(n_1042),
.Y(n_11328)
);

A2O1A1Ixp33_ASAP7_75t_L g11329 ( 
.A1(n_10732),
.A2(n_1045),
.B(n_1043),
.C(n_1044),
.Y(n_11329)
);

INVx1_ASAP7_75t_L g11330 ( 
.A(n_10542),
.Y(n_11330)
);

A2O1A1Ixp33_ASAP7_75t_L g11331 ( 
.A1(n_10776),
.A2(n_1046),
.B(n_1044),
.C(n_1045),
.Y(n_11331)
);

AO21x1_ASAP7_75t_L g11332 ( 
.A1(n_10482),
.A2(n_1046),
.B(n_1047),
.Y(n_11332)
);

O2A1O1Ixp33_ASAP7_75t_L g11333 ( 
.A1(n_10260),
.A2(n_1049),
.B(n_1047),
.C(n_1048),
.Y(n_11333)
);

INVx5_ASAP7_75t_L g11334 ( 
.A(n_10555),
.Y(n_11334)
);

BUFx2_ASAP7_75t_L g11335 ( 
.A(n_10202),
.Y(n_11335)
);

CKINVDCx5p33_ASAP7_75t_R g11336 ( 
.A(n_10451),
.Y(n_11336)
);

NAND2xp5_ASAP7_75t_SL g11337 ( 
.A(n_10413),
.B(n_1049),
.Y(n_11337)
);

CKINVDCx6p67_ASAP7_75t_R g11338 ( 
.A(n_10569),
.Y(n_11338)
);

NAND2x1p5_ASAP7_75t_L g11339 ( 
.A(n_10249),
.B(n_1050),
.Y(n_11339)
);

NAND2xp5_ASAP7_75t_L g11340 ( 
.A(n_10444),
.B(n_1050),
.Y(n_11340)
);

OAI22xp5_ASAP7_75t_L g11341 ( 
.A1(n_10233),
.A2(n_1054),
.B1(n_1051),
.B2(n_1053),
.Y(n_11341)
);

INVx2_ASAP7_75t_L g11342 ( 
.A(n_10576),
.Y(n_11342)
);

AOI21xp5_ASAP7_75t_L g11343 ( 
.A1(n_10375),
.A2(n_1051),
.B(n_1053),
.Y(n_11343)
);

AND2x2_ASAP7_75t_L g11344 ( 
.A(n_10447),
.B(n_1054),
.Y(n_11344)
);

INVx2_ASAP7_75t_SL g11345 ( 
.A(n_10583),
.Y(n_11345)
);

INVx1_ASAP7_75t_L g11346 ( 
.A(n_10520),
.Y(n_11346)
);

INVx3_ASAP7_75t_L g11347 ( 
.A(n_10479),
.Y(n_11347)
);

AND2x2_ASAP7_75t_L g11348 ( 
.A(n_10346),
.B(n_1055),
.Y(n_11348)
);

NAND2xp5_ASAP7_75t_L g11349 ( 
.A(n_10235),
.B(n_1056),
.Y(n_11349)
);

OAI22xp5_ASAP7_75t_L g11350 ( 
.A1(n_10240),
.A2(n_1058),
.B1(n_1056),
.B2(n_1057),
.Y(n_11350)
);

AOI21xp5_ASAP7_75t_L g11351 ( 
.A1(n_10376),
.A2(n_1058),
.B(n_1059),
.Y(n_11351)
);

BUFx3_ASAP7_75t_L g11352 ( 
.A(n_10550),
.Y(n_11352)
);

A2O1A1Ixp33_ASAP7_75t_L g11353 ( 
.A1(n_10435),
.A2(n_1061),
.B(n_1059),
.C(n_1060),
.Y(n_11353)
);

OAI22xp5_ASAP7_75t_L g11354 ( 
.A1(n_10241),
.A2(n_1063),
.B1(n_1060),
.B2(n_1061),
.Y(n_11354)
);

BUFx3_ASAP7_75t_L g11355 ( 
.A(n_10553),
.Y(n_11355)
);

O2A1O1Ixp33_ASAP7_75t_L g11356 ( 
.A1(n_10421),
.A2(n_1065),
.B(n_1063),
.C(n_1064),
.Y(n_11356)
);

INVx1_ASAP7_75t_L g11357 ( 
.A(n_10581),
.Y(n_11357)
);

AOI21xp5_ASAP7_75t_L g11358 ( 
.A1(n_10377),
.A2(n_1064),
.B(n_1065),
.Y(n_11358)
);

A2O1A1Ixp33_ASAP7_75t_L g11359 ( 
.A1(n_10440),
.A2(n_1068),
.B(n_1066),
.C(n_1067),
.Y(n_11359)
);

INVx1_ASAP7_75t_L g11360 ( 
.A(n_10181),
.Y(n_11360)
);

AOI21xp5_ASAP7_75t_L g11361 ( 
.A1(n_10389),
.A2(n_1066),
.B(n_1067),
.Y(n_11361)
);

NAND2xp5_ASAP7_75t_L g11362 ( 
.A(n_10244),
.B(n_1068),
.Y(n_11362)
);

AOI21x1_ASAP7_75t_L g11363 ( 
.A1(n_10125),
.A2(n_1069),
.B(n_1070),
.Y(n_11363)
);

OAI22xp5_ASAP7_75t_L g11364 ( 
.A1(n_10255),
.A2(n_1072),
.B1(n_1070),
.B2(n_1071),
.Y(n_11364)
);

NAND2xp5_ASAP7_75t_L g11365 ( 
.A(n_10256),
.B(n_1071),
.Y(n_11365)
);

NAND2xp5_ASAP7_75t_SL g11366 ( 
.A(n_10411),
.B(n_1072),
.Y(n_11366)
);

NOR2xp33_ASAP7_75t_L g11367 ( 
.A(n_10519),
.B(n_10209),
.Y(n_11367)
);

BUFx2_ASAP7_75t_L g11368 ( 
.A(n_10468),
.Y(n_11368)
);

AOI21x1_ASAP7_75t_L g11369 ( 
.A1(n_10144),
.A2(n_1073),
.B(n_1074),
.Y(n_11369)
);

AOI22xp33_ASAP7_75t_SL g11370 ( 
.A1(n_10134),
.A2(n_1077),
.B1(n_1073),
.B2(n_1075),
.Y(n_11370)
);

AOI21xp5_ASAP7_75t_L g11371 ( 
.A1(n_10393),
.A2(n_1075),
.B(n_1077),
.Y(n_11371)
);

BUFx6f_ASAP7_75t_L g11372 ( 
.A(n_10545),
.Y(n_11372)
);

AOI21xp5_ASAP7_75t_L g11373 ( 
.A1(n_10401),
.A2(n_1078),
.B(n_1080),
.Y(n_11373)
);

AOI21xp5_ASAP7_75t_L g11374 ( 
.A1(n_10286),
.A2(n_1078),
.B(n_1080),
.Y(n_11374)
);

AOI21xp5_ASAP7_75t_L g11375 ( 
.A1(n_10293),
.A2(n_1081),
.B(n_1082),
.Y(n_11375)
);

A2O1A1Ixp33_ASAP7_75t_SL g11376 ( 
.A1(n_10438),
.A2(n_10339),
.B(n_10469),
.C(n_10467),
.Y(n_11376)
);

AND2x2_ASAP7_75t_L g11377 ( 
.A(n_10556),
.B(n_1081),
.Y(n_11377)
);

NOR2xp33_ASAP7_75t_L g11378 ( 
.A(n_10484),
.B(n_10305),
.Y(n_11378)
);

NAND2xp5_ASAP7_75t_L g11379 ( 
.A(n_10177),
.B(n_1082),
.Y(n_11379)
);

NOR3xp33_ASAP7_75t_SL g11380 ( 
.A(n_10472),
.B(n_10476),
.C(n_10251),
.Y(n_11380)
);

NAND2x1p5_ASAP7_75t_L g11381 ( 
.A(n_10278),
.B(n_1083),
.Y(n_11381)
);

INVx1_ASAP7_75t_L g11382 ( 
.A(n_10405),
.Y(n_11382)
);

BUFx2_ASAP7_75t_L g11383 ( 
.A(n_10558),
.Y(n_11383)
);

INVx6_ASAP7_75t_L g11384 ( 
.A(n_10596),
.Y(n_11384)
);

NAND2xp5_ASAP7_75t_SL g11385 ( 
.A(n_10359),
.B(n_1083),
.Y(n_11385)
);

AND2x2_ASAP7_75t_L g11386 ( 
.A(n_10562),
.B(n_10496),
.Y(n_11386)
);

INVx2_ASAP7_75t_L g11387 ( 
.A(n_10283),
.Y(n_11387)
);

NAND2xp5_ASAP7_75t_L g11388 ( 
.A(n_10104),
.B(n_1084),
.Y(n_11388)
);

OR2x4_ASAP7_75t_L g11389 ( 
.A(n_10714),
.B(n_1084),
.Y(n_11389)
);

O2A1O1Ixp5_ASAP7_75t_SL g11390 ( 
.A1(n_10298),
.A2(n_1087),
.B(n_1085),
.C(n_1086),
.Y(n_11390)
);

NAND2xp5_ASAP7_75t_L g11391 ( 
.A(n_10331),
.B(n_1085),
.Y(n_11391)
);

NAND2xp5_ASAP7_75t_L g11392 ( 
.A(n_10239),
.B(n_1086),
.Y(n_11392)
);

OAI22xp5_ASAP7_75t_L g11393 ( 
.A1(n_10753),
.A2(n_1091),
.B1(n_1089),
.B2(n_1090),
.Y(n_11393)
);

OR2x6_ASAP7_75t_L g11394 ( 
.A(n_10432),
.B(n_1089),
.Y(n_11394)
);

A2O1A1Ixp33_ASAP7_75t_L g11395 ( 
.A1(n_10442),
.A2(n_1092),
.B(n_1090),
.C(n_1091),
.Y(n_11395)
);

AOI21xp5_ASAP7_75t_L g11396 ( 
.A1(n_10296),
.A2(n_1093),
.B(n_1094),
.Y(n_11396)
);

AOI21xp5_ASAP7_75t_L g11397 ( 
.A1(n_10308),
.A2(n_1093),
.B(n_1094),
.Y(n_11397)
);

AOI21xp5_ASAP7_75t_L g11398 ( 
.A1(n_10332),
.A2(n_1095),
.B(n_1096),
.Y(n_11398)
);

AND2x2_ASAP7_75t_L g11399 ( 
.A(n_10551),
.B(n_10578),
.Y(n_11399)
);

BUFx6f_ASAP7_75t_L g11400 ( 
.A(n_10598),
.Y(n_11400)
);

AOI21xp5_ASAP7_75t_L g11401 ( 
.A1(n_10446),
.A2(n_1095),
.B(n_1096),
.Y(n_11401)
);

A2O1A1Ixp33_ASAP7_75t_SL g11402 ( 
.A1(n_10253),
.A2(n_1099),
.B(n_1097),
.C(n_1098),
.Y(n_11402)
);

NAND2xp5_ASAP7_75t_L g11403 ( 
.A(n_10257),
.B(n_1097),
.Y(n_11403)
);

INVxp67_ASAP7_75t_L g11404 ( 
.A(n_10218),
.Y(n_11404)
);

INVx2_ASAP7_75t_L g11405 ( 
.A(n_10327),
.Y(n_11405)
);

INVx2_ASAP7_75t_L g11406 ( 
.A(n_10366),
.Y(n_11406)
);

NAND2xp5_ASAP7_75t_L g11407 ( 
.A(n_10072),
.B(n_1098),
.Y(n_11407)
);

BUFx6f_ASAP7_75t_L g11408 ( 
.A(n_10590),
.Y(n_11408)
);

AOI21xp5_ASAP7_75t_L g11409 ( 
.A1(n_10452),
.A2(n_1100),
.B(n_1101),
.Y(n_11409)
);

INVx4_ASAP7_75t_L g11410 ( 
.A(n_10225),
.Y(n_11410)
);

INVx5_ASAP7_75t_L g11411 ( 
.A(n_10774),
.Y(n_11411)
);

NOR2xp33_ASAP7_75t_L g11412 ( 
.A(n_10738),
.B(n_1100),
.Y(n_11412)
);

O2A1O1Ixp33_ASAP7_75t_L g11413 ( 
.A1(n_10303),
.A2(n_1104),
.B(n_1102),
.C(n_1103),
.Y(n_11413)
);

NAND2xp5_ASAP7_75t_SL g11414 ( 
.A(n_10420),
.B(n_1103),
.Y(n_11414)
);

AND2x4_ASAP7_75t_L g11415 ( 
.A(n_10314),
.B(n_1104),
.Y(n_11415)
);

OAI21xp33_ASAP7_75t_L g11416 ( 
.A1(n_10477),
.A2(n_1105),
.B(n_1106),
.Y(n_11416)
);

INVx2_ASAP7_75t_L g11417 ( 
.A(n_10318),
.Y(n_11417)
);

OAI22xp5_ASAP7_75t_L g11418 ( 
.A1(n_10571),
.A2(n_1108),
.B1(n_1106),
.B2(n_1107),
.Y(n_11418)
);

INVx2_ASAP7_75t_L g11419 ( 
.A(n_10518),
.Y(n_11419)
);

OAI21x1_ASAP7_75t_L g11420 ( 
.A1(n_10414),
.A2(n_1107),
.B(n_1108),
.Y(n_11420)
);

INVx1_ASAP7_75t_L g11421 ( 
.A(n_10417),
.Y(n_11421)
);

AO21x1_ASAP7_75t_L g11422 ( 
.A1(n_10116),
.A2(n_1109),
.B(n_1110),
.Y(n_11422)
);

A2O1A1Ixp33_ASAP7_75t_L g11423 ( 
.A1(n_10200),
.A2(n_1111),
.B(n_1109),
.C(n_1110),
.Y(n_11423)
);

OAI221xp5_ASAP7_75t_L g11424 ( 
.A1(n_10502),
.A2(n_1114),
.B1(n_1111),
.B2(n_1112),
.C(n_1115),
.Y(n_11424)
);

NAND2xp5_ASAP7_75t_L g11425 ( 
.A(n_10739),
.B(n_10757),
.Y(n_11425)
);

O2A1O1Ixp5_ASAP7_75t_L g11426 ( 
.A1(n_10152),
.A2(n_1115),
.B(n_1112),
.C(n_1114),
.Y(n_11426)
);

AOI22xp5_ASAP7_75t_SL g11427 ( 
.A1(n_10560),
.A2(n_10565),
.B1(n_10176),
.B2(n_10548),
.Y(n_11427)
);

NOR2xp33_ASAP7_75t_L g11428 ( 
.A(n_10775),
.B(n_1116),
.Y(n_11428)
);

AND2x2_ASAP7_75t_L g11429 ( 
.A(n_10276),
.B(n_1116),
.Y(n_11429)
);

A2O1A1Ixp33_ASAP7_75t_L g11430 ( 
.A1(n_10159),
.A2(n_1119),
.B(n_1117),
.C(n_1118),
.Y(n_11430)
);

BUFx6f_ASAP7_75t_L g11431 ( 
.A(n_10096),
.Y(n_11431)
);

INVx2_ASAP7_75t_L g11432 ( 
.A(n_10430),
.Y(n_11432)
);

INVx6_ASAP7_75t_L g11433 ( 
.A(n_10487),
.Y(n_11433)
);

NAND2xp5_ASAP7_75t_L g11434 ( 
.A(n_10779),
.B(n_1117),
.Y(n_11434)
);

NOR2xp33_ASAP7_75t_L g11435 ( 
.A(n_10780),
.B(n_1118),
.Y(n_11435)
);

NOR2xp33_ASAP7_75t_L g11436 ( 
.A(n_10101),
.B(n_1119),
.Y(n_11436)
);

AOI21xp5_ASAP7_75t_L g11437 ( 
.A1(n_10160),
.A2(n_1120),
.B(n_1121),
.Y(n_11437)
);

NOR2xp33_ASAP7_75t_R g11438 ( 
.A(n_10168),
.B(n_1121),
.Y(n_11438)
);

OAI21xp5_ASAP7_75t_L g11439 ( 
.A1(n_10426),
.A2(n_1122),
.B(n_1123),
.Y(n_11439)
);

NOR2xp33_ASAP7_75t_L g11440 ( 
.A(n_10575),
.B(n_1124),
.Y(n_11440)
);

INVx2_ASAP7_75t_SL g11441 ( 
.A(n_10196),
.Y(n_11441)
);

AOI21xp5_ASAP7_75t_L g11442 ( 
.A1(n_10173),
.A2(n_1125),
.B(n_1126),
.Y(n_11442)
);

OAI22xp5_ASAP7_75t_L g11443 ( 
.A1(n_10530),
.A2(n_1127),
.B1(n_1125),
.B2(n_1126),
.Y(n_11443)
);

INVx3_ASAP7_75t_L g11444 ( 
.A(n_10537),
.Y(n_11444)
);

O2A1O1Ixp33_ASAP7_75t_SL g11445 ( 
.A1(n_10052),
.A2(n_1129),
.B(n_1127),
.C(n_1128),
.Y(n_11445)
);

O2A1O1Ixp33_ASAP7_75t_L g11446 ( 
.A1(n_10612),
.A2(n_1131),
.B(n_1128),
.C(n_1129),
.Y(n_11446)
);

CKINVDCx5p33_ASAP7_75t_R g11447 ( 
.A(n_10149),
.Y(n_11447)
);

NAND2xp5_ASAP7_75t_L g11448 ( 
.A(n_10491),
.B(n_1131),
.Y(n_11448)
);

OAI22xp5_ASAP7_75t_L g11449 ( 
.A1(n_10574),
.A2(n_1134),
.B1(n_1132),
.B2(n_1133),
.Y(n_11449)
);

INVx2_ASAP7_75t_L g11450 ( 
.A(n_10619),
.Y(n_11450)
);

INVx1_ASAP7_75t_L g11451 ( 
.A(n_10121),
.Y(n_11451)
);

OAI21xp5_ASAP7_75t_L g11452 ( 
.A1(n_10174),
.A2(n_10194),
.B(n_10189),
.Y(n_11452)
);

A2O1A1Ixp33_ASAP7_75t_L g11453 ( 
.A1(n_10486),
.A2(n_1135),
.B(n_1132),
.C(n_1134),
.Y(n_11453)
);

INVx2_ASAP7_75t_L g11454 ( 
.A(n_10718),
.Y(n_11454)
);

INVx1_ASAP7_75t_L g11455 ( 
.A(n_10197),
.Y(n_11455)
);

A2O1A1Ixp33_ASAP7_75t_L g11456 ( 
.A1(n_10503),
.A2(n_1137),
.B(n_1135),
.C(n_1136),
.Y(n_11456)
);

NAND2xp5_ASAP7_75t_SL g11457 ( 
.A(n_10543),
.B(n_1136),
.Y(n_11457)
);

AOI22xp33_ASAP7_75t_SL g11458 ( 
.A1(n_10728),
.A2(n_1140),
.B1(n_1137),
.B2(n_1138),
.Y(n_11458)
);

AOI21xp5_ASAP7_75t_L g11459 ( 
.A1(n_10546),
.A2(n_1138),
.B(n_1140),
.Y(n_11459)
);

NAND3xp33_ASAP7_75t_SL g11460 ( 
.A(n_10601),
.B(n_1141),
.C(n_1142),
.Y(n_11460)
);

AND2x2_ASAP7_75t_L g11461 ( 
.A(n_10557),
.B(n_1141),
.Y(n_11461)
);

NAND2xp5_ASAP7_75t_L g11462 ( 
.A(n_10506),
.B(n_10510),
.Y(n_11462)
);

O2A1O1Ixp33_ASAP7_75t_L g11463 ( 
.A1(n_10741),
.A2(n_10788),
.B(n_10511),
.C(n_10515),
.Y(n_11463)
);

O2A1O1Ixp33_ASAP7_75t_L g11464 ( 
.A1(n_10604),
.A2(n_1145),
.B(n_1143),
.C(n_1144),
.Y(n_11464)
);

OAI21x1_ASAP7_75t_L g11465 ( 
.A1(n_10592),
.A2(n_10599),
.B(n_10234),
.Y(n_11465)
);

INVx4_ASAP7_75t_L g11466 ( 
.A(n_10573),
.Y(n_11466)
);

O2A1O1Ixp33_ASAP7_75t_L g11467 ( 
.A1(n_10580),
.A2(n_1145),
.B(n_1143),
.C(n_1144),
.Y(n_11467)
);

INVx1_ASAP7_75t_L g11468 ( 
.A(n_10584),
.Y(n_11468)
);

NAND2xp5_ASAP7_75t_L g11469 ( 
.A(n_10586),
.B(n_1146),
.Y(n_11469)
);

INVx1_ASAP7_75t_L g11470 ( 
.A(n_10563),
.Y(n_11470)
);

BUFx12f_ASAP7_75t_L g11471 ( 
.A(n_10232),
.Y(n_11471)
);

BUFx6f_ASAP7_75t_L g11472 ( 
.A(n_10155),
.Y(n_11472)
);

AOI21xp5_ASAP7_75t_L g11473 ( 
.A1(n_10103),
.A2(n_1146),
.B(n_1147),
.Y(n_11473)
);

A2O1A1Ixp33_ASAP7_75t_L g11474 ( 
.A1(n_10091),
.A2(n_1149),
.B(n_1147),
.C(n_1148),
.Y(n_11474)
);

AOI21xp5_ASAP7_75t_L g11475 ( 
.A1(n_10103),
.A2(n_1149),
.B(n_1150),
.Y(n_11475)
);

HB1xp67_ASAP7_75t_L g11476 ( 
.A(n_10213),
.Y(n_11476)
);

INVx2_ASAP7_75t_L g11477 ( 
.A(n_10336),
.Y(n_11477)
);

AOI21x1_ASAP7_75t_L g11478 ( 
.A1(n_10103),
.A2(n_1150),
.B(n_1151),
.Y(n_11478)
);

NAND2xp5_ASAP7_75t_L g11479 ( 
.A(n_10082),
.B(n_1151),
.Y(n_11479)
);

CKINVDCx5p33_ASAP7_75t_R g11480 ( 
.A(n_10114),
.Y(n_11480)
);

NOR2xp33_ASAP7_75t_L g11481 ( 
.A(n_10724),
.B(n_1152),
.Y(n_11481)
);

NAND2xp5_ASAP7_75t_L g11482 ( 
.A(n_10082),
.B(n_1152),
.Y(n_11482)
);

OAI22xp5_ASAP7_75t_L g11483 ( 
.A1(n_10091),
.A2(n_1157),
.B1(n_1155),
.B2(n_1156),
.Y(n_11483)
);

NAND2xp5_ASAP7_75t_L g11484 ( 
.A(n_10082),
.B(n_1155),
.Y(n_11484)
);

BUFx4f_ASAP7_75t_SL g11485 ( 
.A(n_10706),
.Y(n_11485)
);

AND2x4_ASAP7_75t_L g11486 ( 
.A(n_10385),
.B(n_1157),
.Y(n_11486)
);

INVx1_ASAP7_75t_L g11487 ( 
.A(n_10053),
.Y(n_11487)
);

NAND2xp5_ASAP7_75t_L g11488 ( 
.A(n_10082),
.B(n_1158),
.Y(n_11488)
);

OAI22xp5_ASAP7_75t_L g11489 ( 
.A1(n_10091),
.A2(n_1162),
.B1(n_1160),
.B2(n_1161),
.Y(n_11489)
);

OAI22xp5_ASAP7_75t_L g11490 ( 
.A1(n_10091),
.A2(n_1163),
.B1(n_1161),
.B2(n_1162),
.Y(n_11490)
);

OAI22x1_ASAP7_75t_L g11491 ( 
.A1(n_10243),
.A2(n_1165),
.B1(n_1163),
.B2(n_1164),
.Y(n_11491)
);

AOI21xp5_ASAP7_75t_L g11492 ( 
.A1(n_10103),
.A2(n_1164),
.B(n_1166),
.Y(n_11492)
);

INVx5_ASAP7_75t_L g11493 ( 
.A(n_10706),
.Y(n_11493)
);

O2A1O1Ixp33_ASAP7_75t_L g11494 ( 
.A1(n_10068),
.A2(n_1168),
.B(n_1166),
.C(n_1167),
.Y(n_11494)
);

AOI21xp5_ASAP7_75t_L g11495 ( 
.A1(n_10103),
.A2(n_1167),
.B(n_1168),
.Y(n_11495)
);

A2O1A1Ixp33_ASAP7_75t_L g11496 ( 
.A1(n_10091),
.A2(n_1171),
.B(n_1169),
.C(n_1170),
.Y(n_11496)
);

HB1xp67_ASAP7_75t_L g11497 ( 
.A(n_10213),
.Y(n_11497)
);

OAI22xp5_ASAP7_75t_L g11498 ( 
.A1(n_10091),
.A2(n_1171),
.B1(n_1169),
.B2(n_1170),
.Y(n_11498)
);

A2O1A1Ixp33_ASAP7_75t_L g11499 ( 
.A1(n_10091),
.A2(n_1175),
.B(n_1173),
.C(n_1174),
.Y(n_11499)
);

AND2x6_ASAP7_75t_L g11500 ( 
.A(n_10245),
.B(n_1174),
.Y(n_11500)
);

INVx1_ASAP7_75t_SL g11501 ( 
.A(n_10724),
.Y(n_11501)
);

O2A1O1Ixp5_ASAP7_75t_L g11502 ( 
.A1(n_10094),
.A2(n_1177),
.B(n_1175),
.C(n_1176),
.Y(n_11502)
);

NAND2xp5_ASAP7_75t_L g11503 ( 
.A(n_10082),
.B(n_1177),
.Y(n_11503)
);

NAND2xp5_ASAP7_75t_L g11504 ( 
.A(n_10082),
.B(n_1178),
.Y(n_11504)
);

INVx1_ASAP7_75t_L g11505 ( 
.A(n_10053),
.Y(n_11505)
);

NOR2xp33_ASAP7_75t_L g11506 ( 
.A(n_10724),
.B(n_1178),
.Y(n_11506)
);

NAND2xp5_ASAP7_75t_L g11507 ( 
.A(n_10082),
.B(n_1179),
.Y(n_11507)
);

A2O1A1Ixp33_ASAP7_75t_L g11508 ( 
.A1(n_10091),
.A2(n_1181),
.B(n_1179),
.C(n_1180),
.Y(n_11508)
);

AOI21xp5_ASAP7_75t_L g11509 ( 
.A1(n_10103),
.A2(n_1180),
.B(n_1182),
.Y(n_11509)
);

AND2x4_ASAP7_75t_L g11510 ( 
.A(n_10385),
.B(n_1182),
.Y(n_11510)
);

NOR2xp33_ASAP7_75t_SL g11511 ( 
.A(n_10169),
.B(n_1183),
.Y(n_11511)
);

A2O1A1Ixp33_ASAP7_75t_L g11512 ( 
.A1(n_10091),
.A2(n_1186),
.B(n_1184),
.C(n_1185),
.Y(n_11512)
);

CKINVDCx5p33_ASAP7_75t_R g11513 ( 
.A(n_10114),
.Y(n_11513)
);

INVxp67_ASAP7_75t_SL g11514 ( 
.A(n_10213),
.Y(n_11514)
);

OR2x6_ASAP7_75t_L g11515 ( 
.A(n_10204),
.B(n_1184),
.Y(n_11515)
);

NAND2x1p5_ASAP7_75t_L g11516 ( 
.A(n_10207),
.B(n_1185),
.Y(n_11516)
);

AOI21xp5_ASAP7_75t_L g11517 ( 
.A1(n_10103),
.A2(n_1186),
.B(n_1187),
.Y(n_11517)
);

OAI21x1_ASAP7_75t_L g11518 ( 
.A1(n_10787),
.A2(n_1187),
.B(n_1188),
.Y(n_11518)
);

NOR2xp33_ASAP7_75t_L g11519 ( 
.A(n_10724),
.B(n_1189),
.Y(n_11519)
);

NOR2x1_ASAP7_75t_L g11520 ( 
.A(n_10082),
.B(n_1189),
.Y(n_11520)
);

NAND2xp5_ASAP7_75t_L g11521 ( 
.A(n_10082),
.B(n_1190),
.Y(n_11521)
);

INVx2_ASAP7_75t_L g11522 ( 
.A(n_10336),
.Y(n_11522)
);

O2A1O1Ixp5_ASAP7_75t_L g11523 ( 
.A1(n_10094),
.A2(n_1192),
.B(n_1190),
.C(n_1191),
.Y(n_11523)
);

INVx4_ASAP7_75t_L g11524 ( 
.A(n_10532),
.Y(n_11524)
);

AOI21x1_ASAP7_75t_L g11525 ( 
.A1(n_10103),
.A2(n_1192),
.B(n_1193),
.Y(n_11525)
);

OAI21x1_ASAP7_75t_L g11526 ( 
.A1(n_10787),
.A2(n_1193),
.B(n_1194),
.Y(n_11526)
);

BUFx6f_ASAP7_75t_L g11527 ( 
.A(n_10155),
.Y(n_11527)
);

NAND2xp5_ASAP7_75t_L g11528 ( 
.A(n_10082),
.B(n_1194),
.Y(n_11528)
);

NAND2xp5_ASAP7_75t_L g11529 ( 
.A(n_10082),
.B(n_1195),
.Y(n_11529)
);

AND2x2_ASAP7_75t_L g11530 ( 
.A(n_10089),
.B(n_1195),
.Y(n_11530)
);

BUFx6f_ASAP7_75t_L g11531 ( 
.A(n_10155),
.Y(n_11531)
);

INVx2_ASAP7_75t_L g11532 ( 
.A(n_10336),
.Y(n_11532)
);

NAND2xp5_ASAP7_75t_L g11533 ( 
.A(n_10082),
.B(n_1196),
.Y(n_11533)
);

AOI21xp5_ASAP7_75t_L g11534 ( 
.A1(n_10103),
.A2(n_1197),
.B(n_1198),
.Y(n_11534)
);

AOI21xp5_ASAP7_75t_L g11535 ( 
.A1(n_10103),
.A2(n_1197),
.B(n_1198),
.Y(n_11535)
);

NAND2xp5_ASAP7_75t_L g11536 ( 
.A(n_10082),
.B(n_1199),
.Y(n_11536)
);

NAND2xp5_ASAP7_75t_L g11537 ( 
.A(n_10082),
.B(n_1199),
.Y(n_11537)
);

INVx1_ASAP7_75t_L g11538 ( 
.A(n_10053),
.Y(n_11538)
);

AOI21xp5_ASAP7_75t_L g11539 ( 
.A1(n_10103),
.A2(n_1200),
.B(n_1201),
.Y(n_11539)
);

INVx1_ASAP7_75t_L g11540 ( 
.A(n_10053),
.Y(n_11540)
);

NAND3xp33_ASAP7_75t_L g11541 ( 
.A(n_10091),
.B(n_1200),
.C(n_1201),
.Y(n_11541)
);

NAND2xp5_ASAP7_75t_SL g11542 ( 
.A(n_10103),
.B(n_1202),
.Y(n_11542)
);

NAND2xp5_ASAP7_75t_L g11543 ( 
.A(n_10082),
.B(n_1203),
.Y(n_11543)
);

NAND2xp5_ASAP7_75t_L g11544 ( 
.A(n_10082),
.B(n_1203),
.Y(n_11544)
);

HB1xp67_ASAP7_75t_L g11545 ( 
.A(n_10213),
.Y(n_11545)
);

NAND2xp5_ASAP7_75t_SL g11546 ( 
.A(n_10103),
.B(n_1204),
.Y(n_11546)
);

NAND2xp5_ASAP7_75t_L g11547 ( 
.A(n_10082),
.B(n_1204),
.Y(n_11547)
);

NAND2xp5_ASAP7_75t_SL g11548 ( 
.A(n_10103),
.B(n_1205),
.Y(n_11548)
);

NAND2xp5_ASAP7_75t_L g11549 ( 
.A(n_10082),
.B(n_1205),
.Y(n_11549)
);

NAND2xp5_ASAP7_75t_L g11550 ( 
.A(n_10082),
.B(n_1206),
.Y(n_11550)
);

NAND2xp5_ASAP7_75t_SL g11551 ( 
.A(n_10103),
.B(n_1206),
.Y(n_11551)
);

INVx3_ASAP7_75t_L g11552 ( 
.A(n_10532),
.Y(n_11552)
);

INVx1_ASAP7_75t_L g11553 ( 
.A(n_10053),
.Y(n_11553)
);

AOI21xp5_ASAP7_75t_L g11554 ( 
.A1(n_10103),
.A2(n_1207),
.B(n_1208),
.Y(n_11554)
);

BUFx6f_ASAP7_75t_L g11555 ( 
.A(n_10155),
.Y(n_11555)
);

AOI21x1_ASAP7_75t_L g11556 ( 
.A1(n_10103),
.A2(n_1207),
.B(n_1208),
.Y(n_11556)
);

AOI21xp5_ASAP7_75t_L g11557 ( 
.A1(n_10103),
.A2(n_1209),
.B(n_1210),
.Y(n_11557)
);

AOI21xp5_ASAP7_75t_L g11558 ( 
.A1(n_10103),
.A2(n_1209),
.B(n_1210),
.Y(n_11558)
);

BUFx2_ASAP7_75t_L g11559 ( 
.A(n_10385),
.Y(n_11559)
);

A2O1A1Ixp33_ASAP7_75t_L g11560 ( 
.A1(n_10091),
.A2(n_1213),
.B(n_1211),
.C(n_1212),
.Y(n_11560)
);

OAI22xp33_ASAP7_75t_L g11561 ( 
.A1(n_10099),
.A2(n_1214),
.B1(n_1211),
.B2(n_1213),
.Y(n_11561)
);

INVx1_ASAP7_75t_L g11562 ( 
.A(n_10906),
.Y(n_11562)
);

AO21x1_ASAP7_75t_L g11563 ( 
.A1(n_10795),
.A2(n_1214),
.B(n_1215),
.Y(n_11563)
);

OAI22xp5_ASAP7_75t_L g11564 ( 
.A1(n_10897),
.A2(n_1217),
.B1(n_1215),
.B2(n_1216),
.Y(n_11564)
);

BUFx6f_ASAP7_75t_SL g11565 ( 
.A(n_11076),
.Y(n_11565)
);

AND2x2_ASAP7_75t_L g11566 ( 
.A(n_11559),
.B(n_1216),
.Y(n_11566)
);

OAI21xp33_ASAP7_75t_L g11567 ( 
.A1(n_10896),
.A2(n_1217),
.B(n_1218),
.Y(n_11567)
);

AO21x2_ASAP7_75t_L g11568 ( 
.A1(n_11136),
.A2(n_1219),
.B(n_1220),
.Y(n_11568)
);

OAI22xp5_ASAP7_75t_L g11569 ( 
.A1(n_11139),
.A2(n_1222),
.B1(n_1220),
.B2(n_1221),
.Y(n_11569)
);

O2A1O1Ixp5_ASAP7_75t_L g11570 ( 
.A1(n_10898),
.A2(n_1223),
.B(n_1221),
.C(n_1222),
.Y(n_11570)
);

AND2x4_ASAP7_75t_L g11571 ( 
.A(n_10816),
.B(n_1223),
.Y(n_11571)
);

INVx2_ASAP7_75t_L g11572 ( 
.A(n_10910),
.Y(n_11572)
);

NAND2xp5_ASAP7_75t_L g11573 ( 
.A(n_11132),
.B(n_1224),
.Y(n_11573)
);

INVx3_ASAP7_75t_L g11574 ( 
.A(n_10792),
.Y(n_11574)
);

AOI21xp5_ASAP7_75t_L g11575 ( 
.A1(n_10839),
.A2(n_11010),
.B(n_10986),
.Y(n_11575)
);

NAND2xp5_ASAP7_75t_SL g11576 ( 
.A(n_11520),
.B(n_10832),
.Y(n_11576)
);

OAI21x1_ASAP7_75t_L g11577 ( 
.A1(n_10860),
.A2(n_1224),
.B(n_1225),
.Y(n_11577)
);

OAI21xp5_ASAP7_75t_L g11578 ( 
.A1(n_10888),
.A2(n_11473),
.B(n_10794),
.Y(n_11578)
);

NOR2x1_ASAP7_75t_SL g11579 ( 
.A(n_11515),
.B(n_1225),
.Y(n_11579)
);

OAI21xp5_ASAP7_75t_L g11580 ( 
.A1(n_11475),
.A2(n_1226),
.B(n_1227),
.Y(n_11580)
);

AOI21xp5_ASAP7_75t_L g11581 ( 
.A1(n_10820),
.A2(n_1226),
.B(n_1228),
.Y(n_11581)
);

OR2x2_ASAP7_75t_L g11582 ( 
.A(n_11476),
.B(n_1228),
.Y(n_11582)
);

OAI21x1_ASAP7_75t_L g11583 ( 
.A1(n_11175),
.A2(n_1229),
.B(n_1231),
.Y(n_11583)
);

NAND2xp5_ASAP7_75t_SL g11584 ( 
.A(n_10832),
.B(n_1229),
.Y(n_11584)
);

AND2x2_ASAP7_75t_L g11585 ( 
.A(n_10891),
.B(n_1232),
.Y(n_11585)
);

AOI21xp33_ASAP7_75t_L g11586 ( 
.A1(n_10845),
.A2(n_11376),
.B(n_11462),
.Y(n_11586)
);

OAI21x1_ASAP7_75t_L g11587 ( 
.A1(n_11465),
.A2(n_11311),
.B(n_11305),
.Y(n_11587)
);

OAI21x1_ASAP7_75t_L g11588 ( 
.A1(n_11342),
.A2(n_1232),
.B(n_1233),
.Y(n_11588)
);

NAND2xp5_ASAP7_75t_L g11589 ( 
.A(n_11152),
.B(n_11497),
.Y(n_11589)
);

OAI21x1_ASAP7_75t_L g11590 ( 
.A1(n_11184),
.A2(n_11294),
.B(n_11382),
.Y(n_11590)
);

OAI21x1_ASAP7_75t_L g11591 ( 
.A1(n_11421),
.A2(n_1233),
.B(n_1234),
.Y(n_11591)
);

NAND2xp5_ASAP7_75t_L g11592 ( 
.A(n_11545),
.B(n_1234),
.Y(n_11592)
);

INVx1_ASAP7_75t_L g11593 ( 
.A(n_10920),
.Y(n_11593)
);

AOI22xp5_ASAP7_75t_L g11594 ( 
.A1(n_10840),
.A2(n_10823),
.B1(n_10805),
.B2(n_11062),
.Y(n_11594)
);

A2O1A1Ixp33_ASAP7_75t_L g11595 ( 
.A1(n_11141),
.A2(n_11091),
.B(n_11017),
.C(n_11059),
.Y(n_11595)
);

AO21x2_ASAP7_75t_L g11596 ( 
.A1(n_11330),
.A2(n_11246),
.B(n_11346),
.Y(n_11596)
);

AND2x2_ASAP7_75t_L g11597 ( 
.A(n_10858),
.B(n_1235),
.Y(n_11597)
);

AOI21xp5_ASAP7_75t_L g11598 ( 
.A1(n_10983),
.A2(n_1235),
.B(n_1236),
.Y(n_11598)
);

AOI21xp5_ASAP7_75t_L g11599 ( 
.A1(n_11452),
.A2(n_1236),
.B(n_1237),
.Y(n_11599)
);

AOI21xp5_ASAP7_75t_L g11600 ( 
.A1(n_11123),
.A2(n_11217),
.B(n_10964),
.Y(n_11600)
);

CKINVDCx20_ASAP7_75t_R g11601 ( 
.A(n_10826),
.Y(n_11601)
);

AOI21xp5_ASAP7_75t_L g11602 ( 
.A1(n_10946),
.A2(n_1237),
.B(n_1238),
.Y(n_11602)
);

AOI21xp5_ASAP7_75t_L g11603 ( 
.A1(n_10977),
.A2(n_1238),
.B(n_1239),
.Y(n_11603)
);

OAI21xp5_ASAP7_75t_L g11604 ( 
.A1(n_11492),
.A2(n_1240),
.B(n_1241),
.Y(n_11604)
);

NAND2xp5_ASAP7_75t_L g11605 ( 
.A(n_11514),
.B(n_1240),
.Y(n_11605)
);

OAI21x1_ASAP7_75t_L g11606 ( 
.A1(n_11451),
.A2(n_1241),
.B(n_1242),
.Y(n_11606)
);

INVx1_ASAP7_75t_L g11607 ( 
.A(n_10944),
.Y(n_11607)
);

NOR2x1_ASAP7_75t_R g11608 ( 
.A(n_11471),
.B(n_1243),
.Y(n_11608)
);

OAI21xp5_ASAP7_75t_SL g11609 ( 
.A1(n_11030),
.A2(n_1243),
.B(n_1244),
.Y(n_11609)
);

OAI21x1_ASAP7_75t_L g11610 ( 
.A1(n_11347),
.A2(n_1245),
.B(n_1246),
.Y(n_11610)
);

NAND2xp5_ASAP7_75t_L g11611 ( 
.A(n_10863),
.B(n_1245),
.Y(n_11611)
);

AOI22xp33_ASAP7_75t_L g11612 ( 
.A1(n_11130),
.A2(n_1248),
.B1(n_1246),
.B2(n_1247),
.Y(n_11612)
);

NAND2xp5_ASAP7_75t_L g11613 ( 
.A(n_10893),
.B(n_1247),
.Y(n_11613)
);

OAI21x1_ASAP7_75t_L g11614 ( 
.A1(n_11254),
.A2(n_1248),
.B(n_1249),
.Y(n_11614)
);

AOI21xp5_ASAP7_75t_L g11615 ( 
.A1(n_10852),
.A2(n_1249),
.B(n_1250),
.Y(n_11615)
);

AOI21xp5_ASAP7_75t_L g11616 ( 
.A1(n_11542),
.A2(n_1250),
.B(n_1251),
.Y(n_11616)
);

AOI21x1_ASAP7_75t_SL g11617 ( 
.A1(n_11479),
.A2(n_1252),
.B(n_1253),
.Y(n_11617)
);

NOR2xp33_ASAP7_75t_L g11618 ( 
.A(n_11324),
.B(n_1252),
.Y(n_11618)
);

AOI21xp33_ASAP7_75t_L g11619 ( 
.A1(n_10981),
.A2(n_1253),
.B(n_1254),
.Y(n_11619)
);

OAI21x1_ASAP7_75t_L g11620 ( 
.A1(n_11357),
.A2(n_1255),
.B(n_1256),
.Y(n_11620)
);

AO31x2_ASAP7_75t_L g11621 ( 
.A1(n_10892),
.A2(n_1258),
.A3(n_1256),
.B(n_1257),
.Y(n_11621)
);

OAI21x1_ASAP7_75t_L g11622 ( 
.A1(n_11478),
.A2(n_1257),
.B(n_1258),
.Y(n_11622)
);

AOI21xp5_ASAP7_75t_L g11623 ( 
.A1(n_11546),
.A2(n_11551),
.B(n_11548),
.Y(n_11623)
);

AOI221x1_ASAP7_75t_L g11624 ( 
.A1(n_11491),
.A2(n_1261),
.B1(n_1259),
.B2(n_1260),
.C(n_1262),
.Y(n_11624)
);

AOI21xp5_ASAP7_75t_L g11625 ( 
.A1(n_10899),
.A2(n_1259),
.B(n_1260),
.Y(n_11625)
);

AND2x2_ASAP7_75t_L g11626 ( 
.A(n_11040),
.B(n_1261),
.Y(n_11626)
);

OAI21xp5_ASAP7_75t_L g11627 ( 
.A1(n_11495),
.A2(n_11517),
.B(n_11509),
.Y(n_11627)
);

NAND2xp5_ASAP7_75t_L g11628 ( 
.A(n_11109),
.B(n_1262),
.Y(n_11628)
);

OA21x2_ASAP7_75t_L g11629 ( 
.A1(n_11550),
.A2(n_1263),
.B(n_1264),
.Y(n_11629)
);

BUFx10_ASAP7_75t_L g11630 ( 
.A(n_10804),
.Y(n_11630)
);

AND2x2_ASAP7_75t_L g11631 ( 
.A(n_11383),
.B(n_1263),
.Y(n_11631)
);

NAND2xp5_ASAP7_75t_SL g11632 ( 
.A(n_10833),
.B(n_1265),
.Y(n_11632)
);

NAND2xp5_ASAP7_75t_L g11633 ( 
.A(n_11110),
.B(n_1265),
.Y(n_11633)
);

AO32x2_ASAP7_75t_L g11634 ( 
.A1(n_11306),
.A2(n_1268),
.A3(n_1266),
.B1(n_1267),
.B2(n_1269),
.Y(n_11634)
);

CKINVDCx16_ASAP7_75t_R g11635 ( 
.A(n_11038),
.Y(n_11635)
);

A2O1A1Ixp33_ASAP7_75t_L g11636 ( 
.A1(n_11066),
.A2(n_1268),
.B(n_1266),
.C(n_1267),
.Y(n_11636)
);

AOI21xp5_ASAP7_75t_L g11637 ( 
.A1(n_10842),
.A2(n_1269),
.B(n_1270),
.Y(n_11637)
);

AOI21xp5_ASAP7_75t_L g11638 ( 
.A1(n_10846),
.A2(n_1270),
.B(n_1271),
.Y(n_11638)
);

A2O1A1Ixp33_ASAP7_75t_L g11639 ( 
.A1(n_11078),
.A2(n_1273),
.B(n_1271),
.C(n_1272),
.Y(n_11639)
);

INVx2_ASAP7_75t_L g11640 ( 
.A(n_10912),
.Y(n_11640)
);

O2A1O1Ixp5_ASAP7_75t_L g11641 ( 
.A1(n_11197),
.A2(n_1276),
.B(n_1272),
.C(n_1275),
.Y(n_11641)
);

OAI21x1_ASAP7_75t_L g11642 ( 
.A1(n_11525),
.A2(n_1275),
.B(n_1276),
.Y(n_11642)
);

NAND2x1_ASAP7_75t_L g11643 ( 
.A(n_11384),
.B(n_1277),
.Y(n_11643)
);

NOR3xp33_ASAP7_75t_L g11644 ( 
.A(n_10961),
.B(n_1277),
.C(n_1278),
.Y(n_11644)
);

AND2x2_ASAP7_75t_L g11645 ( 
.A(n_11334),
.B(n_1278),
.Y(n_11645)
);

INVxp67_ASAP7_75t_SL g11646 ( 
.A(n_11056),
.Y(n_11646)
);

OAI21x1_ASAP7_75t_L g11647 ( 
.A1(n_11556),
.A2(n_11161),
.B(n_11122),
.Y(n_11647)
);

AOI21x1_ASAP7_75t_L g11648 ( 
.A1(n_10908),
.A2(n_1279),
.B(n_1280),
.Y(n_11648)
);

NAND2xp5_ASAP7_75t_L g11649 ( 
.A(n_11223),
.B(n_1279),
.Y(n_11649)
);

AO31x2_ASAP7_75t_L g11650 ( 
.A1(n_11422),
.A2(n_10932),
.A3(n_10927),
.B(n_11332),
.Y(n_11650)
);

NOR2xp33_ASAP7_75t_L g11651 ( 
.A(n_11266),
.B(n_1281),
.Y(n_11651)
);

OAI21x1_ASAP7_75t_L g11652 ( 
.A1(n_11178),
.A2(n_1282),
.B(n_1283),
.Y(n_11652)
);

AOI21xp5_ASAP7_75t_L g11653 ( 
.A1(n_10985),
.A2(n_1282),
.B(n_1283),
.Y(n_11653)
);

AOI21xp5_ASAP7_75t_L g11654 ( 
.A1(n_10992),
.A2(n_11011),
.B(n_11008),
.Y(n_11654)
);

OAI21x1_ASAP7_75t_L g11655 ( 
.A1(n_11179),
.A2(n_1284),
.B(n_1285),
.Y(n_11655)
);

INVx5_ASAP7_75t_L g11656 ( 
.A(n_10880),
.Y(n_11656)
);

NAND3xp33_ASAP7_75t_SL g11657 ( 
.A(n_11080),
.B(n_11292),
.C(n_10995),
.Y(n_11657)
);

AND2x2_ASAP7_75t_L g11658 ( 
.A(n_11334),
.B(n_1284),
.Y(n_11658)
);

NOR2xp67_ASAP7_75t_L g11659 ( 
.A(n_11493),
.B(n_1285),
.Y(n_11659)
);

INVx1_ASAP7_75t_L g11660 ( 
.A(n_10953),
.Y(n_11660)
);

OAI21xp5_ASAP7_75t_L g11661 ( 
.A1(n_11534),
.A2(n_1286),
.B(n_1287),
.Y(n_11661)
);

AOI22xp5_ASAP7_75t_L g11662 ( 
.A1(n_11143),
.A2(n_1289),
.B1(n_1286),
.B2(n_1288),
.Y(n_11662)
);

NOR2xp33_ASAP7_75t_L g11663 ( 
.A(n_11431),
.B(n_1289),
.Y(n_11663)
);

NAND2xp5_ASAP7_75t_L g11664 ( 
.A(n_11262),
.B(n_1290),
.Y(n_11664)
);

OAI21x1_ASAP7_75t_L g11665 ( 
.A1(n_10830),
.A2(n_1290),
.B(n_1291),
.Y(n_11665)
);

AOI21xp5_ASAP7_75t_L g11666 ( 
.A1(n_10797),
.A2(n_10984),
.B(n_10838),
.Y(n_11666)
);

INVx1_ASAP7_75t_L g11667 ( 
.A(n_10791),
.Y(n_11667)
);

AO31x2_ASAP7_75t_L g11668 ( 
.A1(n_10837),
.A2(n_1294),
.A3(n_1292),
.B(n_1293),
.Y(n_11668)
);

OAI21x1_ASAP7_75t_L g11669 ( 
.A1(n_10921),
.A2(n_1292),
.B(n_1293),
.Y(n_11669)
);

OAI21xp5_ASAP7_75t_L g11670 ( 
.A1(n_11535),
.A2(n_1294),
.B(n_1295),
.Y(n_11670)
);

O2A1O1Ixp5_ASAP7_75t_L g11671 ( 
.A1(n_10882),
.A2(n_1298),
.B(n_1296),
.C(n_1297),
.Y(n_11671)
);

AO31x2_ASAP7_75t_L g11672 ( 
.A1(n_11195),
.A2(n_1300),
.A3(n_1297),
.B(n_1299),
.Y(n_11672)
);

NAND2xp5_ASAP7_75t_L g11673 ( 
.A(n_11300),
.B(n_1299),
.Y(n_11673)
);

NAND2xp5_ASAP7_75t_L g11674 ( 
.A(n_11146),
.B(n_10874),
.Y(n_11674)
);

AOI21xp5_ASAP7_75t_L g11675 ( 
.A1(n_10870),
.A2(n_1300),
.B(n_1301),
.Y(n_11675)
);

OAI21x1_ASAP7_75t_L g11676 ( 
.A1(n_10950),
.A2(n_1302),
.B(n_1303),
.Y(n_11676)
);

INVx3_ASAP7_75t_L g11677 ( 
.A(n_10812),
.Y(n_11677)
);

OAI21x1_ASAP7_75t_L g11678 ( 
.A1(n_11518),
.A2(n_1302),
.B(n_1303),
.Y(n_11678)
);

OAI21xp5_ASAP7_75t_L g11679 ( 
.A1(n_11539),
.A2(n_1304),
.B(n_1305),
.Y(n_11679)
);

INVx1_ASAP7_75t_L g11680 ( 
.A(n_10796),
.Y(n_11680)
);

NAND2xp5_ASAP7_75t_L g11681 ( 
.A(n_10909),
.B(n_1304),
.Y(n_11681)
);

OR2x6_ASAP7_75t_L g11682 ( 
.A(n_11515),
.B(n_1305),
.Y(n_11682)
);

NAND2xp5_ASAP7_75t_L g11683 ( 
.A(n_11243),
.B(n_1306),
.Y(n_11683)
);

A2O1A1Ixp33_ASAP7_75t_L g11684 ( 
.A1(n_10844),
.A2(n_1308),
.B(n_1306),
.C(n_1307),
.Y(n_11684)
);

AOI21xp5_ASAP7_75t_L g11685 ( 
.A1(n_10831),
.A2(n_1308),
.B(n_1309),
.Y(n_11685)
);

OAI21x1_ASAP7_75t_L g11686 ( 
.A1(n_11526),
.A2(n_1309),
.B(n_1310),
.Y(n_11686)
);

NAND2xp5_ASAP7_75t_L g11687 ( 
.A(n_11248),
.B(n_1311),
.Y(n_11687)
);

BUFx3_ASAP7_75t_L g11688 ( 
.A(n_10976),
.Y(n_11688)
);

NAND2xp5_ASAP7_75t_L g11689 ( 
.A(n_11253),
.B(n_1312),
.Y(n_11689)
);

INVx2_ASAP7_75t_L g11690 ( 
.A(n_10930),
.Y(n_11690)
);

NOR2xp67_ASAP7_75t_L g11691 ( 
.A(n_11493),
.B(n_1312),
.Y(n_11691)
);

AO31x2_ASAP7_75t_L g11692 ( 
.A1(n_11212),
.A2(n_1315),
.A3(n_1313),
.B(n_1314),
.Y(n_11692)
);

NAND2xp5_ASAP7_75t_L g11693 ( 
.A(n_11264),
.B(n_1313),
.Y(n_11693)
);

INVx4_ASAP7_75t_L g11694 ( 
.A(n_10941),
.Y(n_11694)
);

INVx2_ASAP7_75t_L g11695 ( 
.A(n_10933),
.Y(n_11695)
);

INVx1_ASAP7_75t_L g11696 ( 
.A(n_10809),
.Y(n_11696)
);

AOI21x1_ASAP7_75t_L g11697 ( 
.A1(n_11482),
.A2(n_1314),
.B(n_1315),
.Y(n_11697)
);

AO21x1_ASAP7_75t_L g11698 ( 
.A1(n_11231),
.A2(n_1316),
.B(n_1318),
.Y(n_11698)
);

HB1xp67_ASAP7_75t_L g11699 ( 
.A(n_10966),
.Y(n_11699)
);

NAND2xp5_ASAP7_75t_SL g11700 ( 
.A(n_10833),
.B(n_1318),
.Y(n_11700)
);

OAI22xp5_ASAP7_75t_L g11701 ( 
.A1(n_10824),
.A2(n_1322),
.B1(n_1320),
.B2(n_1321),
.Y(n_11701)
);

OAI21xp5_ASAP7_75t_L g11702 ( 
.A1(n_11554),
.A2(n_1321),
.B(n_1322),
.Y(n_11702)
);

NOR2xp33_ASAP7_75t_L g11703 ( 
.A(n_11431),
.B(n_1323),
.Y(n_11703)
);

AOI21xp5_ASAP7_75t_L g11704 ( 
.A1(n_10883),
.A2(n_1323),
.B(n_1324),
.Y(n_11704)
);

NAND2xp5_ASAP7_75t_L g11705 ( 
.A(n_11272),
.B(n_1325),
.Y(n_11705)
);

CKINVDCx20_ASAP7_75t_R g11706 ( 
.A(n_10916),
.Y(n_11706)
);

INVx2_ASAP7_75t_L g11707 ( 
.A(n_10975),
.Y(n_11707)
);

NAND2xp5_ASAP7_75t_L g11708 ( 
.A(n_11299),
.B(n_1325),
.Y(n_11708)
);

INVx2_ASAP7_75t_L g11709 ( 
.A(n_10991),
.Y(n_11709)
);

NAND2xp5_ASAP7_75t_L g11710 ( 
.A(n_11188),
.B(n_1327),
.Y(n_11710)
);

NAND2xp5_ASAP7_75t_L g11711 ( 
.A(n_11203),
.B(n_1327),
.Y(n_11711)
);

INVx1_ASAP7_75t_L g11712 ( 
.A(n_10818),
.Y(n_11712)
);

NAND3x1_ASAP7_75t_L g11713 ( 
.A(n_11169),
.B(n_1328),
.C(n_1329),
.Y(n_11713)
);

NAND2xp5_ASAP7_75t_SL g11714 ( 
.A(n_11260),
.B(n_1328),
.Y(n_11714)
);

AOI21xp5_ASAP7_75t_L g11715 ( 
.A1(n_11494),
.A2(n_1329),
.B(n_1330),
.Y(n_11715)
);

AND2x4_ASAP7_75t_L g11716 ( 
.A(n_11067),
.B(n_1330),
.Y(n_11716)
);

NAND2xp5_ASAP7_75t_L g11717 ( 
.A(n_11242),
.B(n_1331),
.Y(n_11717)
);

OAI21x1_ASAP7_75t_L g11718 ( 
.A1(n_11468),
.A2(n_1331),
.B(n_1332),
.Y(n_11718)
);

AOI21xp5_ASAP7_75t_L g11719 ( 
.A1(n_11533),
.A2(n_11488),
.B(n_11484),
.Y(n_11719)
);

NAND2xp5_ASAP7_75t_L g11720 ( 
.A(n_10996),
.B(n_1332),
.Y(n_11720)
);

BUFx2_ASAP7_75t_L g11721 ( 
.A(n_11285),
.Y(n_11721)
);

BUFx6f_ASAP7_75t_L g11722 ( 
.A(n_10817),
.Y(n_11722)
);

AO31x2_ASAP7_75t_L g11723 ( 
.A1(n_11213),
.A2(n_1335),
.A3(n_1333),
.B(n_1334),
.Y(n_11723)
);

OAI21x1_ASAP7_75t_L g11724 ( 
.A1(n_11060),
.A2(n_11470),
.B(n_11444),
.Y(n_11724)
);

OAI21x1_ASAP7_75t_L g11725 ( 
.A1(n_11249),
.A2(n_1333),
.B(n_1334),
.Y(n_11725)
);

INVx1_ASAP7_75t_L g11726 ( 
.A(n_10828),
.Y(n_11726)
);

INVx1_ASAP7_75t_L g11727 ( 
.A(n_10836),
.Y(n_11727)
);

AOI21xp5_ASAP7_75t_L g11728 ( 
.A1(n_11504),
.A2(n_1335),
.B(n_1336),
.Y(n_11728)
);

OAI21x1_ASAP7_75t_L g11729 ( 
.A1(n_11455),
.A2(n_1337),
.B(n_1338),
.Y(n_11729)
);

INVx1_ASAP7_75t_L g11730 ( 
.A(n_10841),
.Y(n_11730)
);

NAND2xp5_ASAP7_75t_L g11731 ( 
.A(n_11007),
.B(n_1337),
.Y(n_11731)
);

BUFx8_ASAP7_75t_L g11732 ( 
.A(n_11020),
.Y(n_11732)
);

INVx4_ASAP7_75t_L g11733 ( 
.A(n_11480),
.Y(n_11733)
);

OAI21xp5_ASAP7_75t_L g11734 ( 
.A1(n_11557),
.A2(n_11558),
.B(n_10850),
.Y(n_11734)
);

BUFx6f_ASAP7_75t_L g11735 ( 
.A(n_10817),
.Y(n_11735)
);

AOI21xp5_ASAP7_75t_L g11736 ( 
.A1(n_11503),
.A2(n_1338),
.B(n_1339),
.Y(n_11736)
);

BUFx3_ASAP7_75t_L g11737 ( 
.A(n_11014),
.Y(n_11737)
);

AND2x2_ASAP7_75t_L g11738 ( 
.A(n_11335),
.B(n_1339),
.Y(n_11738)
);

OAI21x1_ASAP7_75t_L g11739 ( 
.A1(n_10965),
.A2(n_1340),
.B(n_1341),
.Y(n_11739)
);

OAI21x1_ASAP7_75t_SL g11740 ( 
.A1(n_11322),
.A2(n_1341),
.B(n_1342),
.Y(n_11740)
);

INVx2_ASAP7_75t_L g11741 ( 
.A(n_11012),
.Y(n_11741)
);

AOI221xp5_ASAP7_75t_L g11742 ( 
.A1(n_10798),
.A2(n_1344),
.B1(n_1342),
.B2(n_1343),
.C(n_1345),
.Y(n_11742)
);

NAND2x1_ASAP7_75t_L g11743 ( 
.A(n_11384),
.B(n_1343),
.Y(n_11743)
);

AOI21xp5_ASAP7_75t_L g11744 ( 
.A1(n_11528),
.A2(n_1344),
.B(n_1346),
.Y(n_11744)
);

NAND2xp5_ASAP7_75t_L g11745 ( 
.A(n_11015),
.B(n_1346),
.Y(n_11745)
);

INVx2_ASAP7_75t_SL g11746 ( 
.A(n_11194),
.Y(n_11746)
);

OAI21x1_ASAP7_75t_L g11747 ( 
.A1(n_11133),
.A2(n_1347),
.B(n_1348),
.Y(n_11747)
);

AOI21xp5_ASAP7_75t_L g11748 ( 
.A1(n_11507),
.A2(n_1348),
.B(n_1349),
.Y(n_11748)
);

OAI22xp5_ASAP7_75t_L g11749 ( 
.A1(n_10886),
.A2(n_1351),
.B1(n_1349),
.B2(n_1350),
.Y(n_11749)
);

INVx4_ASAP7_75t_L g11750 ( 
.A(n_11513),
.Y(n_11750)
);

NAND2xp5_ASAP7_75t_L g11751 ( 
.A(n_11021),
.B(n_1350),
.Y(n_11751)
);

OAI21xp5_ASAP7_75t_L g11752 ( 
.A1(n_10945),
.A2(n_1351),
.B(n_1352),
.Y(n_11752)
);

NOR2xp67_ASAP7_75t_SL g11753 ( 
.A(n_11541),
.B(n_1353),
.Y(n_11753)
);

INVx2_ASAP7_75t_L g11754 ( 
.A(n_10875),
.Y(n_11754)
);

AOI21xp5_ASAP7_75t_L g11755 ( 
.A1(n_11544),
.A2(n_1353),
.B(n_1354),
.Y(n_11755)
);

NAND2xp5_ASAP7_75t_L g11756 ( 
.A(n_11259),
.B(n_1354),
.Y(n_11756)
);

NAND3xp33_ASAP7_75t_SL g11757 ( 
.A(n_11241),
.B(n_1355),
.C(n_1356),
.Y(n_11757)
);

AOI21xp5_ASAP7_75t_L g11758 ( 
.A1(n_11521),
.A2(n_1357),
.B(n_1358),
.Y(n_11758)
);

OA21x2_ASAP7_75t_L g11759 ( 
.A1(n_11536),
.A2(n_1357),
.B(n_1358),
.Y(n_11759)
);

AO31x2_ASAP7_75t_L g11760 ( 
.A1(n_10864),
.A2(n_1361),
.A3(n_1359),
.B(n_1360),
.Y(n_11760)
);

NAND2xp5_ASAP7_75t_L g11761 ( 
.A(n_11307),
.B(n_1360),
.Y(n_11761)
);

AO21x2_ASAP7_75t_L g11762 ( 
.A1(n_11543),
.A2(n_1361),
.B(n_1362),
.Y(n_11762)
);

OA22x2_ASAP7_75t_L g11763 ( 
.A1(n_10960),
.A2(n_1364),
.B1(n_1362),
.B2(n_1363),
.Y(n_11763)
);

OAI21x1_ASAP7_75t_L g11764 ( 
.A1(n_11529),
.A2(n_1363),
.B(n_1365),
.Y(n_11764)
);

INVx2_ASAP7_75t_L g11765 ( 
.A(n_10843),
.Y(n_11765)
);

NAND2xp5_ASAP7_75t_SL g11766 ( 
.A(n_11411),
.B(n_1366),
.Y(n_11766)
);

NAND2xp5_ASAP7_75t_L g11767 ( 
.A(n_11309),
.B(n_1366),
.Y(n_11767)
);

AND2x6_ASAP7_75t_L g11768 ( 
.A(n_11419),
.B(n_1367),
.Y(n_11768)
);

OAI22xp5_ASAP7_75t_L g11769 ( 
.A1(n_11024),
.A2(n_1370),
.B1(n_1368),
.B2(n_1369),
.Y(n_11769)
);

AND3x4_ASAP7_75t_L g11770 ( 
.A(n_11267),
.B(n_1368),
.C(n_1369),
.Y(n_11770)
);

NOR2x1_ASAP7_75t_L g11771 ( 
.A(n_11003),
.B(n_1370),
.Y(n_11771)
);

HB1xp67_ASAP7_75t_L g11772 ( 
.A(n_10853),
.Y(n_11772)
);

NAND2xp5_ASAP7_75t_L g11773 ( 
.A(n_11368),
.B(n_1371),
.Y(n_11773)
);

INVx1_ASAP7_75t_L g11774 ( 
.A(n_10859),
.Y(n_11774)
);

AND2x2_ASAP7_75t_L g11775 ( 
.A(n_11312),
.B(n_1371),
.Y(n_11775)
);

INVx4_ASAP7_75t_L g11776 ( 
.A(n_10971),
.Y(n_11776)
);

OAI21x1_ASAP7_75t_L g11777 ( 
.A1(n_11537),
.A2(n_1372),
.B(n_1373),
.Y(n_11777)
);

INVx1_ASAP7_75t_L g11778 ( 
.A(n_10876),
.Y(n_11778)
);

OAI21x1_ASAP7_75t_L g11779 ( 
.A1(n_11547),
.A2(n_1372),
.B(n_1374),
.Y(n_11779)
);

AOI21xp5_ASAP7_75t_L g11780 ( 
.A1(n_11549),
.A2(n_1374),
.B(n_1375),
.Y(n_11780)
);

NAND2xp5_ASAP7_75t_L g11781 ( 
.A(n_11314),
.B(n_1375),
.Y(n_11781)
);

NOR2x1_ASAP7_75t_SL g11782 ( 
.A(n_11177),
.B(n_1376),
.Y(n_11782)
);

INVx2_ASAP7_75t_SL g11783 ( 
.A(n_11220),
.Y(n_11783)
);

AOI21xp5_ASAP7_75t_L g11784 ( 
.A1(n_10847),
.A2(n_1377),
.B(n_1378),
.Y(n_11784)
);

INVx2_ASAP7_75t_L g11785 ( 
.A(n_10889),
.Y(n_11785)
);

NAND2x1_ASAP7_75t_L g11786 ( 
.A(n_11298),
.B(n_1377),
.Y(n_11786)
);

NOR2xp67_ASAP7_75t_L g11787 ( 
.A(n_11228),
.B(n_1378),
.Y(n_11787)
);

NOR2xp33_ASAP7_75t_L g11788 ( 
.A(n_11336),
.B(n_1379),
.Y(n_11788)
);

OAI21x1_ASAP7_75t_L g11789 ( 
.A1(n_10877),
.A2(n_1380),
.B(n_1381),
.Y(n_11789)
);

AOI21x1_ASAP7_75t_SL g11790 ( 
.A1(n_11392),
.A2(n_1380),
.B(n_1381),
.Y(n_11790)
);

OAI21x1_ASAP7_75t_L g11791 ( 
.A1(n_11420),
.A2(n_1382),
.B(n_1383),
.Y(n_11791)
);

AO31x2_ASAP7_75t_L g11792 ( 
.A1(n_11126),
.A2(n_1384),
.A3(n_1382),
.B(n_1383),
.Y(n_11792)
);

OAI21x1_ASAP7_75t_L g11793 ( 
.A1(n_11193),
.A2(n_1385),
.B(n_1386),
.Y(n_11793)
);

OAI21xp33_ASAP7_75t_L g11794 ( 
.A1(n_11380),
.A2(n_1385),
.B(n_1387),
.Y(n_11794)
);

OAI22xp5_ASAP7_75t_L g11795 ( 
.A1(n_11103),
.A2(n_1389),
.B1(n_1387),
.B2(n_1388),
.Y(n_11795)
);

NAND3xp33_ASAP7_75t_L g11796 ( 
.A(n_11148),
.B(n_1388),
.C(n_1389),
.Y(n_11796)
);

OAI21x1_ASAP7_75t_L g11797 ( 
.A1(n_10947),
.A2(n_1390),
.B(n_1391),
.Y(n_11797)
);

INVx2_ASAP7_75t_SL g11798 ( 
.A(n_11247),
.Y(n_11798)
);

OAI21xp33_ASAP7_75t_L g11799 ( 
.A1(n_10884),
.A2(n_1391),
.B(n_1392),
.Y(n_11799)
);

AO31x2_ASAP7_75t_L g11800 ( 
.A1(n_10958),
.A2(n_1394),
.A3(n_1392),
.B(n_1393),
.Y(n_11800)
);

NAND3xp33_ASAP7_75t_L g11801 ( 
.A(n_11353),
.B(n_11395),
.C(n_11359),
.Y(n_11801)
);

OAI21x1_ASAP7_75t_L g11802 ( 
.A1(n_10955),
.A2(n_1393),
.B(n_1395),
.Y(n_11802)
);

AO31x2_ASAP7_75t_L g11803 ( 
.A1(n_10974),
.A2(n_1397),
.A3(n_1395),
.B(n_1396),
.Y(n_11803)
);

AO21x2_ASAP7_75t_L g11804 ( 
.A1(n_11258),
.A2(n_1396),
.B(n_1398),
.Y(n_11804)
);

OAI21xp33_ASAP7_75t_L g11805 ( 
.A1(n_11416),
.A2(n_1398),
.B(n_1400),
.Y(n_11805)
);

AOI21xp5_ASAP7_75t_L g11806 ( 
.A1(n_10867),
.A2(n_1400),
.B(n_1401),
.Y(n_11806)
);

A2O1A1Ixp33_ASAP7_75t_L g11807 ( 
.A1(n_10922),
.A2(n_1403),
.B(n_1401),
.C(n_1402),
.Y(n_11807)
);

NAND2xp5_ASAP7_75t_L g11808 ( 
.A(n_11303),
.B(n_1402),
.Y(n_11808)
);

AO31x2_ASAP7_75t_L g11809 ( 
.A1(n_11074),
.A2(n_1405),
.A3(n_1403),
.B(n_1404),
.Y(n_11809)
);

INVx2_ASAP7_75t_L g11810 ( 
.A(n_10890),
.Y(n_11810)
);

OAI22xp5_ASAP7_75t_L g11811 ( 
.A1(n_11142),
.A2(n_1407),
.B1(n_1404),
.B2(n_1406),
.Y(n_11811)
);

NAND2xp5_ASAP7_75t_L g11812 ( 
.A(n_11043),
.B(n_1406),
.Y(n_11812)
);

BUFx8_ASAP7_75t_SL g11813 ( 
.A(n_10806),
.Y(n_11813)
);

AOI21xp5_ASAP7_75t_L g11814 ( 
.A1(n_11439),
.A2(n_1408),
.B(n_1409),
.Y(n_11814)
);

BUFx6f_ASAP7_75t_L g11815 ( 
.A(n_10871),
.Y(n_11815)
);

OAI21x1_ASAP7_75t_L g11816 ( 
.A1(n_10811),
.A2(n_1408),
.B(n_1409),
.Y(n_11816)
);

OAI21xp5_ASAP7_75t_L g11817 ( 
.A1(n_11013),
.A2(n_1410),
.B(n_1411),
.Y(n_11817)
);

OAI21x1_ASAP7_75t_L g11818 ( 
.A1(n_10943),
.A2(n_1410),
.B(n_1411),
.Y(n_11818)
);

AND2x2_ASAP7_75t_L g11819 ( 
.A(n_11222),
.B(n_1412),
.Y(n_11819)
);

A2O1A1Ixp33_ASAP7_75t_L g11820 ( 
.A1(n_10938),
.A2(n_10952),
.B(n_11093),
.C(n_11129),
.Y(n_11820)
);

NAND2xp5_ASAP7_75t_L g11821 ( 
.A(n_11057),
.B(n_1412),
.Y(n_11821)
);

NAND2xp5_ASAP7_75t_L g11822 ( 
.A(n_11063),
.B(n_1413),
.Y(n_11822)
);

AOI21xp5_ASAP7_75t_L g11823 ( 
.A1(n_11385),
.A2(n_1413),
.B(n_1414),
.Y(n_11823)
);

AOI22xp5_ASAP7_75t_L g11824 ( 
.A1(n_11032),
.A2(n_1416),
.B1(n_1414),
.B2(n_1415),
.Y(n_11824)
);

NAND2xp5_ASAP7_75t_L g11825 ( 
.A(n_11085),
.B(n_1415),
.Y(n_11825)
);

BUFx3_ASAP7_75t_L g11826 ( 
.A(n_11082),
.Y(n_11826)
);

NAND2xp5_ASAP7_75t_L g11827 ( 
.A(n_11096),
.B(n_1416),
.Y(n_11827)
);

INVx2_ASAP7_75t_L g11828 ( 
.A(n_10904),
.Y(n_11828)
);

BUFx3_ASAP7_75t_L g11829 ( 
.A(n_11100),
.Y(n_11829)
);

AOI21xp5_ASAP7_75t_L g11830 ( 
.A1(n_11414),
.A2(n_1417),
.B(n_1419),
.Y(n_11830)
);

AO31x2_ASAP7_75t_L g11831 ( 
.A1(n_11106),
.A2(n_1422),
.A3(n_1419),
.B(n_1421),
.Y(n_11831)
);

NAND2x1_ASAP7_75t_L g11832 ( 
.A(n_11037),
.B(n_11051),
.Y(n_11832)
);

INVx2_ASAP7_75t_L g11833 ( 
.A(n_10914),
.Y(n_11833)
);

INVx1_ASAP7_75t_L g11834 ( 
.A(n_10942),
.Y(n_11834)
);

AOI21x1_ASAP7_75t_L g11835 ( 
.A1(n_10939),
.A2(n_1421),
.B(n_1422),
.Y(n_11835)
);

AOI21x1_ASAP7_75t_L g11836 ( 
.A1(n_11209),
.A2(n_1423),
.B(n_1424),
.Y(n_11836)
);

CKINVDCx5p33_ASAP7_75t_R g11837 ( 
.A(n_11028),
.Y(n_11837)
);

OAI21x1_ASAP7_75t_L g11838 ( 
.A1(n_11025),
.A2(n_10799),
.B(n_10814),
.Y(n_11838)
);

OAI21x1_ASAP7_75t_SL g11839 ( 
.A1(n_11044),
.A2(n_11369),
.B(n_11363),
.Y(n_11839)
);

A2O1A1Ixp33_ASAP7_75t_L g11840 ( 
.A1(n_11134),
.A2(n_11427),
.B(n_11464),
.C(n_11321),
.Y(n_11840)
);

OAI21x1_ASAP7_75t_L g11841 ( 
.A1(n_11374),
.A2(n_1423),
.B(n_1424),
.Y(n_11841)
);

OAI21x1_ASAP7_75t_L g11842 ( 
.A1(n_11375),
.A2(n_1425),
.B(n_1426),
.Y(n_11842)
);

OAI21xp5_ASAP7_75t_L g11843 ( 
.A1(n_11295),
.A2(n_1426),
.B(n_1427),
.Y(n_11843)
);

NAND2xp5_ASAP7_75t_SL g11844 ( 
.A(n_11411),
.B(n_1427),
.Y(n_11844)
);

BUFx2_ASAP7_75t_L g11845 ( 
.A(n_11211),
.Y(n_11845)
);

OAI21x1_ASAP7_75t_L g11846 ( 
.A1(n_11396),
.A2(n_11398),
.B(n_11397),
.Y(n_11846)
);

OAI21x1_ASAP7_75t_L g11847 ( 
.A1(n_11401),
.A2(n_1428),
.B(n_1429),
.Y(n_11847)
);

AOI221x1_ASAP7_75t_L g11848 ( 
.A1(n_11230),
.A2(n_1430),
.B1(n_1428),
.B2(n_1429),
.C(n_1431),
.Y(n_11848)
);

AOI21x1_ASAP7_75t_L g11849 ( 
.A1(n_11238),
.A2(n_1432),
.B(n_1434),
.Y(n_11849)
);

NAND2xp5_ASAP7_75t_L g11850 ( 
.A(n_11097),
.B(n_1434),
.Y(n_11850)
);

OAI21x1_ASAP7_75t_L g11851 ( 
.A1(n_11409),
.A2(n_1435),
.B(n_1436),
.Y(n_11851)
);

OAI21xp5_ASAP7_75t_L g11852 ( 
.A1(n_11315),
.A2(n_1437),
.B(n_1438),
.Y(n_11852)
);

INVx2_ASAP7_75t_L g11853 ( 
.A(n_10954),
.Y(n_11853)
);

OA21x2_ASAP7_75t_L g11854 ( 
.A1(n_10887),
.A2(n_1437),
.B(n_1438),
.Y(n_11854)
);

OAI21x1_ASAP7_75t_L g11855 ( 
.A1(n_11343),
.A2(n_1439),
.B(n_1440),
.Y(n_11855)
);

OAI21xp33_ASAP7_75t_L g11856 ( 
.A1(n_10902),
.A2(n_1439),
.B(n_1440),
.Y(n_11856)
);

NAND2xp5_ASAP7_75t_L g11857 ( 
.A(n_10970),
.B(n_1441),
.Y(n_11857)
);

NAND2xp5_ASAP7_75t_L g11858 ( 
.A(n_10979),
.B(n_1442),
.Y(n_11858)
);

AOI21xp5_ASAP7_75t_L g11859 ( 
.A1(n_11502),
.A2(n_1443),
.B(n_1444),
.Y(n_11859)
);

BUFx2_ASAP7_75t_L g11860 ( 
.A(n_10969),
.Y(n_11860)
);

OAI21x1_ASAP7_75t_L g11861 ( 
.A1(n_11351),
.A2(n_1443),
.B(n_1444),
.Y(n_11861)
);

NAND2xp5_ASAP7_75t_L g11862 ( 
.A(n_10987),
.B(n_1445),
.Y(n_11862)
);

NAND2xp5_ASAP7_75t_L g11863 ( 
.A(n_11000),
.B(n_1445),
.Y(n_11863)
);

AOI21xp5_ASAP7_75t_L g11864 ( 
.A1(n_11523),
.A2(n_1446),
.B(n_1447),
.Y(n_11864)
);

NAND2xp5_ASAP7_75t_L g11865 ( 
.A(n_11022),
.B(n_1446),
.Y(n_11865)
);

OAI21x1_ASAP7_75t_L g11866 ( 
.A1(n_11358),
.A2(n_11371),
.B(n_11361),
.Y(n_11866)
);

OAI21xp5_ASAP7_75t_L g11867 ( 
.A1(n_11373),
.A2(n_1447),
.B(n_1448),
.Y(n_11867)
);

CKINVDCx5p33_ASAP7_75t_R g11868 ( 
.A(n_10999),
.Y(n_11868)
);

BUFx12f_ASAP7_75t_L g11869 ( 
.A(n_11081),
.Y(n_11869)
);

A2O1A1Ixp33_ASAP7_75t_L g11870 ( 
.A1(n_11119),
.A2(n_1451),
.B(n_1449),
.C(n_1450),
.Y(n_11870)
);

NAND2xp5_ASAP7_75t_L g11871 ( 
.A(n_11487),
.B(n_11505),
.Y(n_11871)
);

OAI22xp5_ASAP7_75t_L g11872 ( 
.A1(n_10873),
.A2(n_1452),
.B1(n_1449),
.B2(n_1451),
.Y(n_11872)
);

OAI22xp5_ASAP7_75t_L g11873 ( 
.A1(n_10905),
.A2(n_1454),
.B1(n_1452),
.B2(n_1453),
.Y(n_11873)
);

AO21x2_ASAP7_75t_L g11874 ( 
.A1(n_10895),
.A2(n_1453),
.B(n_1454),
.Y(n_11874)
);

NAND2xp5_ASAP7_75t_L g11875 ( 
.A(n_11538),
.B(n_1455),
.Y(n_11875)
);

NAND2xp5_ASAP7_75t_L g11876 ( 
.A(n_11540),
.B(n_1455),
.Y(n_11876)
);

A2O1A1Ixp33_ASAP7_75t_L g11877 ( 
.A1(n_10936),
.A2(n_1458),
.B(n_1456),
.C(n_1457),
.Y(n_11877)
);

NAND2xp5_ASAP7_75t_L g11878 ( 
.A(n_11553),
.B(n_1457),
.Y(n_11878)
);

NOR2xp33_ASAP7_75t_L g11879 ( 
.A(n_11425),
.B(n_1458),
.Y(n_11879)
);

INVx1_ASAP7_75t_L g11880 ( 
.A(n_10834),
.Y(n_11880)
);

INVx2_ASAP7_75t_L g11881 ( 
.A(n_10868),
.Y(n_11881)
);

INVx1_ASAP7_75t_L g11882 ( 
.A(n_11477),
.Y(n_11882)
);

NAND2xp5_ASAP7_75t_L g11883 ( 
.A(n_11004),
.B(n_1459),
.Y(n_11883)
);

OAI21x1_ASAP7_75t_L g11884 ( 
.A1(n_11273),
.A2(n_1459),
.B(n_1460),
.Y(n_11884)
);

NAND2xp5_ASAP7_75t_SL g11885 ( 
.A(n_11408),
.B(n_1460),
.Y(n_11885)
);

NAND2x1_ASAP7_75t_L g11886 ( 
.A(n_11061),
.B(n_1461),
.Y(n_11886)
);

INVx2_ASAP7_75t_L g11887 ( 
.A(n_11522),
.Y(n_11887)
);

NAND2xp5_ASAP7_75t_L g11888 ( 
.A(n_11532),
.B(n_1461),
.Y(n_11888)
);

OAI21x1_ASAP7_75t_L g11889 ( 
.A1(n_11437),
.A2(n_1462),
.B(n_1463),
.Y(n_11889)
);

AO31x2_ASAP7_75t_L g11890 ( 
.A1(n_11114),
.A2(n_1465),
.A3(n_1463),
.B(n_1464),
.Y(n_11890)
);

A2O1A1Ixp33_ASAP7_75t_L g11891 ( 
.A1(n_11463),
.A2(n_1466),
.B(n_1464),
.C(n_1465),
.Y(n_11891)
);

AOI21xp5_ASAP7_75t_L g11892 ( 
.A1(n_10990),
.A2(n_1466),
.B(n_1467),
.Y(n_11892)
);

INVx1_ASAP7_75t_L g11893 ( 
.A(n_11068),
.Y(n_11893)
);

NAND2xp5_ASAP7_75t_L g11894 ( 
.A(n_11280),
.B(n_1467),
.Y(n_11894)
);

INVx1_ASAP7_75t_L g11895 ( 
.A(n_10825),
.Y(n_11895)
);

OAI21x1_ASAP7_75t_L g11896 ( 
.A1(n_11442),
.A2(n_1468),
.B(n_1469),
.Y(n_11896)
);

NAND2xp5_ASAP7_75t_L g11897 ( 
.A(n_11302),
.B(n_1468),
.Y(n_11897)
);

OAI21x1_ASAP7_75t_SL g11898 ( 
.A1(n_11289),
.A2(n_1469),
.B(n_1470),
.Y(n_11898)
);

NAND2xp5_ASAP7_75t_L g11899 ( 
.A(n_11201),
.B(n_1470),
.Y(n_11899)
);

O2A1O1Ixp5_ASAP7_75t_L g11900 ( 
.A1(n_10919),
.A2(n_11117),
.B(n_10926),
.C(n_11018),
.Y(n_11900)
);

INVx1_ASAP7_75t_L g11901 ( 
.A(n_10790),
.Y(n_11901)
);

OAI21x1_ASAP7_75t_L g11902 ( 
.A1(n_11426),
.A2(n_1471),
.B(n_1472),
.Y(n_11902)
);

NOR2xp33_ASAP7_75t_L g11903 ( 
.A(n_11501),
.B(n_1471),
.Y(n_11903)
);

BUFx6f_ASAP7_75t_L g11904 ( 
.A(n_10871),
.Y(n_11904)
);

AND2x2_ASAP7_75t_L g11905 ( 
.A(n_11338),
.B(n_1472),
.Y(n_11905)
);

NAND2xp5_ASAP7_75t_L g11906 ( 
.A(n_11200),
.B(n_1473),
.Y(n_11906)
);

AND2x2_ASAP7_75t_L g11907 ( 
.A(n_10872),
.B(n_1473),
.Y(n_11907)
);

AO31x2_ASAP7_75t_L g11908 ( 
.A1(n_10998),
.A2(n_1476),
.A3(n_1474),
.B(n_1475),
.Y(n_11908)
);

OAI21x1_ASAP7_75t_L g11909 ( 
.A1(n_11308),
.A2(n_1475),
.B(n_1476),
.Y(n_11909)
);

OAI21x1_ASAP7_75t_L g11910 ( 
.A1(n_11297),
.A2(n_1477),
.B(n_1478),
.Y(n_11910)
);

AOI21xp5_ASAP7_75t_L g11911 ( 
.A1(n_10925),
.A2(n_1477),
.B(n_1478),
.Y(n_11911)
);

INVx1_ASAP7_75t_SL g11912 ( 
.A(n_10988),
.Y(n_11912)
);

AO21x1_ASAP7_75t_L g11913 ( 
.A1(n_11274),
.A2(n_1479),
.B(n_1480),
.Y(n_11913)
);

BUFx6f_ASAP7_75t_L g11914 ( 
.A(n_10937),
.Y(n_11914)
);

AO31x2_ASAP7_75t_L g11915 ( 
.A1(n_11029),
.A2(n_1482),
.A3(n_1480),
.B(n_1481),
.Y(n_11915)
);

AOI21xp5_ASAP7_75t_L g11916 ( 
.A1(n_11318),
.A2(n_1481),
.B(n_1482),
.Y(n_11916)
);

AOI21xp5_ASAP7_75t_L g11917 ( 
.A1(n_11402),
.A2(n_1483),
.B(n_1484),
.Y(n_11917)
);

INVx1_ASAP7_75t_L g11918 ( 
.A(n_10827),
.Y(n_11918)
);

OAI21xp5_ASAP7_75t_L g11919 ( 
.A1(n_11459),
.A2(n_1483),
.B(n_1484),
.Y(n_11919)
);

OAI21x1_ASAP7_75t_L g11920 ( 
.A1(n_11387),
.A2(n_11417),
.B(n_11124),
.Y(n_11920)
);

NAND2xp5_ASAP7_75t_L g11921 ( 
.A(n_10801),
.B(n_1485),
.Y(n_11921)
);

OAI21xp33_ASAP7_75t_L g11922 ( 
.A1(n_10951),
.A2(n_1486),
.B(n_1487),
.Y(n_11922)
);

HB1xp67_ASAP7_75t_L g11923 ( 
.A(n_11360),
.Y(n_11923)
);

NOR2xp33_ASAP7_75t_L g11924 ( 
.A(n_11404),
.B(n_1486),
.Y(n_11924)
);

INVx3_ASAP7_75t_L g11925 ( 
.A(n_10971),
.Y(n_11925)
);

AOI221x1_ASAP7_75t_L g11926 ( 
.A1(n_10901),
.A2(n_1489),
.B1(n_1487),
.B2(n_1488),
.C(n_1490),
.Y(n_11926)
);

NAND2xp5_ASAP7_75t_L g11927 ( 
.A(n_10819),
.B(n_1488),
.Y(n_11927)
);

NAND2xp5_ASAP7_75t_L g11928 ( 
.A(n_10829),
.B(n_1489),
.Y(n_11928)
);

AOI211x1_ASAP7_75t_L g11929 ( 
.A1(n_11561),
.A2(n_1493),
.B(n_1491),
.C(n_1492),
.Y(n_11929)
);

INVx1_ASAP7_75t_L g11930 ( 
.A(n_10815),
.Y(n_11930)
);

AOI21x1_ASAP7_75t_L g11931 ( 
.A1(n_11281),
.A2(n_1491),
.B(n_1493),
.Y(n_11931)
);

NOR2xp33_ASAP7_75t_L g11932 ( 
.A(n_11378),
.B(n_1494),
.Y(n_11932)
);

AO31x2_ASAP7_75t_L g11933 ( 
.A1(n_11474),
.A2(n_11496),
.A3(n_11508),
.B(n_11499),
.Y(n_11933)
);

OAI22xp5_ASAP7_75t_L g11934 ( 
.A1(n_11111),
.A2(n_1496),
.B1(n_1494),
.B2(n_1495),
.Y(n_11934)
);

CKINVDCx5p33_ASAP7_75t_R g11935 ( 
.A(n_10928),
.Y(n_11935)
);

AOI21xp33_ASAP7_75t_L g11936 ( 
.A1(n_11403),
.A2(n_1496),
.B(n_1497),
.Y(n_11936)
);

OAI21xp5_ASAP7_75t_L g11937 ( 
.A1(n_11083),
.A2(n_1497),
.B(n_1498),
.Y(n_11937)
);

OAI21x1_ASAP7_75t_L g11938 ( 
.A1(n_11087),
.A2(n_1498),
.B(n_1499),
.Y(n_11938)
);

INVx5_ASAP7_75t_L g11939 ( 
.A(n_11076),
.Y(n_11939)
);

OAI21x1_ASAP7_75t_L g11940 ( 
.A1(n_11135),
.A2(n_1499),
.B(n_1500),
.Y(n_11940)
);

NAND2xp5_ASAP7_75t_L g11941 ( 
.A(n_11345),
.B(n_1500),
.Y(n_11941)
);

AOI21xp5_ASAP7_75t_L g11942 ( 
.A1(n_11457),
.A2(n_1501),
.B(n_1502),
.Y(n_11942)
);

BUFx10_ASAP7_75t_L g11943 ( 
.A(n_11145),
.Y(n_11943)
);

NAND2xp5_ASAP7_75t_L g11944 ( 
.A(n_10885),
.B(n_1501),
.Y(n_11944)
);

AOI21xp5_ASAP7_75t_L g11945 ( 
.A1(n_11327),
.A2(n_1502),
.B(n_1503),
.Y(n_11945)
);

INVx2_ASAP7_75t_L g11946 ( 
.A(n_10862),
.Y(n_11946)
);

BUFx3_ASAP7_75t_L g11947 ( 
.A(n_10810),
.Y(n_11947)
);

AO31x2_ASAP7_75t_L g11948 ( 
.A1(n_11512),
.A2(n_11560),
.A3(n_11102),
.B(n_11430),
.Y(n_11948)
);

AOI21xp5_ASAP7_75t_L g11949 ( 
.A1(n_11316),
.A2(n_1504),
.B(n_1506),
.Y(n_11949)
);

OAI21x1_ASAP7_75t_L g11950 ( 
.A1(n_11138),
.A2(n_1506),
.B(n_1507),
.Y(n_11950)
);

NAND2xp5_ASAP7_75t_L g11951 ( 
.A(n_10865),
.B(n_1508),
.Y(n_11951)
);

AND2x2_ASAP7_75t_L g11952 ( 
.A(n_11372),
.B(n_1508),
.Y(n_11952)
);

OAI21x1_ASAP7_75t_L g11953 ( 
.A1(n_11153),
.A2(n_1509),
.B(n_1510),
.Y(n_11953)
);

AOI21xp33_ASAP7_75t_L g11954 ( 
.A1(n_11448),
.A2(n_1509),
.B(n_1510),
.Y(n_11954)
);

NAND2xp5_ASAP7_75t_L g11955 ( 
.A(n_11399),
.B(n_11386),
.Y(n_11955)
);

BUFx3_ASAP7_75t_L g11956 ( 
.A(n_10924),
.Y(n_11956)
);

OAI21x1_ASAP7_75t_L g11957 ( 
.A1(n_11163),
.A2(n_1511),
.B(n_1512),
.Y(n_11957)
);

OAI21x1_ASAP7_75t_L g11958 ( 
.A1(n_11166),
.A2(n_1512),
.B(n_1513),
.Y(n_11958)
);

INVx1_ASAP7_75t_SL g11959 ( 
.A(n_11221),
.Y(n_11959)
);

OAI21x1_ASAP7_75t_SL g11960 ( 
.A1(n_11333),
.A2(n_1513),
.B(n_1514),
.Y(n_11960)
);

NAND2xp5_ASAP7_75t_L g11961 ( 
.A(n_11352),
.B(n_1515),
.Y(n_11961)
);

AOI21xp5_ASAP7_75t_L g11962 ( 
.A1(n_11328),
.A2(n_1515),
.B(n_1516),
.Y(n_11962)
);

OAI21x1_ASAP7_75t_L g11963 ( 
.A1(n_11176),
.A2(n_11187),
.B(n_11180),
.Y(n_11963)
);

OAI21x1_ASAP7_75t_L g11964 ( 
.A1(n_11190),
.A2(n_1516),
.B(n_1517),
.Y(n_11964)
);

AND2x2_ASAP7_75t_L g11965 ( 
.A(n_11372),
.B(n_1517),
.Y(n_11965)
);

AOI21xp5_ASAP7_75t_L g11966 ( 
.A1(n_11467),
.A2(n_1518),
.B(n_1519),
.Y(n_11966)
);

AND2x2_ASAP7_75t_L g11967 ( 
.A(n_11355),
.B(n_1520),
.Y(n_11967)
);

NAND2xp5_ASAP7_75t_L g11968 ( 
.A(n_10989),
.B(n_1520),
.Y(n_11968)
);

OAI21x1_ASAP7_75t_L g11969 ( 
.A1(n_11214),
.A2(n_1521),
.B(n_1522),
.Y(n_11969)
);

OAI21x1_ASAP7_75t_L g11970 ( 
.A1(n_11215),
.A2(n_1521),
.B(n_1522),
.Y(n_11970)
);

OAI21xp5_ASAP7_75t_L g11971 ( 
.A1(n_11216),
.A2(n_1523),
.B(n_1524),
.Y(n_11971)
);

NAND2xp5_ASAP7_75t_L g11972 ( 
.A(n_10835),
.B(n_1523),
.Y(n_11972)
);

AOI22xp5_ASAP7_75t_L g11973 ( 
.A1(n_11460),
.A2(n_1526),
.B1(n_1524),
.B2(n_1525),
.Y(n_11973)
);

AO21x2_ASAP7_75t_L g11974 ( 
.A1(n_11469),
.A2(n_1526),
.B(n_1527),
.Y(n_11974)
);

AOI21xp5_ASAP7_75t_L g11975 ( 
.A1(n_11466),
.A2(n_1527),
.B(n_1528),
.Y(n_11975)
);

INVx3_ASAP7_75t_L g11976 ( 
.A(n_11027),
.Y(n_11976)
);

AOI22xp5_ASAP7_75t_L g11977 ( 
.A1(n_11026),
.A2(n_1530),
.B1(n_1528),
.B2(n_1529),
.Y(n_11977)
);

INVx1_ASAP7_75t_L g11978 ( 
.A(n_10894),
.Y(n_11978)
);

OAI21xp5_ASAP7_75t_L g11979 ( 
.A1(n_11224),
.A2(n_1530),
.B(n_1531),
.Y(n_11979)
);

BUFx3_ASAP7_75t_L g11980 ( 
.A(n_10924),
.Y(n_11980)
);

INVx2_ASAP7_75t_L g11981 ( 
.A(n_10913),
.Y(n_11981)
);

NOR4xp25_ASAP7_75t_L g11982 ( 
.A(n_11356),
.B(n_1534),
.C(n_1532),
.D(n_1533),
.Y(n_11982)
);

BUFx10_ASAP7_75t_L g11983 ( 
.A(n_11182),
.Y(n_11983)
);

INVx1_ASAP7_75t_L g11984 ( 
.A(n_10911),
.Y(n_11984)
);

HB1xp67_ASAP7_75t_L g11985 ( 
.A(n_11405),
.Y(n_11985)
);

AND2x2_ASAP7_75t_L g11986 ( 
.A(n_11050),
.B(n_1532),
.Y(n_11986)
);

AOI21xp5_ASAP7_75t_L g11987 ( 
.A1(n_11198),
.A2(n_1533),
.B(n_1534),
.Y(n_11987)
);

INVx2_ASAP7_75t_SL g11988 ( 
.A(n_11172),
.Y(n_11988)
);

NAND2xp5_ASAP7_75t_L g11989 ( 
.A(n_10821),
.B(n_1535),
.Y(n_11989)
);

NAND2x1p5_ASAP7_75t_L g11990 ( 
.A(n_11237),
.B(n_1537),
.Y(n_11990)
);

AOI22xp33_ASAP7_75t_L g11991 ( 
.A1(n_10878),
.A2(n_1539),
.B1(n_1537),
.B2(n_1538),
.Y(n_11991)
);

NAND2xp5_ASAP7_75t_L g11992 ( 
.A(n_11406),
.B(n_1539),
.Y(n_11992)
);

INVx2_ASAP7_75t_L g11993 ( 
.A(n_11310),
.Y(n_11993)
);

NAND2xp5_ASAP7_75t_L g11994 ( 
.A(n_11137),
.B(n_1540),
.Y(n_11994)
);

OAI21x1_ASAP7_75t_L g11995 ( 
.A1(n_11227),
.A2(n_1540),
.B(n_1541),
.Y(n_11995)
);

INVx1_ASAP7_75t_L g11996 ( 
.A(n_10918),
.Y(n_11996)
);

BUFx6f_ASAP7_75t_L g11997 ( 
.A(n_10937),
.Y(n_11997)
);

NAND2xp5_ASAP7_75t_SL g11998 ( 
.A(n_11408),
.B(n_11400),
.Y(n_11998)
);

OAI21x1_ASAP7_75t_L g11999 ( 
.A1(n_11229),
.A2(n_1541),
.B(n_1542),
.Y(n_11999)
);

INVx1_ASAP7_75t_SL g12000 ( 
.A(n_11244),
.Y(n_12000)
);

OAI21x1_ASAP7_75t_SL g12001 ( 
.A1(n_10948),
.A2(n_1542),
.B(n_1543),
.Y(n_12001)
);

NAND2xp5_ASAP7_75t_L g12002 ( 
.A(n_11150),
.B(n_1544),
.Y(n_12002)
);

AOI22xp5_ASAP7_75t_L g12003 ( 
.A1(n_11144),
.A2(n_1546),
.B1(n_1544),
.B2(n_1545),
.Y(n_12003)
);

AND2x2_ASAP7_75t_L g12004 ( 
.A(n_11290),
.B(n_1545),
.Y(n_12004)
);

NAND2xp5_ASAP7_75t_L g12005 ( 
.A(n_11151),
.B(n_1546),
.Y(n_12005)
);

AOI21xp5_ASAP7_75t_L g12006 ( 
.A1(n_11234),
.A2(n_1547),
.B(n_1548),
.Y(n_12006)
);

OAI21xp33_ASAP7_75t_L g12007 ( 
.A1(n_10994),
.A2(n_1549),
.B(n_1550),
.Y(n_12007)
);

CKINVDCx6p67_ASAP7_75t_R g12008 ( 
.A(n_11192),
.Y(n_12008)
);

OAI21xp5_ASAP7_75t_L g12009 ( 
.A1(n_11268),
.A2(n_1550),
.B(n_1551),
.Y(n_12009)
);

INVx2_ASAP7_75t_L g12010 ( 
.A(n_11310),
.Y(n_12010)
);

OAI21x1_ASAP7_75t_L g12011 ( 
.A1(n_10929),
.A2(n_1551),
.B(n_1552),
.Y(n_12011)
);

NAND2xp5_ASAP7_75t_L g12012 ( 
.A(n_11155),
.B(n_1552),
.Y(n_12012)
);

OAI21x1_ASAP7_75t_L g12013 ( 
.A1(n_10931),
.A2(n_1553),
.B(n_1554),
.Y(n_12013)
);

OAI21x1_ASAP7_75t_L g12014 ( 
.A1(n_10935),
.A2(n_1553),
.B(n_1554),
.Y(n_12014)
);

AOI21xp5_ASAP7_75t_L g12015 ( 
.A1(n_11165),
.A2(n_1555),
.B(n_1556),
.Y(n_12015)
);

CKINVDCx5p33_ASAP7_75t_R g12016 ( 
.A(n_11485),
.Y(n_12016)
);

NAND2xp5_ASAP7_75t_L g12017 ( 
.A(n_11159),
.B(n_1555),
.Y(n_12017)
);

OAI21x1_ASAP7_75t_L g12018 ( 
.A1(n_10957),
.A2(n_1556),
.B(n_1557),
.Y(n_12018)
);

AOI21xp5_ASAP7_75t_L g12019 ( 
.A1(n_11323),
.A2(n_1557),
.B(n_1559),
.Y(n_12019)
);

AO31x2_ASAP7_75t_L g12020 ( 
.A1(n_11423),
.A2(n_1561),
.A3(n_1559),
.B(n_1560),
.Y(n_12020)
);

OAI21x1_ASAP7_75t_L g12021 ( 
.A1(n_10962),
.A2(n_1561),
.B(n_1562),
.Y(n_12021)
);

AO31x2_ASAP7_75t_L g12022 ( 
.A1(n_11453),
.A2(n_1564),
.A3(n_1562),
.B(n_1563),
.Y(n_12022)
);

AND2x2_ASAP7_75t_L g12023 ( 
.A(n_11293),
.B(n_1564),
.Y(n_12023)
);

AND2x4_ASAP7_75t_L g12024 ( 
.A(n_11149),
.B(n_11049),
.Y(n_12024)
);

OAI21xp5_ASAP7_75t_L g12025 ( 
.A1(n_11456),
.A2(n_11156),
.B(n_11154),
.Y(n_12025)
);

NAND2x1_ASAP7_75t_L g12026 ( 
.A(n_11433),
.B(n_11410),
.Y(n_12026)
);

AOI21xp33_ASAP7_75t_L g12027 ( 
.A1(n_11440),
.A2(n_11424),
.B(n_10915),
.Y(n_12027)
);

CKINVDCx5p33_ASAP7_75t_R g12028 ( 
.A(n_10973),
.Y(n_12028)
);

AND2x2_ASAP7_75t_L g12029 ( 
.A(n_11275),
.B(n_1565),
.Y(n_12029)
);

AOI21x1_ASAP7_75t_L g12030 ( 
.A1(n_11034),
.A2(n_1566),
.B(n_1567),
.Y(n_12030)
);

AOI21xp5_ASAP7_75t_L g12031 ( 
.A1(n_11337),
.A2(n_1566),
.B(n_1567),
.Y(n_12031)
);

NAND2xp5_ASAP7_75t_L g12032 ( 
.A(n_11160),
.B(n_1568),
.Y(n_12032)
);

INVx2_ASAP7_75t_L g12033 ( 
.A(n_11310),
.Y(n_12033)
);

NAND2xp5_ASAP7_75t_SL g12034 ( 
.A(n_11400),
.B(n_1568),
.Y(n_12034)
);

OAI21x1_ASAP7_75t_L g12035 ( 
.A1(n_11006),
.A2(n_1569),
.B(n_1570),
.Y(n_12035)
);

NAND2xp5_ASAP7_75t_L g12036 ( 
.A(n_11167),
.B(n_1569),
.Y(n_12036)
);

OA22x2_ASAP7_75t_L g12037 ( 
.A1(n_10960),
.A2(n_1572),
.B1(n_1570),
.B2(n_1571),
.Y(n_12037)
);

AOI211x1_ASAP7_75t_L g12038 ( 
.A1(n_11069),
.A2(n_1573),
.B(n_1571),
.C(n_1572),
.Y(n_12038)
);

OAI21x1_ASAP7_75t_L g12039 ( 
.A1(n_11016),
.A2(n_1573),
.B(n_1574),
.Y(n_12039)
);

AOI21xp5_ASAP7_75t_L g12040 ( 
.A1(n_11329),
.A2(n_1574),
.B(n_1575),
.Y(n_12040)
);

NAND2xp5_ASAP7_75t_SL g12041 ( 
.A(n_11045),
.B(n_1575),
.Y(n_12041)
);

AOI21x1_ASAP7_75t_L g12042 ( 
.A1(n_11086),
.A2(n_1576),
.B(n_1577),
.Y(n_12042)
);

INVx3_ASAP7_75t_L g12043 ( 
.A(n_11027),
.Y(n_12043)
);

INVx1_ASAP7_75t_L g12044 ( 
.A(n_11033),
.Y(n_12044)
);

AND2x2_ASAP7_75t_L g12045 ( 
.A(n_11287),
.B(n_1576),
.Y(n_12045)
);

OAI21x1_ASAP7_75t_L g12046 ( 
.A1(n_11039),
.A2(n_1577),
.B(n_1578),
.Y(n_12046)
);

AOI21xp5_ASAP7_75t_L g12047 ( 
.A1(n_11331),
.A2(n_1578),
.B(n_1579),
.Y(n_12047)
);

OAI21x1_ASAP7_75t_L g12048 ( 
.A1(n_11054),
.A2(n_1579),
.B(n_1580),
.Y(n_12048)
);

NAND2xp5_ASAP7_75t_L g12049 ( 
.A(n_11173),
.B(n_1580),
.Y(n_12049)
);

AOI21xp33_ASAP7_75t_L g12050 ( 
.A1(n_11075),
.A2(n_1581),
.B(n_1582),
.Y(n_12050)
);

OAI21x1_ASAP7_75t_L g12051 ( 
.A1(n_11095),
.A2(n_1581),
.B(n_1582),
.Y(n_12051)
);

OAI21x1_ASAP7_75t_L g12052 ( 
.A1(n_11099),
.A2(n_1583),
.B(n_1584),
.Y(n_12052)
);

AOI21xp5_ASAP7_75t_L g12053 ( 
.A1(n_11002),
.A2(n_1583),
.B(n_1584),
.Y(n_12053)
);

INVx1_ASAP7_75t_L g12054 ( 
.A(n_10963),
.Y(n_12054)
);

OAI21x1_ASAP7_75t_L g12055 ( 
.A1(n_11390),
.A2(n_1585),
.B(n_1586),
.Y(n_12055)
);

OAI21x1_ASAP7_75t_L g12056 ( 
.A1(n_11189),
.A2(n_1585),
.B(n_1586),
.Y(n_12056)
);

AOI21xp5_ASAP7_75t_L g12057 ( 
.A1(n_11394),
.A2(n_1587),
.B(n_1588),
.Y(n_12057)
);

OAI21xp33_ASAP7_75t_L g12058 ( 
.A1(n_11084),
.A2(n_1587),
.B(n_1588),
.Y(n_12058)
);

AND2x4_ASAP7_75t_L g12059 ( 
.A(n_10869),
.B(n_1589),
.Y(n_12059)
);

A2O1A1Ixp33_ASAP7_75t_L g12060 ( 
.A1(n_11157),
.A2(n_1591),
.B(n_1589),
.C(n_1590),
.Y(n_12060)
);

A2O1A1Ixp33_ASAP7_75t_L g12061 ( 
.A1(n_11162),
.A2(n_1592),
.B(n_1590),
.C(n_1591),
.Y(n_12061)
);

NAND2xp5_ASAP7_75t_L g12062 ( 
.A(n_11174),
.B(n_1592),
.Y(n_12062)
);

CKINVDCx16_ASAP7_75t_R g12063 ( 
.A(n_11042),
.Y(n_12063)
);

INVx1_ASAP7_75t_L g12064 ( 
.A(n_10963),
.Y(n_12064)
);

AOI221x1_ASAP7_75t_L g12065 ( 
.A1(n_11239),
.A2(n_1595),
.B1(n_1593),
.B2(n_1594),
.C(n_1596),
.Y(n_12065)
);

OAI21xp5_ASAP7_75t_L g12066 ( 
.A1(n_11170),
.A2(n_1593),
.B(n_1595),
.Y(n_12066)
);

OAI21x1_ASAP7_75t_L g12067 ( 
.A1(n_11432),
.A2(n_1596),
.B(n_1597),
.Y(n_12067)
);

HB1xp67_ASAP7_75t_L g12068 ( 
.A(n_10949),
.Y(n_12068)
);

BUFx2_ASAP7_75t_SL g12069 ( 
.A(n_11158),
.Y(n_12069)
);

OAI21x1_ASAP7_75t_L g12070 ( 
.A1(n_11449),
.A2(n_1597),
.B(n_1598),
.Y(n_12070)
);

AOI31xp67_ASAP7_75t_L g12071 ( 
.A1(n_10861),
.A2(n_11454),
.A3(n_11450),
.B(n_11098),
.Y(n_12071)
);

NAND2xp5_ASAP7_75t_L g12072 ( 
.A(n_11183),
.B(n_1598),
.Y(n_12072)
);

BUFx2_ASAP7_75t_SL g12073 ( 
.A(n_11206),
.Y(n_12073)
);

NAND2xp5_ASAP7_75t_L g12074 ( 
.A(n_10848),
.B(n_1599),
.Y(n_12074)
);

OAI22xp5_ASAP7_75t_L g12075 ( 
.A1(n_11058),
.A2(n_1602),
.B1(n_1600),
.B2(n_1601),
.Y(n_12075)
);

OAI21x1_ASAP7_75t_SL g12076 ( 
.A1(n_10900),
.A2(n_1600),
.B(n_1601),
.Y(n_12076)
);

INVx1_ASAP7_75t_L g12077 ( 
.A(n_11310),
.Y(n_12077)
);

AOI21xp5_ASAP7_75t_L g12078 ( 
.A1(n_11394),
.A2(n_1602),
.B(n_1603),
.Y(n_12078)
);

AO31x2_ASAP7_75t_L g12079 ( 
.A1(n_11233),
.A2(n_1605),
.A3(n_1603),
.B(n_1604),
.Y(n_12079)
);

NAND3xp33_ASAP7_75t_L g12080 ( 
.A(n_11236),
.B(n_1604),
.C(n_1605),
.Y(n_12080)
);

AOI21xp5_ASAP7_75t_L g12081 ( 
.A1(n_11191),
.A2(n_1606),
.B(n_1607),
.Y(n_12081)
);

OAI21x1_ASAP7_75t_L g12082 ( 
.A1(n_11443),
.A2(n_1606),
.B(n_1607),
.Y(n_12082)
);

AOI21xp5_ASAP7_75t_L g12083 ( 
.A1(n_11250),
.A2(n_1608),
.B(n_1609),
.Y(n_12083)
);

INVx3_ASAP7_75t_L g12084 ( 
.A(n_11036),
.Y(n_12084)
);

OAI21x1_ASAP7_75t_L g12085 ( 
.A1(n_11418),
.A2(n_1608),
.B(n_1609),
.Y(n_12085)
);

INVx4_ASAP7_75t_L g12086 ( 
.A(n_11036),
.Y(n_12086)
);

OAI21x1_ASAP7_75t_L g12087 ( 
.A1(n_11199),
.A2(n_1610),
.B(n_1611),
.Y(n_12087)
);

NAND2xp5_ASAP7_75t_L g12088 ( 
.A(n_11113),
.B(n_1610),
.Y(n_12088)
);

AOI21xp5_ASAP7_75t_L g12089 ( 
.A1(n_11263),
.A2(n_1611),
.B(n_1612),
.Y(n_12089)
);

OAI21x1_ASAP7_75t_L g12090 ( 
.A1(n_11461),
.A2(n_1612),
.B(n_1613),
.Y(n_12090)
);

NAND2xp5_ASAP7_75t_L g12091 ( 
.A(n_11092),
.B(n_1613),
.Y(n_12091)
);

INVx1_ASAP7_75t_L g12092 ( 
.A(n_10851),
.Y(n_12092)
);

NAND2xp5_ASAP7_75t_L g12093 ( 
.A(n_11186),
.B(n_11412),
.Y(n_12093)
);

OAI21x1_ASAP7_75t_L g12094 ( 
.A1(n_11261),
.A2(n_1614),
.B(n_1615),
.Y(n_12094)
);

INVx1_ASAP7_75t_L g12095 ( 
.A(n_10854),
.Y(n_12095)
);

AOI21xp5_ASAP7_75t_L g12096 ( 
.A1(n_11276),
.A2(n_1615),
.B(n_1616),
.Y(n_12096)
);

AOI211x1_ASAP7_75t_L g12097 ( 
.A1(n_11090),
.A2(n_1618),
.B(n_1616),
.C(n_1617),
.Y(n_12097)
);

A2O1A1Ixp33_ASAP7_75t_L g12098 ( 
.A1(n_11413),
.A2(n_1619),
.B(n_1617),
.C(n_1618),
.Y(n_12098)
);

NAND2xp5_ASAP7_75t_SL g12099 ( 
.A(n_11317),
.B(n_1619),
.Y(n_12099)
);

NAND2xp5_ASAP7_75t_L g12100 ( 
.A(n_11428),
.B(n_11435),
.Y(n_12100)
);

AOI21xp5_ASAP7_75t_L g12101 ( 
.A1(n_11255),
.A2(n_1620),
.B(n_1621),
.Y(n_12101)
);

OAI21x1_ASAP7_75t_L g12102 ( 
.A1(n_11271),
.A2(n_1620),
.B(n_1621),
.Y(n_12102)
);

AND2x2_ASAP7_75t_L g12103 ( 
.A(n_11244),
.B(n_1622),
.Y(n_12103)
);

AOI21xp5_ASAP7_75t_L g12104 ( 
.A1(n_11366),
.A2(n_1622),
.B(n_1623),
.Y(n_12104)
);

AOI21xp5_ASAP7_75t_L g12105 ( 
.A1(n_11446),
.A2(n_1623),
.B(n_1624),
.Y(n_12105)
);

OAI22xp5_ASAP7_75t_L g12106 ( 
.A1(n_11447),
.A2(n_1626),
.B1(n_1624),
.B2(n_1625),
.Y(n_12106)
);

OAI21x1_ASAP7_75t_L g12107 ( 
.A1(n_10856),
.A2(n_10866),
.B(n_11304),
.Y(n_12107)
);

OAI21x1_ASAP7_75t_L g12108 ( 
.A1(n_11339),
.A2(n_1625),
.B(n_1626),
.Y(n_12108)
);

AO31x2_ASAP7_75t_L g12109 ( 
.A1(n_10802),
.A2(n_1629),
.A3(n_1627),
.B(n_1628),
.Y(n_12109)
);

AO31x2_ASAP7_75t_L g12110 ( 
.A1(n_11483),
.A2(n_1629),
.A3(n_1627),
.B(n_1628),
.Y(n_12110)
);

AND2x4_ASAP7_75t_L g12111 ( 
.A(n_10879),
.B(n_1630),
.Y(n_12111)
);

AND2x4_ASAP7_75t_L g12112 ( 
.A(n_11052),
.B(n_1630),
.Y(n_12112)
);

OAI22xp5_ASAP7_75t_L g12113 ( 
.A1(n_11320),
.A2(n_1633),
.B1(n_1631),
.B2(n_1632),
.Y(n_12113)
);

NAND2xp5_ASAP7_75t_L g12114 ( 
.A(n_11367),
.B(n_1632),
.Y(n_12114)
);

AO31x2_ASAP7_75t_L g12115 ( 
.A1(n_11489),
.A2(n_1635),
.A3(n_1633),
.B(n_1634),
.Y(n_12115)
);

AOI21xp5_ASAP7_75t_L g12116 ( 
.A1(n_11048),
.A2(n_11116),
.B(n_11104),
.Y(n_12116)
);

INVx3_ASAP7_75t_SL g12117 ( 
.A(n_11172),
.Y(n_12117)
);

NAND2x1_ASAP7_75t_L g12118 ( 
.A(n_11433),
.B(n_1636),
.Y(n_12118)
);

AOI21xp5_ASAP7_75t_L g12119 ( 
.A1(n_11121),
.A2(n_11140),
.B(n_11131),
.Y(n_12119)
);

BUFx2_ASAP7_75t_L g12120 ( 
.A(n_11047),
.Y(n_12120)
);

AOI21xp5_ASAP7_75t_L g12121 ( 
.A1(n_11445),
.A2(n_1636),
.B(n_1637),
.Y(n_12121)
);

OAI21x1_ASAP7_75t_L g12122 ( 
.A1(n_11381),
.A2(n_1637),
.B(n_1638),
.Y(n_12122)
);

BUFx12f_ASAP7_75t_L g12123 ( 
.A(n_11524),
.Y(n_12123)
);

OAI21xp5_ASAP7_75t_L g12124 ( 
.A1(n_11490),
.A2(n_1639),
.B(n_1640),
.Y(n_12124)
);

INVx2_ASAP7_75t_L g12125 ( 
.A(n_11047),
.Y(n_12125)
);

AOI21xp5_ASAP7_75t_L g12126 ( 
.A1(n_10855),
.A2(n_1640),
.B(n_1641),
.Y(n_12126)
);

BUFx2_ASAP7_75t_L g12127 ( 
.A(n_11064),
.Y(n_12127)
);

INVxp67_ASAP7_75t_L g12128 ( 
.A(n_11226),
.Y(n_12128)
);

OAI21xp5_ASAP7_75t_L g12129 ( 
.A1(n_11498),
.A2(n_11065),
.B(n_11005),
.Y(n_12129)
);

BUFx2_ASAP7_75t_SL g12130 ( 
.A(n_10967),
.Y(n_12130)
);

AND2x2_ASAP7_75t_L g12131 ( 
.A(n_11073),
.B(n_1641),
.Y(n_12131)
);

HB1xp67_ASAP7_75t_L g12132 ( 
.A(n_11064),
.Y(n_12132)
);

OAI21x1_ASAP7_75t_L g12133 ( 
.A1(n_11204),
.A2(n_1642),
.B(n_1643),
.Y(n_12133)
);

BUFx3_ASAP7_75t_L g12134 ( 
.A(n_10808),
.Y(n_12134)
);

AOI21x1_ASAP7_75t_L g12135 ( 
.A1(n_11278),
.A2(n_1643),
.B(n_1644),
.Y(n_12135)
);

AND2x2_ASAP7_75t_L g12136 ( 
.A(n_10813),
.B(n_1644),
.Y(n_12136)
);

OAI22xp5_ASAP7_75t_L g12137 ( 
.A1(n_11171),
.A2(n_11269),
.B1(n_10980),
.B2(n_11370),
.Y(n_12137)
);

NOR2xp33_ASAP7_75t_L g12138 ( 
.A(n_11389),
.B(n_1645),
.Y(n_12138)
);

NAND2xp5_ASAP7_75t_L g12139 ( 
.A(n_11379),
.B(n_11208),
.Y(n_12139)
);

OAI21x1_ASAP7_75t_L g12140 ( 
.A1(n_11210),
.A2(n_1646),
.B(n_1647),
.Y(n_12140)
);

O2A1O1Ixp33_ASAP7_75t_L g12141 ( 
.A1(n_10982),
.A2(n_1648),
.B(n_1646),
.C(n_1647),
.Y(n_12141)
);

AOI21xp5_ASAP7_75t_L g12142 ( 
.A1(n_10849),
.A2(n_1648),
.B(n_1649),
.Y(n_12142)
);

AO22x2_ASAP7_75t_L g12143 ( 
.A1(n_11283),
.A2(n_1651),
.B1(n_1649),
.B2(n_1650),
.Y(n_12143)
);

NAND2xp5_ASAP7_75t_SL g12144 ( 
.A(n_11127),
.B(n_10881),
.Y(n_12144)
);

AOI211x1_ASAP7_75t_L g12145 ( 
.A1(n_11391),
.A2(n_1652),
.B(n_1650),
.C(n_1651),
.Y(n_12145)
);

AOI21xp33_ASAP7_75t_L g12146 ( 
.A1(n_11105),
.A2(n_11279),
.B(n_11341),
.Y(n_12146)
);

OAI21x1_ASAP7_75t_L g12147 ( 
.A1(n_11225),
.A2(n_1652),
.B(n_1653),
.Y(n_12147)
);

AOI21x1_ASAP7_75t_L g12148 ( 
.A1(n_11350),
.A2(n_1653),
.B(n_1654),
.Y(n_12148)
);

AOI21xp5_ASAP7_75t_L g12149 ( 
.A1(n_10822),
.A2(n_1654),
.B(n_1655),
.Y(n_12149)
);

OAI21xp5_ASAP7_75t_L g12150 ( 
.A1(n_11354),
.A2(n_1655),
.B(n_1656),
.Y(n_12150)
);

NAND2xp5_ASAP7_75t_L g12151 ( 
.A(n_11232),
.B(n_1656),
.Y(n_12151)
);

NAND2xp5_ASAP7_75t_L g12152 ( 
.A(n_11240),
.B(n_11245),
.Y(n_12152)
);

OAI21xp5_ASAP7_75t_L g12153 ( 
.A1(n_11364),
.A2(n_1657),
.B(n_1658),
.Y(n_12153)
);

BUFx6f_ASAP7_75t_L g12154 ( 
.A(n_10940),
.Y(n_12154)
);

INVxp67_ASAP7_75t_SL g12155 ( 
.A(n_11070),
.Y(n_12155)
);

NAND2xp5_ASAP7_75t_L g12156 ( 
.A(n_11256),
.B(n_1657),
.Y(n_12156)
);

NOR2xp67_ASAP7_75t_L g12157 ( 
.A(n_11277),
.B(n_1658),
.Y(n_12157)
);

AOI211x1_ASAP7_75t_L g12158 ( 
.A1(n_11340),
.A2(n_1661),
.B(n_1659),
.C(n_1660),
.Y(n_12158)
);

AO31x2_ASAP7_75t_L g12159 ( 
.A1(n_10917),
.A2(n_1662),
.A3(n_1659),
.B(n_1660),
.Y(n_12159)
);

OAI21x1_ASAP7_75t_L g12160 ( 
.A1(n_11282),
.A2(n_1662),
.B(n_1663),
.Y(n_12160)
);

BUFx2_ASAP7_75t_L g12161 ( 
.A(n_11070),
.Y(n_12161)
);

OAI21x1_ASAP7_75t_L g12162 ( 
.A1(n_11286),
.A2(n_1664),
.B(n_1665),
.Y(n_12162)
);

AO31x2_ASAP7_75t_L g12163 ( 
.A1(n_11164),
.A2(n_1667),
.A3(n_1665),
.B(n_1666),
.Y(n_12163)
);

OAI21x1_ASAP7_75t_SL g12164 ( 
.A1(n_11441),
.A2(n_1666),
.B(n_1667),
.Y(n_12164)
);

AOI211x1_ASAP7_75t_L g12165 ( 
.A1(n_11407),
.A2(n_1670),
.B(n_1668),
.C(n_1669),
.Y(n_12165)
);

OAI21x1_ASAP7_75t_L g12166 ( 
.A1(n_11301),
.A2(n_1668),
.B(n_1669),
.Y(n_12166)
);

INVx1_ASAP7_75t_L g12167 ( 
.A(n_10956),
.Y(n_12167)
);

AOI21xp5_ASAP7_75t_L g12168 ( 
.A1(n_10972),
.A2(n_1670),
.B(n_1672),
.Y(n_12168)
);

INVx4_ASAP7_75t_L g12169 ( 
.A(n_11072),
.Y(n_12169)
);

NAND2xp5_ASAP7_75t_L g12170 ( 
.A(n_11313),
.B(n_1672),
.Y(n_12170)
);

INVxp67_ASAP7_75t_SL g12171 ( 
.A(n_11072),
.Y(n_12171)
);

INVx4_ASAP7_75t_L g12172 ( 
.A(n_11077),
.Y(n_12172)
);

NAND2xp5_ASAP7_75t_L g12173 ( 
.A(n_10793),
.B(n_1673),
.Y(n_12173)
);

OAI21x1_ASAP7_75t_L g12174 ( 
.A1(n_11516),
.A2(n_1673),
.B(n_1674),
.Y(n_12174)
);

NAND2xp5_ASAP7_75t_L g12175 ( 
.A(n_11481),
.B(n_1674),
.Y(n_12175)
);

BUFx6f_ASAP7_75t_L g12176 ( 
.A(n_10940),
.Y(n_12176)
);

INVx5_ASAP7_75t_L g12177 ( 
.A(n_11055),
.Y(n_12177)
);

OAI21x1_ASAP7_75t_L g12178 ( 
.A1(n_11393),
.A2(n_1675),
.B(n_1677),
.Y(n_12178)
);

OAI21x1_ASAP7_75t_L g12179 ( 
.A1(n_11349),
.A2(n_1675),
.B(n_1677),
.Y(n_12179)
);

AND2x2_ASAP7_75t_L g12180 ( 
.A(n_11530),
.B(n_1678),
.Y(n_12180)
);

NAND2xp5_ASAP7_75t_L g12181 ( 
.A(n_11506),
.B(n_1678),
.Y(n_12181)
);

INVx1_ASAP7_75t_L g12182 ( 
.A(n_11001),
.Y(n_12182)
);

NAND2xp5_ASAP7_75t_L g12183 ( 
.A(n_11519),
.B(n_11053),
.Y(n_12183)
);

OAI21x1_ASAP7_75t_L g12184 ( 
.A1(n_11362),
.A2(n_1679),
.B(n_1680),
.Y(n_12184)
);

OAI21x1_ASAP7_75t_L g12185 ( 
.A1(n_11365),
.A2(n_1679),
.B(n_1680),
.Y(n_12185)
);

AND2x2_ASAP7_75t_L g12186 ( 
.A(n_10800),
.B(n_1681),
.Y(n_12186)
);

INVx1_ASAP7_75t_L g12187 ( 
.A(n_10968),
.Y(n_12187)
);

BUFx2_ASAP7_75t_L g12188 ( 
.A(n_11077),
.Y(n_12188)
);

NAND2x1p5_ASAP7_75t_L g12189 ( 
.A(n_11088),
.B(n_1681),
.Y(n_12189)
);

BUFx2_ASAP7_75t_SL g12190 ( 
.A(n_11656),
.Y(n_12190)
);

BUFx3_ASAP7_75t_L g12191 ( 
.A(n_11813),
.Y(n_12191)
);

INVx1_ASAP7_75t_L g12192 ( 
.A(n_11772),
.Y(n_12192)
);

BUFx6f_ASAP7_75t_L g12193 ( 
.A(n_11722),
.Y(n_12193)
);

INVxp67_ASAP7_75t_SL g12194 ( 
.A(n_11832),
.Y(n_12194)
);

INVx2_ASAP7_75t_SL g12195 ( 
.A(n_11737),
.Y(n_12195)
);

OAI21x1_ASAP7_75t_L g12196 ( 
.A1(n_11587),
.A2(n_10997),
.B(n_11196),
.Y(n_12196)
);

BUFx12f_ASAP7_75t_L g12197 ( 
.A(n_12016),
.Y(n_12197)
);

OAI21x1_ASAP7_75t_L g12198 ( 
.A1(n_11647),
.A2(n_11202),
.B(n_11434),
.Y(n_12198)
);

AND2x4_ASAP7_75t_L g12199 ( 
.A(n_11845),
.B(n_11207),
.Y(n_12199)
);

OAI21x1_ASAP7_75t_L g12200 ( 
.A1(n_11590),
.A2(n_11388),
.B(n_11118),
.Y(n_12200)
);

INVx1_ASAP7_75t_L g12201 ( 
.A(n_11667),
.Y(n_12201)
);

INVx1_ASAP7_75t_SL g12202 ( 
.A(n_12117),
.Y(n_12202)
);

CKINVDCx14_ASAP7_75t_R g12203 ( 
.A(n_11601),
.Y(n_12203)
);

BUFx2_ASAP7_75t_SL g12204 ( 
.A(n_11656),
.Y(n_12204)
);

NAND2x1p5_ASAP7_75t_L g12205 ( 
.A(n_12177),
.B(n_11486),
.Y(n_12205)
);

INVx3_ASAP7_75t_L g12206 ( 
.A(n_12026),
.Y(n_12206)
);

BUFx6f_ASAP7_75t_L g12207 ( 
.A(n_11722),
.Y(n_12207)
);

INVx4_ASAP7_75t_L g12208 ( 
.A(n_11868),
.Y(n_12208)
);

INVx2_ASAP7_75t_L g12209 ( 
.A(n_11721),
.Y(n_12209)
);

INVx1_ASAP7_75t_L g12210 ( 
.A(n_11680),
.Y(n_12210)
);

OAI21x1_ASAP7_75t_SL g12211 ( 
.A1(n_11575),
.A2(n_11108),
.B(n_11055),
.Y(n_12211)
);

AO21x2_ASAP7_75t_L g12212 ( 
.A1(n_12077),
.A2(n_12064),
.B(n_12054),
.Y(n_12212)
);

OAI21x1_ASAP7_75t_L g12213 ( 
.A1(n_11724),
.A2(n_11019),
.B(n_10993),
.Y(n_12213)
);

BUFx3_ASAP7_75t_L g12214 ( 
.A(n_11732),
.Y(n_12214)
);

BUFx2_ASAP7_75t_SL g12215 ( 
.A(n_11565),
.Y(n_12215)
);

OAI21xp5_ASAP7_75t_L g12216 ( 
.A1(n_11595),
.A2(n_11291),
.B(n_10978),
.Y(n_12216)
);

INVx1_ASAP7_75t_SL g12217 ( 
.A(n_11912),
.Y(n_12217)
);

BUFx3_ASAP7_75t_L g12218 ( 
.A(n_11688),
.Y(n_12218)
);

INVx1_ASAP7_75t_L g12219 ( 
.A(n_11696),
.Y(n_12219)
);

INVx1_ASAP7_75t_L g12220 ( 
.A(n_11712),
.Y(n_12220)
);

OA21x2_ASAP7_75t_L g12221 ( 
.A1(n_11920),
.A2(n_11436),
.B(n_11325),
.Y(n_12221)
);

BUFx2_ASAP7_75t_L g12222 ( 
.A(n_11646),
.Y(n_12222)
);

INVx1_ASAP7_75t_L g12223 ( 
.A(n_11726),
.Y(n_12223)
);

INVx2_ASAP7_75t_R g12224 ( 
.A(n_12177),
.Y(n_12224)
);

AO21x2_ASAP7_75t_L g12225 ( 
.A1(n_11586),
.A2(n_11438),
.B(n_10923),
.Y(n_12225)
);

INVx1_ASAP7_75t_SL g12226 ( 
.A(n_11959),
.Y(n_12226)
);

INVx1_ASAP7_75t_L g12227 ( 
.A(n_11727),
.Y(n_12227)
);

INVx4_ASAP7_75t_L g12228 ( 
.A(n_11869),
.Y(n_12228)
);

INVx4_ASAP7_75t_L g12229 ( 
.A(n_11694),
.Y(n_12229)
);

NAND2xp5_ASAP7_75t_L g12230 ( 
.A(n_11589),
.B(n_11429),
.Y(n_12230)
);

INVx5_ASAP7_75t_L g12231 ( 
.A(n_11768),
.Y(n_12231)
);

BUFx2_ASAP7_75t_SL g12232 ( 
.A(n_11706),
.Y(n_12232)
);

AND2x4_ASAP7_75t_L g12233 ( 
.A(n_11985),
.B(n_11207),
.Y(n_12233)
);

BUFx6f_ASAP7_75t_L g12234 ( 
.A(n_11735),
.Y(n_12234)
);

INVx1_ASAP7_75t_L g12235 ( 
.A(n_11730),
.Y(n_12235)
);

CKINVDCx8_ASAP7_75t_R g12236 ( 
.A(n_11635),
.Y(n_12236)
);

BUFx3_ASAP7_75t_L g12237 ( 
.A(n_11630),
.Y(n_12237)
);

BUFx3_ASAP7_75t_L g12238 ( 
.A(n_11943),
.Y(n_12238)
);

AOI22x1_ASAP7_75t_L g12239 ( 
.A1(n_11654),
.A2(n_11415),
.B1(n_11344),
.B2(n_10903),
.Y(n_12239)
);

BUFx2_ASAP7_75t_R g12240 ( 
.A(n_11935),
.Y(n_12240)
);

BUFx6f_ASAP7_75t_L g12241 ( 
.A(n_11735),
.Y(n_12241)
);

INVx1_ASAP7_75t_L g12242 ( 
.A(n_11774),
.Y(n_12242)
);

OR2x2_ASAP7_75t_L g12243 ( 
.A(n_11562),
.B(n_11510),
.Y(n_12243)
);

AOI22xp33_ASAP7_75t_L g12244 ( 
.A1(n_11644),
.A2(n_11120),
.B1(n_11168),
.B2(n_11055),
.Y(n_12244)
);

INVx1_ASAP7_75t_L g12245 ( 
.A(n_11778),
.Y(n_12245)
);

AND2x4_ASAP7_75t_L g12246 ( 
.A(n_12155),
.B(n_12171),
.Y(n_12246)
);

INVx1_ASAP7_75t_L g12247 ( 
.A(n_11834),
.Y(n_12247)
);

BUFx12f_ASAP7_75t_L g12248 ( 
.A(n_11837),
.Y(n_12248)
);

BUFx3_ASAP7_75t_L g12249 ( 
.A(n_11983),
.Y(n_12249)
);

AO21x2_ASAP7_75t_L g12250 ( 
.A1(n_11993),
.A2(n_11101),
.B(n_11348),
.Y(n_12250)
);

AO21x2_ASAP7_75t_L g12251 ( 
.A1(n_12010),
.A2(n_11377),
.B(n_11257),
.Y(n_12251)
);

BUFx3_ASAP7_75t_L g12252 ( 
.A(n_11947),
.Y(n_12252)
);

NAND2x1p5_ASAP7_75t_L g12253 ( 
.A(n_11939),
.B(n_11088),
.Y(n_12253)
);

AOI22x1_ASAP7_75t_L g12254 ( 
.A1(n_11599),
.A2(n_11009),
.B1(n_11319),
.B2(n_11031),
.Y(n_12254)
);

NOR2x1_ASAP7_75t_SL g12255 ( 
.A(n_11576),
.B(n_11094),
.Y(n_12255)
);

OAI21x1_ASAP7_75t_L g12256 ( 
.A1(n_11600),
.A2(n_11552),
.B(n_10934),
.Y(n_12256)
);

AOI22x1_ASAP7_75t_L g12257 ( 
.A1(n_11581),
.A2(n_11023),
.B1(n_11035),
.B2(n_11205),
.Y(n_12257)
);

BUFx8_ASAP7_75t_L g12258 ( 
.A(n_11819),
.Y(n_12258)
);

AND2x2_ASAP7_75t_L g12259 ( 
.A(n_11895),
.B(n_11296),
.Y(n_12259)
);

BUFx4f_ASAP7_75t_SL g12260 ( 
.A(n_12123),
.Y(n_12260)
);

INVx1_ASAP7_75t_L g12261 ( 
.A(n_11699),
.Y(n_12261)
);

AND2x4_ASAP7_75t_L g12262 ( 
.A(n_11593),
.B(n_11218),
.Y(n_12262)
);

BUFx12f_ASAP7_75t_L g12263 ( 
.A(n_12028),
.Y(n_12263)
);

BUFx3_ASAP7_75t_L g12264 ( 
.A(n_11826),
.Y(n_12264)
);

INVx2_ASAP7_75t_L g12265 ( 
.A(n_11765),
.Y(n_12265)
);

NAND2xp5_ASAP7_75t_L g12266 ( 
.A(n_11923),
.B(n_11674),
.Y(n_12266)
);

INVx1_ASAP7_75t_L g12267 ( 
.A(n_11785),
.Y(n_12267)
);

INVx4_ASAP7_75t_L g12268 ( 
.A(n_11733),
.Y(n_12268)
);

AOI21x1_ASAP7_75t_L g12269 ( 
.A1(n_11719),
.A2(n_11089),
.B(n_11071),
.Y(n_12269)
);

OR2x6_ASAP7_75t_L g12270 ( 
.A(n_12073),
.B(n_11296),
.Y(n_12270)
);

AND2x2_ASAP7_75t_L g12271 ( 
.A(n_11946),
.B(n_11218),
.Y(n_12271)
);

NAND2x1p5_ASAP7_75t_L g12272 ( 
.A(n_11939),
.B(n_11094),
.Y(n_12272)
);

HB1xp67_ASAP7_75t_L g12273 ( 
.A(n_11607),
.Y(n_12273)
);

OAI21x1_ASAP7_75t_L g12274 ( 
.A1(n_12033),
.A2(n_11838),
.B(n_11846),
.Y(n_12274)
);

AO21x2_ASAP7_75t_L g12275 ( 
.A1(n_11596),
.A2(n_11251),
.B(n_11125),
.Y(n_12275)
);

OR2x6_ASAP7_75t_L g12276 ( 
.A(n_12069),
.B(n_11107),
.Y(n_12276)
);

INVx6_ASAP7_75t_L g12277 ( 
.A(n_11750),
.Y(n_12277)
);

CKINVDCx20_ASAP7_75t_R g12278 ( 
.A(n_12008),
.Y(n_12278)
);

NAND2x1p5_ASAP7_75t_L g12279 ( 
.A(n_11574),
.B(n_11677),
.Y(n_12279)
);

OAI21x1_ASAP7_75t_L g12280 ( 
.A1(n_11866),
.A2(n_11115),
.B(n_11112),
.Y(n_12280)
);

INVx2_ASAP7_75t_L g12281 ( 
.A(n_11810),
.Y(n_12281)
);

OAI21x1_ASAP7_75t_L g12282 ( 
.A1(n_11963),
.A2(n_11181),
.B(n_11128),
.Y(n_12282)
);

NAND2xp5_ASAP7_75t_L g12283 ( 
.A(n_11660),
.B(n_11219),
.Y(n_12283)
);

NAND2xp5_ASAP7_75t_L g12284 ( 
.A(n_11930),
.B(n_11235),
.Y(n_12284)
);

BUFx3_ASAP7_75t_L g12285 ( 
.A(n_11829),
.Y(n_12285)
);

INVx4_ASAP7_75t_L g12286 ( 
.A(n_11815),
.Y(n_12286)
);

BUFx6f_ASAP7_75t_L g12287 ( 
.A(n_11815),
.Y(n_12287)
);

INVx1_ASAP7_75t_L g12288 ( 
.A(n_11828),
.Y(n_12288)
);

BUFx8_ASAP7_75t_L g12289 ( 
.A(n_11905),
.Y(n_12289)
);

INVx1_ASAP7_75t_L g12290 ( 
.A(n_11833),
.Y(n_12290)
);

INVx1_ASAP7_75t_SL g12291 ( 
.A(n_12000),
.Y(n_12291)
);

BUFx3_ASAP7_75t_L g12292 ( 
.A(n_11956),
.Y(n_12292)
);

CKINVDCx5p33_ASAP7_75t_R g12293 ( 
.A(n_12063),
.Y(n_12293)
);

AND2x4_ASAP7_75t_L g12294 ( 
.A(n_11981),
.B(n_11107),
.Y(n_12294)
);

OA21x2_ASAP7_75t_L g12295 ( 
.A1(n_11871),
.A2(n_11270),
.B(n_11265),
.Y(n_12295)
);

INVx5_ASAP7_75t_SL g12296 ( 
.A(n_11904),
.Y(n_12296)
);

BUFx2_ASAP7_75t_L g12297 ( 
.A(n_12132),
.Y(n_12297)
);

AND2x4_ASAP7_75t_L g12298 ( 
.A(n_12120),
.B(n_12127),
.Y(n_12298)
);

INVx1_ASAP7_75t_L g12299 ( 
.A(n_11853),
.Y(n_12299)
);

INVx2_ASAP7_75t_L g12300 ( 
.A(n_11572),
.Y(n_12300)
);

BUFx6f_ASAP7_75t_L g12301 ( 
.A(n_11904),
.Y(n_12301)
);

AO21x2_ASAP7_75t_L g12302 ( 
.A1(n_11605),
.A2(n_10907),
.B(n_11284),
.Y(n_12302)
);

OAI21x1_ASAP7_75t_L g12303 ( 
.A1(n_11578),
.A2(n_11326),
.B(n_11288),
.Y(n_12303)
);

OAI21x1_ASAP7_75t_L g12304 ( 
.A1(n_11734),
.A2(n_11627),
.B(n_11577),
.Y(n_12304)
);

INVx1_ASAP7_75t_L g12305 ( 
.A(n_11640),
.Y(n_12305)
);

NAND2x1p5_ASAP7_75t_L g12306 ( 
.A(n_11998),
.B(n_11147),
.Y(n_12306)
);

CKINVDCx5p33_ASAP7_75t_R g12307 ( 
.A(n_11980),
.Y(n_12307)
);

AO21x2_ASAP7_75t_L g12308 ( 
.A1(n_11857),
.A2(n_11500),
.B(n_11168),
.Y(n_12308)
);

OAI21xp5_ASAP7_75t_L g12309 ( 
.A1(n_11594),
.A2(n_11500),
.B(n_11168),
.Y(n_12309)
);

NAND2xp5_ASAP7_75t_SL g12310 ( 
.A(n_11746),
.B(n_10807),
.Y(n_12310)
);

AO21x2_ASAP7_75t_L g12311 ( 
.A1(n_11858),
.A2(n_11500),
.B(n_11041),
.Y(n_12311)
);

NAND2x1p5_ASAP7_75t_L g12312 ( 
.A(n_11643),
.B(n_11743),
.Y(n_12312)
);

BUFx3_ASAP7_75t_L g12313 ( 
.A(n_12134),
.Y(n_12313)
);

AO21x2_ASAP7_75t_L g12314 ( 
.A1(n_11862),
.A2(n_11046),
.B(n_11252),
.Y(n_12314)
);

OAI21x1_ASAP7_75t_L g12315 ( 
.A1(n_11622),
.A2(n_11079),
.B(n_10857),
.Y(n_12315)
);

AOI22xp33_ASAP7_75t_L g12316 ( 
.A1(n_11657),
.A2(n_11458),
.B1(n_10959),
.B2(n_10803),
.Y(n_12316)
);

AO21x2_ASAP7_75t_L g12317 ( 
.A1(n_11863),
.A2(n_11511),
.B(n_11185),
.Y(n_12317)
);

INVx2_ASAP7_75t_L g12318 ( 
.A(n_11690),
.Y(n_12318)
);

NAND2x1p5_ASAP7_75t_L g12319 ( 
.A(n_12161),
.B(n_11147),
.Y(n_12319)
);

BUFx12f_ASAP7_75t_L g12320 ( 
.A(n_12059),
.Y(n_12320)
);

INVx1_ASAP7_75t_L g12321 ( 
.A(n_11695),
.Y(n_12321)
);

OAI21xp5_ASAP7_75t_L g12322 ( 
.A1(n_11840),
.A2(n_1682),
.B(n_1684),
.Y(n_12322)
);

OR3x4_ASAP7_75t_SL g12323 ( 
.A(n_11608),
.B(n_1684),
.C(n_1685),
.Y(n_12323)
);

AND2x2_ASAP7_75t_L g12324 ( 
.A(n_12068),
.B(n_11185),
.Y(n_12324)
);

INVx2_ASAP7_75t_SL g12325 ( 
.A(n_11783),
.Y(n_12325)
);

INVx1_ASAP7_75t_L g12326 ( 
.A(n_11707),
.Y(n_12326)
);

AND2x4_ASAP7_75t_L g12327 ( 
.A(n_12188),
.B(n_11472),
.Y(n_12327)
);

NOR2xp33_ASAP7_75t_L g12328 ( 
.A(n_12152),
.B(n_11472),
.Y(n_12328)
);

NAND2x1p5_ASAP7_75t_L g12329 ( 
.A(n_12024),
.B(n_11527),
.Y(n_12329)
);

OAI21xp5_ASAP7_75t_L g12330 ( 
.A1(n_11814),
.A2(n_1685),
.B(n_1686),
.Y(n_12330)
);

OAI21xp5_ASAP7_75t_L g12331 ( 
.A1(n_11666),
.A2(n_1686),
.B(n_1687),
.Y(n_12331)
);

OAI21x1_ASAP7_75t_L g12332 ( 
.A1(n_11642),
.A2(n_11531),
.B(n_11527),
.Y(n_12332)
);

AO21x2_ASAP7_75t_L g12333 ( 
.A1(n_11865),
.A2(n_11555),
.B(n_11531),
.Y(n_12333)
);

INVx1_ASAP7_75t_L g12334 ( 
.A(n_11709),
.Y(n_12334)
);

BUFx12f_ASAP7_75t_L g12335 ( 
.A(n_12111),
.Y(n_12335)
);

AND2x2_ASAP7_75t_SL g12336 ( 
.A(n_11982),
.B(n_11555),
.Y(n_12336)
);

AO21x2_ASAP7_75t_L g12337 ( 
.A1(n_11875),
.A2(n_1687),
.B(n_1688),
.Y(n_12337)
);

OAI21x1_ASAP7_75t_L g12338 ( 
.A1(n_11839),
.A2(n_1689),
.B(n_1690),
.Y(n_12338)
);

INVx2_ASAP7_75t_L g12339 ( 
.A(n_11741),
.Y(n_12339)
);

OAI21xp5_ASAP7_75t_L g12340 ( 
.A1(n_11728),
.A2(n_1689),
.B(n_1691),
.Y(n_12340)
);

INVx1_ASAP7_75t_L g12341 ( 
.A(n_11754),
.Y(n_12341)
);

HB1xp67_ASAP7_75t_L g12342 ( 
.A(n_11881),
.Y(n_12342)
);

BUFx2_ASAP7_75t_L g12343 ( 
.A(n_11901),
.Y(n_12343)
);

OAI21x1_ASAP7_75t_L g12344 ( 
.A1(n_11591),
.A2(n_1691),
.B(n_1692),
.Y(n_12344)
);

BUFx12f_ASAP7_75t_L g12345 ( 
.A(n_12112),
.Y(n_12345)
);

OAI21x1_ASAP7_75t_L g12346 ( 
.A1(n_11606),
.A2(n_1692),
.B(n_1693),
.Y(n_12346)
);

INVx1_ASAP7_75t_SL g12347 ( 
.A(n_11798),
.Y(n_12347)
);

INVx2_ASAP7_75t_SL g12348 ( 
.A(n_11988),
.Y(n_12348)
);

INVxp67_ASAP7_75t_SL g12349 ( 
.A(n_11880),
.Y(n_12349)
);

NAND2x1p5_ASAP7_75t_L g12350 ( 
.A(n_11776),
.B(n_1693),
.Y(n_12350)
);

AO21x2_ASAP7_75t_L g12351 ( 
.A1(n_11876),
.A2(n_1694),
.B(n_1695),
.Y(n_12351)
);

AND2x2_ASAP7_75t_L g12352 ( 
.A(n_11918),
.B(n_1694),
.Y(n_12352)
);

BUFx6f_ASAP7_75t_L g12353 ( 
.A(n_11914),
.Y(n_12353)
);

OAI21x1_ASAP7_75t_L g12354 ( 
.A1(n_11718),
.A2(n_1696),
.B(n_1697),
.Y(n_12354)
);

INVx1_ASAP7_75t_SL g12355 ( 
.A(n_11955),
.Y(n_12355)
);

OR2x6_ASAP7_75t_L g12356 ( 
.A(n_12130),
.B(n_1696),
.Y(n_12356)
);

AO21x2_ASAP7_75t_L g12357 ( 
.A1(n_11878),
.A2(n_11563),
.B(n_11592),
.Y(n_12357)
);

INVx1_ASAP7_75t_L g12358 ( 
.A(n_11882),
.Y(n_12358)
);

OAI21x1_ASAP7_75t_L g12359 ( 
.A1(n_11729),
.A2(n_1697),
.B(n_1698),
.Y(n_12359)
);

NAND2xp5_ASAP7_75t_L g12360 ( 
.A(n_11996),
.B(n_12044),
.Y(n_12360)
);

AO21x2_ASAP7_75t_L g12361 ( 
.A1(n_11720),
.A2(n_1698),
.B(n_1699),
.Y(n_12361)
);

INVx2_ASAP7_75t_L g12362 ( 
.A(n_11887),
.Y(n_12362)
);

INVx2_ASAP7_75t_L g12363 ( 
.A(n_11893),
.Y(n_12363)
);

OA21x2_ASAP7_75t_L g12364 ( 
.A1(n_12107),
.A2(n_1699),
.B(n_1700),
.Y(n_12364)
);

BUFx3_ASAP7_75t_L g12365 ( 
.A(n_11860),
.Y(n_12365)
);

BUFx2_ASAP7_75t_SL g12366 ( 
.A(n_11659),
.Y(n_12366)
);

OAI21x1_ASAP7_75t_L g12367 ( 
.A1(n_11610),
.A2(n_1700),
.B(n_1701),
.Y(n_12367)
);

CKINVDCx5p33_ASAP7_75t_R g12368 ( 
.A(n_11914),
.Y(n_12368)
);

OAI21xp5_ASAP7_75t_L g12369 ( 
.A1(n_11736),
.A2(n_1701),
.B(n_1702),
.Y(n_12369)
);

INVx1_ASAP7_75t_SL g12370 ( 
.A(n_11997),
.Y(n_12370)
);

OAI21xp5_ASAP7_75t_L g12371 ( 
.A1(n_11744),
.A2(n_1703),
.B(n_1704),
.Y(n_12371)
);

AO21x2_ASAP7_75t_L g12372 ( 
.A1(n_11731),
.A2(n_1703),
.B(n_1705),
.Y(n_12372)
);

INVx1_ASAP7_75t_SL g12373 ( 
.A(n_11997),
.Y(n_12373)
);

AND2x2_ASAP7_75t_L g12374 ( 
.A(n_12167),
.B(n_1705),
.Y(n_12374)
);

AO21x2_ASAP7_75t_L g12375 ( 
.A1(n_11745),
.A2(n_1706),
.B(n_1707),
.Y(n_12375)
);

OR2x6_ASAP7_75t_L g12376 ( 
.A(n_11682),
.B(n_1706),
.Y(n_12376)
);

BUFx3_ASAP7_75t_L g12377 ( 
.A(n_12154),
.Y(n_12377)
);

AOI22xp33_ASAP7_75t_SL g12378 ( 
.A1(n_12137),
.A2(n_1709),
.B1(n_1707),
.B2(n_1708),
.Y(n_12378)
);

INVx1_ASAP7_75t_L g12379 ( 
.A(n_11978),
.Y(n_12379)
);

NAND2x1p5_ASAP7_75t_L g12380 ( 
.A(n_12086),
.B(n_1708),
.Y(n_12380)
);

AND2x4_ASAP7_75t_L g12381 ( 
.A(n_12125),
.B(n_1709),
.Y(n_12381)
);

INVx2_ASAP7_75t_SL g12382 ( 
.A(n_12154),
.Y(n_12382)
);

NAND2xp5_ASAP7_75t_L g12383 ( 
.A(n_11984),
.B(n_1710),
.Y(n_12383)
);

BUFx3_ASAP7_75t_L g12384 ( 
.A(n_12176),
.Y(n_12384)
);

CKINVDCx11_ASAP7_75t_R g12385 ( 
.A(n_12176),
.Y(n_12385)
);

BUFx4f_ASAP7_75t_SL g12386 ( 
.A(n_12169),
.Y(n_12386)
);

CKINVDCx20_ASAP7_75t_R g12387 ( 
.A(n_12139),
.Y(n_12387)
);

BUFx2_ASAP7_75t_L g12388 ( 
.A(n_12128),
.Y(n_12388)
);

OAI21xp5_ASAP7_75t_L g12389 ( 
.A1(n_11748),
.A2(n_11758),
.B(n_11755),
.Y(n_12389)
);

HB1xp67_ASAP7_75t_L g12390 ( 
.A(n_11582),
.Y(n_12390)
);

BUFx3_ASAP7_75t_L g12391 ( 
.A(n_11925),
.Y(n_12391)
);

OAI21x1_ASAP7_75t_L g12392 ( 
.A1(n_11739),
.A2(n_1710),
.B(n_1711),
.Y(n_12392)
);

CKINVDCx8_ASAP7_75t_R g12393 ( 
.A(n_11768),
.Y(n_12393)
);

OAI21x1_ASAP7_75t_L g12394 ( 
.A1(n_11747),
.A2(n_1711),
.B(n_1712),
.Y(n_12394)
);

AO21x2_ASAP7_75t_L g12395 ( 
.A1(n_11751),
.A2(n_1712),
.B(n_1713),
.Y(n_12395)
);

OR2x6_ASAP7_75t_L g12396 ( 
.A(n_11682),
.B(n_1713),
.Y(n_12396)
);

AND2x2_ASAP7_75t_L g12397 ( 
.A(n_12092),
.B(n_1714),
.Y(n_12397)
);

INVx3_ASAP7_75t_L g12398 ( 
.A(n_12172),
.Y(n_12398)
);

INVx1_ASAP7_75t_L g12399 ( 
.A(n_12095),
.Y(n_12399)
);

BUFx3_ASAP7_75t_L g12400 ( 
.A(n_11976),
.Y(n_12400)
);

OAI21xp5_ASAP7_75t_L g12401 ( 
.A1(n_11780),
.A2(n_1715),
.B(n_1716),
.Y(n_12401)
);

INVx1_ASAP7_75t_L g12402 ( 
.A(n_11812),
.Y(n_12402)
);

INVx1_ASAP7_75t_L g12403 ( 
.A(n_11821),
.Y(n_12403)
);

BUFx6f_ASAP7_75t_L g12404 ( 
.A(n_12043),
.Y(n_12404)
);

OAI21x1_ASAP7_75t_L g12405 ( 
.A1(n_11793),
.A2(n_1715),
.B(n_1716),
.Y(n_12405)
);

INVx1_ASAP7_75t_L g12406 ( 
.A(n_11822),
.Y(n_12406)
);

BUFx2_ASAP7_75t_L g12407 ( 
.A(n_12084),
.Y(n_12407)
);

OA21x2_ASAP7_75t_L g12408 ( 
.A1(n_11573),
.A2(n_1717),
.B(n_1718),
.Y(n_12408)
);

INVx8_ASAP7_75t_L g12409 ( 
.A(n_11571),
.Y(n_12409)
);

OAI21x1_ASAP7_75t_L g12410 ( 
.A1(n_11665),
.A2(n_1717),
.B(n_1718),
.Y(n_12410)
);

INVx1_ASAP7_75t_L g12411 ( 
.A(n_11825),
.Y(n_12411)
);

AOI22x1_ASAP7_75t_L g12412 ( 
.A1(n_12015),
.A2(n_1721),
.B1(n_1719),
.B2(n_1720),
.Y(n_12412)
);

INVx2_ASAP7_75t_L g12413 ( 
.A(n_12182),
.Y(n_12413)
);

NAND2xp5_ASAP7_75t_L g12414 ( 
.A(n_12187),
.B(n_1719),
.Y(n_12414)
);

BUFx2_ASAP7_75t_L g12415 ( 
.A(n_11716),
.Y(n_12415)
);

OA21x2_ASAP7_75t_L g12416 ( 
.A1(n_11649),
.A2(n_1721),
.B(n_1722),
.Y(n_12416)
);

INVx2_ASAP7_75t_SL g12417 ( 
.A(n_11952),
.Y(n_12417)
);

OAI21x1_ASAP7_75t_L g12418 ( 
.A1(n_11669),
.A2(n_1722),
.B(n_1723),
.Y(n_12418)
);

INVx1_ASAP7_75t_L g12419 ( 
.A(n_11827),
.Y(n_12419)
);

AO21x2_ASAP7_75t_L g12420 ( 
.A1(n_11628),
.A2(n_1724),
.B(n_1725),
.Y(n_12420)
);

INVx2_ASAP7_75t_L g12421 ( 
.A(n_11850),
.Y(n_12421)
);

INVx2_ASAP7_75t_L g12422 ( 
.A(n_11585),
.Y(n_12422)
);

OR2x2_ASAP7_75t_L g12423 ( 
.A(n_11673),
.B(n_1724),
.Y(n_12423)
);

INVx2_ASAP7_75t_L g12424 ( 
.A(n_11681),
.Y(n_12424)
);

INVx1_ASAP7_75t_L g12425 ( 
.A(n_11672),
.Y(n_12425)
);

BUFx3_ASAP7_75t_L g12426 ( 
.A(n_11965),
.Y(n_12426)
);

OAI21x1_ASAP7_75t_L g12427 ( 
.A1(n_11676),
.A2(n_1726),
.B(n_1727),
.Y(n_12427)
);

INVx2_ASAP7_75t_SL g12428 ( 
.A(n_11566),
.Y(n_12428)
);

OAI21x1_ASAP7_75t_L g12429 ( 
.A1(n_11678),
.A2(n_1726),
.B(n_1727),
.Y(n_12429)
);

BUFx2_ASAP7_75t_R g12430 ( 
.A(n_12144),
.Y(n_12430)
);

INVx1_ASAP7_75t_L g12431 ( 
.A(n_11672),
.Y(n_12431)
);

INVx2_ASAP7_75t_L g12432 ( 
.A(n_11888),
.Y(n_12432)
);

INVx2_ASAP7_75t_L g12433 ( 
.A(n_11629),
.Y(n_12433)
);

INVx1_ASAP7_75t_L g12434 ( 
.A(n_11692),
.Y(n_12434)
);

AO21x2_ASAP7_75t_L g12435 ( 
.A1(n_11664),
.A2(n_1728),
.B(n_1730),
.Y(n_12435)
);

BUFx4_ASAP7_75t_SL g12436 ( 
.A(n_11796),
.Y(n_12436)
);

BUFx5_ASAP7_75t_L g12437 ( 
.A(n_11768),
.Y(n_12437)
);

OR2x6_ASAP7_75t_L g12438 ( 
.A(n_12116),
.B(n_1728),
.Y(n_12438)
);

NAND2x1p5_ASAP7_75t_L g12439 ( 
.A(n_11771),
.B(n_1731),
.Y(n_12439)
);

INVx1_ASAP7_75t_L g12440 ( 
.A(n_11692),
.Y(n_12440)
);

INVx4_ASAP7_75t_L g12441 ( 
.A(n_12103),
.Y(n_12441)
);

AND2x2_ASAP7_75t_L g12442 ( 
.A(n_11597),
.B(n_1732),
.Y(n_12442)
);

AOI22xp33_ASAP7_75t_L g12443 ( 
.A1(n_12027),
.A2(n_1734),
.B1(n_1732),
.B2(n_1733),
.Y(n_12443)
);

INVx2_ASAP7_75t_L g12444 ( 
.A(n_11759),
.Y(n_12444)
);

OAI21xp5_ASAP7_75t_L g12445 ( 
.A1(n_11653),
.A2(n_1735),
.B(n_1736),
.Y(n_12445)
);

INVx1_ASAP7_75t_L g12446 ( 
.A(n_11723),
.Y(n_12446)
);

BUFx6f_ASAP7_75t_L g12447 ( 
.A(n_12131),
.Y(n_12447)
);

BUFx3_ASAP7_75t_L g12448 ( 
.A(n_11907),
.Y(n_12448)
);

AOI21x1_ASAP7_75t_L g12449 ( 
.A1(n_11697),
.A2(n_1735),
.B(n_1736),
.Y(n_12449)
);

BUFx2_ASAP7_75t_L g12450 ( 
.A(n_11645),
.Y(n_12450)
);

NAND2x1p5_ASAP7_75t_L g12451 ( 
.A(n_11658),
.B(n_1737),
.Y(n_12451)
);

NOR2xp33_ASAP7_75t_L g12452 ( 
.A(n_12114),
.B(n_12183),
.Y(n_12452)
);

INVx1_ASAP7_75t_L g12453 ( 
.A(n_11723),
.Y(n_12453)
);

OAI21xp5_ASAP7_75t_L g12454 ( 
.A1(n_11820),
.A2(n_1737),
.B(n_1738),
.Y(n_12454)
);

INVx3_ASAP7_75t_SL g12455 ( 
.A(n_11986),
.Y(n_12455)
);

INVx2_ASAP7_75t_L g12456 ( 
.A(n_11611),
.Y(n_12456)
);

OAI21x1_ASAP7_75t_L g12457 ( 
.A1(n_11686),
.A2(n_1739),
.B(n_1740),
.Y(n_12457)
);

INVx1_ASAP7_75t_L g12458 ( 
.A(n_11633),
.Y(n_12458)
);

BUFx3_ASAP7_75t_L g12459 ( 
.A(n_12029),
.Y(n_12459)
);

NOR2xp33_ASAP7_75t_L g12460 ( 
.A(n_12093),
.B(n_1741),
.Y(n_12460)
);

AOI22x1_ASAP7_75t_L g12461 ( 
.A1(n_12019),
.A2(n_1743),
.B1(n_1741),
.B2(n_1742),
.Y(n_12461)
);

OAI21x1_ASAP7_75t_L g12462 ( 
.A1(n_11614),
.A2(n_1742),
.B(n_1743),
.Y(n_12462)
);

INVx3_ASAP7_75t_L g12463 ( 
.A(n_12023),
.Y(n_12463)
);

INVx1_ASAP7_75t_SL g12464 ( 
.A(n_11738),
.Y(n_12464)
);

OAI21x1_ASAP7_75t_L g12465 ( 
.A1(n_11583),
.A2(n_1744),
.B(n_1746),
.Y(n_12465)
);

INVx1_ASAP7_75t_L g12466 ( 
.A(n_11683),
.Y(n_12466)
);

BUFx2_ASAP7_75t_L g12467 ( 
.A(n_11631),
.Y(n_12467)
);

NAND2xp5_ASAP7_75t_L g12468 ( 
.A(n_11613),
.B(n_1744),
.Y(n_12468)
);

AO21x2_ASAP7_75t_L g12469 ( 
.A1(n_11698),
.A2(n_1746),
.B(n_1747),
.Y(n_12469)
);

INVx1_ASAP7_75t_L g12470 ( 
.A(n_11687),
.Y(n_12470)
);

INVx2_ASAP7_75t_L g12471 ( 
.A(n_11762),
.Y(n_12471)
);

INVx2_ASAP7_75t_SL g12472 ( 
.A(n_11773),
.Y(n_12472)
);

AO21x2_ASAP7_75t_L g12473 ( 
.A1(n_11883),
.A2(n_1747),
.B(n_1749),
.Y(n_12473)
);

INVx1_ASAP7_75t_L g12474 ( 
.A(n_11689),
.Y(n_12474)
);

AO21x2_ASAP7_75t_L g12475 ( 
.A1(n_11568),
.A2(n_1749),
.B(n_1750),
.Y(n_12475)
);

NAND2x1p5_ASAP7_75t_L g12476 ( 
.A(n_11584),
.B(n_1750),
.Y(n_12476)
);

BUFx3_ASAP7_75t_L g12477 ( 
.A(n_12045),
.Y(n_12477)
);

NOR2x1_ASAP7_75t_R g12478 ( 
.A(n_11766),
.B(n_1751),
.Y(n_12478)
);

BUFx6f_ASAP7_75t_L g12479 ( 
.A(n_12118),
.Y(n_12479)
);

INVx3_ASAP7_75t_L g12480 ( 
.A(n_11775),
.Y(n_12480)
);

INVx1_ASAP7_75t_SL g12481 ( 
.A(n_11967),
.Y(n_12481)
);

INVx1_ASAP7_75t_L g12482 ( 
.A(n_11693),
.Y(n_12482)
);

AO21x1_ASAP7_75t_L g12483 ( 
.A1(n_12121),
.A2(n_1751),
.B(n_1752),
.Y(n_12483)
);

OR2x2_ASAP7_75t_L g12484 ( 
.A(n_11906),
.B(n_11961),
.Y(n_12484)
);

INVx1_ASAP7_75t_L g12485 ( 
.A(n_11705),
.Y(n_12485)
);

OAI21x1_ASAP7_75t_L g12486 ( 
.A1(n_11789),
.A2(n_1752),
.B(n_1753),
.Y(n_12486)
);

INVx1_ASAP7_75t_SL g12487 ( 
.A(n_11921),
.Y(n_12487)
);

AO21x2_ASAP7_75t_L g12488 ( 
.A1(n_11787),
.A2(n_1754),
.B(n_1755),
.Y(n_12488)
);

INVx1_ASAP7_75t_L g12489 ( 
.A(n_11708),
.Y(n_12489)
);

AO21x2_ASAP7_75t_L g12490 ( 
.A1(n_11992),
.A2(n_1754),
.B(n_1755),
.Y(n_12490)
);

BUFx10_ASAP7_75t_L g12491 ( 
.A(n_11903),
.Y(n_12491)
);

OAI21x1_ASAP7_75t_L g12492 ( 
.A1(n_11802),
.A2(n_1756),
.B(n_1757),
.Y(n_12492)
);

OA21x2_ASAP7_75t_L g12493 ( 
.A1(n_11655),
.A2(n_1758),
.B(n_1759),
.Y(n_12493)
);

INVx1_ASAP7_75t_SL g12494 ( 
.A(n_11808),
.Y(n_12494)
);

AND2x4_ASAP7_75t_L g12495 ( 
.A(n_12090),
.B(n_11579),
.Y(n_12495)
);

BUFx3_ASAP7_75t_L g12496 ( 
.A(n_12186),
.Y(n_12496)
);

BUFx12f_ASAP7_75t_L g12497 ( 
.A(n_12189),
.Y(n_12497)
);

AO21x2_ASAP7_75t_L g12498 ( 
.A1(n_11756),
.A2(n_1758),
.B(n_1760),
.Y(n_12498)
);

OAI21xp33_ASAP7_75t_SL g12499 ( 
.A1(n_11763),
.A2(n_1761),
.B(n_1762),
.Y(n_12499)
);

OAI21x1_ASAP7_75t_L g12500 ( 
.A1(n_11623),
.A2(n_1762),
.B(n_1763),
.Y(n_12500)
);

OA21x2_ASAP7_75t_L g12501 ( 
.A1(n_11620),
.A2(n_1763),
.B(n_1764),
.Y(n_12501)
);

CKINVDCx11_ASAP7_75t_R g12502 ( 
.A(n_12106),
.Y(n_12502)
);

HB1xp67_ASAP7_75t_L g12503 ( 
.A(n_11974),
.Y(n_12503)
);

OR2x2_ASAP7_75t_L g12504 ( 
.A(n_11941),
.B(n_1764),
.Y(n_12504)
);

INVxp67_ASAP7_75t_SL g12505 ( 
.A(n_11710),
.Y(n_12505)
);

INVx6_ASAP7_75t_L g12506 ( 
.A(n_12004),
.Y(n_12506)
);

INVx1_ASAP7_75t_SL g12507 ( 
.A(n_11951),
.Y(n_12507)
);

OAI21xp5_ASAP7_75t_L g12508 ( 
.A1(n_11609),
.A2(n_1765),
.B(n_1766),
.Y(n_12508)
);

INVx3_ASAP7_75t_L g12509 ( 
.A(n_11886),
.Y(n_12509)
);

BUFx2_ASAP7_75t_L g12510 ( 
.A(n_11990),
.Y(n_12510)
);

AND2x4_ASAP7_75t_L g12511 ( 
.A(n_11652),
.B(n_1766),
.Y(n_12511)
);

INVx1_ASAP7_75t_L g12512 ( 
.A(n_11711),
.Y(n_12512)
);

AND2x2_ASAP7_75t_L g12513 ( 
.A(n_11626),
.B(n_1767),
.Y(n_12513)
);

BUFx3_ASAP7_75t_L g12514 ( 
.A(n_11663),
.Y(n_12514)
);

AO21x2_ASAP7_75t_L g12515 ( 
.A1(n_11761),
.A2(n_1767),
.B(n_1768),
.Y(n_12515)
);

INVx1_ASAP7_75t_L g12516 ( 
.A(n_11717),
.Y(n_12516)
);

OAI21xp5_ASAP7_75t_L g12517 ( 
.A1(n_11801),
.A2(n_1769),
.B(n_1770),
.Y(n_12517)
);

BUFx6f_ASAP7_75t_L g12518 ( 
.A(n_11770),
.Y(n_12518)
);

INVx2_ASAP7_75t_L g12519 ( 
.A(n_12071),
.Y(n_12519)
);

OA21x2_ASAP7_75t_L g12520 ( 
.A1(n_11767),
.A2(n_1769),
.B(n_1770),
.Y(n_12520)
);

INVx2_ASAP7_75t_L g12521 ( 
.A(n_11781),
.Y(n_12521)
);

BUFx5_ASAP7_75t_L g12522 ( 
.A(n_12136),
.Y(n_12522)
);

OAI21x1_ASAP7_75t_L g12523 ( 
.A1(n_11902),
.A2(n_1771),
.B(n_1773),
.Y(n_12523)
);

INVx8_ASAP7_75t_L g12524 ( 
.A(n_12180),
.Y(n_12524)
);

INVx2_ASAP7_75t_L g12525 ( 
.A(n_11764),
.Y(n_12525)
);

HB1xp67_ASAP7_75t_L g12526 ( 
.A(n_11777),
.Y(n_12526)
);

BUFx4f_ASAP7_75t_SL g12527 ( 
.A(n_11844),
.Y(n_12527)
);

OAI21x1_ASAP7_75t_L g12528 ( 
.A1(n_11910),
.A2(n_1771),
.B(n_1773),
.Y(n_12528)
);

OAI21x1_ASAP7_75t_L g12529 ( 
.A1(n_11791),
.A2(n_1774),
.B(n_1775),
.Y(n_12529)
);

INVx5_ASAP7_75t_SL g12530 ( 
.A(n_11804),
.Y(n_12530)
);

BUFx6f_ASAP7_75t_L g12531 ( 
.A(n_11786),
.Y(n_12531)
);

OAI21x1_ASAP7_75t_L g12532 ( 
.A1(n_11588),
.A2(n_1774),
.B(n_1775),
.Y(n_12532)
);

INVx1_ASAP7_75t_L g12533 ( 
.A(n_11621),
.Y(n_12533)
);

CKINVDCx16_ASAP7_75t_R g12534 ( 
.A(n_11618),
.Y(n_12534)
);

BUFx2_ASAP7_75t_L g12535 ( 
.A(n_11779),
.Y(n_12535)
);

AND2x2_ASAP7_75t_L g12536 ( 
.A(n_11703),
.B(n_1776),
.Y(n_12536)
);

INVx2_ASAP7_75t_L g12537 ( 
.A(n_11909),
.Y(n_12537)
);

INVx1_ASAP7_75t_L g12538 ( 
.A(n_11621),
.Y(n_12538)
);

BUFx3_ASAP7_75t_L g12539 ( 
.A(n_11788),
.Y(n_12539)
);

OR2x2_ASAP7_75t_L g12540 ( 
.A(n_12091),
.B(n_1777),
.Y(n_12540)
);

AO21x2_ASAP7_75t_L g12541 ( 
.A1(n_11859),
.A2(n_1778),
.B(n_1779),
.Y(n_12541)
);

INVx3_ASAP7_75t_L g12542 ( 
.A(n_12011),
.Y(n_12542)
);

AO21x2_ASAP7_75t_L g12543 ( 
.A1(n_11864),
.A2(n_1778),
.B(n_1780),
.Y(n_12543)
);

BUFx6f_ASAP7_75t_L g12544 ( 
.A(n_11899),
.Y(n_12544)
);

OAI21x1_ASAP7_75t_L g12545 ( 
.A1(n_11797),
.A2(n_1780),
.B(n_1781),
.Y(n_12545)
);

AND2x4_ASAP7_75t_L g12546 ( 
.A(n_12013),
.B(n_1781),
.Y(n_12546)
);

INVx2_ASAP7_75t_SL g12547 ( 
.A(n_11989),
.Y(n_12547)
);

INVx3_ASAP7_75t_L g12548 ( 
.A(n_12014),
.Y(n_12548)
);

INVx2_ASAP7_75t_L g12549 ( 
.A(n_12018),
.Y(n_12549)
);

NAND2xp5_ASAP7_75t_SL g12550 ( 
.A(n_12119),
.B(n_1782),
.Y(n_12550)
);

AOI21x1_ASAP7_75t_L g12551 ( 
.A1(n_11753),
.A2(n_1782),
.B(n_1783),
.Y(n_12551)
);

BUFx3_ASAP7_75t_L g12552 ( 
.A(n_11924),
.Y(n_12552)
);

NOR2xp33_ASAP7_75t_L g12553 ( 
.A(n_11932),
.B(n_1783),
.Y(n_12553)
);

AO21x2_ASAP7_75t_L g12554 ( 
.A1(n_11987),
.A2(n_1784),
.B(n_1786),
.Y(n_12554)
);

BUFx4f_ASAP7_75t_L g12555 ( 
.A(n_11854),
.Y(n_12555)
);

INVx2_ASAP7_75t_SL g12556 ( 
.A(n_12074),
.Y(n_12556)
);

INVx1_ASAP7_75t_L g12557 ( 
.A(n_11760),
.Y(n_12557)
);

AND2x4_ASAP7_75t_L g12558 ( 
.A(n_12021),
.B(n_12035),
.Y(n_12558)
);

NAND2xp5_ASAP7_75t_L g12559 ( 
.A(n_11879),
.B(n_1784),
.Y(n_12559)
);

NAND2xp5_ASAP7_75t_L g12560 ( 
.A(n_11894),
.B(n_1786),
.Y(n_12560)
);

NAND2xp5_ASAP7_75t_L g12561 ( 
.A(n_11897),
.B(n_1787),
.Y(n_12561)
);

INVx2_ASAP7_75t_SL g12562 ( 
.A(n_11972),
.Y(n_12562)
);

HB1xp67_ASAP7_75t_L g12563 ( 
.A(n_11650),
.Y(n_12563)
);

INVx1_ASAP7_75t_L g12564 ( 
.A(n_11760),
.Y(n_12564)
);

BUFx4f_ASAP7_75t_L g12565 ( 
.A(n_11782),
.Y(n_12565)
);

BUFx6f_ASAP7_75t_L g12566 ( 
.A(n_12174),
.Y(n_12566)
);

INVx1_ASAP7_75t_L g12567 ( 
.A(n_11650),
.Y(n_12567)
);

AO21x2_ASAP7_75t_L g12568 ( 
.A1(n_11740),
.A2(n_1787),
.B(n_1788),
.Y(n_12568)
);

AOI22x1_ASAP7_75t_L g12569 ( 
.A1(n_12143),
.A2(n_1790),
.B1(n_1788),
.B2(n_1789),
.Y(n_12569)
);

AND2x4_ASAP7_75t_L g12570 ( 
.A(n_12039),
.B(n_1789),
.Y(n_12570)
);

INVx2_ASAP7_75t_L g12571 ( 
.A(n_12046),
.Y(n_12571)
);

AOI22xp33_ASAP7_75t_SL g12572 ( 
.A1(n_12025),
.A2(n_1792),
.B1(n_1790),
.B2(n_1791),
.Y(n_12572)
);

INVx2_ASAP7_75t_SL g12573 ( 
.A(n_11994),
.Y(n_12573)
);

BUFx3_ASAP7_75t_L g12574 ( 
.A(n_12173),
.Y(n_12574)
);

NOR2xp33_ASAP7_75t_L g12575 ( 
.A(n_12100),
.B(n_1791),
.Y(n_12575)
);

INVx2_ASAP7_75t_L g12576 ( 
.A(n_12048),
.Y(n_12576)
);

INVx2_ASAP7_75t_SL g12577 ( 
.A(n_12002),
.Y(n_12577)
);

INVx3_ASAP7_75t_L g12578 ( 
.A(n_12051),
.Y(n_12578)
);

INVx1_ASAP7_75t_L g12579 ( 
.A(n_12179),
.Y(n_12579)
);

AOI22xp33_ASAP7_75t_L g12580 ( 
.A1(n_12129),
.A2(n_1794),
.B1(n_1792),
.B2(n_1793),
.Y(n_12580)
);

INVx8_ASAP7_75t_L g12581 ( 
.A(n_11691),
.Y(n_12581)
);

INVx2_ASAP7_75t_SL g12582 ( 
.A(n_12005),
.Y(n_12582)
);

OAI21x1_ASAP7_75t_L g12583 ( 
.A1(n_11816),
.A2(n_1793),
.B(n_1794),
.Y(n_12583)
);

BUFx2_ASAP7_75t_L g12584 ( 
.A(n_12052),
.Y(n_12584)
);

INVx2_ASAP7_75t_L g12585 ( 
.A(n_11725),
.Y(n_12585)
);

BUFx6f_ASAP7_75t_L g12586 ( 
.A(n_12087),
.Y(n_12586)
);

AOI22x1_ASAP7_75t_L g12587 ( 
.A1(n_12143),
.A2(n_1797),
.B1(n_1795),
.B2(n_1796),
.Y(n_12587)
);

AO21x2_ASAP7_75t_L g12588 ( 
.A1(n_12053),
.A2(n_1795),
.B(n_1797),
.Y(n_12588)
);

AND2x4_ASAP7_75t_L g12589 ( 
.A(n_12102),
.B(n_1798),
.Y(n_12589)
);

NAND2x1p5_ASAP7_75t_L g12590 ( 
.A(n_11632),
.B(n_1798),
.Y(n_12590)
);

AOI22x1_ASAP7_75t_L g12591 ( 
.A1(n_11685),
.A2(n_1801),
.B1(n_1799),
.B2(n_1800),
.Y(n_12591)
);

BUFx6f_ASAP7_75t_L g12592 ( 
.A(n_12012),
.Y(n_12592)
);

AND2x2_ASAP7_75t_L g12593 ( 
.A(n_12138),
.B(n_1799),
.Y(n_12593)
);

AND2x4_ASAP7_75t_L g12594 ( 
.A(n_12140),
.B(n_1800),
.Y(n_12594)
);

AOI22x1_ASAP7_75t_L g12595 ( 
.A1(n_11598),
.A2(n_1804),
.B1(n_1802),
.B2(n_1803),
.Y(n_12595)
);

BUFx3_ASAP7_75t_L g12596 ( 
.A(n_12175),
.Y(n_12596)
);

AO21x1_ASAP7_75t_L g12597 ( 
.A1(n_11700),
.A2(n_1802),
.B(n_1803),
.Y(n_12597)
);

AO21x2_ASAP7_75t_L g12598 ( 
.A1(n_11580),
.A2(n_11661),
.B(n_11604),
.Y(n_12598)
);

INVx1_ASAP7_75t_L g12599 ( 
.A(n_12184),
.Y(n_12599)
);

BUFx3_ASAP7_75t_L g12600 ( 
.A(n_12181),
.Y(n_12600)
);

OAI21x1_ASAP7_75t_L g12601 ( 
.A1(n_11648),
.A2(n_1804),
.B(n_1805),
.Y(n_12601)
);

BUFx2_ASAP7_75t_SL g12602 ( 
.A(n_12157),
.Y(n_12602)
);

INVx2_ASAP7_75t_L g12603 ( 
.A(n_12147),
.Y(n_12603)
);

INVx3_ASAP7_75t_L g12604 ( 
.A(n_12185),
.Y(n_12604)
);

INVx2_ASAP7_75t_L g12605 ( 
.A(n_12160),
.Y(n_12605)
);

AO21x2_ASAP7_75t_L g12606 ( 
.A1(n_11670),
.A2(n_1805),
.B(n_1806),
.Y(n_12606)
);

AND2x4_ASAP7_75t_L g12607 ( 
.A(n_12162),
.B(n_1807),
.Y(n_12607)
);

NAND2x1p5_ASAP7_75t_L g12608 ( 
.A(n_11885),
.B(n_1807),
.Y(n_12608)
);

BUFx3_ASAP7_75t_L g12609 ( 
.A(n_12017),
.Y(n_12609)
);

INVx1_ASAP7_75t_SL g12610 ( 
.A(n_12032),
.Y(n_12610)
);

CKINVDCx16_ASAP7_75t_R g12611 ( 
.A(n_11651),
.Y(n_12611)
);

AND2x2_ASAP7_75t_L g12612 ( 
.A(n_12166),
.B(n_1808),
.Y(n_12612)
);

INVx3_ASAP7_75t_L g12613 ( 
.A(n_12133),
.Y(n_12613)
);

INVx2_ASAP7_75t_L g12614 ( 
.A(n_12067),
.Y(n_12614)
);

AOI22x1_ASAP7_75t_L g12615 ( 
.A1(n_11784),
.A2(n_1810),
.B1(n_1808),
.B2(n_1809),
.Y(n_12615)
);

INVx1_ASAP7_75t_L g12616 ( 
.A(n_11634),
.Y(n_12616)
);

OAI21x1_ASAP7_75t_L g12617 ( 
.A1(n_11938),
.A2(n_1809),
.B(n_1811),
.Y(n_12617)
);

INVx2_ASAP7_75t_L g12618 ( 
.A(n_12056),
.Y(n_12618)
);

BUFx2_ASAP7_75t_L g12619 ( 
.A(n_11634),
.Y(n_12619)
);

INVx1_ASAP7_75t_L g12620 ( 
.A(n_11913),
.Y(n_12620)
);

NAND2xp5_ASAP7_75t_L g12621 ( 
.A(n_11944),
.B(n_1811),
.Y(n_12621)
);

INVx2_ASAP7_75t_SL g12622 ( 
.A(n_12036),
.Y(n_12622)
);

CKINVDCx20_ASAP7_75t_R g12623 ( 
.A(n_11968),
.Y(n_12623)
);

BUFx3_ASAP7_75t_L g12624 ( 
.A(n_12049),
.Y(n_12624)
);

OAI21x1_ASAP7_75t_L g12625 ( 
.A1(n_11940),
.A2(n_1812),
.B(n_1813),
.Y(n_12625)
);

OAI21x1_ASAP7_75t_L g12626 ( 
.A1(n_11950),
.A2(n_11957),
.B(n_11953),
.Y(n_12626)
);

OAI21xp5_ASAP7_75t_L g12627 ( 
.A1(n_11892),
.A2(n_1812),
.B(n_1814),
.Y(n_12627)
);

INVxp67_ASAP7_75t_SL g12628 ( 
.A(n_12034),
.Y(n_12628)
);

NOR2xp33_ASAP7_75t_L g12629 ( 
.A(n_11927),
.B(n_1815),
.Y(n_12629)
);

BUFx3_ASAP7_75t_L g12630 ( 
.A(n_12062),
.Y(n_12630)
);

AND2x4_ASAP7_75t_L g12631 ( 
.A(n_11874),
.B(n_1815),
.Y(n_12631)
);

INVx4_ASAP7_75t_L g12632 ( 
.A(n_12037),
.Y(n_12632)
);

OAI21x1_ASAP7_75t_L g12633 ( 
.A1(n_11958),
.A2(n_1816),
.B(n_1817),
.Y(n_12633)
);

AOI21xp33_ASAP7_75t_L g12634 ( 
.A1(n_11794),
.A2(n_1816),
.B(n_1818),
.Y(n_12634)
);

NAND3xp33_ASAP7_75t_SL g12635 ( 
.A(n_11679),
.B(n_1818),
.C(n_1819),
.Y(n_12635)
);

INVx3_ASAP7_75t_L g12636 ( 
.A(n_11713),
.Y(n_12636)
);

INVx1_ASAP7_75t_SL g12637 ( 
.A(n_12072),
.Y(n_12637)
);

OAI21x1_ASAP7_75t_SL g12638 ( 
.A1(n_12135),
.A2(n_1819),
.B(n_1821),
.Y(n_12638)
);

BUFx2_ASAP7_75t_SL g12639 ( 
.A(n_12099),
.Y(n_12639)
);

INVx3_ASAP7_75t_SL g12640 ( 
.A(n_12041),
.Y(n_12640)
);

OAI21x1_ASAP7_75t_L g12641 ( 
.A1(n_11964),
.A2(n_1821),
.B(n_1822),
.Y(n_12641)
);

AO21x2_ASAP7_75t_L g12642 ( 
.A1(n_11702),
.A2(n_11615),
.B(n_11817),
.Y(n_12642)
);

INVx5_ASAP7_75t_L g12643 ( 
.A(n_11790),
.Y(n_12643)
);

OAI21x1_ASAP7_75t_SL g12644 ( 
.A1(n_12066),
.A2(n_12164),
.B(n_11849),
.Y(n_12644)
);

INVx2_ASAP7_75t_L g12645 ( 
.A(n_12333),
.Y(n_12645)
);

OAI21x1_ASAP7_75t_L g12646 ( 
.A1(n_12274),
.A2(n_11931),
.B(n_11836),
.Y(n_12646)
);

OAI21x1_ASAP7_75t_L g12647 ( 
.A1(n_12304),
.A2(n_12213),
.B(n_12567),
.Y(n_12647)
);

INVx1_ASAP7_75t_L g12648 ( 
.A(n_12349),
.Y(n_12648)
);

CKINVDCx16_ASAP7_75t_R g12649 ( 
.A(n_12323),
.Y(n_12649)
);

BUFx2_ASAP7_75t_L g12650 ( 
.A(n_12253),
.Y(n_12650)
);

NAND2xp5_ASAP7_75t_L g12651 ( 
.A(n_12505),
.B(n_11928),
.Y(n_12651)
);

AND2x4_ASAP7_75t_L g12652 ( 
.A(n_12206),
.B(n_11841),
.Y(n_12652)
);

INVx1_ASAP7_75t_L g12653 ( 
.A(n_12201),
.Y(n_12653)
);

OA21x2_ASAP7_75t_L g12654 ( 
.A1(n_12519),
.A2(n_11624),
.B(n_11641),
.Y(n_12654)
);

OAI21x1_ASAP7_75t_L g12655 ( 
.A1(n_12256),
.A2(n_11617),
.B(n_11969),
.Y(n_12655)
);

INVx2_ASAP7_75t_L g12656 ( 
.A(n_12280),
.Y(n_12656)
);

INVx1_ASAP7_75t_L g12657 ( 
.A(n_12210),
.Y(n_12657)
);

INVx2_ASAP7_75t_L g12658 ( 
.A(n_12282),
.Y(n_12658)
);

INVx1_ASAP7_75t_L g12659 ( 
.A(n_12219),
.Y(n_12659)
);

OAI21x1_ASAP7_75t_L g12660 ( 
.A1(n_12433),
.A2(n_11995),
.B(n_11970),
.Y(n_12660)
);

NOR3xp33_ASAP7_75t_L g12661 ( 
.A(n_12322),
.B(n_11619),
.C(n_12146),
.Y(n_12661)
);

OAI22xp5_ASAP7_75t_L g12662 ( 
.A1(n_12430),
.A2(n_11891),
.B1(n_12003),
.B2(n_11824),
.Y(n_12662)
);

OAI21x1_ASAP7_75t_L g12663 ( 
.A1(n_12444),
.A2(n_11999),
.B(n_11847),
.Y(n_12663)
);

INVx1_ASAP7_75t_L g12664 ( 
.A(n_12220),
.Y(n_12664)
);

AO21x2_ASAP7_75t_L g12665 ( 
.A1(n_12563),
.A2(n_11945),
.B(n_11757),
.Y(n_12665)
);

INVx3_ASAP7_75t_L g12666 ( 
.A(n_12246),
.Y(n_12666)
);

OAI21x1_ASAP7_75t_L g12667 ( 
.A1(n_12542),
.A2(n_11851),
.B(n_11842),
.Y(n_12667)
);

OAI21x1_ASAP7_75t_L g12668 ( 
.A1(n_12548),
.A2(n_11861),
.B(n_11855),
.Y(n_12668)
);

O2A1O1Ixp33_ASAP7_75t_L g12669 ( 
.A1(n_12454),
.A2(n_11639),
.B(n_11636),
.C(n_11684),
.Y(n_12669)
);

O2A1O1Ixp33_ASAP7_75t_L g12670 ( 
.A1(n_12331),
.A2(n_12309),
.B(n_12550),
.C(n_12636),
.Y(n_12670)
);

BUFx2_ASAP7_75t_L g12671 ( 
.A(n_12272),
.Y(n_12671)
);

INVx1_ASAP7_75t_L g12672 ( 
.A(n_12223),
.Y(n_12672)
);

INVx3_ASAP7_75t_L g12673 ( 
.A(n_12298),
.Y(n_12673)
);

AND4x1_ASAP7_75t_L g12674 ( 
.A(n_12244),
.B(n_11926),
.C(n_12065),
.D(n_11742),
.Y(n_12674)
);

OAI21x1_ASAP7_75t_L g12675 ( 
.A1(n_12578),
.A2(n_11889),
.B(n_11884),
.Y(n_12675)
);

OAI21x1_ASAP7_75t_L g12676 ( 
.A1(n_12604),
.A2(n_11896),
.B(n_11818),
.Y(n_12676)
);

OAI22xp5_ASAP7_75t_L g12677 ( 
.A1(n_12632),
.A2(n_11807),
.B1(n_11662),
.B2(n_11973),
.Y(n_12677)
);

INVx1_ASAP7_75t_L g12678 ( 
.A(n_12227),
.Y(n_12678)
);

INVx3_ASAP7_75t_L g12679 ( 
.A(n_12365),
.Y(n_12679)
);

AOI21xp5_ASAP7_75t_L g12680 ( 
.A1(n_12389),
.A2(n_11852),
.B(n_11843),
.Y(n_12680)
);

CKINVDCx5p33_ASAP7_75t_R g12681 ( 
.A(n_12203),
.Y(n_12681)
);

NAND3xp33_ASAP7_75t_L g12682 ( 
.A(n_12216),
.B(n_11638),
.C(n_11637),
.Y(n_12682)
);

OAI21x1_ASAP7_75t_L g12683 ( 
.A1(n_12471),
.A2(n_11975),
.B(n_12030),
.Y(n_12683)
);

A2O1A1Ixp33_ASAP7_75t_L g12684 ( 
.A1(n_12508),
.A2(n_12330),
.B(n_12565),
.C(n_12517),
.Y(n_12684)
);

BUFx8_ASAP7_75t_L g12685 ( 
.A(n_12197),
.Y(n_12685)
);

OAI221xp5_ASAP7_75t_L g12686 ( 
.A1(n_12378),
.A2(n_12153),
.B1(n_12150),
.B2(n_11919),
.C(n_11867),
.Y(n_12686)
);

INVx2_ASAP7_75t_L g12687 ( 
.A(n_12363),
.Y(n_12687)
);

AOI21xp5_ASAP7_75t_L g12688 ( 
.A1(n_12642),
.A2(n_12598),
.B(n_12555),
.Y(n_12688)
);

AND2x4_ASAP7_75t_L g12689 ( 
.A(n_12233),
.B(n_12022),
.Y(n_12689)
);

OAI21x1_ASAP7_75t_L g12690 ( 
.A1(n_12613),
.A2(n_12042),
.B(n_11835),
.Y(n_12690)
);

INVx3_ASAP7_75t_L g12691 ( 
.A(n_12264),
.Y(n_12691)
);

INVx1_ASAP7_75t_L g12692 ( 
.A(n_12235),
.Y(n_12692)
);

OAI21x1_ASAP7_75t_L g12693 ( 
.A1(n_12425),
.A2(n_12122),
.B(n_12108),
.Y(n_12693)
);

INVx1_ASAP7_75t_L g12694 ( 
.A(n_12242),
.Y(n_12694)
);

INVx2_ASAP7_75t_L g12695 ( 
.A(n_12297),
.Y(n_12695)
);

INVx1_ASAP7_75t_L g12696 ( 
.A(n_12245),
.Y(n_12696)
);

BUFx2_ASAP7_75t_L g12697 ( 
.A(n_12222),
.Y(n_12697)
);

HB1xp67_ASAP7_75t_L g12698 ( 
.A(n_12603),
.Y(n_12698)
);

NOR2xp33_ASAP7_75t_L g12699 ( 
.A(n_12236),
.B(n_12088),
.Y(n_12699)
);

INVx2_ASAP7_75t_L g12700 ( 
.A(n_12192),
.Y(n_12700)
);

AOI22xp33_ASAP7_75t_SL g12701 ( 
.A1(n_12530),
.A2(n_12619),
.B1(n_12611),
.B2(n_12527),
.Y(n_12701)
);

BUFx6f_ASAP7_75t_L g12702 ( 
.A(n_12191),
.Y(n_12702)
);

INVx1_ASAP7_75t_L g12703 ( 
.A(n_12247),
.Y(n_12703)
);

NAND2xp5_ASAP7_75t_L g12704 ( 
.A(n_12458),
.B(n_12151),
.Y(n_12704)
);

INVx2_ASAP7_75t_SL g12705 ( 
.A(n_12277),
.Y(n_12705)
);

INVx2_ASAP7_75t_L g12706 ( 
.A(n_12265),
.Y(n_12706)
);

AO31x2_ASAP7_75t_L g12707 ( 
.A1(n_12255),
.A2(n_12434),
.A3(n_12440),
.B(n_12431),
.Y(n_12707)
);

A2O1A1Ixp33_ASAP7_75t_L g12708 ( 
.A1(n_12499),
.A2(n_11856),
.B(n_11567),
.C(n_11799),
.Y(n_12708)
);

OAI21xp5_ASAP7_75t_L g12709 ( 
.A1(n_12627),
.A2(n_11900),
.B(n_11715),
.Y(n_12709)
);

AO31x2_ASAP7_75t_L g12710 ( 
.A1(n_12446),
.A2(n_11848),
.A3(n_11917),
.B(n_11873),
.Y(n_12710)
);

INVx6_ASAP7_75t_L g12711 ( 
.A(n_12248),
.Y(n_12711)
);

OAI22xp5_ASAP7_75t_L g12712 ( 
.A1(n_12640),
.A2(n_12080),
.B1(n_11612),
.B2(n_11877),
.Y(n_12712)
);

BUFx8_ASAP7_75t_L g12713 ( 
.A(n_12263),
.Y(n_12713)
);

OAI21x1_ASAP7_75t_L g12714 ( 
.A1(n_12453),
.A2(n_12078),
.B(n_12057),
.Y(n_12714)
);

INVx1_ASAP7_75t_L g12715 ( 
.A(n_12273),
.Y(n_12715)
);

OAI21x1_ASAP7_75t_L g12716 ( 
.A1(n_12585),
.A2(n_11704),
.B(n_12178),
.Y(n_12716)
);

NOR2x1_ASAP7_75t_SL g12717 ( 
.A(n_12275),
.B(n_11714),
.Y(n_12717)
);

INVx1_ASAP7_75t_L g12718 ( 
.A(n_12358),
.Y(n_12718)
);

INVx1_ASAP7_75t_L g12719 ( 
.A(n_12267),
.Y(n_12719)
);

BUFx2_ASAP7_75t_L g12720 ( 
.A(n_12495),
.Y(n_12720)
);

NAND2xp5_ASAP7_75t_L g12721 ( 
.A(n_12466),
.B(n_12156),
.Y(n_12721)
);

INVx2_ASAP7_75t_L g12722 ( 
.A(n_12281),
.Y(n_12722)
);

INVx1_ASAP7_75t_L g12723 ( 
.A(n_12288),
.Y(n_12723)
);

INVx2_ASAP7_75t_L g12724 ( 
.A(n_12261),
.Y(n_12724)
);

OAI21x1_ASAP7_75t_L g12725 ( 
.A1(n_12557),
.A2(n_12148),
.B(n_12006),
.Y(n_12725)
);

OAI21x1_ASAP7_75t_SL g12726 ( 
.A1(n_12269),
.A2(n_11752),
.B(n_11806),
.Y(n_12726)
);

OAI21x1_ASAP7_75t_L g12727 ( 
.A1(n_12564),
.A2(n_12082),
.B(n_12070),
.Y(n_12727)
);

BUFx6f_ASAP7_75t_L g12728 ( 
.A(n_12385),
.Y(n_12728)
);

HB1xp67_ASAP7_75t_L g12729 ( 
.A(n_12605),
.Y(n_12729)
);

NOR2xp33_ASAP7_75t_SL g12730 ( 
.A(n_12240),
.B(n_12058),
.Y(n_12730)
);

OAI22xp5_ASAP7_75t_L g12731 ( 
.A1(n_12231),
.A2(n_12061),
.B1(n_12060),
.B2(n_12098),
.Y(n_12731)
);

OAI21x1_ASAP7_75t_L g12732 ( 
.A1(n_12618),
.A2(n_12085),
.B(n_12094),
.Y(n_12732)
);

CKINVDCx8_ASAP7_75t_R g12733 ( 
.A(n_12232),
.Y(n_12733)
);

OAI21xp5_ASAP7_75t_L g12734 ( 
.A1(n_12200),
.A2(n_11625),
.B(n_11937),
.Y(n_12734)
);

INVx1_ASAP7_75t_L g12735 ( 
.A(n_12290),
.Y(n_12735)
);

INVx1_ASAP7_75t_L g12736 ( 
.A(n_12299),
.Y(n_12736)
);

OAI21x1_ASAP7_75t_L g12737 ( 
.A1(n_12537),
.A2(n_11962),
.B(n_11949),
.Y(n_12737)
);

OA21x2_ASAP7_75t_L g12738 ( 
.A1(n_12194),
.A2(n_12170),
.B(n_12055),
.Y(n_12738)
);

OAI21xp5_ASAP7_75t_L g12739 ( 
.A1(n_12340),
.A2(n_11979),
.B(n_11971),
.Y(n_12739)
);

OAI21x1_ASAP7_75t_L g12740 ( 
.A1(n_12614),
.A2(n_12571),
.B(n_12549),
.Y(n_12740)
);

INVx1_ASAP7_75t_L g12741 ( 
.A(n_12379),
.Y(n_12741)
);

NAND2x1p5_ASAP7_75t_L g12742 ( 
.A(n_12217),
.B(n_12226),
.Y(n_12742)
);

NAND2xp5_ASAP7_75t_L g12743 ( 
.A(n_12470),
.B(n_12145),
.Y(n_12743)
);

INVx1_ASAP7_75t_L g12744 ( 
.A(n_12399),
.Y(n_12744)
);

OAI21xp33_ASAP7_75t_SL g12745 ( 
.A1(n_12616),
.A2(n_11977),
.B(n_12050),
.Y(n_12745)
);

OAI21x1_ASAP7_75t_L g12746 ( 
.A1(n_12576),
.A2(n_12538),
.B(n_12533),
.Y(n_12746)
);

INVx1_ASAP7_75t_L g12747 ( 
.A(n_12343),
.Y(n_12747)
);

CKINVDCx5p33_ASAP7_75t_R g12748 ( 
.A(n_12278),
.Y(n_12748)
);

A2O1A1Ixp33_ASAP7_75t_L g12749 ( 
.A1(n_12369),
.A2(n_12401),
.B(n_12371),
.C(n_12553),
.Y(n_12749)
);

NOR2xp33_ASAP7_75t_L g12750 ( 
.A(n_12208),
.B(n_12007),
.Y(n_12750)
);

OAI21x1_ASAP7_75t_L g12751 ( 
.A1(n_12525),
.A2(n_11916),
.B(n_11616),
.Y(n_12751)
);

OAI21x1_ASAP7_75t_L g12752 ( 
.A1(n_12198),
.A2(n_11830),
.B(n_11823),
.Y(n_12752)
);

AOI22x1_ASAP7_75t_L g12753 ( 
.A1(n_12503),
.A2(n_11675),
.B1(n_12047),
.B2(n_12040),
.Y(n_12753)
);

HB1xp67_ASAP7_75t_L g12754 ( 
.A(n_12579),
.Y(n_12754)
);

AOI21x1_ASAP7_75t_L g12755 ( 
.A1(n_12620),
.A2(n_11966),
.B(n_12105),
.Y(n_12755)
);

OAI21xp5_ASAP7_75t_L g12756 ( 
.A1(n_12196),
.A2(n_12009),
.B(n_12101),
.Y(n_12756)
);

O2A1O1Ixp33_ASAP7_75t_SL g12757 ( 
.A1(n_12310),
.A2(n_11870),
.B(n_12124),
.C(n_11569),
.Y(n_12757)
);

OAI21x1_ASAP7_75t_L g12758 ( 
.A1(n_12626),
.A2(n_12332),
.B(n_12599),
.Y(n_12758)
);

INVx2_ASAP7_75t_L g12759 ( 
.A(n_12212),
.Y(n_12759)
);

INVx1_ASAP7_75t_L g12760 ( 
.A(n_12305),
.Y(n_12760)
);

INVx1_ASAP7_75t_L g12761 ( 
.A(n_12321),
.Y(n_12761)
);

AOI221xp5_ASAP7_75t_L g12762 ( 
.A1(n_12635),
.A2(n_11564),
.B1(n_11936),
.B2(n_11954),
.C(n_11749),
.Y(n_12762)
);

AOI22xp33_ASAP7_75t_L g12763 ( 
.A1(n_12502),
.A2(n_11922),
.B1(n_11805),
.B2(n_11811),
.Y(n_12763)
);

OAI21xp5_ASAP7_75t_L g12764 ( 
.A1(n_12445),
.A2(n_11603),
.B(n_11602),
.Y(n_12764)
);

NAND2xp5_ASAP7_75t_L g12765 ( 
.A(n_12474),
.B(n_12158),
.Y(n_12765)
);

AOI22xp33_ASAP7_75t_SL g12766 ( 
.A1(n_12211),
.A2(n_11795),
.B1(n_12075),
.B2(n_11934),
.Y(n_12766)
);

NAND2xp5_ASAP7_75t_SL g12767 ( 
.A(n_12231),
.B(n_12165),
.Y(n_12767)
);

NAND2xp33_ASAP7_75t_L g12768 ( 
.A(n_12437),
.B(n_11991),
.Y(n_12768)
);

CKINVDCx20_ASAP7_75t_R g12769 ( 
.A(n_12260),
.Y(n_12769)
);

AND2x2_ASAP7_75t_L g12770 ( 
.A(n_12209),
.B(n_12020),
.Y(n_12770)
);

NOR2xp33_ASAP7_75t_L g12771 ( 
.A(n_12190),
.B(n_12031),
.Y(n_12771)
);

INVx1_ASAP7_75t_L g12772 ( 
.A(n_12326),
.Y(n_12772)
);

NOR2xp67_ASAP7_75t_L g12773 ( 
.A(n_12228),
.B(n_12268),
.Y(n_12773)
);

BUFx2_ASAP7_75t_L g12774 ( 
.A(n_12279),
.Y(n_12774)
);

CKINVDCx5p33_ASAP7_75t_R g12775 ( 
.A(n_12293),
.Y(n_12775)
);

OAI21x1_ASAP7_75t_SL g12776 ( 
.A1(n_12597),
.A2(n_11960),
.B(n_11898),
.Y(n_12776)
);

AOI22x1_ASAP7_75t_L g12777 ( 
.A1(n_12204),
.A2(n_12083),
.B1(n_12089),
.B2(n_12081),
.Y(n_12777)
);

AO21x2_ASAP7_75t_L g12778 ( 
.A1(n_12526),
.A2(n_12360),
.B(n_12402),
.Y(n_12778)
);

INVx1_ASAP7_75t_L g12779 ( 
.A(n_12334),
.Y(n_12779)
);

INVx1_ASAP7_75t_L g12780 ( 
.A(n_12341),
.Y(n_12780)
);

AOI21xp5_ASAP7_75t_L g12781 ( 
.A1(n_12634),
.A2(n_12096),
.B(n_12141),
.Y(n_12781)
);

OAI21xp5_ASAP7_75t_L g12782 ( 
.A1(n_12221),
.A2(n_11570),
.B(n_11671),
.Y(n_12782)
);

INVx1_ASAP7_75t_L g12783 ( 
.A(n_12342),
.Y(n_12783)
);

NAND3xp33_ASAP7_75t_L g12784 ( 
.A(n_12591),
.B(n_12142),
.C(n_11942),
.Y(n_12784)
);

AOI22xp33_ASAP7_75t_L g12785 ( 
.A1(n_12225),
.A2(n_11769),
.B1(n_12113),
.B2(n_12126),
.Y(n_12785)
);

INVx1_ASAP7_75t_L g12786 ( 
.A(n_12413),
.Y(n_12786)
);

AOI21xp5_ASAP7_75t_L g12787 ( 
.A1(n_12483),
.A2(n_11911),
.B(n_12168),
.Y(n_12787)
);

AOI22xp5_ASAP7_75t_L g12788 ( 
.A1(n_12311),
.A2(n_11701),
.B1(n_11872),
.B2(n_12149),
.Y(n_12788)
);

NOR2xp33_ASAP7_75t_L g12789 ( 
.A(n_12229),
.B(n_12104),
.Y(n_12789)
);

NAND2xp5_ASAP7_75t_L g12790 ( 
.A(n_12482),
.B(n_11668),
.Y(n_12790)
);

NAND3xp33_ASAP7_75t_L g12791 ( 
.A(n_12412),
.B(n_11929),
.C(n_12038),
.Y(n_12791)
);

NOR2xp33_ASAP7_75t_L g12792 ( 
.A(n_12202),
.B(n_1822),
.Y(n_12792)
);

OAI21xp5_ASAP7_75t_L g12793 ( 
.A1(n_12460),
.A2(n_11948),
.B(n_11933),
.Y(n_12793)
);

OAI21x1_ASAP7_75t_L g12794 ( 
.A1(n_12303),
.A2(n_12076),
.B(n_12001),
.Y(n_12794)
);

AOI21x1_ASAP7_75t_L g12795 ( 
.A1(n_12584),
.A2(n_12097),
.B(n_11668),
.Y(n_12795)
);

INVx1_ASAP7_75t_L g12796 ( 
.A(n_12300),
.Y(n_12796)
);

OAI21x1_ASAP7_75t_L g12797 ( 
.A1(n_12306),
.A2(n_12022),
.B(n_12020),
.Y(n_12797)
);

INVx1_ASAP7_75t_L g12798 ( 
.A(n_12318),
.Y(n_12798)
);

OAI21x1_ASAP7_75t_L g12799 ( 
.A1(n_12338),
.A2(n_12319),
.B(n_12315),
.Y(n_12799)
);

OAI21x1_ASAP7_75t_L g12800 ( 
.A1(n_12329),
.A2(n_12079),
.B(n_11800),
.Y(n_12800)
);

OAI21x1_ASAP7_75t_L g12801 ( 
.A1(n_12521),
.A2(n_12079),
.B(n_11800),
.Y(n_12801)
);

OAI21x1_ASAP7_75t_L g12802 ( 
.A1(n_12432),
.A2(n_11803),
.B(n_11792),
.Y(n_12802)
);

INVx2_ASAP7_75t_SL g12803 ( 
.A(n_12409),
.Y(n_12803)
);

INVx1_ASAP7_75t_L g12804 ( 
.A(n_12339),
.Y(n_12804)
);

OAI21x1_ASAP7_75t_L g12805 ( 
.A1(n_12266),
.A2(n_12421),
.B(n_12362),
.Y(n_12805)
);

AND2x4_ASAP7_75t_L g12806 ( 
.A(n_12199),
.B(n_11792),
.Y(n_12806)
);

OAI22xp5_ASAP7_75t_L g12807 ( 
.A1(n_12393),
.A2(n_11948),
.B1(n_11933),
.B2(n_11809),
.Y(n_12807)
);

OAI21x1_ASAP7_75t_L g12808 ( 
.A1(n_12424),
.A2(n_12489),
.B(n_12485),
.Y(n_12808)
);

AOI21x1_ASAP7_75t_L g12809 ( 
.A1(n_12535),
.A2(n_11809),
.B(n_11803),
.Y(n_12809)
);

INVx1_ASAP7_75t_L g12810 ( 
.A(n_12390),
.Y(n_12810)
);

NAND2xp5_ASAP7_75t_L g12811 ( 
.A(n_12512),
.B(n_11831),
.Y(n_12811)
);

NAND3xp33_ASAP7_75t_L g12812 ( 
.A(n_12461),
.B(n_12110),
.C(n_12109),
.Y(n_12812)
);

NAND2xp5_ASAP7_75t_L g12813 ( 
.A(n_12516),
.B(n_11831),
.Y(n_12813)
);

INVx2_ASAP7_75t_L g12814 ( 
.A(n_12447),
.Y(n_12814)
);

INVx2_ASAP7_75t_L g12815 ( 
.A(n_12447),
.Y(n_12815)
);

BUFx2_ASAP7_75t_L g12816 ( 
.A(n_12450),
.Y(n_12816)
);

AOI22x1_ASAP7_75t_L g12817 ( 
.A1(n_12366),
.A2(n_12110),
.B1(n_12115),
.B2(n_12109),
.Y(n_12817)
);

NAND2xp5_ASAP7_75t_L g12818 ( 
.A(n_12403),
.B(n_11890),
.Y(n_12818)
);

AOI22xp33_ASAP7_75t_L g12819 ( 
.A1(n_12606),
.A2(n_12615),
.B1(n_12595),
.B2(n_12554),
.Y(n_12819)
);

INVx2_ASAP7_75t_SL g12820 ( 
.A(n_12214),
.Y(n_12820)
);

INVx1_ASAP7_75t_L g12821 ( 
.A(n_12406),
.Y(n_12821)
);

OAI21x1_ASAP7_75t_L g12822 ( 
.A1(n_12411),
.A2(n_11890),
.B(n_12159),
.Y(n_12822)
);

NAND2xp5_ASAP7_75t_L g12823 ( 
.A(n_12419),
.B(n_12115),
.Y(n_12823)
);

INVx2_ASAP7_75t_L g12824 ( 
.A(n_12250),
.Y(n_12824)
);

AO21x2_ASAP7_75t_L g12825 ( 
.A1(n_12638),
.A2(n_11915),
.B(n_11908),
.Y(n_12825)
);

OAI22xp5_ASAP7_75t_L g12826 ( 
.A1(n_12336),
.A2(n_11915),
.B1(n_11908),
.B2(n_12159),
.Y(n_12826)
);

AO21x2_ASAP7_75t_L g12827 ( 
.A1(n_12383),
.A2(n_12163),
.B(n_1823),
.Y(n_12827)
);

INVx1_ASAP7_75t_L g12828 ( 
.A(n_12295),
.Y(n_12828)
);

AOI22xp33_ASAP7_75t_L g12829 ( 
.A1(n_12541),
.A2(n_12163),
.B1(n_1825),
.B2(n_1823),
.Y(n_12829)
);

INVx1_ASAP7_75t_L g12830 ( 
.A(n_12283),
.Y(n_12830)
);

OAI21x1_ASAP7_75t_L g12831 ( 
.A1(n_12509),
.A2(n_1824),
.B(n_1825),
.Y(n_12831)
);

AOI211xp5_ASAP7_75t_L g12832 ( 
.A1(n_12478),
.A2(n_1828),
.B(n_1826),
.C(n_1827),
.Y(n_12832)
);

AOI22xp33_ASAP7_75t_L g12833 ( 
.A1(n_12543),
.A2(n_1830),
.B1(n_1827),
.B2(n_1829),
.Y(n_12833)
);

OAI21x1_ASAP7_75t_L g12834 ( 
.A1(n_12523),
.A2(n_1829),
.B(n_1832),
.Y(n_12834)
);

AND2x4_ASAP7_75t_SL g12835 ( 
.A(n_12270),
.B(n_1832),
.Y(n_12835)
);

AND2x4_ASAP7_75t_L g12836 ( 
.A(n_12327),
.B(n_1833),
.Y(n_12836)
);

INVx2_ASAP7_75t_SL g12837 ( 
.A(n_12238),
.Y(n_12837)
);

OAI21x1_ASAP7_75t_L g12838 ( 
.A1(n_12528),
.A2(n_1833),
.B(n_1834),
.Y(n_12838)
);

INVx1_ASAP7_75t_L g12839 ( 
.A(n_12456),
.Y(n_12839)
);

AO21x2_ASAP7_75t_L g12840 ( 
.A1(n_12475),
.A2(n_1834),
.B(n_1835),
.Y(n_12840)
);

BUFx12f_ASAP7_75t_L g12841 ( 
.A(n_12307),
.Y(n_12841)
);

O2A1O1Ixp33_ASAP7_75t_SL g12842 ( 
.A1(n_12559),
.A2(n_1837),
.B(n_1835),
.C(n_1836),
.Y(n_12842)
);

INVx1_ASAP7_75t_L g12843 ( 
.A(n_12243),
.Y(n_12843)
);

AND2x2_ASAP7_75t_L g12844 ( 
.A(n_12388),
.B(n_1836),
.Y(n_12844)
);

AOI22xp33_ASAP7_75t_L g12845 ( 
.A1(n_12438),
.A2(n_1840),
.B1(n_1838),
.B2(n_1839),
.Y(n_12845)
);

OAI21x1_ASAP7_75t_L g12846 ( 
.A1(n_12449),
.A2(n_12346),
.B(n_12344),
.Y(n_12846)
);

AND2x2_ASAP7_75t_L g12847 ( 
.A(n_12407),
.B(n_1838),
.Y(n_12847)
);

NAND3xp33_ASAP7_75t_L g12848 ( 
.A(n_12572),
.B(n_1839),
.C(n_1841),
.Y(n_12848)
);

NAND2xp5_ASAP7_75t_L g12849 ( 
.A(n_12355),
.B(n_1841),
.Y(n_12849)
);

OA21x2_ASAP7_75t_L g12850 ( 
.A1(n_12628),
.A2(n_1842),
.B(n_1843),
.Y(n_12850)
);

OAI21x1_ASAP7_75t_L g12851 ( 
.A1(n_12354),
.A2(n_1842),
.B(n_1843),
.Y(n_12851)
);

OAI21x1_ASAP7_75t_L g12852 ( 
.A1(n_12359),
.A2(n_1844),
.B(n_1845),
.Y(n_12852)
);

AO21x2_ASAP7_75t_L g12853 ( 
.A1(n_12414),
.A2(n_1844),
.B(n_1847),
.Y(n_12853)
);

INVx1_ASAP7_75t_SL g12854 ( 
.A(n_12602),
.Y(n_12854)
);

OAI21x1_ASAP7_75t_L g12855 ( 
.A1(n_12239),
.A2(n_1847),
.B(n_1848),
.Y(n_12855)
);

INVx1_ASAP7_75t_L g12856 ( 
.A(n_12558),
.Y(n_12856)
);

A2O1A1Ixp33_ASAP7_75t_L g12857 ( 
.A1(n_12316),
.A2(n_12575),
.B(n_12629),
.C(n_12643),
.Y(n_12857)
);

INVx1_ASAP7_75t_L g12858 ( 
.A(n_12284),
.Y(n_12858)
);

AND2x2_ASAP7_75t_L g12859 ( 
.A(n_12467),
.B(n_1848),
.Y(n_12859)
);

INVx1_ASAP7_75t_L g12860 ( 
.A(n_12259),
.Y(n_12860)
);

INVx3_ASAP7_75t_L g12861 ( 
.A(n_12285),
.Y(n_12861)
);

AOI21xp5_ASAP7_75t_L g12862 ( 
.A1(n_12588),
.A2(n_1849),
.B(n_1850),
.Y(n_12862)
);

AOI22xp33_ASAP7_75t_L g12863 ( 
.A1(n_12308),
.A2(n_12254),
.B1(n_12587),
.B2(n_12569),
.Y(n_12863)
);

HB1xp67_ASAP7_75t_L g12864 ( 
.A(n_12251),
.Y(n_12864)
);

INVx2_ASAP7_75t_L g12865 ( 
.A(n_12522),
.Y(n_12865)
);

INVx1_ASAP7_75t_SL g12866 ( 
.A(n_12455),
.Y(n_12866)
);

NAND2xp5_ASAP7_75t_L g12867 ( 
.A(n_12472),
.B(n_1850),
.Y(n_12867)
);

AOI21xp33_ASAP7_75t_L g12868 ( 
.A1(n_12644),
.A2(n_1851),
.B(n_1852),
.Y(n_12868)
);

OA21x2_ASAP7_75t_L g12869 ( 
.A1(n_12230),
.A2(n_1851),
.B(n_1853),
.Y(n_12869)
);

INVx1_ASAP7_75t_L g12870 ( 
.A(n_12422),
.Y(n_12870)
);

OA21x2_ASAP7_75t_L g12871 ( 
.A1(n_12415),
.A2(n_1853),
.B(n_1854),
.Y(n_12871)
);

NAND2xp5_ASAP7_75t_L g12872 ( 
.A(n_12494),
.B(n_1854),
.Y(n_12872)
);

INVx2_ASAP7_75t_L g12873 ( 
.A(n_12522),
.Y(n_12873)
);

INVx3_ASAP7_75t_L g12874 ( 
.A(n_12218),
.Y(n_12874)
);

AOI22xp33_ASAP7_75t_L g12875 ( 
.A1(n_12566),
.A2(n_1857),
.B1(n_1855),
.B2(n_1856),
.Y(n_12875)
);

INVx1_ASAP7_75t_L g12876 ( 
.A(n_12271),
.Y(n_12876)
);

INVx1_ASAP7_75t_L g12877 ( 
.A(n_12364),
.Y(n_12877)
);

INVx2_ASAP7_75t_L g12878 ( 
.A(n_12522),
.Y(n_12878)
);

A2O1A1Ixp33_ASAP7_75t_L g12879 ( 
.A1(n_12643),
.A2(n_1859),
.B(n_1857),
.C(n_1858),
.Y(n_12879)
);

INVx1_ASAP7_75t_L g12880 ( 
.A(n_12352),
.Y(n_12880)
);

OAI21x1_ASAP7_75t_L g12881 ( 
.A1(n_12410),
.A2(n_1858),
.B(n_1859),
.Y(n_12881)
);

OAI21xp5_ASAP7_75t_L g12882 ( 
.A1(n_12500),
.A2(n_12452),
.B(n_12621),
.Y(n_12882)
);

AO21x2_ASAP7_75t_L g12883 ( 
.A1(n_12468),
.A2(n_12561),
.B(n_12560),
.Y(n_12883)
);

OAI21xp5_ASAP7_75t_L g12884 ( 
.A1(n_12312),
.A2(n_1860),
.B(n_1861),
.Y(n_12884)
);

NAND2xp5_ASAP7_75t_L g12885 ( 
.A(n_12547),
.B(n_1860),
.Y(n_12885)
);

BUFx3_ASAP7_75t_L g12886 ( 
.A(n_12313),
.Y(n_12886)
);

OAI21x1_ASAP7_75t_L g12887 ( 
.A1(n_12418),
.A2(n_1861),
.B(n_1862),
.Y(n_12887)
);

A2O1A1Ixp33_ASAP7_75t_L g12888 ( 
.A1(n_12639),
.A2(n_1864),
.B(n_1862),
.C(n_1863),
.Y(n_12888)
);

AOI22x1_ASAP7_75t_L g12889 ( 
.A1(n_12518),
.A2(n_1866),
.B1(n_1863),
.B2(n_1865),
.Y(n_12889)
);

OR2x2_ASAP7_75t_L g12890 ( 
.A(n_12484),
.B(n_1866),
.Y(n_12890)
);

OAI21x1_ASAP7_75t_L g12891 ( 
.A1(n_12427),
.A2(n_1867),
.B(n_1868),
.Y(n_12891)
);

INVx2_ASAP7_75t_L g12892 ( 
.A(n_12586),
.Y(n_12892)
);

INVx1_ASAP7_75t_L g12893 ( 
.A(n_12294),
.Y(n_12893)
);

OAI21x1_ASAP7_75t_L g12894 ( 
.A1(n_12429),
.A2(n_1867),
.B(n_1868),
.Y(n_12894)
);

CKINVDCx20_ASAP7_75t_R g12895 ( 
.A(n_12386),
.Y(n_12895)
);

INVx1_ASAP7_75t_SL g12896 ( 
.A(n_12215),
.Y(n_12896)
);

INVx1_ASAP7_75t_L g12897 ( 
.A(n_12463),
.Y(n_12897)
);

OA21x2_ASAP7_75t_L g12898 ( 
.A1(n_12324),
.A2(n_1869),
.B(n_1870),
.Y(n_12898)
);

AOI22xp33_ASAP7_75t_L g12899 ( 
.A1(n_12566),
.A2(n_1872),
.B1(n_1870),
.B2(n_1871),
.Y(n_12899)
);

INVx2_ASAP7_75t_L g12900 ( 
.A(n_12586),
.Y(n_12900)
);

INVxp67_ASAP7_75t_L g12901 ( 
.A(n_12408),
.Y(n_12901)
);

INVx2_ASAP7_75t_L g12902 ( 
.A(n_12426),
.Y(n_12902)
);

INVx1_ASAP7_75t_L g12903 ( 
.A(n_12556),
.Y(n_12903)
);

CKINVDCx8_ASAP7_75t_R g12904 ( 
.A(n_12518),
.Y(n_12904)
);

OAI21x1_ASAP7_75t_L g12905 ( 
.A1(n_12457),
.A2(n_1871),
.B(n_1873),
.Y(n_12905)
);

INVx1_ASAP7_75t_L g12906 ( 
.A(n_12562),
.Y(n_12906)
);

INVx3_ASAP7_75t_L g12907 ( 
.A(n_12276),
.Y(n_12907)
);

OAI21x1_ASAP7_75t_L g12908 ( 
.A1(n_12465),
.A2(n_1873),
.B(n_1874),
.Y(n_12908)
);

A2O1A1Ixp33_ASAP7_75t_L g12909 ( 
.A1(n_12580),
.A2(n_1876),
.B(n_1874),
.C(n_1875),
.Y(n_12909)
);

AND2x4_ASAP7_75t_L g12910 ( 
.A(n_12398),
.B(n_1875),
.Y(n_12910)
);

INVx2_ASAP7_75t_SL g12911 ( 
.A(n_12249),
.Y(n_12911)
);

OAI21x1_ASAP7_75t_L g12912 ( 
.A1(n_12392),
.A2(n_1876),
.B(n_1877),
.Y(n_12912)
);

OAI21x1_ASAP7_75t_L g12913 ( 
.A1(n_12394),
.A2(n_1877),
.B(n_1878),
.Y(n_12913)
);

BUFx4f_ASAP7_75t_L g12914 ( 
.A(n_12376),
.Y(n_12914)
);

OAI21x1_ASAP7_75t_L g12915 ( 
.A1(n_12529),
.A2(n_1879),
.B(n_1880),
.Y(n_12915)
);

BUFx12f_ASAP7_75t_L g12916 ( 
.A(n_12356),
.Y(n_12916)
);

AO21x2_ASAP7_75t_L g12917 ( 
.A1(n_12397),
.A2(n_1879),
.B(n_1880),
.Y(n_12917)
);

INVx1_ASAP7_75t_L g12918 ( 
.A(n_12357),
.Y(n_12918)
);

BUFx2_ASAP7_75t_L g12919 ( 
.A(n_12437),
.Y(n_12919)
);

INVx1_ASAP7_75t_L g12920 ( 
.A(n_12573),
.Y(n_12920)
);

OAI21x1_ASAP7_75t_L g12921 ( 
.A1(n_12405),
.A2(n_1881),
.B(n_1882),
.Y(n_12921)
);

OAI21xp5_ASAP7_75t_L g12922 ( 
.A1(n_12439),
.A2(n_1881),
.B(n_1882),
.Y(n_12922)
);

INVx1_ASAP7_75t_L g12923 ( 
.A(n_12577),
.Y(n_12923)
);

NAND2x1_ASAP7_75t_L g12924 ( 
.A(n_12325),
.B(n_1883),
.Y(n_12924)
);

AOI22xp33_ASAP7_75t_L g12925 ( 
.A1(n_12314),
.A2(n_1885),
.B1(n_1883),
.B2(n_1884),
.Y(n_12925)
);

OAI22xp5_ASAP7_75t_L g12926 ( 
.A1(n_12205),
.A2(n_1886),
.B1(n_1884),
.B2(n_1885),
.Y(n_12926)
);

INVx2_ASAP7_75t_L g12927 ( 
.A(n_12262),
.Y(n_12927)
);

OAI21x1_ASAP7_75t_L g12928 ( 
.A1(n_12462),
.A2(n_1886),
.B(n_1887),
.Y(n_12928)
);

INVx1_ASAP7_75t_L g12929 ( 
.A(n_12582),
.Y(n_12929)
);

INVx2_ASAP7_75t_L g12930 ( 
.A(n_12417),
.Y(n_12930)
);

BUFx6f_ASAP7_75t_L g12931 ( 
.A(n_12193),
.Y(n_12931)
);

OA21x2_ASAP7_75t_L g12932 ( 
.A1(n_12328),
.A2(n_1888),
.B(n_1889),
.Y(n_12932)
);

OAI21x1_ASAP7_75t_L g12933 ( 
.A1(n_12367),
.A2(n_1888),
.B(n_1889),
.Y(n_12933)
);

AOI21xp5_ASAP7_75t_L g12934 ( 
.A1(n_12568),
.A2(n_1890),
.B(n_1891),
.Y(n_12934)
);

OAI21x1_ASAP7_75t_L g12935 ( 
.A1(n_12486),
.A2(n_12492),
.B(n_12532),
.Y(n_12935)
);

INVx1_ASAP7_75t_L g12936 ( 
.A(n_12622),
.Y(n_12936)
);

INVx1_ASAP7_75t_L g12937 ( 
.A(n_12416),
.Y(n_12937)
);

OAI21x1_ASAP7_75t_L g12938 ( 
.A1(n_12601),
.A2(n_1891),
.B(n_1892),
.Y(n_12938)
);

NAND3xp33_ASAP7_75t_L g12939 ( 
.A(n_12443),
.B(n_1892),
.C(n_1894),
.Y(n_12939)
);

AOI21x1_ASAP7_75t_L g12940 ( 
.A1(n_12510),
.A2(n_1894),
.B(n_1895),
.Y(n_12940)
);

OAI21x1_ASAP7_75t_L g12941 ( 
.A1(n_12545),
.A2(n_1896),
.B(n_1897),
.Y(n_12941)
);

OAI21xp5_ASAP7_75t_L g12942 ( 
.A1(n_12612),
.A2(n_12617),
.B(n_12583),
.Y(n_12942)
);

A2O1A1Ixp33_ASAP7_75t_L g12943 ( 
.A1(n_12631),
.A2(n_1898),
.B(n_1896),
.C(n_1897),
.Y(n_12943)
);

AOI22x1_ASAP7_75t_L g12944 ( 
.A1(n_12531),
.A2(n_1900),
.B1(n_1898),
.B2(n_1899),
.Y(n_12944)
);

AO21x2_ASAP7_75t_L g12945 ( 
.A1(n_12435),
.A2(n_1899),
.B(n_1900),
.Y(n_12945)
);

INVx1_ASAP7_75t_L g12946 ( 
.A(n_12520),
.Y(n_12946)
);

OAI21x1_ASAP7_75t_L g12947 ( 
.A1(n_12625),
.A2(n_1901),
.B(n_1902),
.Y(n_12947)
);

OAI22xp33_ASAP7_75t_L g12948 ( 
.A1(n_12534),
.A2(n_1903),
.B1(n_1901),
.B2(n_1902),
.Y(n_12948)
);

AOI22xp5_ASAP7_75t_L g12949 ( 
.A1(n_12437),
.A2(n_1905),
.B1(n_1903),
.B2(n_1904),
.Y(n_12949)
);

AO31x2_ASAP7_75t_L g12950 ( 
.A1(n_12286),
.A2(n_1907),
.A3(n_1905),
.B(n_1906),
.Y(n_12950)
);

OR2x2_ASAP7_75t_L g12951 ( 
.A(n_12487),
.B(n_1906),
.Y(n_12951)
);

INVx1_ASAP7_75t_L g12952 ( 
.A(n_12374),
.Y(n_12952)
);

INVx1_ASAP7_75t_SL g12953 ( 
.A(n_12347),
.Y(n_12953)
);

OAI21x1_ASAP7_75t_L g12954 ( 
.A1(n_12633),
.A2(n_1907),
.B(n_1908),
.Y(n_12954)
);

AOI21xp5_ASAP7_75t_L g12955 ( 
.A1(n_12473),
.A2(n_1908),
.B(n_1909),
.Y(n_12955)
);

OAI21x1_ASAP7_75t_L g12956 ( 
.A1(n_12641),
.A2(n_12480),
.B(n_12257),
.Y(n_12956)
);

NAND2xp5_ASAP7_75t_L g12957 ( 
.A(n_12507),
.B(n_1909),
.Y(n_12957)
);

OAI21x1_ASAP7_75t_L g12958 ( 
.A1(n_12493),
.A2(n_1910),
.B(n_1911),
.Y(n_12958)
);

OR2x6_ASAP7_75t_L g12959 ( 
.A(n_12581),
.B(n_12497),
.Y(n_12959)
);

OAI21x1_ASAP7_75t_L g12960 ( 
.A1(n_12501),
.A2(n_1911),
.B(n_1912),
.Y(n_12960)
);

INVx2_ASAP7_75t_L g12961 ( 
.A(n_12459),
.Y(n_12961)
);

INVx4_ASAP7_75t_L g12962 ( 
.A(n_12368),
.Y(n_12962)
);

OAI21xp33_ASAP7_75t_SL g12963 ( 
.A1(n_12428),
.A2(n_1914),
.B(n_1915),
.Y(n_12963)
);

OAI21xp5_ASAP7_75t_L g12964 ( 
.A1(n_12551),
.A2(n_1914),
.B(n_1915),
.Y(n_12964)
);

AND2x2_ASAP7_75t_L g12965 ( 
.A(n_12464),
.B(n_1916),
.Y(n_12965)
);

NAND2xp5_ASAP7_75t_L g12966 ( 
.A(n_12610),
.B(n_1916),
.Y(n_12966)
);

NAND2xp5_ASAP7_75t_L g12967 ( 
.A(n_12637),
.B(n_1917),
.Y(n_12967)
);

BUFx2_ASAP7_75t_SL g12968 ( 
.A(n_12237),
.Y(n_12968)
);

OAI21x1_ASAP7_75t_SL g12969 ( 
.A1(n_12348),
.A2(n_1917),
.B(n_1918),
.Y(n_12969)
);

OAI211xp5_ASAP7_75t_L g12970 ( 
.A1(n_12436),
.A2(n_12423),
.B(n_12504),
.C(n_12593),
.Y(n_12970)
);

A2O1A1Ixp33_ASAP7_75t_L g12971 ( 
.A1(n_12589),
.A2(n_1920),
.B(n_1918),
.C(n_1919),
.Y(n_12971)
);

INVx1_ASAP7_75t_L g12972 ( 
.A(n_12337),
.Y(n_12972)
);

OAI21x1_ASAP7_75t_L g12973 ( 
.A1(n_12451),
.A2(n_1919),
.B(n_1920),
.Y(n_12973)
);

NAND2x1p5_ASAP7_75t_L g12974 ( 
.A(n_12291),
.B(n_1921),
.Y(n_12974)
);

OAI21x1_ASAP7_75t_L g12975 ( 
.A1(n_12224),
.A2(n_1922),
.B(n_1923),
.Y(n_12975)
);

NOR2x1_ASAP7_75t_SL g12976 ( 
.A(n_12317),
.B(n_1922),
.Y(n_12976)
);

HB1xp67_ASAP7_75t_L g12977 ( 
.A(n_12481),
.Y(n_12977)
);

O2A1O1Ixp33_ASAP7_75t_L g12978 ( 
.A1(n_12396),
.A2(n_1925),
.B(n_1923),
.C(n_1924),
.Y(n_12978)
);

CKINVDCx5p33_ASAP7_75t_R g12979 ( 
.A(n_12252),
.Y(n_12979)
);

NAND2xp5_ASAP7_75t_L g12980 ( 
.A(n_12544),
.B(n_1924),
.Y(n_12980)
);

INVx1_ASAP7_75t_L g12981 ( 
.A(n_12351),
.Y(n_12981)
);

OAI21x1_ASAP7_75t_L g12982 ( 
.A1(n_12350),
.A2(n_1925),
.B(n_1926),
.Y(n_12982)
);

INVx2_ASAP7_75t_L g12983 ( 
.A(n_12477),
.Y(n_12983)
);

OAI21x1_ASAP7_75t_L g12984 ( 
.A1(n_12380),
.A2(n_1926),
.B(n_1927),
.Y(n_12984)
);

AND2x4_ASAP7_75t_L g12985 ( 
.A(n_12391),
.B(n_1927),
.Y(n_12985)
);

BUFx3_ASAP7_75t_L g12986 ( 
.A(n_12292),
.Y(n_12986)
);

INVx1_ASAP7_75t_L g12987 ( 
.A(n_12544),
.Y(n_12987)
);

OAI21x1_ASAP7_75t_L g12988 ( 
.A1(n_12476),
.A2(n_12590),
.B(n_12608),
.Y(n_12988)
);

OAI21x1_ASAP7_75t_L g12989 ( 
.A1(n_12540),
.A2(n_1928),
.B(n_1929),
.Y(n_12989)
);

BUFx3_ASAP7_75t_L g12990 ( 
.A(n_12345),
.Y(n_12990)
);

INVx2_ASAP7_75t_L g12991 ( 
.A(n_12592),
.Y(n_12991)
);

AND2x4_ASAP7_75t_L g12992 ( 
.A(n_12400),
.B(n_1928),
.Y(n_12992)
);

OAI21xp33_ASAP7_75t_SL g12993 ( 
.A1(n_12195),
.A2(n_1930),
.B(n_1931),
.Y(n_12993)
);

OR2x2_ASAP7_75t_L g12994 ( 
.A(n_12609),
.B(n_1931),
.Y(n_12994)
);

OAI21xp5_ASAP7_75t_L g12995 ( 
.A1(n_12594),
.A2(n_1932),
.B(n_1933),
.Y(n_12995)
);

INVx1_ASAP7_75t_L g12996 ( 
.A(n_12592),
.Y(n_12996)
);

BUFx3_ASAP7_75t_L g12997 ( 
.A(n_12320),
.Y(n_12997)
);

NAND2xp5_ASAP7_75t_L g12998 ( 
.A(n_12624),
.B(n_1933),
.Y(n_12998)
);

INVx3_ASAP7_75t_L g12999 ( 
.A(n_12404),
.Y(n_12999)
);

AND2x2_ASAP7_75t_L g13000 ( 
.A(n_12448),
.B(n_1934),
.Y(n_13000)
);

AND2x4_ASAP7_75t_L g13001 ( 
.A(n_12377),
.B(n_1935),
.Y(n_13001)
);

O2A1O1Ixp33_ASAP7_75t_L g13002 ( 
.A1(n_12420),
.A2(n_1937),
.B(n_1935),
.C(n_1936),
.Y(n_13002)
);

BUFx6f_ASAP7_75t_L g13003 ( 
.A(n_12193),
.Y(n_13003)
);

OAI21xp5_ASAP7_75t_L g13004 ( 
.A1(n_12607),
.A2(n_1937),
.B(n_1938),
.Y(n_13004)
);

OAI21x1_ASAP7_75t_L g13005 ( 
.A1(n_12536),
.A2(n_12513),
.B(n_12442),
.Y(n_13005)
);

OAI21x1_ASAP7_75t_L g13006 ( 
.A1(n_12531),
.A2(n_1938),
.B(n_1939),
.Y(n_13006)
);

AO21x2_ASAP7_75t_L g13007 ( 
.A1(n_12469),
.A2(n_1939),
.B(n_1940),
.Y(n_13007)
);

OA21x2_ASAP7_75t_L g13008 ( 
.A1(n_12370),
.A2(n_1940),
.B(n_1941),
.Y(n_13008)
);

OAI21x1_ASAP7_75t_L g13009 ( 
.A1(n_12302),
.A2(n_1941),
.B(n_1942),
.Y(n_13009)
);

AND2x2_ASAP7_75t_L g13010 ( 
.A(n_12441),
.B(n_1943),
.Y(n_13010)
);

INVx1_ASAP7_75t_L g13011 ( 
.A(n_12361),
.Y(n_13011)
);

O2A1O1Ixp33_ASAP7_75t_SL g13012 ( 
.A1(n_12387),
.A2(n_1945),
.B(n_1943),
.C(n_1944),
.Y(n_13012)
);

NOR2xp33_ASAP7_75t_R g13013 ( 
.A(n_12289),
.B(n_1944),
.Y(n_13013)
);

INVxp67_ASAP7_75t_SL g13014 ( 
.A(n_12630),
.Y(n_13014)
);

BUFx4f_ASAP7_75t_L g13015 ( 
.A(n_12207),
.Y(n_13015)
);

OAI21xp5_ASAP7_75t_L g13016 ( 
.A1(n_12546),
.A2(n_12570),
.B(n_12511),
.Y(n_13016)
);

OA21x2_ASAP7_75t_L g13017 ( 
.A1(n_12373),
.A2(n_1945),
.B(n_1946),
.Y(n_13017)
);

INVx3_ASAP7_75t_L g13018 ( 
.A(n_12404),
.Y(n_13018)
);

OAI21x1_ASAP7_75t_L g13019 ( 
.A1(n_12372),
.A2(n_1946),
.B(n_1947),
.Y(n_13019)
);

OA21x2_ASAP7_75t_L g13020 ( 
.A1(n_12382),
.A2(n_12381),
.B(n_12258),
.Y(n_13020)
);

INVx1_ASAP7_75t_L g13021 ( 
.A(n_12375),
.Y(n_13021)
);

INVx4_ASAP7_75t_SL g13022 ( 
.A(n_12479),
.Y(n_13022)
);

OAI21x1_ASAP7_75t_L g13023 ( 
.A1(n_12395),
.A2(n_1948),
.B(n_1949),
.Y(n_13023)
);

OR2x2_ASAP7_75t_L g13024 ( 
.A(n_12574),
.B(n_1948),
.Y(n_13024)
);

OAI21x1_ASAP7_75t_L g13025 ( 
.A1(n_12488),
.A2(n_12490),
.B(n_12498),
.Y(n_13025)
);

A2O1A1Ixp33_ASAP7_75t_L g13026 ( 
.A1(n_12539),
.A2(n_1951),
.B(n_1949),
.C(n_1950),
.Y(n_13026)
);

OAI21x1_ASAP7_75t_L g13027 ( 
.A1(n_12515),
.A2(n_1950),
.B(n_1951),
.Y(n_13027)
);

INVx1_ASAP7_75t_L g13028 ( 
.A(n_12596),
.Y(n_13028)
);

OAI221xp5_ASAP7_75t_L g13029 ( 
.A1(n_12479),
.A2(n_1954),
.B1(n_1952),
.B2(n_1953),
.C(n_1955),
.Y(n_13029)
);

AOI221xp5_ASAP7_75t_L g13030 ( 
.A1(n_12600),
.A2(n_1956),
.B1(n_1952),
.B2(n_1954),
.C(n_1957),
.Y(n_13030)
);

OR2x2_ASAP7_75t_L g13031 ( 
.A(n_12816),
.B(n_12552),
.Y(n_13031)
);

A2O1A1Ixp33_ASAP7_75t_L g13032 ( 
.A1(n_12670),
.A2(n_12514),
.B(n_12623),
.C(n_12524),
.Y(n_13032)
);

OAI22xp5_ASAP7_75t_L g13033 ( 
.A1(n_12649),
.A2(n_12506),
.B1(n_12384),
.B2(n_12496),
.Y(n_13033)
);

NAND2xp5_ASAP7_75t_L g13034 ( 
.A(n_12883),
.B(n_12207),
.Y(n_13034)
);

NAND2xp5_ASAP7_75t_L g13035 ( 
.A(n_12937),
.B(n_12234),
.Y(n_13035)
);

INVx1_ASAP7_75t_L g13036 ( 
.A(n_12718),
.Y(n_13036)
);

OR2x6_ASAP7_75t_L g13037 ( 
.A(n_12968),
.B(n_12335),
.Y(n_13037)
);

O2A1O1Ixp33_ASAP7_75t_L g13038 ( 
.A1(n_12684),
.A2(n_12491),
.B(n_1959),
.C(n_1956),
.Y(n_13038)
);

NAND2xp5_ASAP7_75t_L g13039 ( 
.A(n_12901),
.B(n_12234),
.Y(n_13039)
);

INVx1_ASAP7_75t_L g13040 ( 
.A(n_12653),
.Y(n_13040)
);

NAND2xp5_ASAP7_75t_SL g13041 ( 
.A(n_12701),
.B(n_12241),
.Y(n_13041)
);

AND2x2_ASAP7_75t_L g13042 ( 
.A(n_12650),
.B(n_12296),
.Y(n_13042)
);

INVx1_ASAP7_75t_L g13043 ( 
.A(n_12657),
.Y(n_13043)
);

OA21x2_ASAP7_75t_L g13044 ( 
.A1(n_12688),
.A2(n_12287),
.B(n_12241),
.Y(n_13044)
);

AND2x2_ASAP7_75t_L g13045 ( 
.A(n_12671),
.B(n_12287),
.Y(n_13045)
);

OAI21x1_ASAP7_75t_L g13046 ( 
.A1(n_12647),
.A2(n_12353),
.B(n_12301),
.Y(n_13046)
);

AO31x2_ASAP7_75t_L g13047 ( 
.A1(n_12717),
.A2(n_12918),
.A3(n_12981),
.B(n_12972),
.Y(n_13047)
);

AO21x2_ASAP7_75t_L g13048 ( 
.A1(n_12759),
.A2(n_12353),
.B(n_12301),
.Y(n_13048)
);

AND2x2_ASAP7_75t_L g13049 ( 
.A(n_12774),
.B(n_12666),
.Y(n_13049)
);

AO21x2_ASAP7_75t_L g13050 ( 
.A1(n_12864),
.A2(n_1958),
.B(n_1959),
.Y(n_13050)
);

OAI21xp33_ASAP7_75t_L g13051 ( 
.A1(n_12745),
.A2(n_1958),
.B(n_1960),
.Y(n_13051)
);

OAI21x1_ASAP7_75t_L g13052 ( 
.A1(n_12758),
.A2(n_1960),
.B(n_1961),
.Y(n_13052)
);

AO31x2_ASAP7_75t_L g13053 ( 
.A1(n_12946),
.A2(n_1963),
.A3(n_1961),
.B(n_1962),
.Y(n_13053)
);

INVx1_ASAP7_75t_SL g13054 ( 
.A(n_12896),
.Y(n_13054)
);

HB1xp67_ASAP7_75t_L g13055 ( 
.A(n_12697),
.Y(n_13055)
);

NOR2x1_ASAP7_75t_SL g13056 ( 
.A(n_12778),
.B(n_1962),
.Y(n_13056)
);

NAND2xp5_ASAP7_75t_L g13057 ( 
.A(n_12858),
.B(n_1963),
.Y(n_13057)
);

AO31x2_ASAP7_75t_L g13058 ( 
.A1(n_13011),
.A2(n_1966),
.A3(n_1964),
.B(n_1965),
.Y(n_13058)
);

AOI21xp5_ASAP7_75t_L g13059 ( 
.A1(n_12680),
.A2(n_1965),
.B(n_1966),
.Y(n_13059)
);

HB1xp67_ASAP7_75t_L g13060 ( 
.A(n_12754),
.Y(n_13060)
);

OAI21x1_ASAP7_75t_L g13061 ( 
.A1(n_12746),
.A2(n_1968),
.B(n_1969),
.Y(n_13061)
);

AOI21xp5_ASAP7_75t_L g13062 ( 
.A1(n_12709),
.A2(n_1969),
.B(n_1970),
.Y(n_13062)
);

INVx2_ASAP7_75t_SL g13063 ( 
.A(n_12728),
.Y(n_13063)
);

OAI21x1_ASAP7_75t_SL g13064 ( 
.A1(n_12976),
.A2(n_1971),
.B(n_1972),
.Y(n_13064)
);

INVx2_ASAP7_75t_L g13065 ( 
.A(n_12707),
.Y(n_13065)
);

HB1xp67_ASAP7_75t_L g13066 ( 
.A(n_13025),
.Y(n_13066)
);

INVx1_ASAP7_75t_L g13067 ( 
.A(n_12659),
.Y(n_13067)
);

AND2x2_ASAP7_75t_L g13068 ( 
.A(n_12673),
.B(n_1972),
.Y(n_13068)
);

BUFx10_ASAP7_75t_L g13069 ( 
.A(n_12728),
.Y(n_13069)
);

OAI21x1_ASAP7_75t_L g13070 ( 
.A1(n_12740),
.A2(n_12808),
.B(n_12805),
.Y(n_13070)
);

HB1xp67_ASAP7_75t_L g13071 ( 
.A(n_12877),
.Y(n_13071)
);

OAI21x1_ASAP7_75t_L g13072 ( 
.A1(n_12822),
.A2(n_1973),
.B(n_1974),
.Y(n_13072)
);

BUFx2_ASAP7_75t_L g13073 ( 
.A(n_12919),
.Y(n_13073)
);

HB1xp67_ASAP7_75t_L g13074 ( 
.A(n_13021),
.Y(n_13074)
);

INVx3_ASAP7_75t_L g13075 ( 
.A(n_12733),
.Y(n_13075)
);

OAI21xp5_ASAP7_75t_L g13076 ( 
.A1(n_12682),
.A2(n_1973),
.B(n_1974),
.Y(n_13076)
);

AND2x4_ASAP7_75t_L g13077 ( 
.A(n_12907),
.B(n_1975),
.Y(n_13077)
);

NAND2xp33_ASAP7_75t_R g13078 ( 
.A(n_13013),
.B(n_1975),
.Y(n_13078)
);

OAI21x1_ASAP7_75t_SL g13079 ( 
.A1(n_13016),
.A2(n_1976),
.B(n_1977),
.Y(n_13079)
);

INVx1_ASAP7_75t_L g13080 ( 
.A(n_12664),
.Y(n_13080)
);

A2O1A1Ixp33_ASAP7_75t_L g13081 ( 
.A1(n_12793),
.A2(n_1979),
.B(n_1977),
.C(n_1978),
.Y(n_13081)
);

AND2x2_ASAP7_75t_L g13082 ( 
.A(n_12720),
.B(n_1978),
.Y(n_13082)
);

HB1xp67_ASAP7_75t_L g13083 ( 
.A(n_12977),
.Y(n_13083)
);

OA21x2_ASAP7_75t_L g13084 ( 
.A1(n_12828),
.A2(n_1980),
.B(n_1981),
.Y(n_13084)
);

INVx2_ASAP7_75t_L g13085 ( 
.A(n_12707),
.Y(n_13085)
);

BUFx8_ASAP7_75t_SL g13086 ( 
.A(n_12769),
.Y(n_13086)
);

OA21x2_ASAP7_75t_L g13087 ( 
.A1(n_12824),
.A2(n_1980),
.B(n_1981),
.Y(n_13087)
);

AND2x2_ASAP7_75t_L g13088 ( 
.A(n_12695),
.B(n_1982),
.Y(n_13088)
);

INVxp67_ASAP7_75t_L g13089 ( 
.A(n_12898),
.Y(n_13089)
);

INVx2_ASAP7_75t_L g13090 ( 
.A(n_12652),
.Y(n_13090)
);

AOI221xp5_ASAP7_75t_L g13091 ( 
.A1(n_12807),
.A2(n_12677),
.B1(n_12826),
.B2(n_12661),
.C(n_12868),
.Y(n_13091)
);

HB1xp67_ASAP7_75t_L g13092 ( 
.A(n_12770),
.Y(n_13092)
);

INVx1_ASAP7_75t_L g13093 ( 
.A(n_12672),
.Y(n_13093)
);

INVx1_ASAP7_75t_L g13094 ( 
.A(n_12678),
.Y(n_13094)
);

AND2x4_ASAP7_75t_L g13095 ( 
.A(n_12773),
.B(n_1983),
.Y(n_13095)
);

INVxp33_ASAP7_75t_SL g13096 ( 
.A(n_12681),
.Y(n_13096)
);

OAI21x1_ASAP7_75t_L g13097 ( 
.A1(n_12801),
.A2(n_12802),
.B(n_12658),
.Y(n_13097)
);

INVx1_ASAP7_75t_L g13098 ( 
.A(n_12692),
.Y(n_13098)
);

OAI21x1_ASAP7_75t_L g13099 ( 
.A1(n_12656),
.A2(n_1984),
.B(n_1985),
.Y(n_13099)
);

BUFx8_ASAP7_75t_SL g13100 ( 
.A(n_12895),
.Y(n_13100)
);

INVx2_ASAP7_75t_L g13101 ( 
.A(n_12892),
.Y(n_13101)
);

NOR2x1_ASAP7_75t_L g13102 ( 
.A(n_12959),
.B(n_1984),
.Y(n_13102)
);

INVxp67_ASAP7_75t_SL g13103 ( 
.A(n_12742),
.Y(n_13103)
);

OAI21x1_ASAP7_75t_L g13104 ( 
.A1(n_12809),
.A2(n_1985),
.B(n_1986),
.Y(n_13104)
);

INVx1_ASAP7_75t_L g13105 ( 
.A(n_12694),
.Y(n_13105)
);

AOI21xp5_ASAP7_75t_L g13106 ( 
.A1(n_12749),
.A2(n_1986),
.B(n_1987),
.Y(n_13106)
);

AOI222xp33_ASAP7_75t_L g13107 ( 
.A1(n_12739),
.A2(n_1990),
.B1(n_1992),
.B2(n_1988),
.C1(n_1989),
.C2(n_1991),
.Y(n_13107)
);

NAND2x1p5_ASAP7_75t_L g13108 ( 
.A(n_12679),
.B(n_1988),
.Y(n_13108)
);

OR2x2_ASAP7_75t_L g13109 ( 
.A(n_12790),
.B(n_1991),
.Y(n_13109)
);

AO31x2_ASAP7_75t_L g13110 ( 
.A1(n_12645),
.A2(n_1995),
.A3(n_1993),
.B(n_1994),
.Y(n_13110)
);

AOI222xp33_ASAP7_75t_L g13111 ( 
.A1(n_12686),
.A2(n_1997),
.B1(n_1999),
.B2(n_1993),
.C1(n_1996),
.C2(n_1998),
.Y(n_13111)
);

OAI21x1_ASAP7_75t_L g13112 ( 
.A1(n_12732),
.A2(n_1997),
.B(n_1998),
.Y(n_13112)
);

AND2x4_ASAP7_75t_L g13113 ( 
.A(n_13022),
.B(n_1999),
.Y(n_13113)
);

NAND2xp5_ASAP7_75t_L g13114 ( 
.A(n_12830),
.B(n_2000),
.Y(n_13114)
);

AND2x4_ASAP7_75t_L g13115 ( 
.A(n_13022),
.B(n_2001),
.Y(n_13115)
);

AOI21x1_ASAP7_75t_L g13116 ( 
.A1(n_12959),
.A2(n_2002),
.B(n_2003),
.Y(n_13116)
);

AOI22xp33_ASAP7_75t_L g13117 ( 
.A1(n_12753),
.A2(n_2005),
.B1(n_2002),
.B2(n_2004),
.Y(n_13117)
);

OA21x2_ASAP7_75t_L g13118 ( 
.A1(n_12865),
.A2(n_12878),
.B(n_12873),
.Y(n_13118)
);

INVx2_ASAP7_75t_L g13119 ( 
.A(n_12900),
.Y(n_13119)
);

NAND2xp5_ASAP7_75t_L g13120 ( 
.A(n_12821),
.B(n_12810),
.Y(n_13120)
);

OAI21xp33_ASAP7_75t_L g13121 ( 
.A1(n_12756),
.A2(n_2004),
.B(n_2005),
.Y(n_13121)
);

INVx1_ASAP7_75t_L g13122 ( 
.A(n_12696),
.Y(n_13122)
);

OA21x2_ASAP7_75t_L g13123 ( 
.A1(n_12856),
.A2(n_2006),
.B(n_2007),
.Y(n_13123)
);

CKINVDCx14_ASAP7_75t_R g13124 ( 
.A(n_12914),
.Y(n_13124)
);

NAND2xp5_ASAP7_75t_L g13125 ( 
.A(n_12823),
.B(n_12715),
.Y(n_13125)
);

NOR2x1_ASAP7_75t_SL g13126 ( 
.A(n_12747),
.B(n_12648),
.Y(n_13126)
);

CKINVDCx5p33_ASAP7_75t_R g13127 ( 
.A(n_12748),
.Y(n_13127)
);

NAND2xp5_ASAP7_75t_L g13128 ( 
.A(n_12818),
.B(n_2006),
.Y(n_13128)
);

AOI21xp5_ASAP7_75t_L g13129 ( 
.A1(n_12734),
.A2(n_2007),
.B(n_2009),
.Y(n_13129)
);

OAI21xp5_ASAP7_75t_L g13130 ( 
.A1(n_12857),
.A2(n_2009),
.B(n_2010),
.Y(n_13130)
);

AO21x2_ASAP7_75t_L g13131 ( 
.A1(n_12698),
.A2(n_2010),
.B(n_2011),
.Y(n_13131)
);

INVx1_ASAP7_75t_L g13132 ( 
.A(n_12703),
.Y(n_13132)
);

HB1xp67_ASAP7_75t_L g13133 ( 
.A(n_12660),
.Y(n_13133)
);

AOI21x1_ASAP7_75t_L g13134 ( 
.A1(n_12940),
.A2(n_2011),
.B(n_2012),
.Y(n_13134)
);

CKINVDCx20_ASAP7_75t_R g13135 ( 
.A(n_12685),
.Y(n_13135)
);

AND2x2_ASAP7_75t_L g13136 ( 
.A(n_12866),
.B(n_2013),
.Y(n_13136)
);

AOI22xp5_ASAP7_75t_L g13137 ( 
.A1(n_12731),
.A2(n_2016),
.B1(n_2014),
.B2(n_2015),
.Y(n_13137)
);

NAND2xp5_ASAP7_75t_L g13138 ( 
.A(n_12811),
.B(n_2014),
.Y(n_13138)
);

OAI21x1_ASAP7_75t_SL g13139 ( 
.A1(n_12882),
.A2(n_2015),
.B(n_2016),
.Y(n_13139)
);

NAND2xp5_ASAP7_75t_L g13140 ( 
.A(n_12813),
.B(n_2017),
.Y(n_13140)
);

NAND2xp5_ASAP7_75t_L g13141 ( 
.A(n_12843),
.B(n_2017),
.Y(n_13141)
);

NOR2xp33_ASAP7_75t_L g13142 ( 
.A(n_12711),
.B(n_2018),
.Y(n_13142)
);

INVx2_ASAP7_75t_L g13143 ( 
.A(n_12689),
.Y(n_13143)
);

NOR2xp67_ASAP7_75t_SL g13144 ( 
.A(n_12711),
.B(n_2018),
.Y(n_13144)
);

BUFx2_ASAP7_75t_L g13145 ( 
.A(n_13020),
.Y(n_13145)
);

INVx6_ASAP7_75t_L g13146 ( 
.A(n_12713),
.Y(n_13146)
);

NAND2xp5_ASAP7_75t_L g13147 ( 
.A(n_12839),
.B(n_2019),
.Y(n_13147)
);

INVx1_ASAP7_75t_L g13148 ( 
.A(n_12741),
.Y(n_13148)
);

OAI21xp5_ASAP7_75t_L g13149 ( 
.A1(n_12737),
.A2(n_2020),
.B(n_2021),
.Y(n_13149)
);

AO21x2_ASAP7_75t_L g13150 ( 
.A1(n_12729),
.A2(n_2020),
.B(n_2021),
.Y(n_13150)
);

AOI21xp5_ASAP7_75t_L g13151 ( 
.A1(n_12787),
.A2(n_2022),
.B(n_2023),
.Y(n_13151)
);

A2O1A1Ixp33_ASAP7_75t_L g13152 ( 
.A1(n_12669),
.A2(n_12832),
.B(n_13002),
.C(n_12788),
.Y(n_13152)
);

OAI21x1_ASAP7_75t_L g13153 ( 
.A1(n_12727),
.A2(n_2022),
.B(n_2023),
.Y(n_13153)
);

AO21x2_ASAP7_75t_L g13154 ( 
.A1(n_12849),
.A2(n_2024),
.B(n_2025),
.Y(n_13154)
);

AND2x2_ASAP7_75t_L g13155 ( 
.A(n_12814),
.B(n_2025),
.Y(n_13155)
);

AOI21xp5_ASAP7_75t_L g13156 ( 
.A1(n_12764),
.A2(n_12781),
.B(n_12757),
.Y(n_13156)
);

AOI21xp5_ASAP7_75t_L g13157 ( 
.A1(n_12782),
.A2(n_2026),
.B(n_2027),
.Y(n_13157)
);

OAI21x1_ASAP7_75t_L g13158 ( 
.A1(n_12667),
.A2(n_2026),
.B(n_2028),
.Y(n_13158)
);

INVx1_ASAP7_75t_L g13159 ( 
.A(n_12744),
.Y(n_13159)
);

NAND2xp5_ASAP7_75t_L g13160 ( 
.A(n_12743),
.B(n_2028),
.Y(n_13160)
);

AND2x2_ASAP7_75t_L g13161 ( 
.A(n_12815),
.B(n_2029),
.Y(n_13161)
);

INVx1_ASAP7_75t_L g13162 ( 
.A(n_12719),
.Y(n_13162)
);

AOI21x1_ASAP7_75t_L g13163 ( 
.A1(n_12767),
.A2(n_2029),
.B(n_2030),
.Y(n_13163)
);

CKINVDCx5p33_ASAP7_75t_R g13164 ( 
.A(n_12775),
.Y(n_13164)
);

OA21x2_ASAP7_75t_L g13165 ( 
.A1(n_12956),
.A2(n_2031),
.B(n_2032),
.Y(n_13165)
);

OAI21xp33_ASAP7_75t_L g13166 ( 
.A1(n_12863),
.A2(n_2031),
.B(n_2032),
.Y(n_13166)
);

AOI21xp5_ASAP7_75t_L g13167 ( 
.A1(n_12726),
.A2(n_2033),
.B(n_2034),
.Y(n_13167)
);

NAND2xp5_ASAP7_75t_L g13168 ( 
.A(n_12765),
.B(n_2034),
.Y(n_13168)
);

BUFx2_ASAP7_75t_L g13169 ( 
.A(n_13014),
.Y(n_13169)
);

NAND2xp5_ASAP7_75t_L g13170 ( 
.A(n_12869),
.B(n_2035),
.Y(n_13170)
);

CKINVDCx20_ASAP7_75t_R g13171 ( 
.A(n_12979),
.Y(n_13171)
);

INVx2_ASAP7_75t_L g13172 ( 
.A(n_12806),
.Y(n_13172)
);

NAND2xp5_ASAP7_75t_L g13173 ( 
.A(n_12651),
.B(n_2035),
.Y(n_13173)
);

OR2x6_ASAP7_75t_L g13174 ( 
.A(n_12924),
.B(n_2036),
.Y(n_13174)
);

INVx1_ASAP7_75t_L g13175 ( 
.A(n_12723),
.Y(n_13175)
);

OR2x2_ASAP7_75t_L g13176 ( 
.A(n_12783),
.B(n_2036),
.Y(n_13176)
);

AOI21xp5_ASAP7_75t_L g13177 ( 
.A1(n_12712),
.A2(n_2037),
.B(n_2038),
.Y(n_13177)
);

OR2x2_ASAP7_75t_L g13178 ( 
.A(n_12724),
.B(n_2038),
.Y(n_13178)
);

BUFx12f_ASAP7_75t_L g13179 ( 
.A(n_12702),
.Y(n_13179)
);

BUFx4f_ASAP7_75t_L g13180 ( 
.A(n_12702),
.Y(n_13180)
);

INVx1_ASAP7_75t_L g13181 ( 
.A(n_12735),
.Y(n_13181)
);

NAND2xp5_ASAP7_75t_L g13182 ( 
.A(n_12903),
.B(n_2040),
.Y(n_13182)
);

AO21x2_ASAP7_75t_L g13183 ( 
.A1(n_12955),
.A2(n_2041),
.B(n_2042),
.Y(n_13183)
);

INVx1_ASAP7_75t_L g13184 ( 
.A(n_12736),
.Y(n_13184)
);

INVx2_ASAP7_75t_SL g13185 ( 
.A(n_13015),
.Y(n_13185)
);

INVx1_ASAP7_75t_L g13186 ( 
.A(n_12760),
.Y(n_13186)
);

INVx3_ASAP7_75t_L g13187 ( 
.A(n_12841),
.Y(n_13187)
);

INVx2_ASAP7_75t_L g13188 ( 
.A(n_12706),
.Y(n_13188)
);

INVx1_ASAP7_75t_L g13189 ( 
.A(n_12761),
.Y(n_13189)
);

INVx1_ASAP7_75t_L g13190 ( 
.A(n_12772),
.Y(n_13190)
);

INVx6_ASAP7_75t_L g13191 ( 
.A(n_12962),
.Y(n_13191)
);

OAI22xp5_ASAP7_75t_L g13192 ( 
.A1(n_12763),
.A2(n_2044),
.B1(n_2041),
.B2(n_2043),
.Y(n_13192)
);

OAI21x1_ASAP7_75t_L g13193 ( 
.A1(n_12668),
.A2(n_2043),
.B(n_2045),
.Y(n_13193)
);

INVx3_ASAP7_75t_L g13194 ( 
.A(n_12990),
.Y(n_13194)
);

INVx3_ASAP7_75t_L g13195 ( 
.A(n_12997),
.Y(n_13195)
);

OA21x2_ASAP7_75t_L g13196 ( 
.A1(n_12799),
.A2(n_2045),
.B(n_2046),
.Y(n_13196)
);

INVx1_ASAP7_75t_L g13197 ( 
.A(n_12779),
.Y(n_13197)
);

A2O1A1Ixp33_ASAP7_75t_L g13198 ( 
.A1(n_12708),
.A2(n_2048),
.B(n_2046),
.C(n_2047),
.Y(n_13198)
);

OAI21x1_ASAP7_75t_L g13199 ( 
.A1(n_12675),
.A2(n_2048),
.B(n_2049),
.Y(n_13199)
);

NAND2xp5_ASAP7_75t_L g13200 ( 
.A(n_12906),
.B(n_2049),
.Y(n_13200)
);

BUFx2_ASAP7_75t_L g13201 ( 
.A(n_12854),
.Y(n_13201)
);

AND3x1_ASAP7_75t_L g13202 ( 
.A(n_12771),
.B(n_2050),
.C(n_2051),
.Y(n_13202)
);

AOI21xp5_ASAP7_75t_L g13203 ( 
.A1(n_12934),
.A2(n_2050),
.B(n_2051),
.Y(n_13203)
);

OR2x6_ASAP7_75t_L g13204 ( 
.A(n_12916),
.B(n_2052),
.Y(n_13204)
);

AND2x4_ASAP7_75t_SL g13205 ( 
.A(n_12691),
.B(n_2052),
.Y(n_13205)
);

INVx2_ASAP7_75t_SL g13206 ( 
.A(n_12820),
.Y(n_13206)
);

AOI21xp5_ASAP7_75t_L g13207 ( 
.A1(n_12768),
.A2(n_2053),
.B(n_2054),
.Y(n_13207)
);

HB1xp67_ASAP7_75t_L g13208 ( 
.A(n_12663),
.Y(n_13208)
);

CKINVDCx20_ASAP7_75t_R g13209 ( 
.A(n_12904),
.Y(n_13209)
);

AO21x2_ASAP7_75t_L g13210 ( 
.A1(n_12966),
.A2(n_2053),
.B(n_2054),
.Y(n_13210)
);

OAI21x1_ASAP7_75t_L g13211 ( 
.A1(n_12676),
.A2(n_2055),
.B(n_2056),
.Y(n_13211)
);

BUFx2_ASAP7_75t_SL g13212 ( 
.A(n_12837),
.Y(n_13212)
);

INVx2_ASAP7_75t_L g13213 ( 
.A(n_12722),
.Y(n_13213)
);

BUFx3_ASAP7_75t_L g13214 ( 
.A(n_12986),
.Y(n_13214)
);

BUFx6f_ASAP7_75t_L g13215 ( 
.A(n_12931),
.Y(n_13215)
);

OAI21x1_ASAP7_75t_SL g13216 ( 
.A1(n_12795),
.A2(n_2055),
.B(n_2056),
.Y(n_13216)
);

OAI21x1_ASAP7_75t_L g13217 ( 
.A1(n_12797),
.A2(n_2057),
.B(n_2058),
.Y(n_13217)
);

INVx2_ASAP7_75t_L g13218 ( 
.A(n_12687),
.Y(n_13218)
);

OAI21xp5_ASAP7_75t_L g13219 ( 
.A1(n_12812),
.A2(n_2057),
.B(n_2058),
.Y(n_13219)
);

OR2x2_ASAP7_75t_L g13220 ( 
.A(n_12704),
.B(n_2059),
.Y(n_13220)
);

AO21x2_ASAP7_75t_L g13221 ( 
.A1(n_12967),
.A2(n_2059),
.B(n_2060),
.Y(n_13221)
);

INVx2_ASAP7_75t_SL g13222 ( 
.A(n_12886),
.Y(n_13222)
);

NAND2xp5_ASAP7_75t_L g13223 ( 
.A(n_12920),
.B(n_2062),
.Y(n_13223)
);

OAI21xp5_ASAP7_75t_L g13224 ( 
.A1(n_12752),
.A2(n_2063),
.B(n_2064),
.Y(n_13224)
);

INVx1_ASAP7_75t_L g13225 ( 
.A(n_12780),
.Y(n_13225)
);

INVx2_ASAP7_75t_SL g13226 ( 
.A(n_12861),
.Y(n_13226)
);

INVx2_ASAP7_75t_L g13227 ( 
.A(n_12700),
.Y(n_13227)
);

AND2x2_ASAP7_75t_L g13228 ( 
.A(n_12991),
.B(n_2063),
.Y(n_13228)
);

OAI21x1_ASAP7_75t_L g13229 ( 
.A1(n_12800),
.A2(n_2064),
.B(n_2065),
.Y(n_13229)
);

CKINVDCx11_ASAP7_75t_R g13230 ( 
.A(n_12931),
.Y(n_13230)
);

AOI21xp5_ASAP7_75t_L g13231 ( 
.A1(n_12662),
.A2(n_2065),
.B(n_2066),
.Y(n_13231)
);

INVx3_ASAP7_75t_L g13232 ( 
.A(n_12874),
.Y(n_13232)
);

AND2x2_ASAP7_75t_L g13233 ( 
.A(n_12987),
.B(n_2066),
.Y(n_13233)
);

INVx2_ASAP7_75t_L g13234 ( 
.A(n_12796),
.Y(n_13234)
);

INVx2_ASAP7_75t_L g13235 ( 
.A(n_12798),
.Y(n_13235)
);

OAI21xp5_ASAP7_75t_L g13236 ( 
.A1(n_12751),
.A2(n_2067),
.B(n_2068),
.Y(n_13236)
);

AND2x2_ASAP7_75t_L g13237 ( 
.A(n_12996),
.B(n_2067),
.Y(n_13237)
);

OR2x2_ASAP7_75t_L g13238 ( 
.A(n_12721),
.B(n_2068),
.Y(n_13238)
);

NAND2xp5_ASAP7_75t_L g13239 ( 
.A(n_12923),
.B(n_2069),
.Y(n_13239)
);

AOI21xp5_ASAP7_75t_L g13240 ( 
.A1(n_12862),
.A2(n_2069),
.B(n_2070),
.Y(n_13240)
);

AOI21xp5_ASAP7_75t_L g13241 ( 
.A1(n_12665),
.A2(n_2071),
.B(n_2072),
.Y(n_13241)
);

AOI21xp5_ASAP7_75t_L g13242 ( 
.A1(n_12819),
.A2(n_2071),
.B(n_2072),
.Y(n_13242)
);

INVx1_ASAP7_75t_L g13243 ( 
.A(n_12786),
.Y(n_13243)
);

AOI21xp5_ASAP7_75t_L g13244 ( 
.A1(n_12964),
.A2(n_2073),
.B(n_2074),
.Y(n_13244)
);

INVx1_ASAP7_75t_L g13245 ( 
.A(n_12804),
.Y(n_13245)
);

OA21x2_ASAP7_75t_L g13246 ( 
.A1(n_12942),
.A2(n_2075),
.B(n_2076),
.Y(n_13246)
);

INVx2_ASAP7_75t_L g13247 ( 
.A(n_12897),
.Y(n_13247)
);

NAND2xp5_ASAP7_75t_L g13248 ( 
.A(n_12929),
.B(n_2075),
.Y(n_13248)
);

AOI21xp5_ASAP7_75t_L g13249 ( 
.A1(n_12879),
.A2(n_12784),
.B(n_12888),
.Y(n_13249)
);

AOI22xp33_ASAP7_75t_L g13250 ( 
.A1(n_12777),
.A2(n_2078),
.B1(n_2076),
.B2(n_2077),
.Y(n_13250)
);

INVx1_ASAP7_75t_SL g13251 ( 
.A(n_12953),
.Y(n_13251)
);

OAI21x1_ASAP7_75t_L g13252 ( 
.A1(n_12693),
.A2(n_2078),
.B(n_2079),
.Y(n_13252)
);

AOI21xp5_ASAP7_75t_L g13253 ( 
.A1(n_12884),
.A2(n_2081),
.B(n_2082),
.Y(n_13253)
);

AOI22xp5_ASAP7_75t_L g13254 ( 
.A1(n_12785),
.A2(n_2083),
.B1(n_2081),
.B2(n_2082),
.Y(n_13254)
);

NAND2xp5_ASAP7_75t_L g13255 ( 
.A(n_12936),
.B(n_12827),
.Y(n_13255)
);

NAND2x1p5_ASAP7_75t_L g13256 ( 
.A(n_12988),
.B(n_2083),
.Y(n_13256)
);

INVx1_ASAP7_75t_L g13257 ( 
.A(n_12870),
.Y(n_13257)
);

INVx1_ASAP7_75t_L g13258 ( 
.A(n_12850),
.Y(n_13258)
);

OR2x2_ASAP7_75t_L g13259 ( 
.A(n_12880),
.B(n_2084),
.Y(n_13259)
);

OAI21x1_ASAP7_75t_L g13260 ( 
.A1(n_12646),
.A2(n_2084),
.B(n_2086),
.Y(n_13260)
);

INVx2_ASAP7_75t_L g13261 ( 
.A(n_12930),
.Y(n_13261)
);

HB1xp67_ASAP7_75t_L g13262 ( 
.A(n_12846),
.Y(n_13262)
);

AND2x2_ASAP7_75t_L g13263 ( 
.A(n_12927),
.B(n_2086),
.Y(n_13263)
);

INVx1_ASAP7_75t_L g13264 ( 
.A(n_12952),
.Y(n_13264)
);

INVx2_ASAP7_75t_L g13265 ( 
.A(n_12893),
.Y(n_13265)
);

INVx1_ASAP7_75t_L g13266 ( 
.A(n_12935),
.Y(n_13266)
);

INVxp67_ASAP7_75t_L g13267 ( 
.A(n_12871),
.Y(n_13267)
);

NAND2xp5_ASAP7_75t_L g13268 ( 
.A(n_12932),
.B(n_2087),
.Y(n_13268)
);

AND2x4_ASAP7_75t_L g13269 ( 
.A(n_12911),
.B(n_2087),
.Y(n_13269)
);

INVx2_ASAP7_75t_L g13270 ( 
.A(n_12876),
.Y(n_13270)
);

OAI21x1_ASAP7_75t_L g13271 ( 
.A1(n_12716),
.A2(n_2088),
.B(n_2089),
.Y(n_13271)
);

OR2x6_ASAP7_75t_L g13272 ( 
.A(n_12974),
.B(n_2089),
.Y(n_13272)
);

NOR2xp33_ASAP7_75t_L g13273 ( 
.A(n_12789),
.B(n_2090),
.Y(n_13273)
);

INVx2_ASAP7_75t_L g13274 ( 
.A(n_12860),
.Y(n_13274)
);

NAND3xp33_ASAP7_75t_L g13275 ( 
.A(n_12674),
.B(n_2090),
.C(n_2091),
.Y(n_13275)
);

OAI21x1_ASAP7_75t_L g13276 ( 
.A1(n_12683),
.A2(n_2091),
.B(n_2092),
.Y(n_13276)
);

AO21x2_ASAP7_75t_L g13277 ( 
.A1(n_12872),
.A2(n_2092),
.B(n_2093),
.Y(n_13277)
);

NAND2xp5_ASAP7_75t_L g13278 ( 
.A(n_13028),
.B(n_2093),
.Y(n_13278)
);

OAI21x1_ASAP7_75t_L g13279 ( 
.A1(n_12690),
.A2(n_2094),
.B(n_2095),
.Y(n_13279)
);

INVx2_ASAP7_75t_L g13280 ( 
.A(n_12902),
.Y(n_13280)
);

OAI21x1_ASAP7_75t_L g13281 ( 
.A1(n_12725),
.A2(n_12817),
.B(n_12655),
.Y(n_13281)
);

AO31x2_ASAP7_75t_L g13282 ( 
.A1(n_12699),
.A2(n_2098),
.A3(n_2096),
.B(n_2097),
.Y(n_13282)
);

INVx1_ASAP7_75t_L g13283 ( 
.A(n_12825),
.Y(n_13283)
);

AOI21x1_ASAP7_75t_L g13284 ( 
.A1(n_12970),
.A2(n_2097),
.B(n_2098),
.Y(n_13284)
);

OAI21x1_ASAP7_75t_L g13285 ( 
.A1(n_12794),
.A2(n_2099),
.B(n_2100),
.Y(n_13285)
);

AOI22xp33_ASAP7_75t_L g13286 ( 
.A1(n_12766),
.A2(n_2102),
.B1(n_2099),
.B2(n_2101),
.Y(n_13286)
);

HB1xp67_ASAP7_75t_L g13287 ( 
.A(n_13009),
.Y(n_13287)
);

OAI21x1_ASAP7_75t_L g13288 ( 
.A1(n_12714),
.A2(n_2101),
.B(n_2102),
.Y(n_13288)
);

AOI21xp5_ASAP7_75t_L g13289 ( 
.A1(n_13012),
.A2(n_2103),
.B(n_2105),
.Y(n_13289)
);

INVx1_ASAP7_75t_L g13290 ( 
.A(n_12890),
.Y(n_13290)
);

OAI21x1_ASAP7_75t_L g13291 ( 
.A1(n_12961),
.A2(n_2105),
.B(n_2106),
.Y(n_13291)
);

AO31x2_ASAP7_75t_L g13292 ( 
.A1(n_13026),
.A2(n_2108),
.A3(n_2106),
.B(n_2107),
.Y(n_13292)
);

AND2x2_ASAP7_75t_L g13293 ( 
.A(n_12999),
.B(n_2107),
.Y(n_13293)
);

BUFx6f_ASAP7_75t_L g13294 ( 
.A(n_13003),
.Y(n_13294)
);

AO21x2_ASAP7_75t_L g13295 ( 
.A1(n_12957),
.A2(n_2108),
.B(n_2110),
.Y(n_13295)
);

A2O1A1Ixp33_ASAP7_75t_L g13296 ( 
.A1(n_12978),
.A2(n_12848),
.B(n_12925),
.C(n_13030),
.Y(n_13296)
);

OAI21x1_ASAP7_75t_L g13297 ( 
.A1(n_12983),
.A2(n_2110),
.B(n_2111),
.Y(n_13297)
);

AND2x2_ASAP7_75t_L g13298 ( 
.A(n_13018),
.B(n_2111),
.Y(n_13298)
);

CKINVDCx14_ASAP7_75t_R g13299 ( 
.A(n_12859),
.Y(n_13299)
);

NAND2xp5_ASAP7_75t_L g13300 ( 
.A(n_12853),
.B(n_2112),
.Y(n_13300)
);

CKINVDCx11_ASAP7_75t_R g13301 ( 
.A(n_13003),
.Y(n_13301)
);

AO21x2_ASAP7_75t_L g13302 ( 
.A1(n_12867),
.A2(n_2112),
.B(n_2113),
.Y(n_13302)
);

NAND2xp5_ASAP7_75t_L g13303 ( 
.A(n_12847),
.B(n_2113),
.Y(n_13303)
);

A2O1A1Ixp33_ASAP7_75t_L g13304 ( 
.A1(n_12922),
.A2(n_2116),
.B(n_2114),
.C(n_2115),
.Y(n_13304)
);

OAI21xp5_ASAP7_75t_L g13305 ( 
.A1(n_12755),
.A2(n_2116),
.B(n_2117),
.Y(n_13305)
);

INVx1_ASAP7_75t_L g13306 ( 
.A(n_12958),
.Y(n_13306)
);

AOI22xp5_ASAP7_75t_L g13307 ( 
.A1(n_12762),
.A2(n_2120),
.B1(n_2118),
.B2(n_2119),
.Y(n_13307)
);

NAND2xp5_ASAP7_75t_L g13308 ( 
.A(n_12844),
.B(n_2118),
.Y(n_13308)
);

INVx1_ASAP7_75t_SL g13309 ( 
.A(n_12951),
.Y(n_13309)
);

AOI21x1_ASAP7_75t_L g13310 ( 
.A1(n_12998),
.A2(n_2119),
.B(n_2120),
.Y(n_13310)
);

INVx1_ASAP7_75t_L g13311 ( 
.A(n_12960),
.Y(n_13311)
);

AND2x2_ASAP7_75t_L g13312 ( 
.A(n_13005),
.B(n_2121),
.Y(n_13312)
);

AO21x2_ASAP7_75t_L g13313 ( 
.A1(n_12885),
.A2(n_2121),
.B(n_2122),
.Y(n_13313)
);

BUFx2_ASAP7_75t_L g13314 ( 
.A(n_12705),
.Y(n_13314)
);

NAND2xp5_ASAP7_75t_L g13315 ( 
.A(n_12965),
.B(n_12917),
.Y(n_13315)
);

INVx2_ASAP7_75t_SL g13316 ( 
.A(n_12803),
.Y(n_13316)
);

AND2x2_ASAP7_75t_L g13317 ( 
.A(n_13010),
.B(n_2122),
.Y(n_13317)
);

AOI22x1_ASAP7_75t_L g13318 ( 
.A1(n_12776),
.A2(n_2125),
.B1(n_2123),
.B2(n_2124),
.Y(n_13318)
);

INVx1_ASAP7_75t_L g13319 ( 
.A(n_12738),
.Y(n_13319)
);

AO21x2_ASAP7_75t_L g13320 ( 
.A1(n_12948),
.A2(n_2123),
.B(n_2124),
.Y(n_13320)
);

INVx1_ASAP7_75t_L g13321 ( 
.A(n_12945),
.Y(n_13321)
);

OAI21x1_ASAP7_75t_L g13322 ( 
.A1(n_12831),
.A2(n_12975),
.B(n_13027),
.Y(n_13322)
);

NAND2xp5_ASAP7_75t_L g13323 ( 
.A(n_12994),
.B(n_2125),
.Y(n_13323)
);

HB1xp67_ASAP7_75t_L g13324 ( 
.A(n_13008),
.Y(n_13324)
);

OA21x2_ASAP7_75t_L g13325 ( 
.A1(n_13019),
.A2(n_2126),
.B(n_2127),
.Y(n_13325)
);

AO21x2_ASAP7_75t_L g13326 ( 
.A1(n_12969),
.A2(n_2126),
.B(n_2128),
.Y(n_13326)
);

AND2x2_ASAP7_75t_L g13327 ( 
.A(n_13000),
.B(n_2129),
.Y(n_13327)
);

OR2x2_ASAP7_75t_L g13328 ( 
.A(n_13024),
.B(n_2129),
.Y(n_13328)
);

AND2x2_ASAP7_75t_L g13329 ( 
.A(n_12836),
.B(n_2130),
.Y(n_13329)
);

NAND2xp5_ASAP7_75t_SL g13330 ( 
.A(n_12750),
.B(n_2130),
.Y(n_13330)
);

INVx2_ASAP7_75t_L g13331 ( 
.A(n_13017),
.Y(n_13331)
);

AO31x2_ASAP7_75t_L g13332 ( 
.A1(n_12943),
.A2(n_2133),
.A3(n_2131),
.B(n_2132),
.Y(n_13332)
);

OAI22xp33_ASAP7_75t_L g13333 ( 
.A1(n_12730),
.A2(n_2133),
.B1(n_2131),
.B2(n_2132),
.Y(n_13333)
);

AO31x2_ASAP7_75t_L g13334 ( 
.A1(n_12971),
.A2(n_2136),
.A3(n_2134),
.B(n_2135),
.Y(n_13334)
);

INVx1_ASAP7_75t_L g13335 ( 
.A(n_12654),
.Y(n_13335)
);

BUFx3_ASAP7_75t_L g13336 ( 
.A(n_12985),
.Y(n_13336)
);

CKINVDCx20_ASAP7_75t_R g13337 ( 
.A(n_12835),
.Y(n_13337)
);

NAND2xp5_ASAP7_75t_L g13338 ( 
.A(n_12980),
.B(n_2134),
.Y(n_13338)
);

AOI21xp5_ASAP7_75t_L g13339 ( 
.A1(n_12842),
.A2(n_2135),
.B(n_2136),
.Y(n_13339)
);

AOI21xp5_ASAP7_75t_L g13340 ( 
.A1(n_12995),
.A2(n_2137),
.B(n_2138),
.Y(n_13340)
);

NAND2x1p5_ASAP7_75t_L g13341 ( 
.A(n_12992),
.B(n_2138),
.Y(n_13341)
);

AOI21xp5_ASAP7_75t_L g13342 ( 
.A1(n_13004),
.A2(n_2139),
.B(n_2140),
.Y(n_13342)
);

AOI21xp5_ASAP7_75t_L g13343 ( 
.A1(n_12840),
.A2(n_2139),
.B(n_2140),
.Y(n_13343)
);

AND2x2_ASAP7_75t_L g13344 ( 
.A(n_12910),
.B(n_2141),
.Y(n_13344)
);

NAND2xp5_ASAP7_75t_L g13345 ( 
.A(n_12989),
.B(n_2141),
.Y(n_13345)
);

AOI21xp5_ASAP7_75t_L g13346 ( 
.A1(n_12829),
.A2(n_2142),
.B(n_2143),
.Y(n_13346)
);

AO21x2_ASAP7_75t_L g13347 ( 
.A1(n_13007),
.A2(n_2143),
.B(n_2144),
.Y(n_13347)
);

AOI22xp5_ASAP7_75t_L g13348 ( 
.A1(n_12939),
.A2(n_2147),
.B1(n_2145),
.B2(n_2146),
.Y(n_13348)
);

OA21x2_ASAP7_75t_L g13349 ( 
.A1(n_13023),
.A2(n_2145),
.B(n_2146),
.Y(n_13349)
);

INVx2_ASAP7_75t_L g13350 ( 
.A(n_12921),
.Y(n_13350)
);

NAND2x1p5_ASAP7_75t_L g13351 ( 
.A(n_12855),
.B(n_2147),
.Y(n_13351)
);

INVx2_ASAP7_75t_SL g13352 ( 
.A(n_13001),
.Y(n_13352)
);

HB1xp67_ASAP7_75t_L g13353 ( 
.A(n_12950),
.Y(n_13353)
);

INVx1_ASAP7_75t_L g13354 ( 
.A(n_12834),
.Y(n_13354)
);

INVx1_ASAP7_75t_L g13355 ( 
.A(n_12838),
.Y(n_13355)
);

INVx1_ASAP7_75t_L g13356 ( 
.A(n_12950),
.Y(n_13356)
);

AND2x2_ASAP7_75t_L g13357 ( 
.A(n_12792),
.B(n_2148),
.Y(n_13357)
);

AOI21xp5_ASAP7_75t_L g13358 ( 
.A1(n_13029),
.A2(n_2148),
.B(n_2149),
.Y(n_13358)
);

CKINVDCx20_ASAP7_75t_R g13359 ( 
.A(n_12889),
.Y(n_13359)
);

OAI21x1_ASAP7_75t_L g13360 ( 
.A1(n_12881),
.A2(n_2149),
.B(n_2150),
.Y(n_13360)
);

NOR2xp33_ASAP7_75t_L g13361 ( 
.A(n_12993),
.B(n_2150),
.Y(n_13361)
);

INVx2_ASAP7_75t_L g13362 ( 
.A(n_12887),
.Y(n_13362)
);

INVx1_ASAP7_75t_L g13363 ( 
.A(n_12938),
.Y(n_13363)
);

OA21x2_ASAP7_75t_L g13364 ( 
.A1(n_12891),
.A2(n_2151),
.B(n_2152),
.Y(n_13364)
);

AND2x4_ASAP7_75t_L g13365 ( 
.A(n_12973),
.B(n_2151),
.Y(n_13365)
);

AO31x2_ASAP7_75t_L g13366 ( 
.A1(n_12926),
.A2(n_2154),
.A3(n_2152),
.B(n_2153),
.Y(n_13366)
);

AOI21xp5_ASAP7_75t_L g13367 ( 
.A1(n_12833),
.A2(n_2154),
.B(n_2155),
.Y(n_13367)
);

INVx1_ASAP7_75t_L g13368 ( 
.A(n_12894),
.Y(n_13368)
);

INVx2_ASAP7_75t_L g13369 ( 
.A(n_12905),
.Y(n_13369)
);

INVx1_ASAP7_75t_L g13370 ( 
.A(n_12915),
.Y(n_13370)
);

AOI21x1_ASAP7_75t_L g13371 ( 
.A1(n_13006),
.A2(n_2156),
.B(n_2157),
.Y(n_13371)
);

BUFx6f_ASAP7_75t_SL g13372 ( 
.A(n_12944),
.Y(n_13372)
);

AND2x4_ASAP7_75t_L g13373 ( 
.A(n_12851),
.B(n_2156),
.Y(n_13373)
);

OR2x2_ASAP7_75t_L g13374 ( 
.A(n_12710),
.B(n_2157),
.Y(n_13374)
);

INVx2_ASAP7_75t_L g13375 ( 
.A(n_12852),
.Y(n_13375)
);

INVx1_ASAP7_75t_L g13376 ( 
.A(n_12912),
.Y(n_13376)
);

OR2x2_ASAP7_75t_L g13377 ( 
.A(n_12710),
.B(n_2158),
.Y(n_13377)
);

NAND2xp5_ASAP7_75t_L g13378 ( 
.A(n_12963),
.B(n_2158),
.Y(n_13378)
);

AND2x4_ASAP7_75t_L g13379 ( 
.A(n_12908),
.B(n_2160),
.Y(n_13379)
);

NAND2x1p5_ASAP7_75t_L g13380 ( 
.A(n_12982),
.B(n_2160),
.Y(n_13380)
);

OAI21x1_ASAP7_75t_L g13381 ( 
.A1(n_12913),
.A2(n_2161),
.B(n_2162),
.Y(n_13381)
);

NAND2xp5_ASAP7_75t_L g13382 ( 
.A(n_12933),
.B(n_2161),
.Y(n_13382)
);

INVx1_ASAP7_75t_L g13383 ( 
.A(n_12928),
.Y(n_13383)
);

CKINVDCx5p33_ASAP7_75t_R g13384 ( 
.A(n_12949),
.Y(n_13384)
);

A2O1A1Ixp33_ASAP7_75t_L g13385 ( 
.A1(n_12791),
.A2(n_2165),
.B(n_2162),
.C(n_2163),
.Y(n_13385)
);

INVx5_ASAP7_75t_L g13386 ( 
.A(n_12984),
.Y(n_13386)
);

OA21x2_ASAP7_75t_L g13387 ( 
.A1(n_12941),
.A2(n_12954),
.B(n_12947),
.Y(n_13387)
);

INVx2_ASAP7_75t_L g13388 ( 
.A(n_12875),
.Y(n_13388)
);

OR2x2_ASAP7_75t_L g13389 ( 
.A(n_12899),
.B(n_2163),
.Y(n_13389)
);

INVx1_ASAP7_75t_L g13390 ( 
.A(n_12909),
.Y(n_13390)
);

OAI21x1_ASAP7_75t_L g13391 ( 
.A1(n_13046),
.A2(n_12845),
.B(n_2165),
.Y(n_13391)
);

OR2x6_ASAP7_75t_L g13392 ( 
.A(n_13037),
.B(n_2166),
.Y(n_13392)
);

NOR2xp33_ASAP7_75t_L g13393 ( 
.A(n_13146),
.B(n_2167),
.Y(n_13393)
);

OR2x2_ASAP7_75t_L g13394 ( 
.A(n_13083),
.B(n_2167),
.Y(n_13394)
);

INVx2_ASAP7_75t_L g13395 ( 
.A(n_13201),
.Y(n_13395)
);

INVx1_ASAP7_75t_L g13396 ( 
.A(n_13036),
.Y(n_13396)
);

INVx1_ASAP7_75t_L g13397 ( 
.A(n_13040),
.Y(n_13397)
);

INVx2_ASAP7_75t_L g13398 ( 
.A(n_13314),
.Y(n_13398)
);

HB1xp67_ASAP7_75t_L g13399 ( 
.A(n_13169),
.Y(n_13399)
);

INVx5_ASAP7_75t_L g13400 ( 
.A(n_13204),
.Y(n_13400)
);

INVx2_ASAP7_75t_L g13401 ( 
.A(n_13232),
.Y(n_13401)
);

INVx2_ASAP7_75t_SL g13402 ( 
.A(n_13069),
.Y(n_13402)
);

INVx1_ASAP7_75t_L g13403 ( 
.A(n_13043),
.Y(n_13403)
);

INVx1_ASAP7_75t_L g13404 ( 
.A(n_13067),
.Y(n_13404)
);

INVx2_ASAP7_75t_L g13405 ( 
.A(n_13206),
.Y(n_13405)
);

AO31x2_ASAP7_75t_L g13406 ( 
.A1(n_13335),
.A2(n_2170),
.A3(n_2168),
.B(n_2169),
.Y(n_13406)
);

HB1xp67_ASAP7_75t_L g13407 ( 
.A(n_13055),
.Y(n_13407)
);

BUFx6f_ASAP7_75t_L g13408 ( 
.A(n_13179),
.Y(n_13408)
);

INVx1_ASAP7_75t_L g13409 ( 
.A(n_13080),
.Y(n_13409)
);

INVx2_ASAP7_75t_SL g13410 ( 
.A(n_13180),
.Y(n_13410)
);

INVx2_ASAP7_75t_L g13411 ( 
.A(n_13031),
.Y(n_13411)
);

HB1xp67_ASAP7_75t_L g13412 ( 
.A(n_13071),
.Y(n_13412)
);

INVx1_ASAP7_75t_L g13413 ( 
.A(n_13093),
.Y(n_13413)
);

NAND2xp5_ASAP7_75t_L g13414 ( 
.A(n_13324),
.B(n_2168),
.Y(n_13414)
);

INVx3_ASAP7_75t_L g13415 ( 
.A(n_13191),
.Y(n_13415)
);

OA21x2_ASAP7_75t_L g13416 ( 
.A1(n_13032),
.A2(n_2169),
.B(n_2170),
.Y(n_13416)
);

HB1xp67_ASAP7_75t_L g13417 ( 
.A(n_13387),
.Y(n_13417)
);

INVx2_ASAP7_75t_L g13418 ( 
.A(n_13226),
.Y(n_13418)
);

INVx3_ASAP7_75t_L g13419 ( 
.A(n_13037),
.Y(n_13419)
);

INVx2_ASAP7_75t_L g13420 ( 
.A(n_13054),
.Y(n_13420)
);

INVx1_ASAP7_75t_L g13421 ( 
.A(n_13094),
.Y(n_13421)
);

INVx2_ASAP7_75t_L g13422 ( 
.A(n_13194),
.Y(n_13422)
);

INVx1_ASAP7_75t_L g13423 ( 
.A(n_13098),
.Y(n_13423)
);

INVx1_ASAP7_75t_SL g13424 ( 
.A(n_13230),
.Y(n_13424)
);

NAND2xp5_ASAP7_75t_L g13425 ( 
.A(n_13331),
.B(n_2171),
.Y(n_13425)
);

OA21x2_ASAP7_75t_L g13426 ( 
.A1(n_13091),
.A2(n_2172),
.B(n_2173),
.Y(n_13426)
);

INVx2_ASAP7_75t_L g13427 ( 
.A(n_13195),
.Y(n_13427)
);

INVx1_ASAP7_75t_L g13428 ( 
.A(n_13105),
.Y(n_13428)
);

BUFx6f_ASAP7_75t_L g13429 ( 
.A(n_13301),
.Y(n_13429)
);

AND2x2_ASAP7_75t_L g13430 ( 
.A(n_13212),
.B(n_2172),
.Y(n_13430)
);

INVx1_ASAP7_75t_L g13431 ( 
.A(n_13122),
.Y(n_13431)
);

INVx2_ASAP7_75t_L g13432 ( 
.A(n_13048),
.Y(n_13432)
);

INVx2_ASAP7_75t_SL g13433 ( 
.A(n_13063),
.Y(n_13433)
);

INVx2_ASAP7_75t_L g13434 ( 
.A(n_13045),
.Y(n_13434)
);

INVx2_ASAP7_75t_L g13435 ( 
.A(n_13049),
.Y(n_13435)
);

INVx2_ASAP7_75t_L g13436 ( 
.A(n_13316),
.Y(n_13436)
);

BUFx3_ASAP7_75t_L g13437 ( 
.A(n_13100),
.Y(n_13437)
);

AND2x2_ASAP7_75t_L g13438 ( 
.A(n_13145),
.B(n_2173),
.Y(n_13438)
);

INVx1_ASAP7_75t_L g13439 ( 
.A(n_13132),
.Y(n_13439)
);

OR2x6_ASAP7_75t_L g13440 ( 
.A(n_13207),
.B(n_2174),
.Y(n_13440)
);

INVx3_ASAP7_75t_L g13441 ( 
.A(n_13214),
.Y(n_13441)
);

OAI21x1_ASAP7_75t_L g13442 ( 
.A1(n_13097),
.A2(n_2174),
.B(n_2175),
.Y(n_13442)
);

AND2x2_ASAP7_75t_L g13443 ( 
.A(n_13103),
.B(n_2175),
.Y(n_13443)
);

NAND2xp5_ASAP7_75t_L g13444 ( 
.A(n_13267),
.B(n_2176),
.Y(n_13444)
);

INVx1_ASAP7_75t_L g13445 ( 
.A(n_13148),
.Y(n_13445)
);

BUFx3_ASAP7_75t_L g13446 ( 
.A(n_13086),
.Y(n_13446)
);

INVx3_ASAP7_75t_L g13447 ( 
.A(n_13187),
.Y(n_13447)
);

AND2x2_ASAP7_75t_L g13448 ( 
.A(n_13042),
.B(n_2176),
.Y(n_13448)
);

OAI21xp33_ASAP7_75t_SL g13449 ( 
.A1(n_13041),
.A2(n_2177),
.B(n_2178),
.Y(n_13449)
);

INVx1_ASAP7_75t_L g13450 ( 
.A(n_13159),
.Y(n_13450)
);

INVx3_ASAP7_75t_L g13451 ( 
.A(n_13336),
.Y(n_13451)
);

INVx2_ASAP7_75t_L g13452 ( 
.A(n_13075),
.Y(n_13452)
);

INVx1_ASAP7_75t_SL g13453 ( 
.A(n_13209),
.Y(n_13453)
);

INVx2_ASAP7_75t_L g13454 ( 
.A(n_13073),
.Y(n_13454)
);

OR2x6_ASAP7_75t_L g13455 ( 
.A(n_13038),
.B(n_2177),
.Y(n_13455)
);

INVx1_ASAP7_75t_L g13456 ( 
.A(n_13162),
.Y(n_13456)
);

INVx1_ASAP7_75t_L g13457 ( 
.A(n_13175),
.Y(n_13457)
);

INVx2_ASAP7_75t_L g13458 ( 
.A(n_13126),
.Y(n_13458)
);

INVx2_ASAP7_75t_L g13459 ( 
.A(n_13215),
.Y(n_13459)
);

AND2x2_ASAP7_75t_L g13460 ( 
.A(n_13172),
.B(n_2178),
.Y(n_13460)
);

INVx1_ASAP7_75t_L g13461 ( 
.A(n_13181),
.Y(n_13461)
);

BUFx6f_ASAP7_75t_L g13462 ( 
.A(n_13113),
.Y(n_13462)
);

INVx2_ASAP7_75t_L g13463 ( 
.A(n_13215),
.Y(n_13463)
);

INVx3_ASAP7_75t_L g13464 ( 
.A(n_13294),
.Y(n_13464)
);

INVx2_ASAP7_75t_L g13465 ( 
.A(n_13294),
.Y(n_13465)
);

INVx1_ASAP7_75t_L g13466 ( 
.A(n_13184),
.Y(n_13466)
);

INVx3_ASAP7_75t_L g13467 ( 
.A(n_13115),
.Y(n_13467)
);

INVx1_ASAP7_75t_L g13468 ( 
.A(n_13186),
.Y(n_13468)
);

NAND2xp5_ASAP7_75t_L g13469 ( 
.A(n_13051),
.B(n_2179),
.Y(n_13469)
);

OR2x2_ASAP7_75t_L g13470 ( 
.A(n_13315),
.B(n_2179),
.Y(n_13470)
);

OA21x2_ASAP7_75t_L g13471 ( 
.A1(n_13089),
.A2(n_2180),
.B(n_2181),
.Y(n_13471)
);

HB1xp67_ASAP7_75t_L g13472 ( 
.A(n_13060),
.Y(n_13472)
);

AND2x4_ASAP7_75t_L g13473 ( 
.A(n_13222),
.B(n_2180),
.Y(n_13473)
);

AND2x2_ASAP7_75t_L g13474 ( 
.A(n_13143),
.B(n_2181),
.Y(n_13474)
);

NOR2x1_ASAP7_75t_R g13475 ( 
.A(n_13095),
.B(n_2182),
.Y(n_13475)
);

AOI222xp33_ASAP7_75t_L g13476 ( 
.A1(n_13275),
.A2(n_2185),
.B1(n_2187),
.B2(n_2182),
.C1(n_2183),
.C2(n_2186),
.Y(n_13476)
);

INVx5_ASAP7_75t_L g13477 ( 
.A(n_13204),
.Y(n_13477)
);

OAI22xp33_ASAP7_75t_L g13478 ( 
.A1(n_13374),
.A2(n_2188),
.B1(n_2185),
.B2(n_2186),
.Y(n_13478)
);

AND2x4_ASAP7_75t_L g13479 ( 
.A(n_13251),
.B(n_2189),
.Y(n_13479)
);

INVx1_ASAP7_75t_L g13480 ( 
.A(n_13189),
.Y(n_13480)
);

INVx1_ASAP7_75t_L g13481 ( 
.A(n_13190),
.Y(n_13481)
);

INVx2_ASAP7_75t_L g13482 ( 
.A(n_13065),
.Y(n_13482)
);

OAI21xp5_ASAP7_75t_L g13483 ( 
.A1(n_13156),
.A2(n_2189),
.B(n_2190),
.Y(n_13483)
);

AND2x2_ASAP7_75t_L g13484 ( 
.A(n_13290),
.B(n_2190),
.Y(n_13484)
);

AND2x2_ASAP7_75t_L g13485 ( 
.A(n_13090),
.B(n_2192),
.Y(n_13485)
);

OA21x2_ASAP7_75t_L g13486 ( 
.A1(n_13085),
.A2(n_2193),
.B(n_2194),
.Y(n_13486)
);

INVx1_ASAP7_75t_L g13487 ( 
.A(n_13197),
.Y(n_13487)
);

HB1xp67_ASAP7_75t_L g13488 ( 
.A(n_13196),
.Y(n_13488)
);

INVx1_ASAP7_75t_L g13489 ( 
.A(n_13225),
.Y(n_13489)
);

INVx2_ASAP7_75t_L g13490 ( 
.A(n_13118),
.Y(n_13490)
);

INVx2_ASAP7_75t_L g13491 ( 
.A(n_13044),
.Y(n_13491)
);

INVx1_ASAP7_75t_L g13492 ( 
.A(n_13243),
.Y(n_13492)
);

INVx3_ASAP7_75t_L g13493 ( 
.A(n_13185),
.Y(n_13493)
);

INVx2_ASAP7_75t_L g13494 ( 
.A(n_13256),
.Y(n_13494)
);

INVx1_ASAP7_75t_L g13495 ( 
.A(n_13264),
.Y(n_13495)
);

HB1xp67_ASAP7_75t_L g13496 ( 
.A(n_13353),
.Y(n_13496)
);

INVx2_ASAP7_75t_L g13497 ( 
.A(n_13101),
.Y(n_13497)
);

INVx1_ASAP7_75t_L g13498 ( 
.A(n_13245),
.Y(n_13498)
);

INVx1_ASAP7_75t_L g13499 ( 
.A(n_13120),
.Y(n_13499)
);

HB1xp67_ASAP7_75t_L g13500 ( 
.A(n_13087),
.Y(n_13500)
);

AND2x2_ASAP7_75t_L g13501 ( 
.A(n_13280),
.B(n_2193),
.Y(n_13501)
);

INVx2_ASAP7_75t_L g13502 ( 
.A(n_13119),
.Y(n_13502)
);

INVx1_ASAP7_75t_SL g13503 ( 
.A(n_13096),
.Y(n_13503)
);

INVx1_ASAP7_75t_L g13504 ( 
.A(n_13074),
.Y(n_13504)
);

NOR2xp67_ASAP7_75t_L g13505 ( 
.A(n_13033),
.B(n_2195),
.Y(n_13505)
);

INVx2_ASAP7_75t_SL g13506 ( 
.A(n_13352),
.Y(n_13506)
);

INVx2_ASAP7_75t_L g13507 ( 
.A(n_13070),
.Y(n_13507)
);

AOI22xp33_ASAP7_75t_SL g13508 ( 
.A1(n_13056),
.A2(n_2197),
.B1(n_2195),
.B2(n_2196),
.Y(n_13508)
);

AND2x2_ASAP7_75t_L g13509 ( 
.A(n_13265),
.B(n_2196),
.Y(n_13509)
);

INVx2_ASAP7_75t_L g13510 ( 
.A(n_13285),
.Y(n_13510)
);

INVx1_ASAP7_75t_L g13511 ( 
.A(n_13257),
.Y(n_13511)
);

INVx1_ASAP7_75t_L g13512 ( 
.A(n_13234),
.Y(n_13512)
);

INVx1_ASAP7_75t_L g13513 ( 
.A(n_13235),
.Y(n_13513)
);

OR2x2_ASAP7_75t_L g13514 ( 
.A(n_13274),
.B(n_13270),
.Y(n_13514)
);

OR2x6_ASAP7_75t_L g13515 ( 
.A(n_13241),
.B(n_2197),
.Y(n_13515)
);

INVx1_ASAP7_75t_L g13516 ( 
.A(n_13084),
.Y(n_13516)
);

NAND3xp33_ASAP7_75t_L g13517 ( 
.A(n_13152),
.B(n_2198),
.C(n_2199),
.Y(n_13517)
);

OAI22xp5_ASAP7_75t_L g13518 ( 
.A1(n_13299),
.A2(n_2200),
.B1(n_2198),
.B2(n_2199),
.Y(n_13518)
);

NOR2xp67_ASAP7_75t_L g13519 ( 
.A(n_13386),
.B(n_2200),
.Y(n_13519)
);

OR2x6_ASAP7_75t_L g13520 ( 
.A(n_13129),
.B(n_2201),
.Y(n_13520)
);

INVxp67_ASAP7_75t_L g13521 ( 
.A(n_13078),
.Y(n_13521)
);

INVx1_ASAP7_75t_L g13522 ( 
.A(n_13227),
.Y(n_13522)
);

INVx2_ASAP7_75t_SL g13523 ( 
.A(n_13077),
.Y(n_13523)
);

OR2x6_ASAP7_75t_L g13524 ( 
.A(n_13157),
.B(n_2201),
.Y(n_13524)
);

BUFx4f_ASAP7_75t_SL g13525 ( 
.A(n_13135),
.Y(n_13525)
);

INVx1_ASAP7_75t_L g13526 ( 
.A(n_13218),
.Y(n_13526)
);

INVx1_ASAP7_75t_L g13527 ( 
.A(n_13188),
.Y(n_13527)
);

INVx2_ASAP7_75t_L g13528 ( 
.A(n_13261),
.Y(n_13528)
);

OAI21x1_ASAP7_75t_L g13529 ( 
.A1(n_13281),
.A2(n_2202),
.B(n_2203),
.Y(n_13529)
);

AND2x4_ASAP7_75t_L g13530 ( 
.A(n_13039),
.B(n_2202),
.Y(n_13530)
);

INVx1_ASAP7_75t_L g13531 ( 
.A(n_13213),
.Y(n_13531)
);

INVx1_ASAP7_75t_L g13532 ( 
.A(n_13377),
.Y(n_13532)
);

AOI21x1_ASAP7_75t_L g13533 ( 
.A1(n_13066),
.A2(n_2203),
.B(n_2204),
.Y(n_13533)
);

INVx1_ASAP7_75t_L g13534 ( 
.A(n_13058),
.Y(n_13534)
);

AND2x4_ASAP7_75t_L g13535 ( 
.A(n_13035),
.B(n_2204),
.Y(n_13535)
);

AND2x2_ASAP7_75t_L g13536 ( 
.A(n_13309),
.B(n_2205),
.Y(n_13536)
);

BUFx2_ASAP7_75t_L g13537 ( 
.A(n_13124),
.Y(n_13537)
);

INVx3_ASAP7_75t_L g13538 ( 
.A(n_13269),
.Y(n_13538)
);

AO21x1_ASAP7_75t_SL g13539 ( 
.A1(n_13034),
.A2(n_2205),
.B(n_2206),
.Y(n_13539)
);

INVx2_ASAP7_75t_L g13540 ( 
.A(n_13288),
.Y(n_13540)
);

INVxp67_ASAP7_75t_SL g13541 ( 
.A(n_13102),
.Y(n_13541)
);

INVx1_ASAP7_75t_L g13542 ( 
.A(n_13058),
.Y(n_13542)
);

INVx2_ASAP7_75t_L g13543 ( 
.A(n_13322),
.Y(n_13543)
);

HB1xp67_ASAP7_75t_L g13544 ( 
.A(n_13165),
.Y(n_13544)
);

AOI21xp5_ASAP7_75t_L g13545 ( 
.A1(n_13249),
.A2(n_2206),
.B(n_2207),
.Y(n_13545)
);

OA21x2_ASAP7_75t_L g13546 ( 
.A1(n_13319),
.A2(n_2207),
.B(n_2208),
.Y(n_13546)
);

AOI22xp33_ASAP7_75t_L g13547 ( 
.A1(n_13130),
.A2(n_2211),
.B1(n_2209),
.B2(n_2210),
.Y(n_13547)
);

INVx1_ASAP7_75t_L g13548 ( 
.A(n_13110),
.Y(n_13548)
);

OAI21x1_ASAP7_75t_L g13549 ( 
.A1(n_13255),
.A2(n_2209),
.B(n_2210),
.Y(n_13549)
);

INVx1_ASAP7_75t_L g13550 ( 
.A(n_13110),
.Y(n_13550)
);

AO21x2_ASAP7_75t_L g13551 ( 
.A1(n_13258),
.A2(n_2211),
.B(n_2212),
.Y(n_13551)
);

OAI22xp5_ASAP7_75t_L g13552 ( 
.A1(n_13202),
.A2(n_13384),
.B1(n_13296),
.B2(n_13231),
.Y(n_13552)
);

INVx2_ASAP7_75t_L g13553 ( 
.A(n_13229),
.Y(n_13553)
);

INVx2_ASAP7_75t_L g13554 ( 
.A(n_13217),
.Y(n_13554)
);

OAI22xp5_ASAP7_75t_L g13555 ( 
.A1(n_13137),
.A2(n_2214),
.B1(n_2212),
.B2(n_2213),
.Y(n_13555)
);

INVx1_ASAP7_75t_L g13556 ( 
.A(n_13178),
.Y(n_13556)
);

INVx1_ASAP7_75t_L g13557 ( 
.A(n_13306),
.Y(n_13557)
);

INVx4_ASAP7_75t_L g13558 ( 
.A(n_13164),
.Y(n_13558)
);

NAND2xp5_ASAP7_75t_L g13559 ( 
.A(n_13356),
.B(n_2213),
.Y(n_13559)
);

INVx1_ASAP7_75t_L g13560 ( 
.A(n_13311),
.Y(n_13560)
);

OA21x2_ASAP7_75t_L g13561 ( 
.A1(n_13283),
.A2(n_2215),
.B(n_2216),
.Y(n_13561)
);

OR2x2_ASAP7_75t_L g13562 ( 
.A(n_13109),
.B(n_13125),
.Y(n_13562)
);

INVx2_ASAP7_75t_L g13563 ( 
.A(n_13052),
.Y(n_13563)
);

AO21x2_ASAP7_75t_L g13564 ( 
.A1(n_13321),
.A2(n_2217),
.B(n_2218),
.Y(n_13564)
);

AND2x2_ASAP7_75t_L g13565 ( 
.A(n_13082),
.B(n_2217),
.Y(n_13565)
);

AND2x2_ASAP7_75t_L g13566 ( 
.A(n_13312),
.B(n_2218),
.Y(n_13566)
);

CKINVDCx20_ASAP7_75t_R g13567 ( 
.A(n_13171),
.Y(n_13567)
);

INVx2_ASAP7_75t_L g13568 ( 
.A(n_13276),
.Y(n_13568)
);

BUFx6f_ASAP7_75t_L g13569 ( 
.A(n_13293),
.Y(n_13569)
);

INVx1_ASAP7_75t_L g13570 ( 
.A(n_13053),
.Y(n_13570)
);

INVx1_ASAP7_75t_L g13571 ( 
.A(n_13053),
.Y(n_13571)
);

INVx2_ASAP7_75t_L g13572 ( 
.A(n_13247),
.Y(n_13572)
);

BUFx4f_ASAP7_75t_SL g13573 ( 
.A(n_13337),
.Y(n_13573)
);

INVx2_ASAP7_75t_L g13574 ( 
.A(n_13271),
.Y(n_13574)
);

INVx1_ASAP7_75t_L g13575 ( 
.A(n_13050),
.Y(n_13575)
);

INVx1_ASAP7_75t_L g13576 ( 
.A(n_13072),
.Y(n_13576)
);

INVx2_ASAP7_75t_SL g13577 ( 
.A(n_13068),
.Y(n_13577)
);

INVx3_ASAP7_75t_L g13578 ( 
.A(n_13127),
.Y(n_13578)
);

INVx1_ASAP7_75t_L g13579 ( 
.A(n_13176),
.Y(n_13579)
);

HB1xp67_ASAP7_75t_L g13580 ( 
.A(n_13092),
.Y(n_13580)
);

INVx1_ASAP7_75t_L g13581 ( 
.A(n_13123),
.Y(n_13581)
);

INVx2_ASAP7_75t_L g13582 ( 
.A(n_13112),
.Y(n_13582)
);

INVx1_ASAP7_75t_L g13583 ( 
.A(n_13131),
.Y(n_13583)
);

NAND2xp5_ASAP7_75t_L g13584 ( 
.A(n_13354),
.B(n_2219),
.Y(n_13584)
);

INVx1_ASAP7_75t_L g13585 ( 
.A(n_13150),
.Y(n_13585)
);

OR2x2_ASAP7_75t_L g13586 ( 
.A(n_13141),
.B(n_13287),
.Y(n_13586)
);

BUFx6f_ASAP7_75t_L g13587 ( 
.A(n_13298),
.Y(n_13587)
);

INVx3_ASAP7_75t_L g13588 ( 
.A(n_13205),
.Y(n_13588)
);

BUFx2_ASAP7_75t_L g13589 ( 
.A(n_13174),
.Y(n_13589)
);

INVx2_ASAP7_75t_L g13590 ( 
.A(n_13252),
.Y(n_13590)
);

INVx1_ASAP7_75t_L g13591 ( 
.A(n_13259),
.Y(n_13591)
);

INVx3_ASAP7_75t_L g13592 ( 
.A(n_13088),
.Y(n_13592)
);

INVx1_ASAP7_75t_L g13593 ( 
.A(n_13363),
.Y(n_13593)
);

NAND2xp5_ASAP7_75t_L g13594 ( 
.A(n_13355),
.B(n_2219),
.Y(n_13594)
);

OAI21x1_ASAP7_75t_L g13595 ( 
.A1(n_13266),
.A2(n_2220),
.B(n_2221),
.Y(n_13595)
);

INVx3_ASAP7_75t_L g13596 ( 
.A(n_13155),
.Y(n_13596)
);

AND2x2_ASAP7_75t_L g13597 ( 
.A(n_13350),
.B(n_13362),
.Y(n_13597)
);

BUFx6f_ASAP7_75t_L g13598 ( 
.A(n_13136),
.Y(n_13598)
);

INVx1_ASAP7_75t_L g13599 ( 
.A(n_13364),
.Y(n_13599)
);

INVx2_ASAP7_75t_L g13600 ( 
.A(n_13158),
.Y(n_13600)
);

INVx2_ASAP7_75t_L g13601 ( 
.A(n_13193),
.Y(n_13601)
);

INVx2_ASAP7_75t_L g13602 ( 
.A(n_13199),
.Y(n_13602)
);

INVxp67_ASAP7_75t_L g13603 ( 
.A(n_13216),
.Y(n_13603)
);

INVx2_ASAP7_75t_L g13604 ( 
.A(n_13211),
.Y(n_13604)
);

INVx1_ASAP7_75t_L g13605 ( 
.A(n_13368),
.Y(n_13605)
);

INVx1_ASAP7_75t_L g13606 ( 
.A(n_13370),
.Y(n_13606)
);

INVx3_ASAP7_75t_L g13607 ( 
.A(n_13161),
.Y(n_13607)
);

INVx3_ASAP7_75t_L g13608 ( 
.A(n_13228),
.Y(n_13608)
);

HB1xp67_ASAP7_75t_L g13609 ( 
.A(n_13376),
.Y(n_13609)
);

AOI22xp33_ASAP7_75t_SL g13610 ( 
.A1(n_13372),
.A2(n_2222),
.B1(n_2220),
.B2(n_2221),
.Y(n_13610)
);

OAI21xp5_ASAP7_75t_L g13611 ( 
.A1(n_13062),
.A2(n_2222),
.B(n_2223),
.Y(n_13611)
);

OAI21x1_ASAP7_75t_L g13612 ( 
.A1(n_13383),
.A2(n_2223),
.B(n_2224),
.Y(n_13612)
);

INVx2_ASAP7_75t_L g13613 ( 
.A(n_13061),
.Y(n_13613)
);

AOI21xp5_ASAP7_75t_L g13614 ( 
.A1(n_13167),
.A2(n_2224),
.B(n_2225),
.Y(n_13614)
);

INVx2_ASAP7_75t_L g13615 ( 
.A(n_13369),
.Y(n_13615)
);

INVx1_ASAP7_75t_L g13616 ( 
.A(n_13325),
.Y(n_13616)
);

OAI21x1_ASAP7_75t_L g13617 ( 
.A1(n_13262),
.A2(n_2225),
.B(n_2226),
.Y(n_13617)
);

BUFx4f_ASAP7_75t_L g13618 ( 
.A(n_13341),
.Y(n_13618)
);

INVx2_ASAP7_75t_L g13619 ( 
.A(n_13375),
.Y(n_13619)
);

INVx3_ASAP7_75t_L g13620 ( 
.A(n_13174),
.Y(n_13620)
);

INVx1_ASAP7_75t_L g13621 ( 
.A(n_13349),
.Y(n_13621)
);

INVx1_ASAP7_75t_L g13622 ( 
.A(n_13147),
.Y(n_13622)
);

INVx2_ASAP7_75t_L g13623 ( 
.A(n_13153),
.Y(n_13623)
);

NOR2xp33_ASAP7_75t_L g13624 ( 
.A(n_13390),
.B(n_2227),
.Y(n_13624)
);

AND2x2_ASAP7_75t_L g13625 ( 
.A(n_13246),
.B(n_2227),
.Y(n_13625)
);

AND2x2_ASAP7_75t_L g13626 ( 
.A(n_13386),
.B(n_2228),
.Y(n_13626)
);

INVx2_ASAP7_75t_L g13627 ( 
.A(n_13279),
.Y(n_13627)
);

INVx1_ASAP7_75t_L g13628 ( 
.A(n_13260),
.Y(n_13628)
);

INVx2_ASAP7_75t_L g13629 ( 
.A(n_13047),
.Y(n_13629)
);

INVx1_ASAP7_75t_L g13630 ( 
.A(n_13104),
.Y(n_13630)
);

INVx1_ASAP7_75t_L g13631 ( 
.A(n_13128),
.Y(n_13631)
);

AND2x2_ASAP7_75t_L g13632 ( 
.A(n_13233),
.B(n_2228),
.Y(n_13632)
);

AND2x2_ASAP7_75t_L g13633 ( 
.A(n_13237),
.B(n_2229),
.Y(n_13633)
);

INVx1_ASAP7_75t_L g13634 ( 
.A(n_13138),
.Y(n_13634)
);

OR2x2_ASAP7_75t_L g13635 ( 
.A(n_13220),
.B(n_2229),
.Y(n_13635)
);

INVx1_ASAP7_75t_L g13636 ( 
.A(n_13140),
.Y(n_13636)
);

INVx1_ASAP7_75t_L g13637 ( 
.A(n_13347),
.Y(n_13637)
);

INVx1_ASAP7_75t_L g13638 ( 
.A(n_13170),
.Y(n_13638)
);

INVx1_ASAP7_75t_L g13639 ( 
.A(n_13057),
.Y(n_13639)
);

OAI22xp5_ASAP7_75t_L g13640 ( 
.A1(n_13286),
.A2(n_2232),
.B1(n_2230),
.B2(n_2231),
.Y(n_13640)
);

NAND3xp33_ASAP7_75t_L g13641 ( 
.A(n_13107),
.B(n_2230),
.C(n_2232),
.Y(n_13641)
);

NAND2xp5_ASAP7_75t_L g13642 ( 
.A(n_13302),
.B(n_2233),
.Y(n_13642)
);

INVx1_ASAP7_75t_SL g13643 ( 
.A(n_13359),
.Y(n_13643)
);

INVx3_ASAP7_75t_L g13644 ( 
.A(n_13108),
.Y(n_13644)
);

NAND2xp5_ASAP7_75t_L g13645 ( 
.A(n_13313),
.B(n_2234),
.Y(n_13645)
);

AND2x2_ASAP7_75t_L g13646 ( 
.A(n_13263),
.B(n_13236),
.Y(n_13646)
);

AND2x2_ASAP7_75t_L g13647 ( 
.A(n_13149),
.B(n_2234),
.Y(n_13647)
);

INVx1_ASAP7_75t_L g13648 ( 
.A(n_13114),
.Y(n_13648)
);

INVx1_ASAP7_75t_L g13649 ( 
.A(n_13268),
.Y(n_13649)
);

OR2x2_ASAP7_75t_L g13650 ( 
.A(n_13238),
.B(n_2235),
.Y(n_13650)
);

INVx3_ASAP7_75t_L g13651 ( 
.A(n_13272),
.Y(n_13651)
);

OAI21x1_ASAP7_75t_L g13652 ( 
.A1(n_13133),
.A2(n_2235),
.B(n_2236),
.Y(n_13652)
);

INVx1_ASAP7_75t_L g13653 ( 
.A(n_13300),
.Y(n_13653)
);

INVx2_ASAP7_75t_L g13654 ( 
.A(n_13047),
.Y(n_13654)
);

INVx2_ASAP7_75t_SL g13655 ( 
.A(n_13344),
.Y(n_13655)
);

INVx1_ASAP7_75t_L g13656 ( 
.A(n_13382),
.Y(n_13656)
);

BUFx3_ASAP7_75t_L g13657 ( 
.A(n_13329),
.Y(n_13657)
);

INVx1_ASAP7_75t_L g13658 ( 
.A(n_13099),
.Y(n_13658)
);

INVx1_ASAP7_75t_L g13659 ( 
.A(n_13360),
.Y(n_13659)
);

BUFx2_ASAP7_75t_L g13660 ( 
.A(n_13272),
.Y(n_13660)
);

INVx1_ASAP7_75t_L g13661 ( 
.A(n_13381),
.Y(n_13661)
);

INVx6_ASAP7_75t_L g13662 ( 
.A(n_13327),
.Y(n_13662)
);

INVx2_ASAP7_75t_L g13663 ( 
.A(n_13064),
.Y(n_13663)
);

INVx3_ASAP7_75t_L g13664 ( 
.A(n_13116),
.Y(n_13664)
);

AND2x2_ASAP7_75t_L g13665 ( 
.A(n_13388),
.B(n_2236),
.Y(n_13665)
);

BUFx2_ASAP7_75t_L g13666 ( 
.A(n_13380),
.Y(n_13666)
);

INVx2_ASAP7_75t_L g13667 ( 
.A(n_13163),
.Y(n_13667)
);

AND2x2_ASAP7_75t_L g13668 ( 
.A(n_13317),
.B(n_2237),
.Y(n_13668)
);

OAI21xp5_ASAP7_75t_L g13669 ( 
.A1(n_13106),
.A2(n_2238),
.B(n_2239),
.Y(n_13669)
);

BUFx2_ASAP7_75t_L g13670 ( 
.A(n_13373),
.Y(n_13670)
);

OAI21xp5_ASAP7_75t_L g13671 ( 
.A1(n_13177),
.A2(n_2240),
.B(n_2241),
.Y(n_13671)
);

INVx1_ASAP7_75t_L g13672 ( 
.A(n_13182),
.Y(n_13672)
);

INVx1_ASAP7_75t_L g13673 ( 
.A(n_13200),
.Y(n_13673)
);

OR2x2_ASAP7_75t_L g13674 ( 
.A(n_13223),
.B(n_2240),
.Y(n_13674)
);

INVx2_ASAP7_75t_L g13675 ( 
.A(n_13379),
.Y(n_13675)
);

INVx1_ASAP7_75t_L g13676 ( 
.A(n_13239),
.Y(n_13676)
);

INVx1_ASAP7_75t_L g13677 ( 
.A(n_13248),
.Y(n_13677)
);

BUFx12f_ASAP7_75t_L g13678 ( 
.A(n_13328),
.Y(n_13678)
);

AND2x4_ASAP7_75t_L g13679 ( 
.A(n_13365),
.B(n_2241),
.Y(n_13679)
);

INVx2_ASAP7_75t_L g13680 ( 
.A(n_13139),
.Y(n_13680)
);

INVx1_ASAP7_75t_L g13681 ( 
.A(n_13134),
.Y(n_13681)
);

INVx1_ASAP7_75t_L g13682 ( 
.A(n_13173),
.Y(n_13682)
);

INVx1_ASAP7_75t_L g13683 ( 
.A(n_13310),
.Y(n_13683)
);

INVx1_ASAP7_75t_L g13684 ( 
.A(n_13345),
.Y(n_13684)
);

BUFx3_ASAP7_75t_L g13685 ( 
.A(n_13142),
.Y(n_13685)
);

AND2x2_ASAP7_75t_L g13686 ( 
.A(n_13224),
.B(n_2242),
.Y(n_13686)
);

INVx2_ASAP7_75t_SL g13687 ( 
.A(n_13154),
.Y(n_13687)
);

INVxp67_ASAP7_75t_L g13688 ( 
.A(n_13326),
.Y(n_13688)
);

INVx1_ASAP7_75t_L g13689 ( 
.A(n_13278),
.Y(n_13689)
);

INVx2_ASAP7_75t_L g13690 ( 
.A(n_13284),
.Y(n_13690)
);

INVx1_ASAP7_75t_L g13691 ( 
.A(n_13210),
.Y(n_13691)
);

INVx2_ASAP7_75t_L g13692 ( 
.A(n_13221),
.Y(n_13692)
);

INVx2_ASAP7_75t_L g13693 ( 
.A(n_13277),
.Y(n_13693)
);

INVx1_ASAP7_75t_L g13694 ( 
.A(n_13295),
.Y(n_13694)
);

INVx2_ASAP7_75t_L g13695 ( 
.A(n_13208),
.Y(n_13695)
);

INVx1_ASAP7_75t_L g13696 ( 
.A(n_13160),
.Y(n_13696)
);

BUFx12f_ASAP7_75t_L g13697 ( 
.A(n_13357),
.Y(n_13697)
);

OA21x2_ASAP7_75t_L g13698 ( 
.A1(n_13168),
.A2(n_2242),
.B(n_2243),
.Y(n_13698)
);

INVx1_ASAP7_75t_SL g13699 ( 
.A(n_13308),
.Y(n_13699)
);

INVx1_ASAP7_75t_L g13700 ( 
.A(n_13323),
.Y(n_13700)
);

BUFx3_ASAP7_75t_L g13701 ( 
.A(n_13303),
.Y(n_13701)
);

INVx2_ASAP7_75t_L g13702 ( 
.A(n_13079),
.Y(n_13702)
);

INVx1_ASAP7_75t_L g13703 ( 
.A(n_13282),
.Y(n_13703)
);

INVx1_ASAP7_75t_L g13704 ( 
.A(n_13282),
.Y(n_13704)
);

AOI21xp5_ASAP7_75t_L g13705 ( 
.A1(n_13151),
.A2(n_2243),
.B(n_2244),
.Y(n_13705)
);

INVx2_ASAP7_75t_L g13706 ( 
.A(n_13351),
.Y(n_13706)
);

INVx1_ASAP7_75t_L g13707 ( 
.A(n_13183),
.Y(n_13707)
);

NAND2xp5_ASAP7_75t_SL g13708 ( 
.A(n_13305),
.B(n_2244),
.Y(n_13708)
);

INVx1_ASAP7_75t_L g13709 ( 
.A(n_13338),
.Y(n_13709)
);

HB1xp67_ASAP7_75t_L g13710 ( 
.A(n_13291),
.Y(n_13710)
);

INVx2_ASAP7_75t_SL g13711 ( 
.A(n_13297),
.Y(n_13711)
);

AND2x2_ASAP7_75t_L g13712 ( 
.A(n_13273),
.B(n_2245),
.Y(n_13712)
);

AND2x2_ASAP7_75t_L g13713 ( 
.A(n_13330),
.B(n_2246),
.Y(n_13713)
);

HB1xp67_ASAP7_75t_L g13714 ( 
.A(n_13320),
.Y(n_13714)
);

INVx2_ASAP7_75t_L g13715 ( 
.A(n_13371),
.Y(n_13715)
);

INVx2_ASAP7_75t_L g13716 ( 
.A(n_13318),
.Y(n_13716)
);

INVx1_ASAP7_75t_L g13717 ( 
.A(n_13343),
.Y(n_13717)
);

BUFx4f_ASAP7_75t_SL g13718 ( 
.A(n_13389),
.Y(n_13718)
);

AND2x2_ASAP7_75t_L g13719 ( 
.A(n_13361),
.B(n_2247),
.Y(n_13719)
);

HB1xp67_ASAP7_75t_L g13720 ( 
.A(n_13366),
.Y(n_13720)
);

INVx1_ASAP7_75t_L g13721 ( 
.A(n_13378),
.Y(n_13721)
);

INVx2_ASAP7_75t_L g13722 ( 
.A(n_13366),
.Y(n_13722)
);

INVx1_ASAP7_75t_L g13723 ( 
.A(n_13332),
.Y(n_13723)
);

INVx2_ASAP7_75t_L g13724 ( 
.A(n_13334),
.Y(n_13724)
);

INVx2_ASAP7_75t_L g13725 ( 
.A(n_13334),
.Y(n_13725)
);

INVx1_ASAP7_75t_L g13726 ( 
.A(n_13332),
.Y(n_13726)
);

INVx1_ASAP7_75t_L g13727 ( 
.A(n_13292),
.Y(n_13727)
);

CKINVDCx5p33_ASAP7_75t_R g13728 ( 
.A(n_13192),
.Y(n_13728)
);

INVx2_ASAP7_75t_L g13729 ( 
.A(n_13292),
.Y(n_13729)
);

OR2x2_ASAP7_75t_L g13730 ( 
.A(n_13244),
.B(n_2247),
.Y(n_13730)
);

INVx1_ASAP7_75t_L g13731 ( 
.A(n_13219),
.Y(n_13731)
);

INVx1_ASAP7_75t_L g13732 ( 
.A(n_13121),
.Y(n_13732)
);

AND2x4_ASAP7_75t_L g13733 ( 
.A(n_13242),
.B(n_2248),
.Y(n_13733)
);

AOI21x1_ASAP7_75t_L g13734 ( 
.A1(n_13144),
.A2(n_13289),
.B(n_13339),
.Y(n_13734)
);

INVx1_ASAP7_75t_L g13735 ( 
.A(n_13254),
.Y(n_13735)
);

OAI21x1_ASAP7_75t_L g13736 ( 
.A1(n_13059),
.A2(n_2249),
.B(n_2250),
.Y(n_13736)
);

INVx1_ASAP7_75t_L g13737 ( 
.A(n_13203),
.Y(n_13737)
);

AND2x4_ASAP7_75t_L g13738 ( 
.A(n_13076),
.B(n_2249),
.Y(n_13738)
);

INVx2_ASAP7_75t_L g13739 ( 
.A(n_13307),
.Y(n_13739)
);

INVx1_ASAP7_75t_L g13740 ( 
.A(n_13240),
.Y(n_13740)
);

AOI22xp33_ASAP7_75t_SL g13741 ( 
.A1(n_13714),
.A2(n_13340),
.B1(n_13342),
.B2(n_13253),
.Y(n_13741)
);

HB1xp67_ASAP7_75t_L g13742 ( 
.A(n_13399),
.Y(n_13742)
);

INVx4_ASAP7_75t_SL g13743 ( 
.A(n_13429),
.Y(n_13743)
);

OAI22xp5_ASAP7_75t_L g13744 ( 
.A1(n_13455),
.A2(n_13081),
.B1(n_13198),
.B2(n_13385),
.Y(n_13744)
);

OAI22xp5_ASAP7_75t_L g13745 ( 
.A1(n_13455),
.A2(n_13117),
.B1(n_13250),
.B2(n_13348),
.Y(n_13745)
);

OAI22xp5_ASAP7_75t_L g13746 ( 
.A1(n_13541),
.A2(n_13304),
.B1(n_13166),
.B2(n_13333),
.Y(n_13746)
);

NAND2xp5_ASAP7_75t_L g13747 ( 
.A(n_13690),
.B(n_13111),
.Y(n_13747)
);

NAND2xp5_ASAP7_75t_SL g13748 ( 
.A(n_13505),
.B(n_13400),
.Y(n_13748)
);

INVx1_ASAP7_75t_L g13749 ( 
.A(n_13412),
.Y(n_13749)
);

AOI21xp5_ASAP7_75t_L g13750 ( 
.A1(n_13552),
.A2(n_13346),
.B(n_13358),
.Y(n_13750)
);

NAND2x1p5_ASAP7_75t_L g13751 ( 
.A(n_13400),
.B(n_13367),
.Y(n_13751)
);

INVxp67_ASAP7_75t_L g13752 ( 
.A(n_13539),
.Y(n_13752)
);

NAND2xp5_ASAP7_75t_SL g13753 ( 
.A(n_13477),
.B(n_2250),
.Y(n_13753)
);

OAI22xp5_ASAP7_75t_L g13754 ( 
.A1(n_13688),
.A2(n_2253),
.B1(n_2251),
.B2(n_2252),
.Y(n_13754)
);

AND2x2_ASAP7_75t_L g13755 ( 
.A(n_13493),
.B(n_2251),
.Y(n_13755)
);

INVx8_ASAP7_75t_L g13756 ( 
.A(n_13429),
.Y(n_13756)
);

OAI22xp5_ASAP7_75t_L g13757 ( 
.A1(n_13731),
.A2(n_2255),
.B1(n_2252),
.B2(n_2254),
.Y(n_13757)
);

AOI222xp33_ASAP7_75t_L g13758 ( 
.A1(n_13641),
.A2(n_2257),
.B1(n_2259),
.B2(n_2254),
.C1(n_2256),
.C2(n_2258),
.Y(n_13758)
);

AOI21xp33_ASAP7_75t_L g13759 ( 
.A1(n_13544),
.A2(n_2257),
.B(n_2258),
.Y(n_13759)
);

HB1xp67_ASAP7_75t_L g13760 ( 
.A(n_13407),
.Y(n_13760)
);

INVxp67_ASAP7_75t_L g13761 ( 
.A(n_13660),
.Y(n_13761)
);

INVx1_ASAP7_75t_L g13762 ( 
.A(n_13472),
.Y(n_13762)
);

NAND2xp5_ASAP7_75t_SL g13763 ( 
.A(n_13477),
.B(n_2259),
.Y(n_13763)
);

AOI22xp33_ASAP7_75t_L g13764 ( 
.A1(n_13739),
.A2(n_2262),
.B1(n_2260),
.B2(n_2261),
.Y(n_13764)
);

AOI22xp33_ASAP7_75t_L g13765 ( 
.A1(n_13419),
.A2(n_2262),
.B1(n_2260),
.B2(n_2261),
.Y(n_13765)
);

AND2x2_ASAP7_75t_L g13766 ( 
.A(n_13447),
.B(n_2263),
.Y(n_13766)
);

AOI221xp5_ASAP7_75t_L g13767 ( 
.A1(n_13517),
.A2(n_13720),
.B1(n_13687),
.B2(n_13707),
.C(n_13545),
.Y(n_13767)
);

AOI22xp33_ASAP7_75t_SL g13768 ( 
.A1(n_13488),
.A2(n_2265),
.B1(n_2263),
.B2(n_2264),
.Y(n_13768)
);

AOI22xp33_ASAP7_75t_L g13769 ( 
.A1(n_13524),
.A2(n_2268),
.B1(n_2266),
.B2(n_2267),
.Y(n_13769)
);

AOI22xp33_ASAP7_75t_SL g13770 ( 
.A1(n_13416),
.A2(n_2269),
.B1(n_2266),
.B2(n_2267),
.Y(n_13770)
);

OAI21xp33_ASAP7_75t_SL g13771 ( 
.A1(n_13516),
.A2(n_2270),
.B(n_2271),
.Y(n_13771)
);

INVx1_ASAP7_75t_L g13772 ( 
.A(n_13496),
.Y(n_13772)
);

OR2x2_ASAP7_75t_L g13773 ( 
.A(n_13395),
.B(n_2270),
.Y(n_13773)
);

OAI22xp33_ASAP7_75t_L g13774 ( 
.A1(n_13524),
.A2(n_2273),
.B1(n_2271),
.B2(n_2272),
.Y(n_13774)
);

OAI22xp33_ASAP7_75t_L g13775 ( 
.A1(n_13520),
.A2(n_2276),
.B1(n_2272),
.B2(n_2274),
.Y(n_13775)
);

AOI22xp33_ASAP7_75t_L g13776 ( 
.A1(n_13735),
.A2(n_13520),
.B1(n_13411),
.B2(n_13537),
.Y(n_13776)
);

INVx3_ASAP7_75t_L g13777 ( 
.A(n_13408),
.Y(n_13777)
);

AOI22xp33_ASAP7_75t_L g13778 ( 
.A1(n_13717),
.A2(n_2278),
.B1(n_2276),
.B2(n_2277),
.Y(n_13778)
);

AOI21xp33_ASAP7_75t_L g13779 ( 
.A1(n_13730),
.A2(n_2277),
.B(n_2279),
.Y(n_13779)
);

CKINVDCx5p33_ASAP7_75t_R g13780 ( 
.A(n_13525),
.Y(n_13780)
);

AOI21xp5_ASAP7_75t_L g13781 ( 
.A1(n_13483),
.A2(n_2280),
.B(n_2281),
.Y(n_13781)
);

OAI22xp5_ASAP7_75t_L g13782 ( 
.A1(n_13575),
.A2(n_2282),
.B1(n_2280),
.B2(n_2281),
.Y(n_13782)
);

NAND3xp33_ASAP7_75t_L g13783 ( 
.A(n_13476),
.B(n_13581),
.C(n_13500),
.Y(n_13783)
);

CKINVDCx5p33_ASAP7_75t_R g13784 ( 
.A(n_13437),
.Y(n_13784)
);

AOI221xp5_ASAP7_75t_L g13785 ( 
.A1(n_13691),
.A2(n_2284),
.B1(n_2282),
.B2(n_2283),
.C(n_2285),
.Y(n_13785)
);

AND2x2_ASAP7_75t_L g13786 ( 
.A(n_13589),
.B(n_2284),
.Y(n_13786)
);

AND2x4_ASAP7_75t_L g13787 ( 
.A(n_13402),
.B(n_2285),
.Y(n_13787)
);

NAND3xp33_ASAP7_75t_L g13788 ( 
.A(n_13610),
.B(n_2286),
.C(n_2288),
.Y(n_13788)
);

INVx3_ASAP7_75t_L g13789 ( 
.A(n_13408),
.Y(n_13789)
);

AOI22xp33_ASAP7_75t_L g13790 ( 
.A1(n_13718),
.A2(n_2289),
.B1(n_2286),
.B2(n_2288),
.Y(n_13790)
);

INVx4_ASAP7_75t_L g13791 ( 
.A(n_13446),
.Y(n_13791)
);

OR2x2_ASAP7_75t_L g13792 ( 
.A(n_13532),
.B(n_2289),
.Y(n_13792)
);

AOI21xp33_ASAP7_75t_L g13793 ( 
.A1(n_13586),
.A2(n_2290),
.B(n_2291),
.Y(n_13793)
);

HB1xp67_ASAP7_75t_L g13794 ( 
.A(n_13519),
.Y(n_13794)
);

NAND3xp33_ASAP7_75t_L g13795 ( 
.A(n_13637),
.B(n_2290),
.C(n_2292),
.Y(n_13795)
);

AOI22xp33_ASAP7_75t_L g13796 ( 
.A1(n_13452),
.A2(n_2294),
.B1(n_2292),
.B2(n_2293),
.Y(n_13796)
);

INVx1_ASAP7_75t_L g13797 ( 
.A(n_13580),
.Y(n_13797)
);

OAI211xp5_ASAP7_75t_L g13798 ( 
.A1(n_13449),
.A2(n_13508),
.B(n_13669),
.C(n_13611),
.Y(n_13798)
);

AOI22xp33_ASAP7_75t_L g13799 ( 
.A1(n_13728),
.A2(n_2297),
.B1(n_2295),
.B2(n_2296),
.Y(n_13799)
);

AOI222xp33_ASAP7_75t_L g13800 ( 
.A1(n_13732),
.A2(n_2297),
.B1(n_2299),
.B2(n_2295),
.C1(n_2296),
.C2(n_2298),
.Y(n_13800)
);

BUFx2_ASAP7_75t_L g13801 ( 
.A(n_13697),
.Y(n_13801)
);

INVx2_ASAP7_75t_L g13802 ( 
.A(n_13462),
.Y(n_13802)
);

NAND3xp33_ASAP7_75t_L g13803 ( 
.A(n_13583),
.B(n_2298),
.C(n_2299),
.Y(n_13803)
);

OAI22xp5_ASAP7_75t_L g13804 ( 
.A1(n_13585),
.A2(n_2302),
.B1(n_2300),
.B2(n_2301),
.Y(n_13804)
);

OAI22xp5_ASAP7_75t_L g13805 ( 
.A1(n_13547),
.A2(n_2302),
.B1(n_2300),
.B2(n_2301),
.Y(n_13805)
);

AOI221xp5_ASAP7_75t_L g13806 ( 
.A1(n_13694),
.A2(n_2305),
.B1(n_2303),
.B2(n_2304),
.C(n_2306),
.Y(n_13806)
);

INVx1_ASAP7_75t_L g13807 ( 
.A(n_13556),
.Y(n_13807)
);

AOI22xp5_ASAP7_75t_L g13808 ( 
.A1(n_13426),
.A2(n_2305),
.B1(n_2303),
.B2(n_2304),
.Y(n_13808)
);

OAI211xp5_ASAP7_75t_L g13809 ( 
.A1(n_13521),
.A2(n_2308),
.B(n_2306),
.C(n_2307),
.Y(n_13809)
);

AOI21xp5_ASAP7_75t_L g13810 ( 
.A1(n_13708),
.A2(n_2307),
.B(n_2308),
.Y(n_13810)
);

OAI211xp5_ASAP7_75t_SL g13811 ( 
.A1(n_13737),
.A2(n_2311),
.B(n_2309),
.C(n_2310),
.Y(n_13811)
);

OAI22xp5_ASAP7_75t_L g13812 ( 
.A1(n_13458),
.A2(n_2313),
.B1(n_2310),
.B2(n_2312),
.Y(n_13812)
);

AOI211xp5_ASAP7_75t_L g13813 ( 
.A1(n_13478),
.A2(n_2315),
.B(n_2312),
.C(n_2314),
.Y(n_13813)
);

INVx1_ASAP7_75t_L g13814 ( 
.A(n_13512),
.Y(n_13814)
);

INVx1_ASAP7_75t_L g13815 ( 
.A(n_13513),
.Y(n_13815)
);

AND2x2_ASAP7_75t_L g13816 ( 
.A(n_13433),
.B(n_2314),
.Y(n_13816)
);

AOI221xp5_ASAP7_75t_L g13817 ( 
.A1(n_13692),
.A2(n_13693),
.B1(n_13740),
.B2(n_13518),
.C(n_13603),
.Y(n_13817)
);

BUFx4f_ASAP7_75t_SL g13818 ( 
.A(n_13567),
.Y(n_13818)
);

INVx1_ASAP7_75t_L g13819 ( 
.A(n_13396),
.Y(n_13819)
);

AOI222xp33_ASAP7_75t_L g13820 ( 
.A1(n_13653),
.A2(n_2317),
.B1(n_2319),
.B2(n_2315),
.C1(n_2316),
.C2(n_2318),
.Y(n_13820)
);

OAI22xp5_ASAP7_75t_L g13821 ( 
.A1(n_13420),
.A2(n_2318),
.B1(n_2316),
.B2(n_2317),
.Y(n_13821)
);

NAND2xp5_ASAP7_75t_L g13822 ( 
.A(n_13716),
.B(n_2319),
.Y(n_13822)
);

AOI22xp5_ASAP7_75t_L g13823 ( 
.A1(n_13506),
.A2(n_2322),
.B1(n_2320),
.B2(n_2321),
.Y(n_13823)
);

AOI22xp33_ASAP7_75t_L g13824 ( 
.A1(n_13434),
.A2(n_2323),
.B1(n_2320),
.B2(n_2321),
.Y(n_13824)
);

AND2x2_ASAP7_75t_L g13825 ( 
.A(n_13451),
.B(n_2324),
.Y(n_13825)
);

INVx1_ASAP7_75t_L g13826 ( 
.A(n_13397),
.Y(n_13826)
);

AOI22xp33_ASAP7_75t_L g13827 ( 
.A1(n_13738),
.A2(n_2326),
.B1(n_2324),
.B2(n_2325),
.Y(n_13827)
);

AOI21xp5_ASAP7_75t_L g13828 ( 
.A1(n_13414),
.A2(n_2325),
.B(n_2326),
.Y(n_13828)
);

AND2x2_ASAP7_75t_L g13829 ( 
.A(n_13422),
.B(n_2327),
.Y(n_13829)
);

INVx1_ASAP7_75t_L g13830 ( 
.A(n_13403),
.Y(n_13830)
);

INVx1_ASAP7_75t_L g13831 ( 
.A(n_13404),
.Y(n_13831)
);

BUFx12f_ASAP7_75t_L g13832 ( 
.A(n_13392),
.Y(n_13832)
);

INVx1_ASAP7_75t_L g13833 ( 
.A(n_13409),
.Y(n_13833)
);

OAI211xp5_ASAP7_75t_L g13834 ( 
.A1(n_13671),
.A2(n_2329),
.B(n_2327),
.C(n_2328),
.Y(n_13834)
);

AO31x2_ASAP7_75t_L g13835 ( 
.A1(n_13629),
.A2(n_2330),
.A3(n_2328),
.B(n_2329),
.Y(n_13835)
);

AOI22xp5_ASAP7_75t_L g13836 ( 
.A1(n_13398),
.A2(n_2332),
.B1(n_2330),
.B2(n_2331),
.Y(n_13836)
);

AOI22xp33_ASAP7_75t_L g13837 ( 
.A1(n_13616),
.A2(n_2333),
.B1(n_2331),
.B2(n_2332),
.Y(n_13837)
);

AOI22xp33_ASAP7_75t_L g13838 ( 
.A1(n_13621),
.A2(n_2336),
.B1(n_2333),
.B2(n_2335),
.Y(n_13838)
);

INVx2_ASAP7_75t_L g13839 ( 
.A(n_13462),
.Y(n_13839)
);

OR2x6_ASAP7_75t_L g13840 ( 
.A(n_13392),
.B(n_2335),
.Y(n_13840)
);

OAI22xp5_ASAP7_75t_L g13841 ( 
.A1(n_13620),
.A2(n_13440),
.B1(n_13436),
.B2(n_13651),
.Y(n_13841)
);

OAI22xp5_ASAP7_75t_L g13842 ( 
.A1(n_13440),
.A2(n_2338),
.B1(n_2336),
.B2(n_2337),
.Y(n_13842)
);

INVx1_ASAP7_75t_L g13843 ( 
.A(n_13413),
.Y(n_13843)
);

AOI22xp33_ASAP7_75t_L g13844 ( 
.A1(n_13733),
.A2(n_2340),
.B1(n_2337),
.B2(n_2339),
.Y(n_13844)
);

INVx3_ASAP7_75t_L g13845 ( 
.A(n_13467),
.Y(n_13845)
);

OAI21xp33_ASAP7_75t_L g13846 ( 
.A1(n_13454),
.A2(n_2339),
.B(n_2340),
.Y(n_13846)
);

BUFx2_ASAP7_75t_L g13847 ( 
.A(n_13678),
.Y(n_13847)
);

OAI22xp5_ASAP7_75t_L g13848 ( 
.A1(n_13435),
.A2(n_2344),
.B1(n_2341),
.B2(n_2343),
.Y(n_13848)
);

INVx2_ASAP7_75t_L g13849 ( 
.A(n_13441),
.Y(n_13849)
);

AOI21xp5_ASAP7_75t_L g13850 ( 
.A1(n_13643),
.A2(n_2341),
.B(n_2343),
.Y(n_13850)
);

AOI21xp33_ASAP7_75t_L g13851 ( 
.A1(n_13543),
.A2(n_2344),
.B(n_2345),
.Y(n_13851)
);

INVx1_ASAP7_75t_L g13852 ( 
.A(n_13421),
.Y(n_13852)
);

AOI221xp5_ASAP7_75t_L g13853 ( 
.A1(n_13683),
.A2(n_2347),
.B1(n_2345),
.B2(n_2346),
.C(n_2348),
.Y(n_13853)
);

AOI21xp5_ASAP7_75t_L g13854 ( 
.A1(n_13444),
.A2(n_2346),
.B(n_2347),
.Y(n_13854)
);

AND2x2_ASAP7_75t_L g13855 ( 
.A(n_13427),
.B(n_2348),
.Y(n_13855)
);

OAI21x1_ASAP7_75t_L g13856 ( 
.A1(n_13490),
.A2(n_13432),
.B(n_13491),
.Y(n_13856)
);

OAI221xp5_ASAP7_75t_L g13857 ( 
.A1(n_13599),
.A2(n_2351),
.B1(n_2349),
.B2(n_2350),
.C(n_2352),
.Y(n_13857)
);

OAI221xp5_ASAP7_75t_L g13858 ( 
.A1(n_13503),
.A2(n_2352),
.B1(n_2349),
.B2(n_2350),
.C(n_2353),
.Y(n_13858)
);

NAND2xp5_ASAP7_75t_L g13859 ( 
.A(n_13438),
.B(n_13663),
.Y(n_13859)
);

OR2x6_ASAP7_75t_L g13860 ( 
.A(n_13410),
.B(n_2353),
.Y(n_13860)
);

AOI21xp5_ASAP7_75t_L g13861 ( 
.A1(n_13642),
.A2(n_2354),
.B(n_2355),
.Y(n_13861)
);

OAI22xp33_ASAP7_75t_L g13862 ( 
.A1(n_13515),
.A2(n_2356),
.B1(n_2354),
.B2(n_2355),
.Y(n_13862)
);

OAI22xp33_ASAP7_75t_L g13863 ( 
.A1(n_13515),
.A2(n_2358),
.B1(n_2356),
.B2(n_2357),
.Y(n_13863)
);

NAND2xp5_ASAP7_75t_L g13864 ( 
.A(n_13721),
.B(n_2357),
.Y(n_13864)
);

INVx1_ASAP7_75t_L g13865 ( 
.A(n_13423),
.Y(n_13865)
);

AOI22xp33_ASAP7_75t_SL g13866 ( 
.A1(n_13666),
.A2(n_2361),
.B1(n_2358),
.B2(n_2360),
.Y(n_13866)
);

AOI221xp5_ASAP7_75t_L g13867 ( 
.A1(n_13722),
.A2(n_2364),
.B1(n_2362),
.B2(n_2363),
.C(n_2365),
.Y(n_13867)
);

OAI221xp5_ASAP7_75t_L g13868 ( 
.A1(n_13734),
.A2(n_2364),
.B1(n_2362),
.B2(n_2363),
.C(n_2365),
.Y(n_13868)
);

AOI22xp33_ASAP7_75t_L g13869 ( 
.A1(n_13701),
.A2(n_2368),
.B1(n_2366),
.B2(n_2367),
.Y(n_13869)
);

AND2x2_ASAP7_75t_L g13870 ( 
.A(n_13415),
.B(n_2366),
.Y(n_13870)
);

AOI221xp5_ASAP7_75t_L g13871 ( 
.A1(n_13727),
.A2(n_2371),
.B1(n_2369),
.B2(n_2370),
.C(n_2372),
.Y(n_13871)
);

AOI22xp33_ASAP7_75t_L g13872 ( 
.A1(n_13696),
.A2(n_2373),
.B1(n_2370),
.B2(n_2372),
.Y(n_13872)
);

INVx2_ASAP7_75t_L g13873 ( 
.A(n_13662),
.Y(n_13873)
);

BUFx12f_ASAP7_75t_L g13874 ( 
.A(n_13558),
.Y(n_13874)
);

AOI222xp33_ASAP7_75t_L g13875 ( 
.A1(n_13649),
.A2(n_2375),
.B1(n_2377),
.B2(n_2373),
.C1(n_2374),
.C2(n_2376),
.Y(n_13875)
);

OAI21xp33_ASAP7_75t_L g13876 ( 
.A1(n_13562),
.A2(n_2374),
.B(n_2375),
.Y(n_13876)
);

INVx1_ASAP7_75t_L g13877 ( 
.A(n_13428),
.Y(n_13877)
);

OAI211xp5_ASAP7_75t_L g13878 ( 
.A1(n_13417),
.A2(n_2379),
.B(n_2377),
.C(n_2378),
.Y(n_13878)
);

AOI22xp33_ASAP7_75t_L g13879 ( 
.A1(n_13401),
.A2(n_2380),
.B1(n_2378),
.B2(n_2379),
.Y(n_13879)
);

NOR2xp33_ASAP7_75t_L g13880 ( 
.A(n_13424),
.B(n_2381),
.Y(n_13880)
);

INVx1_ASAP7_75t_L g13881 ( 
.A(n_13431),
.Y(n_13881)
);

OR2x2_ASAP7_75t_L g13882 ( 
.A(n_13470),
.B(n_2381),
.Y(n_13882)
);

INVx2_ASAP7_75t_L g13883 ( 
.A(n_13464),
.Y(n_13883)
);

AOI22xp5_ASAP7_75t_L g13884 ( 
.A1(n_13418),
.A2(n_2384),
.B1(n_2382),
.B2(n_2383),
.Y(n_13884)
);

A2O1A1Ixp33_ASAP7_75t_L g13885 ( 
.A1(n_13614),
.A2(n_2384),
.B(n_2382),
.C(n_2383),
.Y(n_13885)
);

BUFx3_ASAP7_75t_L g13886 ( 
.A(n_13573),
.Y(n_13886)
);

NAND2xp5_ASAP7_75t_L g13887 ( 
.A(n_13592),
.B(n_2385),
.Y(n_13887)
);

AOI221xp5_ASAP7_75t_L g13888 ( 
.A1(n_13723),
.A2(n_2387),
.B1(n_2385),
.B2(n_2386),
.C(n_2388),
.Y(n_13888)
);

BUFx3_ASAP7_75t_L g13889 ( 
.A(n_13588),
.Y(n_13889)
);

AOI22xp33_ASAP7_75t_L g13890 ( 
.A1(n_13638),
.A2(n_2388),
.B1(n_2386),
.B2(n_2387),
.Y(n_13890)
);

INVx2_ASAP7_75t_L g13891 ( 
.A(n_13569),
.Y(n_13891)
);

AOI22xp33_ASAP7_75t_L g13892 ( 
.A1(n_13670),
.A2(n_13700),
.B1(n_13631),
.B2(n_13636),
.Y(n_13892)
);

AND2x4_ASAP7_75t_L g13893 ( 
.A(n_13657),
.B(n_2389),
.Y(n_13893)
);

OAI221xp5_ASAP7_75t_L g13894 ( 
.A1(n_13469),
.A2(n_2391),
.B1(n_2389),
.B2(n_2390),
.C(n_2392),
.Y(n_13894)
);

OAI22xp33_ASAP7_75t_L g13895 ( 
.A1(n_13703),
.A2(n_2393),
.B1(n_2390),
.B2(n_2391),
.Y(n_13895)
);

OAI22xp5_ASAP7_75t_L g13896 ( 
.A1(n_13664),
.A2(n_2395),
.B1(n_2393),
.B2(n_2394),
.Y(n_13896)
);

AOI21xp5_ASAP7_75t_L g13897 ( 
.A1(n_13645),
.A2(n_2395),
.B(n_2396),
.Y(n_13897)
);

AND2x2_ASAP7_75t_L g13898 ( 
.A(n_13405),
.B(n_2396),
.Y(n_13898)
);

AOI221xp5_ASAP7_75t_L g13899 ( 
.A1(n_13726),
.A2(n_2400),
.B1(n_2397),
.B2(n_2399),
.C(n_2401),
.Y(n_13899)
);

OAI221xp5_ASAP7_75t_L g13900 ( 
.A1(n_13680),
.A2(n_2401),
.B1(n_2397),
.B2(n_2400),
.C(n_2402),
.Y(n_13900)
);

CKINVDCx20_ASAP7_75t_R g13901 ( 
.A(n_13453),
.Y(n_13901)
);

NAND2xp5_ASAP7_75t_L g13902 ( 
.A(n_13698),
.B(n_2402),
.Y(n_13902)
);

AO21x2_ASAP7_75t_L g13903 ( 
.A1(n_13654),
.A2(n_2403),
.B(n_2404),
.Y(n_13903)
);

NAND2xp5_ASAP7_75t_L g13904 ( 
.A(n_13667),
.B(n_2403),
.Y(n_13904)
);

OAI22xp33_ASAP7_75t_L g13905 ( 
.A1(n_13704),
.A2(n_2406),
.B1(n_2404),
.B2(n_2405),
.Y(n_13905)
);

AND2x2_ASAP7_75t_L g13906 ( 
.A(n_13675),
.B(n_2405),
.Y(n_13906)
);

OAI211xp5_ASAP7_75t_L g13907 ( 
.A1(n_13705),
.A2(n_2408),
.B(n_2406),
.C(n_2407),
.Y(n_13907)
);

OAI211xp5_ASAP7_75t_L g13908 ( 
.A1(n_13570),
.A2(n_2409),
.B(n_2407),
.C(n_2408),
.Y(n_13908)
);

BUFx4f_ASAP7_75t_SL g13909 ( 
.A(n_13578),
.Y(n_13909)
);

AOI21xp5_ASAP7_75t_L g13910 ( 
.A1(n_13618),
.A2(n_2409),
.B(n_2410),
.Y(n_13910)
);

BUFx3_ASAP7_75t_L g13911 ( 
.A(n_13473),
.Y(n_13911)
);

A2O1A1Ixp33_ASAP7_75t_L g13912 ( 
.A1(n_13549),
.A2(n_2412),
.B(n_2410),
.C(n_2411),
.Y(n_13912)
);

OR2x6_ASAP7_75t_SL g13913 ( 
.A(n_13702),
.B(n_2412),
.Y(n_13913)
);

AND2x2_ASAP7_75t_L g13914 ( 
.A(n_13459),
.B(n_2413),
.Y(n_13914)
);

AOI32xp33_ASAP7_75t_L g13915 ( 
.A1(n_13686),
.A2(n_2415),
.A3(n_2413),
.B1(n_2414),
.B2(n_2416),
.Y(n_13915)
);

AND2x4_ASAP7_75t_L g13916 ( 
.A(n_13523),
.B(n_2414),
.Y(n_13916)
);

NOR2xp33_ASAP7_75t_L g13917 ( 
.A(n_13598),
.B(n_2415),
.Y(n_13917)
);

INVx2_ASAP7_75t_L g13918 ( 
.A(n_13569),
.Y(n_13918)
);

AOI22xp33_ASAP7_75t_SL g13919 ( 
.A1(n_13644),
.A2(n_2418),
.B1(n_2416),
.B2(n_2417),
.Y(n_13919)
);

OAI22xp5_ASAP7_75t_L g13920 ( 
.A1(n_13534),
.A2(n_2419),
.B1(n_2417),
.B2(n_2418),
.Y(n_13920)
);

AO31x2_ASAP7_75t_L g13921 ( 
.A1(n_13542),
.A2(n_2421),
.A3(n_2419),
.B(n_2420),
.Y(n_13921)
);

OAI22x1_ASAP7_75t_L g13922 ( 
.A1(n_13494),
.A2(n_2422),
.B1(n_2420),
.B2(n_2421),
.Y(n_13922)
);

HB1xp67_ASAP7_75t_L g13923 ( 
.A(n_13598),
.Y(n_13923)
);

CKINVDCx8_ASAP7_75t_R g13924 ( 
.A(n_13479),
.Y(n_13924)
);

OAI22xp5_ASAP7_75t_L g13925 ( 
.A1(n_13571),
.A2(n_2425),
.B1(n_2423),
.B2(n_2424),
.Y(n_13925)
);

AOI21xp33_ASAP7_75t_L g13926 ( 
.A1(n_13656),
.A2(n_13684),
.B(n_13661),
.Y(n_13926)
);

AOI221xp5_ASAP7_75t_L g13927 ( 
.A1(n_13729),
.A2(n_2426),
.B1(n_2423),
.B2(n_2424),
.C(n_2427),
.Y(n_13927)
);

OAI22xp33_ASAP7_75t_L g13928 ( 
.A1(n_13711),
.A2(n_13710),
.B1(n_13554),
.B2(n_13553),
.Y(n_13928)
);

AOI22xp33_ASAP7_75t_L g13929 ( 
.A1(n_13634),
.A2(n_2428),
.B1(n_2426),
.B2(n_2427),
.Y(n_13929)
);

OAI22xp5_ASAP7_75t_L g13930 ( 
.A1(n_13577),
.A2(n_2430),
.B1(n_2428),
.B2(n_2429),
.Y(n_13930)
);

A2O1A1Ixp33_ASAP7_75t_L g13931 ( 
.A1(n_13391),
.A2(n_13625),
.B(n_13626),
.C(n_13624),
.Y(n_13931)
);

INVx1_ASAP7_75t_L g13932 ( 
.A(n_13439),
.Y(n_13932)
);

INVx1_ASAP7_75t_L g13933 ( 
.A(n_13445),
.Y(n_13933)
);

HB1xp67_ASAP7_75t_L g13934 ( 
.A(n_13486),
.Y(n_13934)
);

OAI22xp5_ASAP7_75t_L g13935 ( 
.A1(n_13706),
.A2(n_2431),
.B1(n_2429),
.B2(n_2430),
.Y(n_13935)
);

INVx1_ASAP7_75t_L g13936 ( 
.A(n_13450),
.Y(n_13936)
);

AND2x2_ASAP7_75t_L g13937 ( 
.A(n_13463),
.B(n_2431),
.Y(n_13937)
);

AND2x2_ASAP7_75t_L g13938 ( 
.A(n_13465),
.B(n_2432),
.Y(n_13938)
);

INVx1_ASAP7_75t_L g13939 ( 
.A(n_13456),
.Y(n_13939)
);

AOI22xp5_ASAP7_75t_L g13940 ( 
.A1(n_13555),
.A2(n_2435),
.B1(n_2433),
.B2(n_2434),
.Y(n_13940)
);

OR2x2_ASAP7_75t_L g13941 ( 
.A(n_13579),
.B(n_2434),
.Y(n_13941)
);

AOI221xp5_ASAP7_75t_L g13942 ( 
.A1(n_13724),
.A2(n_2439),
.B1(n_2437),
.B2(n_2438),
.C(n_2440),
.Y(n_13942)
);

AOI22xp33_ASAP7_75t_L g13943 ( 
.A1(n_13682),
.A2(n_2439),
.B1(n_2437),
.B2(n_2438),
.Y(n_13943)
);

AOI22xp33_ASAP7_75t_L g13944 ( 
.A1(n_13681),
.A2(n_2442),
.B1(n_2440),
.B2(n_2441),
.Y(n_13944)
);

HB1xp67_ASAP7_75t_L g13945 ( 
.A(n_13471),
.Y(n_13945)
);

OAI22xp33_ASAP7_75t_L g13946 ( 
.A1(n_13582),
.A2(n_2445),
.B1(n_2443),
.B2(n_2444),
.Y(n_13946)
);

AOI22xp33_ASAP7_75t_SL g13947 ( 
.A1(n_13647),
.A2(n_2446),
.B1(n_2443),
.B2(n_2444),
.Y(n_13947)
);

BUFx6f_ASAP7_75t_L g13948 ( 
.A(n_13430),
.Y(n_13948)
);

OAI22xp5_ASAP7_75t_L g13949 ( 
.A1(n_13658),
.A2(n_2448),
.B1(n_2446),
.B2(n_2447),
.Y(n_13949)
);

AOI22xp33_ASAP7_75t_SL g13950 ( 
.A1(n_13646),
.A2(n_2449),
.B1(n_2447),
.B2(n_2448),
.Y(n_13950)
);

AOI22xp33_ASAP7_75t_L g13951 ( 
.A1(n_13715),
.A2(n_2451),
.B1(n_2449),
.B2(n_2450),
.Y(n_13951)
);

OR2x2_ASAP7_75t_L g13952 ( 
.A(n_13699),
.B(n_2450),
.Y(n_13952)
);

AND2x2_ASAP7_75t_L g13953 ( 
.A(n_13596),
.B(n_2451),
.Y(n_13953)
);

OR2x2_ASAP7_75t_L g13954 ( 
.A(n_13591),
.B(n_13639),
.Y(n_13954)
);

AND2x2_ASAP7_75t_L g13955 ( 
.A(n_13607),
.B(n_2452),
.Y(n_13955)
);

OR2x2_ASAP7_75t_L g13956 ( 
.A(n_13648),
.B(n_2452),
.Y(n_13956)
);

BUFx4f_ASAP7_75t_SL g13957 ( 
.A(n_13448),
.Y(n_13957)
);

OAI21x1_ASAP7_75t_L g13958 ( 
.A1(n_13695),
.A2(n_2453),
.B(n_2454),
.Y(n_13958)
);

HB1xp67_ASAP7_75t_L g13959 ( 
.A(n_13609),
.Y(n_13959)
);

AOI221xp5_ASAP7_75t_L g13960 ( 
.A1(n_13725),
.A2(n_13499),
.B1(n_13504),
.B2(n_13560),
.C(n_13557),
.Y(n_13960)
);

INVx2_ASAP7_75t_L g13961 ( 
.A(n_13587),
.Y(n_13961)
);

AOI22xp33_ASAP7_75t_L g13962 ( 
.A1(n_13709),
.A2(n_2456),
.B1(n_2453),
.B2(n_2455),
.Y(n_13962)
);

AOI22xp33_ASAP7_75t_L g13963 ( 
.A1(n_13655),
.A2(n_13685),
.B1(n_13689),
.B2(n_13608),
.Y(n_13963)
);

BUFx2_ASAP7_75t_L g13964 ( 
.A(n_13587),
.Y(n_13964)
);

AND2x2_ASAP7_75t_L g13965 ( 
.A(n_13538),
.B(n_2455),
.Y(n_13965)
);

AOI22xp33_ASAP7_75t_L g13966 ( 
.A1(n_13672),
.A2(n_2458),
.B1(n_2456),
.B2(n_2457),
.Y(n_13966)
);

NAND3xp33_ASAP7_75t_L g13967 ( 
.A(n_13593),
.B(n_2458),
.C(n_2459),
.Y(n_13967)
);

AOI22xp33_ASAP7_75t_L g13968 ( 
.A1(n_13673),
.A2(n_2461),
.B1(n_2459),
.B2(n_2460),
.Y(n_13968)
);

OR2x2_ASAP7_75t_L g13969 ( 
.A(n_13622),
.B(n_2460),
.Y(n_13969)
);

HB1xp67_ASAP7_75t_L g13970 ( 
.A(n_13561),
.Y(n_13970)
);

AOI221xp5_ASAP7_75t_L g13971 ( 
.A1(n_13425),
.A2(n_2464),
.B1(n_2461),
.B2(n_2463),
.C(n_2465),
.Y(n_13971)
);

AND2x2_ASAP7_75t_L g13972 ( 
.A(n_13676),
.B(n_2463),
.Y(n_13972)
);

AOI22xp33_ASAP7_75t_L g13973 ( 
.A1(n_13677),
.A2(n_2467),
.B1(n_2464),
.B2(n_2465),
.Y(n_13973)
);

OA21x2_ASAP7_75t_L g13974 ( 
.A1(n_13529),
.A2(n_2467),
.B(n_2468),
.Y(n_13974)
);

OA21x2_ASAP7_75t_L g13975 ( 
.A1(n_13507),
.A2(n_13550),
.B(n_13548),
.Y(n_13975)
);

AOI22xp33_ASAP7_75t_L g13976 ( 
.A1(n_13540),
.A2(n_2470),
.B1(n_2468),
.B2(n_2469),
.Y(n_13976)
);

OAI22xp33_ASAP7_75t_L g13977 ( 
.A1(n_13590),
.A2(n_2471),
.B1(n_2469),
.B2(n_2470),
.Y(n_13977)
);

OR2x2_ASAP7_75t_L g13978 ( 
.A(n_13497),
.B(n_2472),
.Y(n_13978)
);

OAI22xp33_ASAP7_75t_L g13979 ( 
.A1(n_13623),
.A2(n_2474),
.B1(n_2472),
.B2(n_2473),
.Y(n_13979)
);

AOI221xp5_ASAP7_75t_L g13980 ( 
.A1(n_13630),
.A2(n_2475),
.B1(n_2473),
.B2(n_2474),
.C(n_2476),
.Y(n_13980)
);

OAI22xp33_ASAP7_75t_L g13981 ( 
.A1(n_13563),
.A2(n_2478),
.B1(n_2476),
.B2(n_2477),
.Y(n_13981)
);

OAI22xp33_ASAP7_75t_L g13982 ( 
.A1(n_13600),
.A2(n_2481),
.B1(n_2479),
.B2(n_2480),
.Y(n_13982)
);

AND2x4_ASAP7_75t_L g13983 ( 
.A(n_13485),
.B(n_13460),
.Y(n_13983)
);

HB1xp67_ASAP7_75t_L g13984 ( 
.A(n_13546),
.Y(n_13984)
);

AND2x4_ASAP7_75t_L g13985 ( 
.A(n_13474),
.B(n_2479),
.Y(n_13985)
);

INVx3_ASAP7_75t_L g13986 ( 
.A(n_13679),
.Y(n_13986)
);

OAI22xp33_ASAP7_75t_L g13987 ( 
.A1(n_13601),
.A2(n_2483),
.B1(n_2480),
.B2(n_2482),
.Y(n_13987)
);

AND2x2_ASAP7_75t_L g13988 ( 
.A(n_13665),
.B(n_2482),
.Y(n_13988)
);

AOI22xp33_ASAP7_75t_L g13989 ( 
.A1(n_13568),
.A2(n_2486),
.B1(n_2484),
.B2(n_2485),
.Y(n_13989)
);

AOI22xp5_ASAP7_75t_L g13990 ( 
.A1(n_13551),
.A2(n_2486),
.B1(n_2484),
.B2(n_2485),
.Y(n_13990)
);

OAI22xp5_ASAP7_75t_L g13991 ( 
.A1(n_13510),
.A2(n_2489),
.B1(n_2487),
.B2(n_2488),
.Y(n_13991)
);

AOI21xp5_ASAP7_75t_L g13992 ( 
.A1(n_13584),
.A2(n_13594),
.B(n_13559),
.Y(n_13992)
);

NAND2xp5_ASAP7_75t_L g13993 ( 
.A(n_13628),
.B(n_2487),
.Y(n_13993)
);

AOI222xp33_ASAP7_75t_L g13994 ( 
.A1(n_13640),
.A2(n_2490),
.B1(n_2492),
.B2(n_2488),
.C1(n_2489),
.C2(n_2491),
.Y(n_13994)
);

A2O1A1Ixp33_ASAP7_75t_L g13995 ( 
.A1(n_13736),
.A2(n_2492),
.B(n_2490),
.C(n_2491),
.Y(n_13995)
);

NAND3xp33_ASAP7_75t_L g13996 ( 
.A(n_13605),
.B(n_2493),
.C(n_2494),
.Y(n_13996)
);

AOI221xp5_ASAP7_75t_L g13997 ( 
.A1(n_13606),
.A2(n_2496),
.B1(n_2493),
.B2(n_2495),
.C(n_2497),
.Y(n_13997)
);

AO31x2_ASAP7_75t_L g13998 ( 
.A1(n_13482),
.A2(n_2497),
.A3(n_2495),
.B(n_2496),
.Y(n_13998)
);

INVx1_ASAP7_75t_L g13999 ( 
.A(n_13457),
.Y(n_13999)
);

INVx2_ASAP7_75t_SL g14000 ( 
.A(n_13756),
.Y(n_14000)
);

NOR2xp67_ASAP7_75t_L g14001 ( 
.A(n_13832),
.B(n_13602),
.Y(n_14001)
);

HB1xp67_ASAP7_75t_L g14002 ( 
.A(n_13794),
.Y(n_14002)
);

AND2x2_ASAP7_75t_L g14003 ( 
.A(n_13801),
.B(n_13443),
.Y(n_14003)
);

HB1xp67_ASAP7_75t_L g14004 ( 
.A(n_13760),
.Y(n_14004)
);

OR2x2_ASAP7_75t_L g14005 ( 
.A(n_13761),
.B(n_13502),
.Y(n_14005)
);

BUFx3_ASAP7_75t_L g14006 ( 
.A(n_13756),
.Y(n_14006)
);

OR2x2_ASAP7_75t_L g14007 ( 
.A(n_13859),
.B(n_13528),
.Y(n_14007)
);

OR2x2_ASAP7_75t_L g14008 ( 
.A(n_13762),
.B(n_13797),
.Y(n_14008)
);

AND2x4_ASAP7_75t_L g14009 ( 
.A(n_13886),
.B(n_13530),
.Y(n_14009)
);

AND2x2_ASAP7_75t_L g14010 ( 
.A(n_13847),
.B(n_13613),
.Y(n_14010)
);

INVx2_ASAP7_75t_L g14011 ( 
.A(n_13777),
.Y(n_14011)
);

INVx1_ASAP7_75t_L g14012 ( 
.A(n_13742),
.Y(n_14012)
);

INVx2_ASAP7_75t_L g14013 ( 
.A(n_13789),
.Y(n_14013)
);

AND2x2_ASAP7_75t_L g14014 ( 
.A(n_13889),
.B(n_13574),
.Y(n_14014)
);

AND2x2_ASAP7_75t_L g14015 ( 
.A(n_13791),
.B(n_13627),
.Y(n_14015)
);

INVx1_ASAP7_75t_L g14016 ( 
.A(n_13959),
.Y(n_14016)
);

OR2x2_ASAP7_75t_L g14017 ( 
.A(n_13923),
.B(n_13749),
.Y(n_14017)
);

INVx2_ASAP7_75t_L g14018 ( 
.A(n_13901),
.Y(n_14018)
);

INVx1_ASAP7_75t_L g14019 ( 
.A(n_13970),
.Y(n_14019)
);

INVx1_ASAP7_75t_L g14020 ( 
.A(n_13772),
.Y(n_14020)
);

AOI22xp33_ASAP7_75t_L g14021 ( 
.A1(n_13783),
.A2(n_13597),
.B1(n_13619),
.B2(n_13615),
.Y(n_14021)
);

INVx1_ASAP7_75t_L g14022 ( 
.A(n_13984),
.Y(n_14022)
);

HB1xp67_ASAP7_75t_L g14023 ( 
.A(n_13948),
.Y(n_14023)
);

CKINVDCx16_ASAP7_75t_R g14024 ( 
.A(n_13913),
.Y(n_14024)
);

INVx1_ASAP7_75t_L g14025 ( 
.A(n_13978),
.Y(n_14025)
);

INVx2_ASAP7_75t_L g14026 ( 
.A(n_13818),
.Y(n_14026)
);

NOR2xp67_ASAP7_75t_L g14027 ( 
.A(n_13752),
.B(n_13604),
.Y(n_14027)
);

INVxp67_ASAP7_75t_L g14028 ( 
.A(n_13748),
.Y(n_14028)
);

HB1xp67_ASAP7_75t_L g14029 ( 
.A(n_13948),
.Y(n_14029)
);

BUFx3_ASAP7_75t_L g14030 ( 
.A(n_13780),
.Y(n_14030)
);

HB1xp67_ASAP7_75t_L g14031 ( 
.A(n_13924),
.Y(n_14031)
);

INVx1_ASAP7_75t_L g14032 ( 
.A(n_13975),
.Y(n_14032)
);

AND2x2_ASAP7_75t_L g14033 ( 
.A(n_13845),
.B(n_13659),
.Y(n_14033)
);

HB1xp67_ASAP7_75t_L g14034 ( 
.A(n_13934),
.Y(n_14034)
);

BUFx6f_ASAP7_75t_L g14035 ( 
.A(n_13874),
.Y(n_14035)
);

BUFx6f_ASAP7_75t_L g14036 ( 
.A(n_13784),
.Y(n_14036)
);

AND2x2_ASAP7_75t_L g14037 ( 
.A(n_13802),
.B(n_13576),
.Y(n_14037)
);

INVx2_ASAP7_75t_L g14038 ( 
.A(n_13911),
.Y(n_14038)
);

INVx2_ASAP7_75t_L g14039 ( 
.A(n_13839),
.Y(n_14039)
);

HB1xp67_ASAP7_75t_L g14040 ( 
.A(n_13945),
.Y(n_14040)
);

INVx1_ASAP7_75t_L g14041 ( 
.A(n_13975),
.Y(n_14041)
);

AND2x2_ASAP7_75t_L g14042 ( 
.A(n_13964),
.B(n_13535),
.Y(n_14042)
);

HB1xp67_ASAP7_75t_L g14043 ( 
.A(n_13860),
.Y(n_14043)
);

AND2x2_ASAP7_75t_L g14044 ( 
.A(n_13849),
.B(n_13484),
.Y(n_14044)
);

INVx1_ASAP7_75t_SL g14045 ( 
.A(n_13743),
.Y(n_14045)
);

AND2x4_ASAP7_75t_L g14046 ( 
.A(n_13743),
.B(n_13536),
.Y(n_14046)
);

INVx2_ASAP7_75t_SL g14047 ( 
.A(n_13916),
.Y(n_14047)
);

INVx2_ASAP7_75t_L g14048 ( 
.A(n_13986),
.Y(n_14048)
);

INVx2_ASAP7_75t_L g14049 ( 
.A(n_13909),
.Y(n_14049)
);

NOR2x1_ASAP7_75t_SL g14050 ( 
.A(n_13840),
.B(n_13564),
.Y(n_14050)
);

INVx3_ASAP7_75t_L g14051 ( 
.A(n_13787),
.Y(n_14051)
);

AND2x2_ASAP7_75t_L g14052 ( 
.A(n_13873),
.B(n_13572),
.Y(n_14052)
);

AND2x2_ASAP7_75t_L g14053 ( 
.A(n_13983),
.B(n_13566),
.Y(n_14053)
);

NOR2x1p5_ASAP7_75t_L g14054 ( 
.A(n_13891),
.B(n_13635),
.Y(n_14054)
);

AND2x2_ASAP7_75t_L g14055 ( 
.A(n_13883),
.B(n_13526),
.Y(n_14055)
);

AND2x2_ASAP7_75t_L g14056 ( 
.A(n_13918),
.B(n_13961),
.Y(n_14056)
);

INVx2_ASAP7_75t_L g14057 ( 
.A(n_13957),
.Y(n_14057)
);

HB1xp67_ASAP7_75t_L g14058 ( 
.A(n_13860),
.Y(n_14058)
);

AND2x2_ASAP7_75t_L g14059 ( 
.A(n_13776),
.B(n_13527),
.Y(n_14059)
);

OR2x2_ASAP7_75t_L g14060 ( 
.A(n_13954),
.B(n_13514),
.Y(n_14060)
);

INVx1_ASAP7_75t_L g14061 ( 
.A(n_13941),
.Y(n_14061)
);

CKINVDCx20_ASAP7_75t_R g14062 ( 
.A(n_13880),
.Y(n_14062)
);

AND2x4_ASAP7_75t_L g14063 ( 
.A(n_13816),
.B(n_13501),
.Y(n_14063)
);

NAND2xp5_ASAP7_75t_L g14064 ( 
.A(n_13741),
.B(n_13719),
.Y(n_14064)
);

INVx1_ASAP7_75t_L g14065 ( 
.A(n_13819),
.Y(n_14065)
);

NAND3xp33_ASAP7_75t_L g14066 ( 
.A(n_13767),
.B(n_13531),
.C(n_13522),
.Y(n_14066)
);

AOI22xp33_ASAP7_75t_L g14067 ( 
.A1(n_13747),
.A2(n_13498),
.B1(n_13511),
.B2(n_13492),
.Y(n_14067)
);

OR2x2_ASAP7_75t_L g14068 ( 
.A(n_13892),
.B(n_13394),
.Y(n_14068)
);

INVx2_ASAP7_75t_L g14069 ( 
.A(n_13856),
.Y(n_14069)
);

BUFx2_ASAP7_75t_L g14070 ( 
.A(n_13771),
.Y(n_14070)
);

NOR2xp33_ASAP7_75t_L g14071 ( 
.A(n_13753),
.B(n_13475),
.Y(n_14071)
);

INVx2_ASAP7_75t_L g14072 ( 
.A(n_13755),
.Y(n_14072)
);

INVxp67_ASAP7_75t_SL g14073 ( 
.A(n_13763),
.Y(n_14073)
);

AND2x2_ASAP7_75t_L g14074 ( 
.A(n_13751),
.B(n_13963),
.Y(n_14074)
);

AND2x2_ASAP7_75t_L g14075 ( 
.A(n_13786),
.B(n_13632),
.Y(n_14075)
);

AND2x2_ASAP7_75t_L g14076 ( 
.A(n_13841),
.B(n_13633),
.Y(n_14076)
);

INVx1_ASAP7_75t_L g14077 ( 
.A(n_13826),
.Y(n_14077)
);

INVx1_ASAP7_75t_L g14078 ( 
.A(n_13830),
.Y(n_14078)
);

INVx2_ASAP7_75t_L g14079 ( 
.A(n_13766),
.Y(n_14079)
);

BUFx6f_ASAP7_75t_L g14080 ( 
.A(n_13893),
.Y(n_14080)
);

AND2x2_ASAP7_75t_L g14081 ( 
.A(n_13870),
.B(n_13565),
.Y(n_14081)
);

INVx2_ASAP7_75t_L g14082 ( 
.A(n_13906),
.Y(n_14082)
);

INVx2_ASAP7_75t_L g14083 ( 
.A(n_13898),
.Y(n_14083)
);

AND2x2_ASAP7_75t_L g14084 ( 
.A(n_13840),
.B(n_13988),
.Y(n_14084)
);

AOI22xp33_ASAP7_75t_SL g14085 ( 
.A1(n_13746),
.A2(n_13713),
.B1(n_13712),
.B2(n_13617),
.Y(n_14085)
);

INVx2_ASAP7_75t_L g14086 ( 
.A(n_13773),
.Y(n_14086)
);

AND2x2_ASAP7_75t_L g14087 ( 
.A(n_13931),
.B(n_13668),
.Y(n_14087)
);

BUFx3_ASAP7_75t_L g14088 ( 
.A(n_13985),
.Y(n_14088)
);

INVx1_ASAP7_75t_L g14089 ( 
.A(n_13831),
.Y(n_14089)
);

INVx1_ASAP7_75t_L g14090 ( 
.A(n_13833),
.Y(n_14090)
);

AND2x4_ASAP7_75t_L g14091 ( 
.A(n_13829),
.B(n_13509),
.Y(n_14091)
);

NAND2xp5_ASAP7_75t_L g14092 ( 
.A(n_13808),
.B(n_13461),
.Y(n_14092)
);

INVx1_ASAP7_75t_L g14093 ( 
.A(n_13843),
.Y(n_14093)
);

INVx1_ASAP7_75t_L g14094 ( 
.A(n_13852),
.Y(n_14094)
);

INVx2_ASAP7_75t_SL g14095 ( 
.A(n_13825),
.Y(n_14095)
);

INVx1_ASAP7_75t_L g14096 ( 
.A(n_13865),
.Y(n_14096)
);

INVx1_ASAP7_75t_L g14097 ( 
.A(n_13877),
.Y(n_14097)
);

INVx1_ASAP7_75t_L g14098 ( 
.A(n_13881),
.Y(n_14098)
);

INVx3_ASAP7_75t_L g14099 ( 
.A(n_13914),
.Y(n_14099)
);

INVx1_ASAP7_75t_L g14100 ( 
.A(n_13932),
.Y(n_14100)
);

INVx2_ASAP7_75t_L g14101 ( 
.A(n_13855),
.Y(n_14101)
);

INVx2_ASAP7_75t_L g14102 ( 
.A(n_13953),
.Y(n_14102)
);

BUFx2_ASAP7_75t_L g14103 ( 
.A(n_13903),
.Y(n_14103)
);

INVx1_ASAP7_75t_L g14104 ( 
.A(n_13933),
.Y(n_14104)
);

AND2x2_ASAP7_75t_L g14105 ( 
.A(n_13965),
.B(n_13393),
.Y(n_14105)
);

INVx2_ASAP7_75t_L g14106 ( 
.A(n_13955),
.Y(n_14106)
);

BUFx6f_ASAP7_75t_L g14107 ( 
.A(n_13937),
.Y(n_14107)
);

INVx1_ASAP7_75t_L g14108 ( 
.A(n_13936),
.Y(n_14108)
);

INVx1_ASAP7_75t_L g14109 ( 
.A(n_13939),
.Y(n_14109)
);

INVx1_ASAP7_75t_L g14110 ( 
.A(n_13999),
.Y(n_14110)
);

INVx1_ASAP7_75t_L g14111 ( 
.A(n_13972),
.Y(n_14111)
);

AND2x2_ASAP7_75t_L g14112 ( 
.A(n_13938),
.B(n_13495),
.Y(n_14112)
);

INVx4_ASAP7_75t_L g14113 ( 
.A(n_13952),
.Y(n_14113)
);

AND2x2_ASAP7_75t_L g14114 ( 
.A(n_13807),
.B(n_13958),
.Y(n_14114)
);

AND2x2_ASAP7_75t_L g14115 ( 
.A(n_13917),
.B(n_13466),
.Y(n_14115)
);

INVx2_ASAP7_75t_L g14116 ( 
.A(n_13998),
.Y(n_14116)
);

HB1xp67_ASAP7_75t_L g14117 ( 
.A(n_13974),
.Y(n_14117)
);

INVx1_ASAP7_75t_L g14118 ( 
.A(n_13814),
.Y(n_14118)
);

INVx1_ASAP7_75t_L g14119 ( 
.A(n_13815),
.Y(n_14119)
);

AND2x4_ASAP7_75t_L g14120 ( 
.A(n_13910),
.B(n_13650),
.Y(n_14120)
);

AND2x4_ASAP7_75t_L g14121 ( 
.A(n_13887),
.B(n_13468),
.Y(n_14121)
);

HB1xp67_ASAP7_75t_L g14122 ( 
.A(n_13974),
.Y(n_14122)
);

INVx1_ASAP7_75t_L g14123 ( 
.A(n_13792),
.Y(n_14123)
);

BUFx3_ASAP7_75t_L g14124 ( 
.A(n_13922),
.Y(n_14124)
);

AOI22xp33_ASAP7_75t_L g14125 ( 
.A1(n_13750),
.A2(n_13481),
.B1(n_13487),
.B2(n_13480),
.Y(n_14125)
);

HB1xp67_ASAP7_75t_L g14126 ( 
.A(n_13835),
.Y(n_14126)
);

INVx2_ASAP7_75t_L g14127 ( 
.A(n_13998),
.Y(n_14127)
);

INVx2_ASAP7_75t_L g14128 ( 
.A(n_13835),
.Y(n_14128)
);

INVx2_ASAP7_75t_L g14129 ( 
.A(n_13882),
.Y(n_14129)
);

OR2x2_ASAP7_75t_L g14130 ( 
.A(n_13904),
.B(n_13489),
.Y(n_14130)
);

INVx1_ASAP7_75t_L g14131 ( 
.A(n_13956),
.Y(n_14131)
);

BUFx2_ASAP7_75t_L g14132 ( 
.A(n_13969),
.Y(n_14132)
);

INVx2_ASAP7_75t_L g14133 ( 
.A(n_13921),
.Y(n_14133)
);

INVx2_ASAP7_75t_L g14134 ( 
.A(n_13921),
.Y(n_14134)
);

AOI21xp33_ASAP7_75t_L g14135 ( 
.A1(n_13928),
.A2(n_13674),
.B(n_13442),
.Y(n_14135)
);

NAND2xp5_ASAP7_75t_L g14136 ( 
.A(n_13861),
.B(n_13652),
.Y(n_14136)
);

AND2x2_ASAP7_75t_L g14137 ( 
.A(n_13992),
.B(n_13612),
.Y(n_14137)
);

INVx1_ASAP7_75t_L g14138 ( 
.A(n_13864),
.Y(n_14138)
);

OR2x2_ASAP7_75t_L g14139 ( 
.A(n_13993),
.B(n_13406),
.Y(n_14139)
);

INVx2_ASAP7_75t_L g14140 ( 
.A(n_13822),
.Y(n_14140)
);

OR2x2_ASAP7_75t_L g14141 ( 
.A(n_13902),
.B(n_13406),
.Y(n_14141)
);

OR2x2_ASAP7_75t_L g14142 ( 
.A(n_13803),
.B(n_13595),
.Y(n_14142)
);

AOI22xp33_ASAP7_75t_SL g14143 ( 
.A1(n_13798),
.A2(n_13533),
.B1(n_2500),
.B2(n_2498),
.Y(n_14143)
);

INVx1_ASAP7_75t_L g14144 ( 
.A(n_13795),
.Y(n_14144)
);

INVx2_ASAP7_75t_L g14145 ( 
.A(n_13868),
.Y(n_14145)
);

AND2x2_ASAP7_75t_L g14146 ( 
.A(n_13817),
.B(n_2498),
.Y(n_14146)
);

INVx1_ASAP7_75t_L g14147 ( 
.A(n_13967),
.Y(n_14147)
);

AND2x2_ASAP7_75t_L g14148 ( 
.A(n_13828),
.B(n_2499),
.Y(n_14148)
);

INVx3_ASAP7_75t_L g14149 ( 
.A(n_13866),
.Y(n_14149)
);

AND2x4_ASAP7_75t_L g14150 ( 
.A(n_13850),
.B(n_2499),
.Y(n_14150)
);

AND2x2_ASAP7_75t_L g14151 ( 
.A(n_13854),
.B(n_2500),
.Y(n_14151)
);

INVx1_ASAP7_75t_L g14152 ( 
.A(n_13996),
.Y(n_14152)
);

INVx2_ASAP7_75t_L g14153 ( 
.A(n_13990),
.Y(n_14153)
);

AND2x4_ASAP7_75t_SL g14154 ( 
.A(n_13823),
.B(n_2501),
.Y(n_14154)
);

AND2x2_ASAP7_75t_L g14155 ( 
.A(n_13897),
.B(n_2501),
.Y(n_14155)
);

BUFx6f_ASAP7_75t_SL g14156 ( 
.A(n_13919),
.Y(n_14156)
);

AND2x2_ASAP7_75t_L g14157 ( 
.A(n_13770),
.B(n_2502),
.Y(n_14157)
);

INVx1_ASAP7_75t_L g14158 ( 
.A(n_13754),
.Y(n_14158)
);

HB1xp67_ASAP7_75t_L g14159 ( 
.A(n_13812),
.Y(n_14159)
);

NAND2xp5_ASAP7_75t_L g14160 ( 
.A(n_13744),
.B(n_2503),
.Y(n_14160)
);

NAND2xp5_ASAP7_75t_L g14161 ( 
.A(n_13915),
.B(n_2503),
.Y(n_14161)
);

INVx1_ASAP7_75t_L g14162 ( 
.A(n_13782),
.Y(n_14162)
);

BUFx3_ASAP7_75t_L g14163 ( 
.A(n_13836),
.Y(n_14163)
);

INVx2_ASAP7_75t_L g14164 ( 
.A(n_13900),
.Y(n_14164)
);

INVx1_ASAP7_75t_L g14165 ( 
.A(n_13804),
.Y(n_14165)
);

AND2x2_ASAP7_75t_L g14166 ( 
.A(n_13779),
.B(n_2504),
.Y(n_14166)
);

NOR2x1_ASAP7_75t_L g14167 ( 
.A(n_13878),
.B(n_2504),
.Y(n_14167)
);

INVxp67_ASAP7_75t_L g14168 ( 
.A(n_13788),
.Y(n_14168)
);

OR2x2_ASAP7_75t_L g14169 ( 
.A(n_13926),
.B(n_2505),
.Y(n_14169)
);

INVx1_ASAP7_75t_L g14170 ( 
.A(n_13949),
.Y(n_14170)
);

INVxp67_ASAP7_75t_L g14171 ( 
.A(n_13809),
.Y(n_14171)
);

INVxp67_ASAP7_75t_SL g14172 ( 
.A(n_13774),
.Y(n_14172)
);

INVx1_ASAP7_75t_L g14173 ( 
.A(n_13896),
.Y(n_14173)
);

CKINVDCx5p33_ASAP7_75t_R g14174 ( 
.A(n_13842),
.Y(n_14174)
);

INVx1_ASAP7_75t_L g14175 ( 
.A(n_13991),
.Y(n_14175)
);

INVx1_ASAP7_75t_L g14176 ( 
.A(n_13920),
.Y(n_14176)
);

INVx1_ASAP7_75t_L g14177 ( 
.A(n_13925),
.Y(n_14177)
);

INVx2_ASAP7_75t_L g14178 ( 
.A(n_13884),
.Y(n_14178)
);

INVx2_ASAP7_75t_L g14179 ( 
.A(n_13935),
.Y(n_14179)
);

AND2x2_ASAP7_75t_L g14180 ( 
.A(n_13947),
.B(n_2505),
.Y(n_14180)
);

INVx2_ASAP7_75t_L g14181 ( 
.A(n_13857),
.Y(n_14181)
);

AND2x2_ASAP7_75t_L g14182 ( 
.A(n_13960),
.B(n_2506),
.Y(n_14182)
);

INVx2_ASAP7_75t_L g14183 ( 
.A(n_13930),
.Y(n_14183)
);

BUFx8_ASAP7_75t_L g14184 ( 
.A(n_13908),
.Y(n_14184)
);

AND2x2_ASAP7_75t_L g14185 ( 
.A(n_13793),
.B(n_2506),
.Y(n_14185)
);

AND2x2_ASAP7_75t_L g14186 ( 
.A(n_13950),
.B(n_2507),
.Y(n_14186)
);

INVx2_ASAP7_75t_L g14187 ( 
.A(n_13894),
.Y(n_14187)
);

NOR2x1_ASAP7_75t_L g14188 ( 
.A(n_13775),
.B(n_2507),
.Y(n_14188)
);

OAI22xp5_ASAP7_75t_L g14189 ( 
.A1(n_13745),
.A2(n_2510),
.B1(n_2508),
.B2(n_2509),
.Y(n_14189)
);

INVx2_ASAP7_75t_L g14190 ( 
.A(n_13848),
.Y(n_14190)
);

INVx1_ASAP7_75t_L g14191 ( 
.A(n_13895),
.Y(n_14191)
);

INVx1_ASAP7_75t_L g14192 ( 
.A(n_13905),
.Y(n_14192)
);

INVx2_ASAP7_75t_L g14193 ( 
.A(n_13858),
.Y(n_14193)
);

BUFx6f_ASAP7_75t_L g14194 ( 
.A(n_13768),
.Y(n_14194)
);

INVx2_ASAP7_75t_L g14195 ( 
.A(n_13821),
.Y(n_14195)
);

OR2x2_ASAP7_75t_L g14196 ( 
.A(n_13912),
.B(n_2509),
.Y(n_14196)
);

INVx2_ASAP7_75t_L g14197 ( 
.A(n_13757),
.Y(n_14197)
);

NAND2xp5_ASAP7_75t_L g14198 ( 
.A(n_13876),
.B(n_2510),
.Y(n_14198)
);

INVx2_ASAP7_75t_L g14199 ( 
.A(n_13940),
.Y(n_14199)
);

AND2x2_ASAP7_75t_L g14200 ( 
.A(n_13846),
.B(n_2511),
.Y(n_14200)
);

INVx2_ASAP7_75t_L g14201 ( 
.A(n_13805),
.Y(n_14201)
);

BUFx6f_ASAP7_75t_L g14202 ( 
.A(n_13862),
.Y(n_14202)
);

INVx1_ASAP7_75t_L g14203 ( 
.A(n_14002),
.Y(n_14203)
);

AND2x2_ASAP7_75t_L g14204 ( 
.A(n_14045),
.B(n_13810),
.Y(n_14204)
);

INVx2_ASAP7_75t_L g14205 ( 
.A(n_14006),
.Y(n_14205)
);

INVx2_ASAP7_75t_L g14206 ( 
.A(n_14046),
.Y(n_14206)
);

NAND2xp5_ASAP7_75t_L g14207 ( 
.A(n_14024),
.B(n_13758),
.Y(n_14207)
);

AND2x2_ASAP7_75t_L g14208 ( 
.A(n_14018),
.B(n_13799),
.Y(n_14208)
);

INVxp67_ASAP7_75t_L g14209 ( 
.A(n_14043),
.Y(n_14209)
);

INVx1_ASAP7_75t_L g14210 ( 
.A(n_14004),
.Y(n_14210)
);

INVxp67_ASAP7_75t_SL g14211 ( 
.A(n_14058),
.Y(n_14211)
);

INVx1_ASAP7_75t_L g14212 ( 
.A(n_14032),
.Y(n_14212)
);

HB1xp67_ASAP7_75t_L g14213 ( 
.A(n_14027),
.Y(n_14213)
);

INVx1_ASAP7_75t_L g14214 ( 
.A(n_14041),
.Y(n_14214)
);

INVx1_ASAP7_75t_L g14215 ( 
.A(n_14040),
.Y(n_14215)
);

INVx2_ASAP7_75t_L g14216 ( 
.A(n_14035),
.Y(n_14216)
);

BUFx3_ASAP7_75t_L g14217 ( 
.A(n_14035),
.Y(n_14217)
);

INVx2_ASAP7_75t_L g14218 ( 
.A(n_14000),
.Y(n_14218)
);

INVx1_ASAP7_75t_L g14219 ( 
.A(n_14034),
.Y(n_14219)
);

INVx2_ASAP7_75t_L g14220 ( 
.A(n_14036),
.Y(n_14220)
);

INVx2_ASAP7_75t_L g14221 ( 
.A(n_14036),
.Y(n_14221)
);

INVx1_ASAP7_75t_L g14222 ( 
.A(n_14012),
.Y(n_14222)
);

OR2x2_ASAP7_75t_L g14223 ( 
.A(n_14017),
.B(n_13759),
.Y(n_14223)
);

AND2x2_ASAP7_75t_L g14224 ( 
.A(n_14003),
.B(n_13844),
.Y(n_14224)
);

INVx1_ASAP7_75t_L g14225 ( 
.A(n_14008),
.Y(n_14225)
);

INVx2_ASAP7_75t_L g14226 ( 
.A(n_14026),
.Y(n_14226)
);

INVx1_ASAP7_75t_L g14227 ( 
.A(n_14016),
.Y(n_14227)
);

INVx1_ASAP7_75t_L g14228 ( 
.A(n_14019),
.Y(n_14228)
);

AND2x2_ASAP7_75t_L g14229 ( 
.A(n_14031),
.B(n_13813),
.Y(n_14229)
);

INVx2_ASAP7_75t_L g14230 ( 
.A(n_14030),
.Y(n_14230)
);

OAI22xp5_ASAP7_75t_L g14231 ( 
.A1(n_14143),
.A2(n_13781),
.B1(n_13769),
.B2(n_13976),
.Y(n_14231)
);

OR2x2_ASAP7_75t_L g14232 ( 
.A(n_14070),
.B(n_13863),
.Y(n_14232)
);

NAND2xp5_ASAP7_75t_L g14233 ( 
.A(n_14047),
.B(n_13800),
.Y(n_14233)
);

INVx1_ASAP7_75t_L g14234 ( 
.A(n_14022),
.Y(n_14234)
);

NAND2xp5_ASAP7_75t_L g14235 ( 
.A(n_14124),
.B(n_13875),
.Y(n_14235)
);

NAND2xp5_ASAP7_75t_L g14236 ( 
.A(n_14149),
.B(n_13820),
.Y(n_14236)
);

INVx1_ASAP7_75t_L g14237 ( 
.A(n_14132),
.Y(n_14237)
);

INVx2_ASAP7_75t_L g14238 ( 
.A(n_14051),
.Y(n_14238)
);

NOR2x1_ASAP7_75t_L g14239 ( 
.A(n_14062),
.B(n_13946),
.Y(n_14239)
);

BUFx3_ASAP7_75t_L g14240 ( 
.A(n_14080),
.Y(n_14240)
);

AND2x2_ASAP7_75t_L g14241 ( 
.A(n_14049),
.B(n_13827),
.Y(n_14241)
);

INVx2_ASAP7_75t_L g14242 ( 
.A(n_14080),
.Y(n_14242)
);

NAND2xp5_ASAP7_75t_L g14243 ( 
.A(n_14073),
.B(n_13971),
.Y(n_14243)
);

NAND2xp5_ASAP7_75t_L g14244 ( 
.A(n_14075),
.B(n_13977),
.Y(n_14244)
);

AND2x2_ASAP7_75t_L g14245 ( 
.A(n_14057),
.B(n_13851),
.Y(n_14245)
);

OR2x2_ASAP7_75t_L g14246 ( 
.A(n_14191),
.B(n_13979),
.Y(n_14246)
);

INVx2_ASAP7_75t_L g14247 ( 
.A(n_14009),
.Y(n_14247)
);

AND2x2_ASAP7_75t_L g14248 ( 
.A(n_14084),
.B(n_13995),
.Y(n_14248)
);

OAI22xp5_ASAP7_75t_L g14249 ( 
.A1(n_14156),
.A2(n_13989),
.B1(n_13837),
.B2(n_13838),
.Y(n_14249)
);

NAND2xp5_ASAP7_75t_L g14250 ( 
.A(n_14157),
.B(n_13981),
.Y(n_14250)
);

AND2x2_ASAP7_75t_L g14251 ( 
.A(n_14076),
.B(n_14042),
.Y(n_14251)
);

AND2x2_ASAP7_75t_L g14252 ( 
.A(n_14014),
.B(n_13765),
.Y(n_14252)
);

AND2x2_ASAP7_75t_L g14253 ( 
.A(n_14011),
.B(n_13790),
.Y(n_14253)
);

INVx1_ASAP7_75t_L g14254 ( 
.A(n_14129),
.Y(n_14254)
);

AND2x2_ASAP7_75t_L g14255 ( 
.A(n_14013),
.B(n_13764),
.Y(n_14255)
);

NAND2xp5_ASAP7_75t_L g14256 ( 
.A(n_14167),
.B(n_13982),
.Y(n_14256)
);

INVx2_ASAP7_75t_L g14257 ( 
.A(n_14088),
.Y(n_14257)
);

INVx1_ASAP7_75t_L g14258 ( 
.A(n_14126),
.Y(n_14258)
);

AND2x2_ASAP7_75t_L g14259 ( 
.A(n_14081),
.B(n_13885),
.Y(n_14259)
);

INVx1_ASAP7_75t_L g14260 ( 
.A(n_14117),
.Y(n_14260)
);

INVx2_ASAP7_75t_L g14261 ( 
.A(n_14107),
.Y(n_14261)
);

AND2x2_ASAP7_75t_L g14262 ( 
.A(n_14105),
.B(n_13778),
.Y(n_14262)
);

HB1xp67_ASAP7_75t_L g14263 ( 
.A(n_14023),
.Y(n_14263)
);

OR2x2_ASAP7_75t_L g14264 ( 
.A(n_14192),
.B(n_13987),
.Y(n_14264)
);

OR2x2_ASAP7_75t_L g14265 ( 
.A(n_14113),
.B(n_13907),
.Y(n_14265)
);

AND2x2_ASAP7_75t_L g14266 ( 
.A(n_14010),
.B(n_13879),
.Y(n_14266)
);

OR2x2_ASAP7_75t_L g14267 ( 
.A(n_14005),
.B(n_13834),
.Y(n_14267)
);

INVx3_ASAP7_75t_L g14268 ( 
.A(n_14107),
.Y(n_14268)
);

NAND2xp5_ASAP7_75t_L g14269 ( 
.A(n_14184),
.B(n_13785),
.Y(n_14269)
);

AND2x2_ASAP7_75t_L g14270 ( 
.A(n_14053),
.B(n_13869),
.Y(n_14270)
);

BUFx2_ASAP7_75t_L g14271 ( 
.A(n_14029),
.Y(n_14271)
);

AOI22xp33_ASAP7_75t_L g14272 ( 
.A1(n_14202),
.A2(n_14163),
.B1(n_14194),
.B2(n_14172),
.Y(n_14272)
);

AND2x2_ASAP7_75t_L g14273 ( 
.A(n_14015),
.B(n_13824),
.Y(n_14273)
);

INVx1_ASAP7_75t_L g14274 ( 
.A(n_14122),
.Y(n_14274)
);

INVx2_ASAP7_75t_L g14275 ( 
.A(n_14038),
.Y(n_14275)
);

INVx2_ASAP7_75t_L g14276 ( 
.A(n_14048),
.Y(n_14276)
);

INVxp67_ASAP7_75t_SL g14277 ( 
.A(n_14050),
.Y(n_14277)
);

INVx1_ASAP7_75t_L g14278 ( 
.A(n_14111),
.Y(n_14278)
);

AND2x2_ASAP7_75t_L g14279 ( 
.A(n_14028),
.B(n_13796),
.Y(n_14279)
);

NAND2xp5_ASAP7_75t_L g14280 ( 
.A(n_14071),
.B(n_13806),
.Y(n_14280)
);

AND2x2_ASAP7_75t_L g14281 ( 
.A(n_14074),
.B(n_13951),
.Y(n_14281)
);

OR2x2_ASAP7_75t_L g14282 ( 
.A(n_14158),
.B(n_13890),
.Y(n_14282)
);

OR2x2_ASAP7_75t_L g14283 ( 
.A(n_14060),
.B(n_13872),
.Y(n_14283)
);

INVx1_ASAP7_75t_L g14284 ( 
.A(n_14061),
.Y(n_14284)
);

NAND2xp5_ASAP7_75t_L g14285 ( 
.A(n_14171),
.B(n_13927),
.Y(n_14285)
);

NAND2xp5_ASAP7_75t_L g14286 ( 
.A(n_14194),
.B(n_13942),
.Y(n_14286)
);

NOR2x1_ASAP7_75t_L g14287 ( 
.A(n_14103),
.B(n_13811),
.Y(n_14287)
);

INVx2_ASAP7_75t_L g14288 ( 
.A(n_14099),
.Y(n_14288)
);

OR2x2_ASAP7_75t_L g14289 ( 
.A(n_14068),
.B(n_13929),
.Y(n_14289)
);

INVx2_ASAP7_75t_L g14290 ( 
.A(n_14044),
.Y(n_14290)
);

BUFx3_ASAP7_75t_L g14291 ( 
.A(n_14063),
.Y(n_14291)
);

INVx1_ASAP7_75t_L g14292 ( 
.A(n_14123),
.Y(n_14292)
);

AOI22xp33_ASAP7_75t_L g14293 ( 
.A1(n_14202),
.A2(n_13853),
.B1(n_13980),
.B2(n_13867),
.Y(n_14293)
);

INVx1_ASAP7_75t_L g14294 ( 
.A(n_14086),
.Y(n_14294)
);

INVx1_ASAP7_75t_L g14295 ( 
.A(n_14025),
.Y(n_14295)
);

AND2x2_ASAP7_75t_L g14296 ( 
.A(n_14056),
.B(n_14054),
.Y(n_14296)
);

INVx2_ASAP7_75t_L g14297 ( 
.A(n_14091),
.Y(n_14297)
);

AND2x2_ASAP7_75t_L g14298 ( 
.A(n_14059),
.B(n_13943),
.Y(n_14298)
);

BUFx3_ASAP7_75t_L g14299 ( 
.A(n_14037),
.Y(n_14299)
);

AOI22xp33_ASAP7_75t_L g14300 ( 
.A1(n_14187),
.A2(n_13888),
.B1(n_13899),
.B2(n_13871),
.Y(n_14300)
);

INVx1_ASAP7_75t_L g14301 ( 
.A(n_14131),
.Y(n_14301)
);

INVx1_ASAP7_75t_L g14302 ( 
.A(n_14020),
.Y(n_14302)
);

INVx1_ASAP7_75t_L g14303 ( 
.A(n_14133),
.Y(n_14303)
);

NAND2xp5_ASAP7_75t_L g14304 ( 
.A(n_14087),
.B(n_13997),
.Y(n_14304)
);

OR2x2_ASAP7_75t_L g14305 ( 
.A(n_14142),
.B(n_13962),
.Y(n_14305)
);

BUFx6f_ASAP7_75t_L g14306 ( 
.A(n_14039),
.Y(n_14306)
);

INVxp67_ASAP7_75t_SL g14307 ( 
.A(n_14001),
.Y(n_14307)
);

AND2x2_ASAP7_75t_L g14308 ( 
.A(n_14120),
.B(n_13966),
.Y(n_14308)
);

AOI22xp33_ASAP7_75t_L g14309 ( 
.A1(n_14153),
.A2(n_13994),
.B1(n_13944),
.B2(n_13973),
.Y(n_14309)
);

AND2x2_ASAP7_75t_L g14310 ( 
.A(n_14095),
.B(n_13968),
.Y(n_14310)
);

INVxp67_ASAP7_75t_L g14311 ( 
.A(n_14188),
.Y(n_14311)
);

NAND2xp5_ASAP7_75t_L g14312 ( 
.A(n_14150),
.B(n_2511),
.Y(n_14312)
);

HB1xp67_ASAP7_75t_L g14313 ( 
.A(n_14128),
.Y(n_14313)
);

AOI22xp33_ASAP7_75t_L g14314 ( 
.A1(n_14181),
.A2(n_2516),
.B1(n_2513),
.B2(n_2515),
.Y(n_14314)
);

NAND2xp5_ASAP7_75t_L g14315 ( 
.A(n_14085),
.B(n_2513),
.Y(n_14315)
);

INVx1_ASAP7_75t_L g14316 ( 
.A(n_14134),
.Y(n_14316)
);

AND2x2_ASAP7_75t_L g14317 ( 
.A(n_14033),
.B(n_2516),
.Y(n_14317)
);

AND2x2_ASAP7_75t_L g14318 ( 
.A(n_14079),
.B(n_2517),
.Y(n_14318)
);

OR2x2_ASAP7_75t_L g14319 ( 
.A(n_14162),
.B(n_2518),
.Y(n_14319)
);

INVxp67_ASAP7_75t_SL g14320 ( 
.A(n_14137),
.Y(n_14320)
);

AND2x2_ASAP7_75t_L g14321 ( 
.A(n_14072),
.B(n_2519),
.Y(n_14321)
);

BUFx2_ASAP7_75t_L g14322 ( 
.A(n_14114),
.Y(n_14322)
);

AND2x2_ASAP7_75t_L g14323 ( 
.A(n_14082),
.B(n_14052),
.Y(n_14323)
);

INVx1_ASAP7_75t_L g14324 ( 
.A(n_14130),
.Y(n_14324)
);

OR2x2_ASAP7_75t_L g14325 ( 
.A(n_14165),
.B(n_14176),
.Y(n_14325)
);

AND2x2_ASAP7_75t_L g14326 ( 
.A(n_14102),
.B(n_2519),
.Y(n_14326)
);

INVx2_ASAP7_75t_L g14327 ( 
.A(n_14101),
.Y(n_14327)
);

INVx1_ASAP7_75t_L g14328 ( 
.A(n_14083),
.Y(n_14328)
);

HB1xp67_ASAP7_75t_L g14329 ( 
.A(n_14069),
.Y(n_14329)
);

AND2x2_ASAP7_75t_L g14330 ( 
.A(n_14106),
.B(n_2521),
.Y(n_14330)
);

NAND2xp5_ASAP7_75t_L g14331 ( 
.A(n_14168),
.B(n_2522),
.Y(n_14331)
);

NAND2xp5_ASAP7_75t_L g14332 ( 
.A(n_14146),
.B(n_2522),
.Y(n_14332)
);

NOR2xp33_ASAP7_75t_L g14333 ( 
.A(n_14193),
.B(n_2523),
.Y(n_14333)
);

INVx1_ASAP7_75t_L g14334 ( 
.A(n_14112),
.Y(n_14334)
);

INVx2_ASAP7_75t_L g14335 ( 
.A(n_14007),
.Y(n_14335)
);

BUFx3_ASAP7_75t_L g14336 ( 
.A(n_14055),
.Y(n_14336)
);

AND2x2_ASAP7_75t_L g14337 ( 
.A(n_14115),
.B(n_14140),
.Y(n_14337)
);

INVx1_ASAP7_75t_L g14338 ( 
.A(n_14118),
.Y(n_14338)
);

NAND2xp5_ASAP7_75t_L g14339 ( 
.A(n_14159),
.B(n_2523),
.Y(n_14339)
);

BUFx2_ASAP7_75t_L g14340 ( 
.A(n_14116),
.Y(n_14340)
);

NAND2x1_ASAP7_75t_L g14341 ( 
.A(n_14127),
.B(n_2524),
.Y(n_14341)
);

HB1xp67_ASAP7_75t_L g14342 ( 
.A(n_14141),
.Y(n_14342)
);

INVx1_ASAP7_75t_L g14343 ( 
.A(n_14119),
.Y(n_14343)
);

INVx1_ASAP7_75t_L g14344 ( 
.A(n_14065),
.Y(n_14344)
);

AND2x2_ASAP7_75t_L g14345 ( 
.A(n_14179),
.B(n_2524),
.Y(n_14345)
);

HB1xp67_ASAP7_75t_L g14346 ( 
.A(n_14144),
.Y(n_14346)
);

AND2x2_ASAP7_75t_L g14347 ( 
.A(n_14183),
.B(n_2525),
.Y(n_14347)
);

INVx1_ASAP7_75t_L g14348 ( 
.A(n_14077),
.Y(n_14348)
);

INVx1_ASAP7_75t_L g14349 ( 
.A(n_14078),
.Y(n_14349)
);

HB1xp67_ASAP7_75t_L g14350 ( 
.A(n_14139),
.Y(n_14350)
);

HB1xp67_ASAP7_75t_L g14351 ( 
.A(n_14136),
.Y(n_14351)
);

INVx1_ASAP7_75t_L g14352 ( 
.A(n_14089),
.Y(n_14352)
);

AND2x2_ASAP7_75t_L g14353 ( 
.A(n_14195),
.B(n_2525),
.Y(n_14353)
);

INVx2_ASAP7_75t_L g14354 ( 
.A(n_14121),
.Y(n_14354)
);

INVx1_ASAP7_75t_L g14355 ( 
.A(n_14090),
.Y(n_14355)
);

INVx1_ASAP7_75t_L g14356 ( 
.A(n_14093),
.Y(n_14356)
);

BUFx3_ASAP7_75t_L g14357 ( 
.A(n_14200),
.Y(n_14357)
);

NOR2xp33_ASAP7_75t_L g14358 ( 
.A(n_14174),
.B(n_2526),
.Y(n_14358)
);

AND2x2_ASAP7_75t_L g14359 ( 
.A(n_14251),
.B(n_14190),
.Y(n_14359)
);

INVx1_ASAP7_75t_L g14360 ( 
.A(n_14211),
.Y(n_14360)
);

AND2x4_ASAP7_75t_L g14361 ( 
.A(n_14217),
.B(n_14206),
.Y(n_14361)
);

OR2x2_ASAP7_75t_L g14362 ( 
.A(n_14232),
.B(n_14177),
.Y(n_14362)
);

INVx1_ASAP7_75t_L g14363 ( 
.A(n_14313),
.Y(n_14363)
);

OR2x2_ASAP7_75t_L g14364 ( 
.A(n_14311),
.B(n_14170),
.Y(n_14364)
);

INVx2_ASAP7_75t_L g14365 ( 
.A(n_14240),
.Y(n_14365)
);

BUFx2_ASAP7_75t_L g14366 ( 
.A(n_14213),
.Y(n_14366)
);

NOR2x1_ASAP7_75t_L g14367 ( 
.A(n_14341),
.B(n_14160),
.Y(n_14367)
);

AND2x2_ASAP7_75t_L g14368 ( 
.A(n_14296),
.B(n_14175),
.Y(n_14368)
);

INVx3_ASAP7_75t_L g14369 ( 
.A(n_14291),
.Y(n_14369)
);

AND2x2_ASAP7_75t_L g14370 ( 
.A(n_14216),
.B(n_14173),
.Y(n_14370)
);

INVx1_ASAP7_75t_L g14371 ( 
.A(n_14340),
.Y(n_14371)
);

AND2x2_ASAP7_75t_L g14372 ( 
.A(n_14247),
.B(n_14147),
.Y(n_14372)
);

INVx2_ASAP7_75t_SL g14373 ( 
.A(n_14271),
.Y(n_14373)
);

INVx1_ASAP7_75t_SL g14374 ( 
.A(n_14322),
.Y(n_14374)
);

INVx2_ASAP7_75t_L g14375 ( 
.A(n_14299),
.Y(n_14375)
);

INVx2_ASAP7_75t_L g14376 ( 
.A(n_14205),
.Y(n_14376)
);

AND2x2_ASAP7_75t_SL g14377 ( 
.A(n_14207),
.B(n_14196),
.Y(n_14377)
);

INVx1_ASAP7_75t_L g14378 ( 
.A(n_14263),
.Y(n_14378)
);

INVx2_ASAP7_75t_L g14379 ( 
.A(n_14336),
.Y(n_14379)
);

INVx2_ASAP7_75t_L g14380 ( 
.A(n_14218),
.Y(n_14380)
);

OR2x2_ASAP7_75t_L g14381 ( 
.A(n_14256),
.B(n_14197),
.Y(n_14381)
);

INVx1_ASAP7_75t_L g14382 ( 
.A(n_14203),
.Y(n_14382)
);

INVx2_ASAP7_75t_SL g14383 ( 
.A(n_14306),
.Y(n_14383)
);

NAND2xp5_ASAP7_75t_L g14384 ( 
.A(n_14209),
.B(n_14182),
.Y(n_14384)
);

AND2x2_ASAP7_75t_L g14385 ( 
.A(n_14204),
.B(n_14152),
.Y(n_14385)
);

INVx2_ASAP7_75t_L g14386 ( 
.A(n_14268),
.Y(n_14386)
);

INVx1_ASAP7_75t_L g14387 ( 
.A(n_14303),
.Y(n_14387)
);

INVx1_ASAP7_75t_L g14388 ( 
.A(n_14316),
.Y(n_14388)
);

AND2x4_ASAP7_75t_L g14389 ( 
.A(n_14257),
.B(n_14138),
.Y(n_14389)
);

INVx2_ASAP7_75t_L g14390 ( 
.A(n_14242),
.Y(n_14390)
);

AND2x2_ASAP7_75t_L g14391 ( 
.A(n_14238),
.B(n_14178),
.Y(n_14391)
);

AND2x4_ASAP7_75t_SL g14392 ( 
.A(n_14220),
.B(n_14180),
.Y(n_14392)
);

INVx2_ASAP7_75t_L g14393 ( 
.A(n_14306),
.Y(n_14393)
);

AND2x2_ASAP7_75t_L g14394 ( 
.A(n_14229),
.B(n_14199),
.Y(n_14394)
);

NOR2xp33_ASAP7_75t_L g14395 ( 
.A(n_14307),
.B(n_14064),
.Y(n_14395)
);

INVx2_ASAP7_75t_L g14396 ( 
.A(n_14297),
.Y(n_14396)
);

INVx2_ASAP7_75t_L g14397 ( 
.A(n_14230),
.Y(n_14397)
);

NAND2xp5_ASAP7_75t_L g14398 ( 
.A(n_14320),
.B(n_14145),
.Y(n_14398)
);

NAND2xp5_ASAP7_75t_L g14399 ( 
.A(n_14272),
.B(n_14164),
.Y(n_14399)
);

AND2x2_ASAP7_75t_L g14400 ( 
.A(n_14323),
.B(n_14201),
.Y(n_14400)
);

AND2x2_ASAP7_75t_L g14401 ( 
.A(n_14226),
.B(n_14125),
.Y(n_14401)
);

INVx1_ASAP7_75t_L g14402 ( 
.A(n_14237),
.Y(n_14402)
);

INVx1_ASAP7_75t_L g14403 ( 
.A(n_14258),
.Y(n_14403)
);

INVx2_ASAP7_75t_L g14404 ( 
.A(n_14221),
.Y(n_14404)
);

NAND2xp5_ASAP7_75t_L g14405 ( 
.A(n_14277),
.B(n_14148),
.Y(n_14405)
);

INVx2_ASAP7_75t_L g14406 ( 
.A(n_14261),
.Y(n_14406)
);

AND2x4_ASAP7_75t_L g14407 ( 
.A(n_14290),
.B(n_14066),
.Y(n_14407)
);

HB1xp67_ASAP7_75t_L g14408 ( 
.A(n_14260),
.Y(n_14408)
);

INVx1_ASAP7_75t_L g14409 ( 
.A(n_14212),
.Y(n_14409)
);

OR2x2_ASAP7_75t_L g14410 ( 
.A(n_14265),
.B(n_14092),
.Y(n_14410)
);

NAND2xp5_ASAP7_75t_L g14411 ( 
.A(n_14224),
.B(n_14189),
.Y(n_14411)
);

AND2x2_ASAP7_75t_L g14412 ( 
.A(n_14248),
.B(n_14021),
.Y(n_14412)
);

NAND2xp5_ASAP7_75t_L g14413 ( 
.A(n_14239),
.B(n_14151),
.Y(n_14413)
);

OR2x2_ASAP7_75t_L g14414 ( 
.A(n_14267),
.B(n_14246),
.Y(n_14414)
);

INVx1_ASAP7_75t_L g14415 ( 
.A(n_14214),
.Y(n_14415)
);

INVx1_ASAP7_75t_L g14416 ( 
.A(n_14210),
.Y(n_14416)
);

INVx2_ASAP7_75t_L g14417 ( 
.A(n_14317),
.Y(n_14417)
);

OR2x2_ASAP7_75t_L g14418 ( 
.A(n_14264),
.B(n_14067),
.Y(n_14418)
);

AND2x2_ASAP7_75t_L g14419 ( 
.A(n_14253),
.B(n_14135),
.Y(n_14419)
);

AND2x2_ASAP7_75t_L g14420 ( 
.A(n_14241),
.B(n_14155),
.Y(n_14420)
);

INVx2_ASAP7_75t_L g14421 ( 
.A(n_14288),
.Y(n_14421)
);

BUFx2_ASAP7_75t_L g14422 ( 
.A(n_14215),
.Y(n_14422)
);

INVx1_ASAP7_75t_L g14423 ( 
.A(n_14274),
.Y(n_14423)
);

NOR2xp33_ASAP7_75t_L g14424 ( 
.A(n_14250),
.B(n_14161),
.Y(n_14424)
);

AND2x2_ASAP7_75t_L g14425 ( 
.A(n_14357),
.B(n_14154),
.Y(n_14425)
);

NAND2xp5_ASAP7_75t_L g14426 ( 
.A(n_14259),
.B(n_14266),
.Y(n_14426)
);

AND2x2_ASAP7_75t_L g14427 ( 
.A(n_14255),
.B(n_14347),
.Y(n_14427)
);

AND2x2_ASAP7_75t_L g14428 ( 
.A(n_14346),
.B(n_14094),
.Y(n_14428)
);

OR2x2_ASAP7_75t_L g14429 ( 
.A(n_14233),
.B(n_14169),
.Y(n_14429)
);

AND2x4_ASAP7_75t_L g14430 ( 
.A(n_14275),
.B(n_14096),
.Y(n_14430)
);

INVx3_ASAP7_75t_L g14431 ( 
.A(n_14276),
.Y(n_14431)
);

AND2x2_ASAP7_75t_L g14432 ( 
.A(n_14345),
.B(n_14097),
.Y(n_14432)
);

AND2x4_ASAP7_75t_L g14433 ( 
.A(n_14354),
.B(n_14098),
.Y(n_14433)
);

HB1xp67_ASAP7_75t_L g14434 ( 
.A(n_14342),
.Y(n_14434)
);

NAND2xp5_ASAP7_75t_L g14435 ( 
.A(n_14308),
.B(n_14186),
.Y(n_14435)
);

NAND2xp5_ASAP7_75t_L g14436 ( 
.A(n_14219),
.B(n_14185),
.Y(n_14436)
);

OR2x2_ASAP7_75t_L g14437 ( 
.A(n_14325),
.B(n_14100),
.Y(n_14437)
);

HB1xp67_ASAP7_75t_L g14438 ( 
.A(n_14350),
.Y(n_14438)
);

OR2x2_ASAP7_75t_L g14439 ( 
.A(n_14244),
.B(n_14104),
.Y(n_14439)
);

NAND2xp5_ASAP7_75t_L g14440 ( 
.A(n_14298),
.B(n_14270),
.Y(n_14440)
);

AND2x2_ASAP7_75t_L g14441 ( 
.A(n_14353),
.B(n_14108),
.Y(n_14441)
);

AND2x2_ASAP7_75t_L g14442 ( 
.A(n_14337),
.B(n_14109),
.Y(n_14442)
);

AND2x4_ASAP7_75t_L g14443 ( 
.A(n_14334),
.B(n_14327),
.Y(n_14443)
);

NAND2xp5_ASAP7_75t_L g14444 ( 
.A(n_14273),
.B(n_14166),
.Y(n_14444)
);

INVx1_ASAP7_75t_L g14445 ( 
.A(n_14329),
.Y(n_14445)
);

INVx1_ASAP7_75t_L g14446 ( 
.A(n_14225),
.Y(n_14446)
);

INVx2_ASAP7_75t_L g14447 ( 
.A(n_14318),
.Y(n_14447)
);

AND2x2_ASAP7_75t_L g14448 ( 
.A(n_14245),
.B(n_14310),
.Y(n_14448)
);

AND2x2_ASAP7_75t_L g14449 ( 
.A(n_14208),
.B(n_14110),
.Y(n_14449)
);

INVx4_ASAP7_75t_L g14450 ( 
.A(n_14321),
.Y(n_14450)
);

AND2x2_ASAP7_75t_L g14451 ( 
.A(n_14252),
.B(n_14198),
.Y(n_14451)
);

NAND2xp5_ASAP7_75t_L g14452 ( 
.A(n_14262),
.B(n_2526),
.Y(n_14452)
);

NAND2xp5_ASAP7_75t_L g14453 ( 
.A(n_14281),
.B(n_2527),
.Y(n_14453)
);

AND2x2_ASAP7_75t_L g14454 ( 
.A(n_14335),
.B(n_2527),
.Y(n_14454)
);

OR2x2_ASAP7_75t_L g14455 ( 
.A(n_14223),
.B(n_2528),
.Y(n_14455)
);

INVx1_ASAP7_75t_L g14456 ( 
.A(n_14326),
.Y(n_14456)
);

AND2x2_ASAP7_75t_L g14457 ( 
.A(n_14279),
.B(n_2528),
.Y(n_14457)
);

AND2x2_ASAP7_75t_L g14458 ( 
.A(n_14294),
.B(n_2529),
.Y(n_14458)
);

AND2x2_ASAP7_75t_L g14459 ( 
.A(n_14254),
.B(n_2530),
.Y(n_14459)
);

INVx2_ASAP7_75t_L g14460 ( 
.A(n_14330),
.Y(n_14460)
);

INVx2_ASAP7_75t_L g14461 ( 
.A(n_14228),
.Y(n_14461)
);

INVx2_ASAP7_75t_L g14462 ( 
.A(n_14234),
.Y(n_14462)
);

NAND2xp5_ASAP7_75t_L g14463 ( 
.A(n_14287),
.B(n_2530),
.Y(n_14463)
);

INVx1_ASAP7_75t_L g14464 ( 
.A(n_14312),
.Y(n_14464)
);

INVx2_ASAP7_75t_L g14465 ( 
.A(n_14222),
.Y(n_14465)
);

NOR2x1_ASAP7_75t_L g14466 ( 
.A(n_14315),
.B(n_14319),
.Y(n_14466)
);

INVx1_ASAP7_75t_L g14467 ( 
.A(n_14227),
.Y(n_14467)
);

BUFx3_ASAP7_75t_L g14468 ( 
.A(n_14328),
.Y(n_14468)
);

AND2x2_ASAP7_75t_L g14469 ( 
.A(n_14358),
.B(n_2531),
.Y(n_14469)
);

HB1xp67_ASAP7_75t_L g14470 ( 
.A(n_14284),
.Y(n_14470)
);

HB1xp67_ASAP7_75t_L g14471 ( 
.A(n_14292),
.Y(n_14471)
);

INVx1_ASAP7_75t_SL g14472 ( 
.A(n_14339),
.Y(n_14472)
);

INVx1_ASAP7_75t_L g14473 ( 
.A(n_14301),
.Y(n_14473)
);

AND2x2_ASAP7_75t_L g14474 ( 
.A(n_14333),
.B(n_2531),
.Y(n_14474)
);

INVx2_ASAP7_75t_L g14475 ( 
.A(n_14295),
.Y(n_14475)
);

INVx1_ASAP7_75t_L g14476 ( 
.A(n_14278),
.Y(n_14476)
);

NAND2xp5_ASAP7_75t_L g14477 ( 
.A(n_14309),
.B(n_2532),
.Y(n_14477)
);

AND2x4_ASAP7_75t_L g14478 ( 
.A(n_14324),
.B(n_2532),
.Y(n_14478)
);

AND2x2_ASAP7_75t_L g14479 ( 
.A(n_14351),
.B(n_2533),
.Y(n_14479)
);

INVx1_ASAP7_75t_L g14480 ( 
.A(n_14302),
.Y(n_14480)
);

NAND2xp5_ASAP7_75t_L g14481 ( 
.A(n_14293),
.B(n_2533),
.Y(n_14481)
);

AND2x2_ASAP7_75t_L g14482 ( 
.A(n_14269),
.B(n_2534),
.Y(n_14482)
);

INVx1_ASAP7_75t_L g14483 ( 
.A(n_14331),
.Y(n_14483)
);

HB1xp67_ASAP7_75t_L g14484 ( 
.A(n_14338),
.Y(n_14484)
);

INVx1_ASAP7_75t_L g14485 ( 
.A(n_14343),
.Y(n_14485)
);

AND2x2_ASAP7_75t_L g14486 ( 
.A(n_14283),
.B(n_2534),
.Y(n_14486)
);

INVx1_ASAP7_75t_L g14487 ( 
.A(n_14344),
.Y(n_14487)
);

AND2x2_ASAP7_75t_L g14488 ( 
.A(n_14332),
.B(n_2535),
.Y(n_14488)
);

AND2x2_ASAP7_75t_L g14489 ( 
.A(n_14282),
.B(n_2535),
.Y(n_14489)
);

AND2x2_ASAP7_75t_L g14490 ( 
.A(n_14235),
.B(n_2536),
.Y(n_14490)
);

HB1xp67_ASAP7_75t_L g14491 ( 
.A(n_14348),
.Y(n_14491)
);

INVx1_ASAP7_75t_L g14492 ( 
.A(n_14366),
.Y(n_14492)
);

INVx1_ASAP7_75t_L g14493 ( 
.A(n_14434),
.Y(n_14493)
);

AOI22xp5_ASAP7_75t_L g14494 ( 
.A1(n_14377),
.A2(n_14249),
.B1(n_14231),
.B2(n_14304),
.Y(n_14494)
);

INVx1_ASAP7_75t_SL g14495 ( 
.A(n_14374),
.Y(n_14495)
);

AOI21xp5_ASAP7_75t_SL g14496 ( 
.A1(n_14373),
.A2(n_14463),
.B(n_14361),
.Y(n_14496)
);

INVx4_ASAP7_75t_L g14497 ( 
.A(n_14369),
.Y(n_14497)
);

AND2x2_ASAP7_75t_L g14498 ( 
.A(n_14359),
.B(n_14300),
.Y(n_14498)
);

NAND3xp33_ASAP7_75t_L g14499 ( 
.A(n_14413),
.B(n_14285),
.C(n_14286),
.Y(n_14499)
);

INVx2_ASAP7_75t_L g14500 ( 
.A(n_14425),
.Y(n_14500)
);

INVx3_ASAP7_75t_L g14501 ( 
.A(n_14443),
.Y(n_14501)
);

INVx2_ASAP7_75t_L g14502 ( 
.A(n_14360),
.Y(n_14502)
);

NAND2xp5_ASAP7_75t_L g14503 ( 
.A(n_14392),
.B(n_14236),
.Y(n_14503)
);

INVx1_ASAP7_75t_L g14504 ( 
.A(n_14438),
.Y(n_14504)
);

INVxp67_ASAP7_75t_SL g14505 ( 
.A(n_14367),
.Y(n_14505)
);

NAND2xp5_ASAP7_75t_L g14506 ( 
.A(n_14395),
.B(n_14289),
.Y(n_14506)
);

NAND2xp5_ASAP7_75t_L g14507 ( 
.A(n_14368),
.B(n_14305),
.Y(n_14507)
);

AOI222xp33_ASAP7_75t_L g14508 ( 
.A1(n_14412),
.A2(n_14243),
.B1(n_14280),
.B2(n_14349),
.C1(n_14355),
.C2(n_14352),
.Y(n_14508)
);

INVx1_ASAP7_75t_L g14509 ( 
.A(n_14408),
.Y(n_14509)
);

INVx3_ASAP7_75t_L g14510 ( 
.A(n_14468),
.Y(n_14510)
);

AND2x2_ASAP7_75t_L g14511 ( 
.A(n_14420),
.B(n_14356),
.Y(n_14511)
);

INVx1_ASAP7_75t_L g14512 ( 
.A(n_14422),
.Y(n_14512)
);

INVx2_ASAP7_75t_L g14513 ( 
.A(n_14370),
.Y(n_14513)
);

NOR2x1_ASAP7_75t_SL g14514 ( 
.A(n_14437),
.B(n_14314),
.Y(n_14514)
);

AND2x2_ASAP7_75t_L g14515 ( 
.A(n_14385),
.B(n_14448),
.Y(n_14515)
);

AO21x2_ASAP7_75t_L g14516 ( 
.A1(n_14477),
.A2(n_2536),
.B(n_2537),
.Y(n_14516)
);

INVx1_ASAP7_75t_L g14517 ( 
.A(n_14372),
.Y(n_14517)
);

HB1xp67_ASAP7_75t_L g14518 ( 
.A(n_14378),
.Y(n_14518)
);

AND2x2_ASAP7_75t_L g14519 ( 
.A(n_14400),
.B(n_2538),
.Y(n_14519)
);

AND2x2_ASAP7_75t_L g14520 ( 
.A(n_14394),
.B(n_2538),
.Y(n_14520)
);

NAND2x1_ASAP7_75t_L g14521 ( 
.A(n_14450),
.B(n_2539),
.Y(n_14521)
);

INVx1_ASAP7_75t_L g14522 ( 
.A(n_14428),
.Y(n_14522)
);

BUFx3_ASAP7_75t_L g14523 ( 
.A(n_14365),
.Y(n_14523)
);

AND2x2_ASAP7_75t_L g14524 ( 
.A(n_14427),
.B(n_2539),
.Y(n_14524)
);

OR2x2_ASAP7_75t_L g14525 ( 
.A(n_14362),
.B(n_2540),
.Y(n_14525)
);

INVx1_ASAP7_75t_L g14526 ( 
.A(n_14442),
.Y(n_14526)
);

INVx2_ASAP7_75t_L g14527 ( 
.A(n_14380),
.Y(n_14527)
);

INVx1_ASAP7_75t_L g14528 ( 
.A(n_14364),
.Y(n_14528)
);

INVxp67_ASAP7_75t_SL g14529 ( 
.A(n_14414),
.Y(n_14529)
);

INVx2_ASAP7_75t_L g14530 ( 
.A(n_14396),
.Y(n_14530)
);

AND2x2_ASAP7_75t_L g14531 ( 
.A(n_14391),
.B(n_2540),
.Y(n_14531)
);

AND2x2_ASAP7_75t_L g14532 ( 
.A(n_14457),
.B(n_2541),
.Y(n_14532)
);

INVx1_ASAP7_75t_L g14533 ( 
.A(n_14470),
.Y(n_14533)
);

AOI22xp33_ASAP7_75t_L g14534 ( 
.A1(n_14419),
.A2(n_2544),
.B1(n_2542),
.B2(n_2543),
.Y(n_14534)
);

NAND2xp5_ASAP7_75t_L g14535 ( 
.A(n_14383),
.B(n_2542),
.Y(n_14535)
);

AND2x2_ASAP7_75t_L g14536 ( 
.A(n_14482),
.B(n_2543),
.Y(n_14536)
);

OAI21x1_ASAP7_75t_L g14537 ( 
.A1(n_14405),
.A2(n_2544),
.B(n_2545),
.Y(n_14537)
);

INVx1_ASAP7_75t_L g14538 ( 
.A(n_14471),
.Y(n_14538)
);

AO21x2_ASAP7_75t_L g14539 ( 
.A1(n_14481),
.A2(n_14479),
.B(n_14490),
.Y(n_14539)
);

INVx2_ASAP7_75t_L g14540 ( 
.A(n_14375),
.Y(n_14540)
);

AND2x2_ASAP7_75t_L g14541 ( 
.A(n_14401),
.B(n_2545),
.Y(n_14541)
);

INVx1_ASAP7_75t_L g14542 ( 
.A(n_14371),
.Y(n_14542)
);

INVx1_ASAP7_75t_L g14543 ( 
.A(n_14449),
.Y(n_14543)
);

NAND2xp5_ASAP7_75t_L g14544 ( 
.A(n_14407),
.B(n_2546),
.Y(n_14544)
);

INVx2_ASAP7_75t_L g14545 ( 
.A(n_14379),
.Y(n_14545)
);

AND2x4_ASAP7_75t_L g14546 ( 
.A(n_14376),
.B(n_2547),
.Y(n_14546)
);

AOI22xp33_ASAP7_75t_L g14547 ( 
.A1(n_14418),
.A2(n_2549),
.B1(n_2547),
.B2(n_2548),
.Y(n_14547)
);

BUFx3_ASAP7_75t_L g14548 ( 
.A(n_14433),
.Y(n_14548)
);

AND2x4_ASAP7_75t_L g14549 ( 
.A(n_14386),
.B(n_2548),
.Y(n_14549)
);

BUFx3_ASAP7_75t_L g14550 ( 
.A(n_14389),
.Y(n_14550)
);

INVx3_ASAP7_75t_L g14551 ( 
.A(n_14430),
.Y(n_14551)
);

INVx2_ASAP7_75t_L g14552 ( 
.A(n_14417),
.Y(n_14552)
);

OAI21xp5_ASAP7_75t_L g14553 ( 
.A1(n_14424),
.A2(n_2549),
.B(n_2550),
.Y(n_14553)
);

INVx1_ASAP7_75t_SL g14554 ( 
.A(n_14381),
.Y(n_14554)
);

AND2x4_ASAP7_75t_L g14555 ( 
.A(n_14393),
.B(n_2550),
.Y(n_14555)
);

OR2x2_ASAP7_75t_L g14556 ( 
.A(n_14440),
.B(n_2551),
.Y(n_14556)
);

INVx2_ASAP7_75t_L g14557 ( 
.A(n_14431),
.Y(n_14557)
);

OR2x2_ASAP7_75t_L g14558 ( 
.A(n_14435),
.B(n_2551),
.Y(n_14558)
);

AO21x2_ASAP7_75t_L g14559 ( 
.A1(n_14453),
.A2(n_2552),
.B(n_2553),
.Y(n_14559)
);

BUFx3_ASAP7_75t_L g14560 ( 
.A(n_14390),
.Y(n_14560)
);

INVx1_ASAP7_75t_L g14561 ( 
.A(n_14445),
.Y(n_14561)
);

OAI22xp5_ASAP7_75t_L g14562 ( 
.A1(n_14410),
.A2(n_2554),
.B1(n_2552),
.B2(n_2553),
.Y(n_14562)
);

AND2x2_ASAP7_75t_L g14563 ( 
.A(n_14486),
.B(n_2555),
.Y(n_14563)
);

HB1xp67_ASAP7_75t_L g14564 ( 
.A(n_14484),
.Y(n_14564)
);

NAND2x1_ASAP7_75t_L g14565 ( 
.A(n_14363),
.B(n_2555),
.Y(n_14565)
);

AOI22xp33_ASAP7_75t_SL g14566 ( 
.A1(n_14411),
.A2(n_2558),
.B1(n_2556),
.B2(n_2557),
.Y(n_14566)
);

INVx2_ASAP7_75t_L g14567 ( 
.A(n_14478),
.Y(n_14567)
);

AND2x2_ASAP7_75t_L g14568 ( 
.A(n_14489),
.B(n_2556),
.Y(n_14568)
);

INVx1_ASAP7_75t_L g14569 ( 
.A(n_14454),
.Y(n_14569)
);

OAI221xp5_ASAP7_75t_SL g14570 ( 
.A1(n_14429),
.A2(n_2560),
.B1(n_2558),
.B2(n_2559),
.C(n_2561),
.Y(n_14570)
);

NAND3xp33_ASAP7_75t_L g14571 ( 
.A(n_14402),
.B(n_2561),
.C(n_2562),
.Y(n_14571)
);

AND2x2_ASAP7_75t_L g14572 ( 
.A(n_14397),
.B(n_2563),
.Y(n_14572)
);

AND2x2_ASAP7_75t_L g14573 ( 
.A(n_14406),
.B(n_2564),
.Y(n_14573)
);

INVx2_ASAP7_75t_L g14574 ( 
.A(n_14447),
.Y(n_14574)
);

OAI22xp5_ASAP7_75t_L g14575 ( 
.A1(n_14426),
.A2(n_2567),
.B1(n_2565),
.B2(n_2566),
.Y(n_14575)
);

OR2x2_ASAP7_75t_L g14576 ( 
.A(n_14398),
.B(n_14384),
.Y(n_14576)
);

INVx1_ASAP7_75t_L g14577 ( 
.A(n_14458),
.Y(n_14577)
);

NOR3xp33_ASAP7_75t_SL g14578 ( 
.A(n_14399),
.B(n_2565),
.C(n_2568),
.Y(n_14578)
);

NAND2xp5_ASAP7_75t_L g14579 ( 
.A(n_14451),
.B(n_2568),
.Y(n_14579)
);

AND2x2_ASAP7_75t_L g14580 ( 
.A(n_14460),
.B(n_2569),
.Y(n_14580)
);

HB1xp67_ASAP7_75t_L g14581 ( 
.A(n_14491),
.Y(n_14581)
);

INVx1_ASAP7_75t_L g14582 ( 
.A(n_14459),
.Y(n_14582)
);

INVxp67_ASAP7_75t_SL g14583 ( 
.A(n_14466),
.Y(n_14583)
);

INVx1_ASAP7_75t_L g14584 ( 
.A(n_14432),
.Y(n_14584)
);

INVx1_ASAP7_75t_L g14585 ( 
.A(n_14441),
.Y(n_14585)
);

AOI211xp5_ASAP7_75t_L g14586 ( 
.A1(n_14382),
.A2(n_2572),
.B(n_2570),
.C(n_2571),
.Y(n_14586)
);

OR2x2_ASAP7_75t_L g14587 ( 
.A(n_14444),
.B(n_14452),
.Y(n_14587)
);

OAI211xp5_ASAP7_75t_SL g14588 ( 
.A1(n_14436),
.A2(n_14472),
.B(n_14439),
.C(n_14483),
.Y(n_14588)
);

INVx1_ASAP7_75t_L g14589 ( 
.A(n_14488),
.Y(n_14589)
);

OR2x2_ASAP7_75t_L g14590 ( 
.A(n_14455),
.B(n_2570),
.Y(n_14590)
);

AOI22xp33_ASAP7_75t_L g14591 ( 
.A1(n_14404),
.A2(n_2573),
.B1(n_2571),
.B2(n_2572),
.Y(n_14591)
);

BUFx2_ASAP7_75t_L g14592 ( 
.A(n_14423),
.Y(n_14592)
);

OR2x2_ASAP7_75t_L g14593 ( 
.A(n_14421),
.B(n_2574),
.Y(n_14593)
);

INVx2_ASAP7_75t_L g14594 ( 
.A(n_14456),
.Y(n_14594)
);

NAND2xp5_ASAP7_75t_L g14595 ( 
.A(n_14474),
.B(n_2574),
.Y(n_14595)
);

INVx1_ASAP7_75t_L g14596 ( 
.A(n_14416),
.Y(n_14596)
);

INVx1_ASAP7_75t_L g14597 ( 
.A(n_14446),
.Y(n_14597)
);

BUFx6f_ASAP7_75t_L g14598 ( 
.A(n_14469),
.Y(n_14598)
);

INVx1_ASAP7_75t_L g14599 ( 
.A(n_14403),
.Y(n_14599)
);

NAND2xp5_ASAP7_75t_L g14600 ( 
.A(n_14464),
.B(n_2575),
.Y(n_14600)
);

NOR2x1_ASAP7_75t_SL g14601 ( 
.A(n_14475),
.B(n_2575),
.Y(n_14601)
);

AO21x2_ASAP7_75t_L g14602 ( 
.A1(n_14409),
.A2(n_2576),
.B(n_2577),
.Y(n_14602)
);

AND2x4_ASAP7_75t_L g14603 ( 
.A(n_14461),
.B(n_2576),
.Y(n_14603)
);

HB1xp67_ASAP7_75t_L g14604 ( 
.A(n_14415),
.Y(n_14604)
);

NAND2x1_ASAP7_75t_L g14605 ( 
.A(n_14462),
.B(n_14465),
.Y(n_14605)
);

AND2x2_ASAP7_75t_L g14606 ( 
.A(n_14473),
.B(n_2577),
.Y(n_14606)
);

INVx2_ASAP7_75t_L g14607 ( 
.A(n_14601),
.Y(n_14607)
);

OR2x6_ASAP7_75t_L g14608 ( 
.A(n_14496),
.B(n_14467),
.Y(n_14608)
);

INVx1_ASAP7_75t_L g14609 ( 
.A(n_14529),
.Y(n_14609)
);

NAND2xp67_ASAP7_75t_L g14610 ( 
.A(n_14515),
.B(n_14387),
.Y(n_14610)
);

INVx1_ASAP7_75t_L g14611 ( 
.A(n_14583),
.Y(n_14611)
);

INVx2_ASAP7_75t_L g14612 ( 
.A(n_14521),
.Y(n_14612)
);

OR2x2_ASAP7_75t_L g14613 ( 
.A(n_14495),
.B(n_14476),
.Y(n_14613)
);

INVx1_ASAP7_75t_L g14614 ( 
.A(n_14505),
.Y(n_14614)
);

NAND2x1p5_ASAP7_75t_L g14615 ( 
.A(n_14497),
.B(n_14480),
.Y(n_14615)
);

INVx1_ASAP7_75t_L g14616 ( 
.A(n_14564),
.Y(n_14616)
);

INVx1_ASAP7_75t_L g14617 ( 
.A(n_14581),
.Y(n_14617)
);

NAND2xp5_ASAP7_75t_L g14618 ( 
.A(n_14501),
.B(n_14388),
.Y(n_14618)
);

AND2x2_ASAP7_75t_SL g14619 ( 
.A(n_14498),
.B(n_14485),
.Y(n_14619)
);

OR2x2_ASAP7_75t_L g14620 ( 
.A(n_14507),
.B(n_14487),
.Y(n_14620)
);

INVx1_ASAP7_75t_L g14621 ( 
.A(n_14518),
.Y(n_14621)
);

AND2x4_ASAP7_75t_L g14622 ( 
.A(n_14548),
.B(n_2578),
.Y(n_14622)
);

INVx1_ASAP7_75t_L g14623 ( 
.A(n_14492),
.Y(n_14623)
);

NAND2xp5_ASAP7_75t_L g14624 ( 
.A(n_14551),
.B(n_2578),
.Y(n_14624)
);

NOR2x1p5_ASAP7_75t_L g14625 ( 
.A(n_14550),
.B(n_2579),
.Y(n_14625)
);

INVx1_ASAP7_75t_L g14626 ( 
.A(n_14524),
.Y(n_14626)
);

AND2x2_ASAP7_75t_L g14627 ( 
.A(n_14500),
.B(n_2579),
.Y(n_14627)
);

NAND2xp5_ASAP7_75t_L g14628 ( 
.A(n_14512),
.B(n_2580),
.Y(n_14628)
);

AND2x2_ASAP7_75t_L g14629 ( 
.A(n_14511),
.B(n_2580),
.Y(n_14629)
);

AND2x4_ASAP7_75t_SL g14630 ( 
.A(n_14510),
.B(n_14598),
.Y(n_14630)
);

AND2x2_ASAP7_75t_L g14631 ( 
.A(n_14523),
.B(n_2581),
.Y(n_14631)
);

INVx2_ASAP7_75t_L g14632 ( 
.A(n_14565),
.Y(n_14632)
);

OR2x2_ASAP7_75t_L g14633 ( 
.A(n_14525),
.B(n_2582),
.Y(n_14633)
);

HB1xp67_ASAP7_75t_L g14634 ( 
.A(n_14602),
.Y(n_14634)
);

AND2x2_ASAP7_75t_L g14635 ( 
.A(n_14520),
.B(n_2582),
.Y(n_14635)
);

INVx1_ASAP7_75t_L g14636 ( 
.A(n_14519),
.Y(n_14636)
);

AND2x2_ASAP7_75t_L g14637 ( 
.A(n_14513),
.B(n_2583),
.Y(n_14637)
);

INVx1_ASAP7_75t_SL g14638 ( 
.A(n_14554),
.Y(n_14638)
);

OR2x2_ASAP7_75t_L g14639 ( 
.A(n_14493),
.B(n_2583),
.Y(n_14639)
);

AND2x4_ASAP7_75t_L g14640 ( 
.A(n_14560),
.B(n_2584),
.Y(n_14640)
);

AND2x2_ASAP7_75t_L g14641 ( 
.A(n_14567),
.B(n_14543),
.Y(n_14641)
);

AND2x4_ASAP7_75t_L g14642 ( 
.A(n_14517),
.B(n_2584),
.Y(n_14642)
);

OR2x2_ASAP7_75t_L g14643 ( 
.A(n_14504),
.B(n_2585),
.Y(n_14643)
);

NAND2xp5_ASAP7_75t_L g14644 ( 
.A(n_14532),
.B(n_2585),
.Y(n_14644)
);

INVx1_ASAP7_75t_L g14645 ( 
.A(n_14531),
.Y(n_14645)
);

AND2x2_ASAP7_75t_L g14646 ( 
.A(n_14526),
.B(n_2586),
.Y(n_14646)
);

OAI22xp5_ASAP7_75t_L g14647 ( 
.A1(n_14494),
.A2(n_2588),
.B1(n_2586),
.B2(n_2587),
.Y(n_14647)
);

INVx2_ASAP7_75t_L g14648 ( 
.A(n_14598),
.Y(n_14648)
);

HB1xp67_ASAP7_75t_L g14649 ( 
.A(n_14559),
.Y(n_14649)
);

OR2x2_ASAP7_75t_L g14650 ( 
.A(n_14503),
.B(n_14522),
.Y(n_14650)
);

AND2x4_ASAP7_75t_L g14651 ( 
.A(n_14584),
.B(n_2589),
.Y(n_14651)
);

INVx1_ASAP7_75t_L g14652 ( 
.A(n_14536),
.Y(n_14652)
);

NAND2xp5_ASAP7_75t_L g14653 ( 
.A(n_14568),
.B(n_2589),
.Y(n_14653)
);

OR2x2_ASAP7_75t_L g14654 ( 
.A(n_14556),
.B(n_2590),
.Y(n_14654)
);

INVx1_ASAP7_75t_L g14655 ( 
.A(n_14563),
.Y(n_14655)
);

AND2x4_ASAP7_75t_SL g14656 ( 
.A(n_14557),
.B(n_2590),
.Y(n_14656)
);

INVx1_ASAP7_75t_L g14657 ( 
.A(n_14541),
.Y(n_14657)
);

AND2x4_ASAP7_75t_L g14658 ( 
.A(n_14585),
.B(n_2591),
.Y(n_14658)
);

INVx1_ASAP7_75t_L g14659 ( 
.A(n_14509),
.Y(n_14659)
);

AND2x4_ASAP7_75t_L g14660 ( 
.A(n_14552),
.B(n_2591),
.Y(n_14660)
);

AND2x2_ASAP7_75t_L g14661 ( 
.A(n_14539),
.B(n_2592),
.Y(n_14661)
);

AND2x2_ASAP7_75t_L g14662 ( 
.A(n_14540),
.B(n_2592),
.Y(n_14662)
);

OR2x2_ASAP7_75t_L g14663 ( 
.A(n_14506),
.B(n_2593),
.Y(n_14663)
);

NAND2xp5_ASAP7_75t_L g14664 ( 
.A(n_14566),
.B(n_2593),
.Y(n_14664)
);

INVx2_ASAP7_75t_L g14665 ( 
.A(n_14590),
.Y(n_14665)
);

NAND2xp5_ASAP7_75t_L g14666 ( 
.A(n_14533),
.B(n_2594),
.Y(n_14666)
);

INVx2_ASAP7_75t_L g14667 ( 
.A(n_14549),
.Y(n_14667)
);

INVx1_ASAP7_75t_L g14668 ( 
.A(n_14592),
.Y(n_14668)
);

INVx2_ASAP7_75t_L g14669 ( 
.A(n_14555),
.Y(n_14669)
);

INVx1_ASAP7_75t_L g14670 ( 
.A(n_14544),
.Y(n_14670)
);

INVx1_ASAP7_75t_L g14671 ( 
.A(n_14573),
.Y(n_14671)
);

AND2x2_ASAP7_75t_L g14672 ( 
.A(n_14545),
.B(n_2594),
.Y(n_14672)
);

NAND2xp5_ASAP7_75t_L g14673 ( 
.A(n_14538),
.B(n_2595),
.Y(n_14673)
);

INVx2_ASAP7_75t_L g14674 ( 
.A(n_14546),
.Y(n_14674)
);

AND2x2_ASAP7_75t_L g14675 ( 
.A(n_14574),
.B(n_2595),
.Y(n_14675)
);

AND2x2_ASAP7_75t_L g14676 ( 
.A(n_14577),
.B(n_2596),
.Y(n_14676)
);

INVx2_ASAP7_75t_L g14677 ( 
.A(n_14593),
.Y(n_14677)
);

INVx2_ASAP7_75t_L g14678 ( 
.A(n_14603),
.Y(n_14678)
);

NAND2xp5_ASAP7_75t_L g14679 ( 
.A(n_14582),
.B(n_2596),
.Y(n_14679)
);

OR2x2_ASAP7_75t_L g14680 ( 
.A(n_14558),
.B(n_2597),
.Y(n_14680)
);

NAND2xp5_ASAP7_75t_L g14681 ( 
.A(n_14569),
.B(n_2597),
.Y(n_14681)
);

INVx1_ASAP7_75t_L g14682 ( 
.A(n_14572),
.Y(n_14682)
);

AND2x4_ASAP7_75t_L g14683 ( 
.A(n_14530),
.B(n_14542),
.Y(n_14683)
);

AND2x2_ASAP7_75t_L g14684 ( 
.A(n_14528),
.B(n_2598),
.Y(n_14684)
);

AND2x4_ASAP7_75t_L g14685 ( 
.A(n_14594),
.B(n_2598),
.Y(n_14685)
);

OR2x2_ASAP7_75t_L g14686 ( 
.A(n_14579),
.B(n_2599),
.Y(n_14686)
);

OR2x2_ASAP7_75t_L g14687 ( 
.A(n_14499),
.B(n_2599),
.Y(n_14687)
);

AND2x2_ASAP7_75t_L g14688 ( 
.A(n_14514),
.B(n_2600),
.Y(n_14688)
);

NAND2xp5_ASAP7_75t_L g14689 ( 
.A(n_14580),
.B(n_2600),
.Y(n_14689)
);

INVx2_ASAP7_75t_L g14690 ( 
.A(n_14537),
.Y(n_14690)
);

OR2x2_ASAP7_75t_L g14691 ( 
.A(n_14502),
.B(n_2601),
.Y(n_14691)
);

AND2x4_ASAP7_75t_L g14692 ( 
.A(n_14527),
.B(n_2601),
.Y(n_14692)
);

NAND2xp5_ASAP7_75t_L g14693 ( 
.A(n_14589),
.B(n_2602),
.Y(n_14693)
);

INVx1_ASAP7_75t_L g14694 ( 
.A(n_14595),
.Y(n_14694)
);

AND2x2_ASAP7_75t_L g14695 ( 
.A(n_14578),
.B(n_2602),
.Y(n_14695)
);

INVx1_ASAP7_75t_L g14696 ( 
.A(n_14604),
.Y(n_14696)
);

AND2x2_ASAP7_75t_L g14697 ( 
.A(n_14508),
.B(n_2603),
.Y(n_14697)
);

INVx1_ASAP7_75t_L g14698 ( 
.A(n_14606),
.Y(n_14698)
);

INVx1_ASAP7_75t_L g14699 ( 
.A(n_14535),
.Y(n_14699)
);

AND2x2_ASAP7_75t_L g14700 ( 
.A(n_14516),
.B(n_2604),
.Y(n_14700)
);

NAND2xp5_ASAP7_75t_L g14701 ( 
.A(n_14534),
.B(n_2604),
.Y(n_14701)
);

INVx1_ASAP7_75t_L g14702 ( 
.A(n_14605),
.Y(n_14702)
);

AND2x2_ASAP7_75t_L g14703 ( 
.A(n_14553),
.B(n_2605),
.Y(n_14703)
);

OR2x2_ASAP7_75t_L g14704 ( 
.A(n_14587),
.B(n_2605),
.Y(n_14704)
);

AND2x2_ASAP7_75t_L g14705 ( 
.A(n_14561),
.B(n_2606),
.Y(n_14705)
);

INVx1_ASAP7_75t_L g14706 ( 
.A(n_14576),
.Y(n_14706)
);

NAND2xp5_ASAP7_75t_L g14707 ( 
.A(n_14547),
.B(n_2606),
.Y(n_14707)
);

NOR2xp33_ASAP7_75t_L g14708 ( 
.A(n_14588),
.B(n_2607),
.Y(n_14708)
);

AND3x2_ASAP7_75t_L g14709 ( 
.A(n_14586),
.B(n_2608),
.C(n_2609),
.Y(n_14709)
);

AND2x2_ASAP7_75t_L g14710 ( 
.A(n_14597),
.B(n_2608),
.Y(n_14710)
);

INVx1_ASAP7_75t_L g14711 ( 
.A(n_14600),
.Y(n_14711)
);

OR2x6_ASAP7_75t_L g14712 ( 
.A(n_14596),
.B(n_14599),
.Y(n_14712)
);

INVx1_ASAP7_75t_L g14713 ( 
.A(n_14571),
.Y(n_14713)
);

INVx1_ASAP7_75t_L g14714 ( 
.A(n_14562),
.Y(n_14714)
);

OR2x2_ASAP7_75t_L g14715 ( 
.A(n_14570),
.B(n_2609),
.Y(n_14715)
);

AND2x2_ASAP7_75t_L g14716 ( 
.A(n_14575),
.B(n_2610),
.Y(n_14716)
);

INVx1_ASAP7_75t_L g14717 ( 
.A(n_14591),
.Y(n_14717)
);

AND2x4_ASAP7_75t_L g14718 ( 
.A(n_14548),
.B(n_2611),
.Y(n_14718)
);

AND2x4_ASAP7_75t_L g14719 ( 
.A(n_14548),
.B(n_2611),
.Y(n_14719)
);

INVxp67_ASAP7_75t_SL g14720 ( 
.A(n_14601),
.Y(n_14720)
);

AND2x4_ASAP7_75t_SL g14721 ( 
.A(n_14497),
.B(n_2612),
.Y(n_14721)
);

AND2x2_ASAP7_75t_L g14722 ( 
.A(n_14515),
.B(n_2612),
.Y(n_14722)
);

NAND2xp5_ASAP7_75t_L g14723 ( 
.A(n_14529),
.B(n_2613),
.Y(n_14723)
);

NAND2xp5_ASAP7_75t_L g14724 ( 
.A(n_14529),
.B(n_2613),
.Y(n_14724)
);

NAND3xp33_ASAP7_75t_L g14725 ( 
.A(n_14494),
.B(n_2614),
.C(n_2615),
.Y(n_14725)
);

INVx1_ASAP7_75t_L g14726 ( 
.A(n_14529),
.Y(n_14726)
);

INVx2_ASAP7_75t_L g14727 ( 
.A(n_14601),
.Y(n_14727)
);

INVx1_ASAP7_75t_L g14728 ( 
.A(n_14529),
.Y(n_14728)
);

INVx2_ASAP7_75t_L g14729 ( 
.A(n_14601),
.Y(n_14729)
);

OR2x2_ASAP7_75t_L g14730 ( 
.A(n_14529),
.B(n_2614),
.Y(n_14730)
);

OR2x6_ASAP7_75t_L g14731 ( 
.A(n_14496),
.B(n_2615),
.Y(n_14731)
);

AND2x4_ASAP7_75t_L g14732 ( 
.A(n_14607),
.B(n_2616),
.Y(n_14732)
);

NAND2xp5_ASAP7_75t_L g14733 ( 
.A(n_14612),
.B(n_2616),
.Y(n_14733)
);

AND2x2_ASAP7_75t_L g14734 ( 
.A(n_14630),
.B(n_2617),
.Y(n_14734)
);

NAND2xp5_ASAP7_75t_L g14735 ( 
.A(n_14632),
.B(n_2618),
.Y(n_14735)
);

NOR2x1p5_ASAP7_75t_L g14736 ( 
.A(n_14720),
.B(n_2619),
.Y(n_14736)
);

NAND2xp5_ASAP7_75t_L g14737 ( 
.A(n_14727),
.B(n_2619),
.Y(n_14737)
);

INVx1_ASAP7_75t_L g14738 ( 
.A(n_14634),
.Y(n_14738)
);

AND2x2_ASAP7_75t_L g14739 ( 
.A(n_14688),
.B(n_2620),
.Y(n_14739)
);

OR2x2_ASAP7_75t_L g14740 ( 
.A(n_14729),
.B(n_2621),
.Y(n_14740)
);

OR2x2_ASAP7_75t_L g14741 ( 
.A(n_14609),
.B(n_2621),
.Y(n_14741)
);

NAND2x1p5_ASAP7_75t_L g14742 ( 
.A(n_14638),
.B(n_2622),
.Y(n_14742)
);

INVx2_ASAP7_75t_L g14743 ( 
.A(n_14625),
.Y(n_14743)
);

AND2x2_ASAP7_75t_L g14744 ( 
.A(n_14619),
.B(n_2622),
.Y(n_14744)
);

AND2x4_ASAP7_75t_L g14745 ( 
.A(n_14726),
.B(n_2624),
.Y(n_14745)
);

AND2x2_ASAP7_75t_L g14746 ( 
.A(n_14641),
.B(n_2624),
.Y(n_14746)
);

NAND2xp5_ASAP7_75t_L g14747 ( 
.A(n_14728),
.B(n_2625),
.Y(n_14747)
);

INVx1_ASAP7_75t_L g14748 ( 
.A(n_14649),
.Y(n_14748)
);

AND2x2_ASAP7_75t_L g14749 ( 
.A(n_14722),
.B(n_14648),
.Y(n_14749)
);

AND2x2_ASAP7_75t_L g14750 ( 
.A(n_14669),
.B(n_14657),
.Y(n_14750)
);

INVx2_ASAP7_75t_L g14751 ( 
.A(n_14731),
.Y(n_14751)
);

OR2x2_ASAP7_75t_L g14752 ( 
.A(n_14615),
.B(n_2625),
.Y(n_14752)
);

OR2x2_ASAP7_75t_L g14753 ( 
.A(n_14730),
.B(n_2626),
.Y(n_14753)
);

OR2x2_ASAP7_75t_L g14754 ( 
.A(n_14613),
.B(n_2626),
.Y(n_14754)
);

OR2x2_ASAP7_75t_L g14755 ( 
.A(n_14715),
.B(n_2627),
.Y(n_14755)
);

INVx2_ASAP7_75t_L g14756 ( 
.A(n_14731),
.Y(n_14756)
);

INVx2_ASAP7_75t_SL g14757 ( 
.A(n_14721),
.Y(n_14757)
);

INVx1_ASAP7_75t_L g14758 ( 
.A(n_14610),
.Y(n_14758)
);

INVx2_ASAP7_75t_L g14759 ( 
.A(n_14608),
.Y(n_14759)
);

AND2x4_ASAP7_75t_L g14760 ( 
.A(n_14667),
.B(n_14626),
.Y(n_14760)
);

HB1xp67_ASAP7_75t_L g14761 ( 
.A(n_14608),
.Y(n_14761)
);

NAND2xp5_ASAP7_75t_L g14762 ( 
.A(n_14629),
.B(n_2627),
.Y(n_14762)
);

BUFx2_ASAP7_75t_L g14763 ( 
.A(n_14661),
.Y(n_14763)
);

NOR2xp33_ASAP7_75t_L g14764 ( 
.A(n_14616),
.B(n_14617),
.Y(n_14764)
);

INVx1_ASAP7_75t_L g14765 ( 
.A(n_14631),
.Y(n_14765)
);

INVx1_ASAP7_75t_L g14766 ( 
.A(n_14700),
.Y(n_14766)
);

NOR2xp33_ASAP7_75t_L g14767 ( 
.A(n_14636),
.B(n_14621),
.Y(n_14767)
);

NAND2xp5_ASAP7_75t_L g14768 ( 
.A(n_14709),
.B(n_2628),
.Y(n_14768)
);

AOI32xp33_ASAP7_75t_L g14769 ( 
.A1(n_14697),
.A2(n_2630),
.A3(n_2628),
.B1(n_2629),
.B2(n_2631),
.Y(n_14769)
);

AND2x2_ASAP7_75t_L g14770 ( 
.A(n_14645),
.B(n_2629),
.Y(n_14770)
);

AND2x2_ASAP7_75t_L g14771 ( 
.A(n_14655),
.B(n_2630),
.Y(n_14771)
);

OR2x2_ASAP7_75t_L g14772 ( 
.A(n_14723),
.B(n_2631),
.Y(n_14772)
);

INVx1_ASAP7_75t_L g14773 ( 
.A(n_14656),
.Y(n_14773)
);

AND2x2_ASAP7_75t_L g14774 ( 
.A(n_14695),
.B(n_2632),
.Y(n_14774)
);

AOI22xp5_ASAP7_75t_L g14775 ( 
.A1(n_14708),
.A2(n_2634),
.B1(n_2632),
.B2(n_2633),
.Y(n_14775)
);

INVx1_ASAP7_75t_L g14776 ( 
.A(n_14627),
.Y(n_14776)
);

AND2x4_ASAP7_75t_L g14777 ( 
.A(n_14674),
.B(n_14678),
.Y(n_14777)
);

INVx1_ASAP7_75t_L g14778 ( 
.A(n_14635),
.Y(n_14778)
);

INVx1_ASAP7_75t_L g14779 ( 
.A(n_14724),
.Y(n_14779)
);

INVx1_ASAP7_75t_L g14780 ( 
.A(n_14646),
.Y(n_14780)
);

INVx2_ASAP7_75t_SL g14781 ( 
.A(n_14622),
.Y(n_14781)
);

NAND2xp5_ASAP7_75t_SL g14782 ( 
.A(n_14668),
.B(n_2633),
.Y(n_14782)
);

OR2x2_ASAP7_75t_L g14783 ( 
.A(n_14624),
.B(n_2634),
.Y(n_14783)
);

AND2x2_ASAP7_75t_L g14784 ( 
.A(n_14652),
.B(n_2635),
.Y(n_14784)
);

INVx1_ASAP7_75t_L g14785 ( 
.A(n_14718),
.Y(n_14785)
);

INVx1_ASAP7_75t_L g14786 ( 
.A(n_14719),
.Y(n_14786)
);

INVx1_ASAP7_75t_L g14787 ( 
.A(n_14684),
.Y(n_14787)
);

INVx1_ASAP7_75t_L g14788 ( 
.A(n_14676),
.Y(n_14788)
);

AND2x2_ASAP7_75t_L g14789 ( 
.A(n_14698),
.B(n_2635),
.Y(n_14789)
);

NAND2xp5_ASAP7_75t_L g14790 ( 
.A(n_14702),
.B(n_2636),
.Y(n_14790)
);

OR2x2_ASAP7_75t_L g14791 ( 
.A(n_14650),
.B(n_2636),
.Y(n_14791)
);

AND2x2_ASAP7_75t_L g14792 ( 
.A(n_14665),
.B(n_2637),
.Y(n_14792)
);

INVxp67_ASAP7_75t_L g14793 ( 
.A(n_14637),
.Y(n_14793)
);

INVx2_ASAP7_75t_L g14794 ( 
.A(n_14633),
.Y(n_14794)
);

INVx1_ASAP7_75t_L g14795 ( 
.A(n_14639),
.Y(n_14795)
);

INVxp67_ASAP7_75t_L g14796 ( 
.A(n_14675),
.Y(n_14796)
);

INVx1_ASAP7_75t_L g14797 ( 
.A(n_14643),
.Y(n_14797)
);

INVxp67_ASAP7_75t_SL g14798 ( 
.A(n_14690),
.Y(n_14798)
);

INVx1_ASAP7_75t_L g14799 ( 
.A(n_14662),
.Y(n_14799)
);

INVx1_ASAP7_75t_L g14800 ( 
.A(n_14672),
.Y(n_14800)
);

OR2x6_ASAP7_75t_L g14801 ( 
.A(n_14618),
.B(n_2637),
.Y(n_14801)
);

NAND2xp5_ASAP7_75t_L g14802 ( 
.A(n_14660),
.B(n_2638),
.Y(n_14802)
);

INVx1_ASAP7_75t_L g14803 ( 
.A(n_14640),
.Y(n_14803)
);

AND2x2_ASAP7_75t_L g14804 ( 
.A(n_14671),
.B(n_2639),
.Y(n_14804)
);

INVx1_ASAP7_75t_L g14805 ( 
.A(n_14705),
.Y(n_14805)
);

NAND2xp5_ASAP7_75t_L g14806 ( 
.A(n_14614),
.B(n_2640),
.Y(n_14806)
);

INVxp67_ASAP7_75t_L g14807 ( 
.A(n_14664),
.Y(n_14807)
);

INVx1_ASAP7_75t_L g14808 ( 
.A(n_14611),
.Y(n_14808)
);

BUFx2_ASAP7_75t_L g14809 ( 
.A(n_14712),
.Y(n_14809)
);

AND2x2_ASAP7_75t_L g14810 ( 
.A(n_14682),
.B(n_2640),
.Y(n_14810)
);

OR2x2_ASAP7_75t_L g14811 ( 
.A(n_14687),
.B(n_2641),
.Y(n_14811)
);

OR2x2_ASAP7_75t_L g14812 ( 
.A(n_14663),
.B(n_2641),
.Y(n_14812)
);

AOI211xp5_ASAP7_75t_L g14813 ( 
.A1(n_14647),
.A2(n_2645),
.B(n_2642),
.C(n_2643),
.Y(n_14813)
);

INVx2_ASAP7_75t_L g14814 ( 
.A(n_14654),
.Y(n_14814)
);

AND2x2_ASAP7_75t_L g14815 ( 
.A(n_14623),
.B(n_2643),
.Y(n_14815)
);

INVx1_ASAP7_75t_L g14816 ( 
.A(n_14651),
.Y(n_14816)
);

OR2x2_ASAP7_75t_L g14817 ( 
.A(n_14704),
.B(n_2645),
.Y(n_14817)
);

INVx1_ASAP7_75t_L g14818 ( 
.A(n_14658),
.Y(n_14818)
);

AND2x2_ASAP7_75t_L g14819 ( 
.A(n_14714),
.B(n_2646),
.Y(n_14819)
);

INVx1_ASAP7_75t_L g14820 ( 
.A(n_14644),
.Y(n_14820)
);

AND2x2_ASAP7_75t_SL g14821 ( 
.A(n_14683),
.B(n_14620),
.Y(n_14821)
);

INVx1_ASAP7_75t_L g14822 ( 
.A(n_14653),
.Y(n_14822)
);

HB1xp67_ASAP7_75t_L g14823 ( 
.A(n_14712),
.Y(n_14823)
);

OR2x2_ASAP7_75t_L g14824 ( 
.A(n_14696),
.B(n_2646),
.Y(n_14824)
);

NAND2xp5_ASAP7_75t_L g14825 ( 
.A(n_14685),
.B(n_2647),
.Y(n_14825)
);

NAND2xp5_ASAP7_75t_L g14826 ( 
.A(n_14692),
.B(n_2647),
.Y(n_14826)
);

AND2x2_ASAP7_75t_L g14827 ( 
.A(n_14706),
.B(n_2648),
.Y(n_14827)
);

INVx1_ASAP7_75t_L g14828 ( 
.A(n_14642),
.Y(n_14828)
);

OR2x2_ASAP7_75t_L g14829 ( 
.A(n_14628),
.B(n_2648),
.Y(n_14829)
);

INVx1_ASAP7_75t_L g14830 ( 
.A(n_14680),
.Y(n_14830)
);

AND2x2_ASAP7_75t_L g14831 ( 
.A(n_14703),
.B(n_2649),
.Y(n_14831)
);

INVx1_ASAP7_75t_L g14832 ( 
.A(n_14710),
.Y(n_14832)
);

INVx1_ASAP7_75t_L g14833 ( 
.A(n_14691),
.Y(n_14833)
);

NAND2xp5_ASAP7_75t_L g14834 ( 
.A(n_14659),
.B(n_2649),
.Y(n_14834)
);

INVx3_ASAP7_75t_L g14835 ( 
.A(n_14677),
.Y(n_14835)
);

INVx1_ASAP7_75t_L g14836 ( 
.A(n_14689),
.Y(n_14836)
);

INVx1_ASAP7_75t_L g14837 ( 
.A(n_14666),
.Y(n_14837)
);

AND2x2_ASAP7_75t_L g14838 ( 
.A(n_14713),
.B(n_14716),
.Y(n_14838)
);

INVx2_ASAP7_75t_L g14839 ( 
.A(n_14686),
.Y(n_14839)
);

NAND2xp5_ASAP7_75t_L g14840 ( 
.A(n_14694),
.B(n_2651),
.Y(n_14840)
);

BUFx2_ASAP7_75t_L g14841 ( 
.A(n_14673),
.Y(n_14841)
);

NAND2xp5_ASAP7_75t_L g14842 ( 
.A(n_14670),
.B(n_2651),
.Y(n_14842)
);

INVx2_ASAP7_75t_L g14843 ( 
.A(n_14699),
.Y(n_14843)
);

AND2x2_ASAP7_75t_L g14844 ( 
.A(n_14717),
.B(n_2652),
.Y(n_14844)
);

INVx1_ASAP7_75t_L g14845 ( 
.A(n_14679),
.Y(n_14845)
);

OR2x6_ASAP7_75t_L g14846 ( 
.A(n_14693),
.B(n_14681),
.Y(n_14846)
);

INVx1_ASAP7_75t_L g14847 ( 
.A(n_14701),
.Y(n_14847)
);

OR2x2_ASAP7_75t_L g14848 ( 
.A(n_14725),
.B(n_2653),
.Y(n_14848)
);

INVx2_ASAP7_75t_SL g14849 ( 
.A(n_14711),
.Y(n_14849)
);

INVx1_ASAP7_75t_L g14850 ( 
.A(n_14707),
.Y(n_14850)
);

NAND5xp2_ASAP7_75t_L g14851 ( 
.A(n_14609),
.B(n_2655),
.C(n_2653),
.D(n_2654),
.E(n_2656),
.Y(n_14851)
);

OR2x2_ASAP7_75t_L g14852 ( 
.A(n_14607),
.B(n_2654),
.Y(n_14852)
);

BUFx2_ASAP7_75t_L g14853 ( 
.A(n_14731),
.Y(n_14853)
);

NAND2xp5_ASAP7_75t_L g14854 ( 
.A(n_14612),
.B(n_2656),
.Y(n_14854)
);

INVx1_ASAP7_75t_L g14855 ( 
.A(n_14634),
.Y(n_14855)
);

OAI22xp5_ASAP7_75t_L g14856 ( 
.A1(n_14638),
.A2(n_2660),
.B1(n_2657),
.B2(n_2658),
.Y(n_14856)
);

INVx2_ASAP7_75t_L g14857 ( 
.A(n_14607),
.Y(n_14857)
);

AND2x2_ASAP7_75t_L g14858 ( 
.A(n_14630),
.B(n_2657),
.Y(n_14858)
);

AND2x2_ASAP7_75t_L g14859 ( 
.A(n_14630),
.B(n_2658),
.Y(n_14859)
);

AND2x2_ASAP7_75t_L g14860 ( 
.A(n_14630),
.B(n_2660),
.Y(n_14860)
);

NOR2xp33_ASAP7_75t_L g14861 ( 
.A(n_14607),
.B(n_2661),
.Y(n_14861)
);

NAND2x1p5_ASAP7_75t_L g14862 ( 
.A(n_14607),
.B(n_2661),
.Y(n_14862)
);

INVx2_ASAP7_75t_L g14863 ( 
.A(n_14607),
.Y(n_14863)
);

AND2x2_ASAP7_75t_L g14864 ( 
.A(n_14630),
.B(n_2663),
.Y(n_14864)
);

NOR2xp33_ASAP7_75t_SL g14865 ( 
.A(n_14720),
.B(n_2663),
.Y(n_14865)
);

NAND2xp5_ASAP7_75t_L g14866 ( 
.A(n_14612),
.B(n_2664),
.Y(n_14866)
);

NAND2xp5_ASAP7_75t_L g14867 ( 
.A(n_14612),
.B(n_2665),
.Y(n_14867)
);

INVx2_ASAP7_75t_L g14868 ( 
.A(n_14607),
.Y(n_14868)
);

INVx1_ASAP7_75t_L g14869 ( 
.A(n_14634),
.Y(n_14869)
);

NAND2xp5_ASAP7_75t_L g14870 ( 
.A(n_14612),
.B(n_2666),
.Y(n_14870)
);

INVx2_ASAP7_75t_L g14871 ( 
.A(n_14607),
.Y(n_14871)
);

NAND3xp33_ASAP7_75t_L g14872 ( 
.A(n_14708),
.B(n_2666),
.C(n_2667),
.Y(n_14872)
);

INVxp67_ASAP7_75t_SL g14873 ( 
.A(n_14634),
.Y(n_14873)
);

AND2x2_ASAP7_75t_L g14874 ( 
.A(n_14630),
.B(n_2667),
.Y(n_14874)
);

INVx1_ASAP7_75t_L g14875 ( 
.A(n_14634),
.Y(n_14875)
);

INVx1_ASAP7_75t_SL g14876 ( 
.A(n_14688),
.Y(n_14876)
);

NAND2xp5_ASAP7_75t_L g14877 ( 
.A(n_14612),
.B(n_2668),
.Y(n_14877)
);

AND2x2_ASAP7_75t_L g14878 ( 
.A(n_14630),
.B(n_2669),
.Y(n_14878)
);

INVxp67_ASAP7_75t_L g14879 ( 
.A(n_14634),
.Y(n_14879)
);

AND2x2_ASAP7_75t_L g14880 ( 
.A(n_14630),
.B(n_2669),
.Y(n_14880)
);

AND2x4_ASAP7_75t_L g14881 ( 
.A(n_14607),
.B(n_2670),
.Y(n_14881)
);

INVx2_ASAP7_75t_L g14882 ( 
.A(n_14742),
.Y(n_14882)
);

OR2x2_ASAP7_75t_L g14883 ( 
.A(n_14862),
.B(n_14853),
.Y(n_14883)
);

INVx2_ASAP7_75t_L g14884 ( 
.A(n_14736),
.Y(n_14884)
);

INVxp67_ASAP7_75t_SL g14885 ( 
.A(n_14823),
.Y(n_14885)
);

OR2x2_ASAP7_75t_L g14886 ( 
.A(n_14757),
.B(n_2670),
.Y(n_14886)
);

CKINVDCx14_ASAP7_75t_R g14887 ( 
.A(n_14809),
.Y(n_14887)
);

INVx1_ASAP7_75t_L g14888 ( 
.A(n_14744),
.Y(n_14888)
);

OR2x2_ASAP7_75t_L g14889 ( 
.A(n_14876),
.B(n_2671),
.Y(n_14889)
);

INVx1_ASAP7_75t_L g14890 ( 
.A(n_14763),
.Y(n_14890)
);

INVx1_ASAP7_75t_L g14891 ( 
.A(n_14739),
.Y(n_14891)
);

INVx1_ASAP7_75t_L g14892 ( 
.A(n_14740),
.Y(n_14892)
);

NAND2xp5_ASAP7_75t_L g14893 ( 
.A(n_14732),
.B(n_2672),
.Y(n_14893)
);

INVx1_ASAP7_75t_L g14894 ( 
.A(n_14852),
.Y(n_14894)
);

AND2x2_ASAP7_75t_L g14895 ( 
.A(n_14749),
.B(n_2672),
.Y(n_14895)
);

NAND2xp5_ASAP7_75t_L g14896 ( 
.A(n_14881),
.B(n_2673),
.Y(n_14896)
);

NAND2xp5_ASAP7_75t_L g14897 ( 
.A(n_14781),
.B(n_14857),
.Y(n_14897)
);

NAND2xp5_ASAP7_75t_L g14898 ( 
.A(n_14863),
.B(n_2674),
.Y(n_14898)
);

NAND2xp5_ASAP7_75t_L g14899 ( 
.A(n_14868),
.B(n_2674),
.Y(n_14899)
);

OR2x2_ASAP7_75t_L g14900 ( 
.A(n_14871),
.B(n_2675),
.Y(n_14900)
);

OR2x2_ASAP7_75t_L g14901 ( 
.A(n_14751),
.B(n_2675),
.Y(n_14901)
);

INVx1_ASAP7_75t_L g14902 ( 
.A(n_14746),
.Y(n_14902)
);

INVx2_ASAP7_75t_L g14903 ( 
.A(n_14821),
.Y(n_14903)
);

INVx1_ASAP7_75t_L g14904 ( 
.A(n_14734),
.Y(n_14904)
);

INVxp67_ASAP7_75t_L g14905 ( 
.A(n_14865),
.Y(n_14905)
);

INVx1_ASAP7_75t_L g14906 ( 
.A(n_14858),
.Y(n_14906)
);

INVx1_ASAP7_75t_L g14907 ( 
.A(n_14859),
.Y(n_14907)
);

INVx2_ASAP7_75t_L g14908 ( 
.A(n_14756),
.Y(n_14908)
);

AND2x2_ASAP7_75t_L g14909 ( 
.A(n_14750),
.B(n_2676),
.Y(n_14909)
);

AND2x2_ASAP7_75t_L g14910 ( 
.A(n_14774),
.B(n_2676),
.Y(n_14910)
);

OR2x2_ASAP7_75t_L g14911 ( 
.A(n_14752),
.B(n_2677),
.Y(n_14911)
);

AND2x2_ASAP7_75t_L g14912 ( 
.A(n_14743),
.B(n_2677),
.Y(n_14912)
);

INVx2_ASAP7_75t_L g14913 ( 
.A(n_14801),
.Y(n_14913)
);

INVx1_ASAP7_75t_SL g14914 ( 
.A(n_14860),
.Y(n_14914)
);

INVxp67_ASAP7_75t_SL g14915 ( 
.A(n_14761),
.Y(n_14915)
);

INVx2_ASAP7_75t_L g14916 ( 
.A(n_14801),
.Y(n_14916)
);

INVx1_ASAP7_75t_L g14917 ( 
.A(n_14864),
.Y(n_14917)
);

OR2x2_ASAP7_75t_L g14918 ( 
.A(n_14754),
.B(n_2678),
.Y(n_14918)
);

INVx1_ASAP7_75t_L g14919 ( 
.A(n_14874),
.Y(n_14919)
);

OR2x2_ASAP7_75t_L g14920 ( 
.A(n_14737),
.B(n_2679),
.Y(n_14920)
);

INVx1_ASAP7_75t_L g14921 ( 
.A(n_14878),
.Y(n_14921)
);

INVx1_ASAP7_75t_L g14922 ( 
.A(n_14880),
.Y(n_14922)
);

AND2x4_ASAP7_75t_L g14923 ( 
.A(n_14760),
.B(n_2679),
.Y(n_14923)
);

INVx2_ASAP7_75t_SL g14924 ( 
.A(n_14745),
.Y(n_14924)
);

NAND2xp5_ASAP7_75t_L g14925 ( 
.A(n_14777),
.B(n_14773),
.Y(n_14925)
);

INVx1_ASAP7_75t_L g14926 ( 
.A(n_14873),
.Y(n_14926)
);

INVx1_ASAP7_75t_L g14927 ( 
.A(n_14753),
.Y(n_14927)
);

INVx2_ASAP7_75t_L g14928 ( 
.A(n_14817),
.Y(n_14928)
);

INVxp67_ASAP7_75t_SL g14929 ( 
.A(n_14879),
.Y(n_14929)
);

AND2x2_ASAP7_75t_L g14930 ( 
.A(n_14819),
.B(n_2681),
.Y(n_14930)
);

INVx2_ASAP7_75t_L g14931 ( 
.A(n_14812),
.Y(n_14931)
);

INVx1_ASAP7_75t_L g14932 ( 
.A(n_14770),
.Y(n_14932)
);

NAND2x1p5_ASAP7_75t_L g14933 ( 
.A(n_14835),
.B(n_2681),
.Y(n_14933)
);

INVx1_ASAP7_75t_L g14934 ( 
.A(n_14771),
.Y(n_14934)
);

OR2x2_ASAP7_75t_SL g14935 ( 
.A(n_14759),
.B(n_2682),
.Y(n_14935)
);

OR2x2_ASAP7_75t_L g14936 ( 
.A(n_14766),
.B(n_2682),
.Y(n_14936)
);

INVxp67_ASAP7_75t_L g14937 ( 
.A(n_14851),
.Y(n_14937)
);

INVx2_ASAP7_75t_L g14938 ( 
.A(n_14791),
.Y(n_14938)
);

INVx1_ASAP7_75t_L g14939 ( 
.A(n_14784),
.Y(n_14939)
);

INVx1_ASAP7_75t_L g14940 ( 
.A(n_14824),
.Y(n_14940)
);

AND2x2_ASAP7_75t_L g14941 ( 
.A(n_14785),
.B(n_2683),
.Y(n_14941)
);

NAND2xp5_ASAP7_75t_L g14942 ( 
.A(n_14786),
.B(n_14861),
.Y(n_14942)
);

AND2x2_ASAP7_75t_L g14943 ( 
.A(n_14803),
.B(n_2683),
.Y(n_14943)
);

INVx1_ASAP7_75t_L g14944 ( 
.A(n_14741),
.Y(n_14944)
);

BUFx2_ASAP7_75t_L g14945 ( 
.A(n_14798),
.Y(n_14945)
);

AND2x2_ASAP7_75t_L g14946 ( 
.A(n_14816),
.B(n_2684),
.Y(n_14946)
);

INVxp67_ASAP7_75t_L g14947 ( 
.A(n_14764),
.Y(n_14947)
);

OR2x2_ASAP7_75t_L g14948 ( 
.A(n_14768),
.B(n_2686),
.Y(n_14948)
);

AND2x2_ASAP7_75t_L g14949 ( 
.A(n_14818),
.B(n_2686),
.Y(n_14949)
);

NOR2x1p5_ASAP7_75t_SL g14950 ( 
.A(n_14738),
.B(n_2687),
.Y(n_14950)
);

NAND2xp5_ASAP7_75t_L g14951 ( 
.A(n_14828),
.B(n_2687),
.Y(n_14951)
);

INVx1_ASAP7_75t_L g14952 ( 
.A(n_14789),
.Y(n_14952)
);

AND2x2_ASAP7_75t_L g14953 ( 
.A(n_14844),
.B(n_2688),
.Y(n_14953)
);

INVx1_ASAP7_75t_L g14954 ( 
.A(n_14815),
.Y(n_14954)
);

NAND2xp5_ASAP7_75t_L g14955 ( 
.A(n_14778),
.B(n_2688),
.Y(n_14955)
);

INVx2_ASAP7_75t_L g14956 ( 
.A(n_14811),
.Y(n_14956)
);

AND2x2_ASAP7_75t_L g14957 ( 
.A(n_14838),
.B(n_2689),
.Y(n_14957)
);

INVx1_ASAP7_75t_L g14958 ( 
.A(n_14827),
.Y(n_14958)
);

A2O1A1Ixp33_ASAP7_75t_L g14959 ( 
.A1(n_14767),
.A2(n_2691),
.B(n_2689),
.C(n_2690),
.Y(n_14959)
);

AND2x2_ASAP7_75t_L g14960 ( 
.A(n_14765),
.B(n_2690),
.Y(n_14960)
);

OAI21xp33_ASAP7_75t_L g14961 ( 
.A1(n_14807),
.A2(n_14788),
.B(n_14780),
.Y(n_14961)
);

INVx2_ASAP7_75t_L g14962 ( 
.A(n_14831),
.Y(n_14962)
);

NOR2x1_ASAP7_75t_L g14963 ( 
.A(n_14855),
.B(n_2691),
.Y(n_14963)
);

AND2x2_ASAP7_75t_L g14964 ( 
.A(n_14787),
.B(n_2692),
.Y(n_14964)
);

NAND2xp5_ASAP7_75t_L g14965 ( 
.A(n_14792),
.B(n_2692),
.Y(n_14965)
);

OAI21xp33_ASAP7_75t_L g14966 ( 
.A1(n_14850),
.A2(n_2693),
.B(n_2694),
.Y(n_14966)
);

INVxp67_ASAP7_75t_SL g14967 ( 
.A(n_14869),
.Y(n_14967)
);

OR2x2_ASAP7_75t_L g14968 ( 
.A(n_14735),
.B(n_2694),
.Y(n_14968)
);

NAND2xp5_ASAP7_75t_L g14969 ( 
.A(n_14804),
.B(n_2695),
.Y(n_14969)
);

OR2x2_ASAP7_75t_L g14970 ( 
.A(n_14755),
.B(n_2696),
.Y(n_14970)
);

INVx1_ASAP7_75t_L g14971 ( 
.A(n_14810),
.Y(n_14971)
);

INVx1_ASAP7_75t_L g14972 ( 
.A(n_14733),
.Y(n_14972)
);

NAND2x1_ASAP7_75t_L g14973 ( 
.A(n_14748),
.B(n_14875),
.Y(n_14973)
);

INVxp67_ASAP7_75t_L g14974 ( 
.A(n_14854),
.Y(n_14974)
);

OR2x2_ASAP7_75t_L g14975 ( 
.A(n_14866),
.B(n_2696),
.Y(n_14975)
);

INVx2_ASAP7_75t_L g14976 ( 
.A(n_14783),
.Y(n_14976)
);

BUFx2_ASAP7_75t_L g14977 ( 
.A(n_14758),
.Y(n_14977)
);

OR2x2_ASAP7_75t_L g14978 ( 
.A(n_14867),
.B(n_2697),
.Y(n_14978)
);

NAND2xp5_ASAP7_75t_L g14979 ( 
.A(n_14769),
.B(n_2697),
.Y(n_14979)
);

INVx2_ASAP7_75t_L g14980 ( 
.A(n_14772),
.Y(n_14980)
);

NAND2xp5_ASAP7_75t_L g14981 ( 
.A(n_14805),
.B(n_2698),
.Y(n_14981)
);

NAND2xp5_ASAP7_75t_L g14982 ( 
.A(n_14832),
.B(n_2698),
.Y(n_14982)
);

NAND2xp5_ASAP7_75t_L g14983 ( 
.A(n_14776),
.B(n_2700),
.Y(n_14983)
);

INVx3_ASAP7_75t_L g14984 ( 
.A(n_14794),
.Y(n_14984)
);

INVx1_ASAP7_75t_L g14985 ( 
.A(n_14870),
.Y(n_14985)
);

NOR2x1p5_ASAP7_75t_L g14986 ( 
.A(n_14762),
.B(n_2700),
.Y(n_14986)
);

CKINVDCx5p33_ASAP7_75t_R g14987 ( 
.A(n_14846),
.Y(n_14987)
);

NAND2x1p5_ASAP7_75t_L g14988 ( 
.A(n_14795),
.B(n_2701),
.Y(n_14988)
);

INVx1_ASAP7_75t_L g14989 ( 
.A(n_14877),
.Y(n_14989)
);

AOI211xp5_ASAP7_75t_L g14990 ( 
.A1(n_14808),
.A2(n_2704),
.B(n_2702),
.C(n_2703),
.Y(n_14990)
);

AND2x2_ASAP7_75t_L g14991 ( 
.A(n_14814),
.B(n_2703),
.Y(n_14991)
);

INVx1_ASAP7_75t_L g14992 ( 
.A(n_14790),
.Y(n_14992)
);

INVxp67_ASAP7_75t_L g14993 ( 
.A(n_14802),
.Y(n_14993)
);

INVx2_ASAP7_75t_L g14994 ( 
.A(n_14829),
.Y(n_14994)
);

INVx1_ASAP7_75t_L g14995 ( 
.A(n_14826),
.Y(n_14995)
);

AND2x2_ASAP7_75t_L g14996 ( 
.A(n_14799),
.B(n_2704),
.Y(n_14996)
);

NAND2xp5_ASAP7_75t_L g14997 ( 
.A(n_14800),
.B(n_14830),
.Y(n_14997)
);

INVx1_ASAP7_75t_L g14998 ( 
.A(n_14825),
.Y(n_14998)
);

AND2x2_ASAP7_75t_L g14999 ( 
.A(n_14793),
.B(n_2705),
.Y(n_14999)
);

AOI22xp5_ASAP7_75t_L g15000 ( 
.A1(n_14796),
.A2(n_2707),
.B1(n_2705),
.B2(n_2706),
.Y(n_15000)
);

INVx1_ASAP7_75t_L g15001 ( 
.A(n_14848),
.Y(n_15001)
);

HB1xp67_ASAP7_75t_L g15002 ( 
.A(n_14856),
.Y(n_15002)
);

INVxp67_ASAP7_75t_L g15003 ( 
.A(n_14782),
.Y(n_15003)
);

AND2x2_ASAP7_75t_L g15004 ( 
.A(n_14797),
.B(n_14839),
.Y(n_15004)
);

INVx1_ASAP7_75t_L g15005 ( 
.A(n_14747),
.Y(n_15005)
);

NAND2xp5_ASAP7_75t_L g15006 ( 
.A(n_14833),
.B(n_2706),
.Y(n_15006)
);

INVx1_ASAP7_75t_L g15007 ( 
.A(n_14806),
.Y(n_15007)
);

AND2x2_ASAP7_75t_L g15008 ( 
.A(n_14846),
.B(n_2707),
.Y(n_15008)
);

AND2x4_ASAP7_75t_SL g15009 ( 
.A(n_14843),
.B(n_2710),
.Y(n_15009)
);

INVx1_ASAP7_75t_L g15010 ( 
.A(n_14834),
.Y(n_15010)
);

OR2x2_ASAP7_75t_L g15011 ( 
.A(n_14840),
.B(n_2711),
.Y(n_15011)
);

NAND2xp5_ASAP7_75t_L g15012 ( 
.A(n_14775),
.B(n_14813),
.Y(n_15012)
);

INVx1_ASAP7_75t_L g15013 ( 
.A(n_14842),
.Y(n_15013)
);

AND2x2_ASAP7_75t_L g15014 ( 
.A(n_14841),
.B(n_2711),
.Y(n_15014)
);

OAI21xp5_ASAP7_75t_L g15015 ( 
.A1(n_14872),
.A2(n_2712),
.B(n_2713),
.Y(n_15015)
);

INVx2_ASAP7_75t_SL g15016 ( 
.A(n_14849),
.Y(n_15016)
);

OR2x2_ASAP7_75t_L g15017 ( 
.A(n_14820),
.B(n_2712),
.Y(n_15017)
);

NAND2xp5_ASAP7_75t_L g15018 ( 
.A(n_14822),
.B(n_2713),
.Y(n_15018)
);

INVx1_ASAP7_75t_L g15019 ( 
.A(n_14836),
.Y(n_15019)
);

INVx1_ASAP7_75t_L g15020 ( 
.A(n_14779),
.Y(n_15020)
);

OR2x2_ASAP7_75t_L g15021 ( 
.A(n_14847),
.B(n_14845),
.Y(n_15021)
);

INVx2_ASAP7_75t_L g15022 ( 
.A(n_14837),
.Y(n_15022)
);

AND2x2_ASAP7_75t_L g15023 ( 
.A(n_14757),
.B(n_2714),
.Y(n_15023)
);

AND2x2_ASAP7_75t_L g15024 ( 
.A(n_14757),
.B(n_2714),
.Y(n_15024)
);

INVx1_ASAP7_75t_L g15025 ( 
.A(n_14950),
.Y(n_15025)
);

OR2x2_ASAP7_75t_L g15026 ( 
.A(n_14935),
.B(n_2715),
.Y(n_15026)
);

AOI22xp33_ASAP7_75t_L g15027 ( 
.A1(n_14887),
.A2(n_2717),
.B1(n_2715),
.B2(n_2716),
.Y(n_15027)
);

INVx1_ASAP7_75t_L g15028 ( 
.A(n_14885),
.Y(n_15028)
);

INVx1_ASAP7_75t_L g15029 ( 
.A(n_14925),
.Y(n_15029)
);

OAI22xp5_ASAP7_75t_L g15030 ( 
.A1(n_14915),
.A2(n_2718),
.B1(n_2716),
.B2(n_2717),
.Y(n_15030)
);

NAND2xp5_ASAP7_75t_L g15031 ( 
.A(n_14923),
.B(n_2718),
.Y(n_15031)
);

INVx1_ASAP7_75t_L g15032 ( 
.A(n_14933),
.Y(n_15032)
);

NAND2xp5_ASAP7_75t_L g15033 ( 
.A(n_15023),
.B(n_2719),
.Y(n_15033)
);

INVx2_ASAP7_75t_L g15034 ( 
.A(n_14988),
.Y(n_15034)
);

INVxp67_ASAP7_75t_L g15035 ( 
.A(n_15024),
.Y(n_15035)
);

AND2x2_ASAP7_75t_L g15036 ( 
.A(n_14903),
.B(n_2719),
.Y(n_15036)
);

NOR3xp33_ASAP7_75t_L g15037 ( 
.A(n_14961),
.B(n_2720),
.C(n_2721),
.Y(n_15037)
);

INVx2_ASAP7_75t_SL g15038 ( 
.A(n_15009),
.Y(n_15038)
);

INVx2_ASAP7_75t_L g15039 ( 
.A(n_14886),
.Y(n_15039)
);

INVx1_ASAP7_75t_L g15040 ( 
.A(n_14895),
.Y(n_15040)
);

HB1xp67_ASAP7_75t_L g15041 ( 
.A(n_14963),
.Y(n_15041)
);

NAND2xp5_ASAP7_75t_L g15042 ( 
.A(n_14914),
.B(n_2720),
.Y(n_15042)
);

NAND3xp33_ASAP7_75t_SL g15043 ( 
.A(n_14987),
.B(n_2721),
.C(n_2722),
.Y(n_15043)
);

AND2x2_ASAP7_75t_L g15044 ( 
.A(n_14884),
.B(n_2722),
.Y(n_15044)
);

INVxp67_ASAP7_75t_L g15045 ( 
.A(n_14909),
.Y(n_15045)
);

INVxp67_ASAP7_75t_L g15046 ( 
.A(n_14945),
.Y(n_15046)
);

INVx1_ASAP7_75t_L g15047 ( 
.A(n_14957),
.Y(n_15047)
);

INVx2_ASAP7_75t_SL g15048 ( 
.A(n_14883),
.Y(n_15048)
);

INVx2_ASAP7_75t_L g15049 ( 
.A(n_14918),
.Y(n_15049)
);

OR2x2_ASAP7_75t_L g15050 ( 
.A(n_14882),
.B(n_2724),
.Y(n_15050)
);

AND3x2_ASAP7_75t_L g15051 ( 
.A(n_14990),
.B(n_2724),
.C(n_2725),
.Y(n_15051)
);

AOI32xp33_ASAP7_75t_L g15052 ( 
.A1(n_14890),
.A2(n_2727),
.A3(n_2725),
.B1(n_2726),
.B2(n_2728),
.Y(n_15052)
);

AOI22xp33_ASAP7_75t_L g15053 ( 
.A1(n_15016),
.A2(n_2731),
.B1(n_2729),
.B2(n_2730),
.Y(n_15053)
);

INVx1_ASAP7_75t_L g15054 ( 
.A(n_14941),
.Y(n_15054)
);

INVx1_ASAP7_75t_L g15055 ( 
.A(n_14943),
.Y(n_15055)
);

INVx2_ASAP7_75t_SL g15056 ( 
.A(n_14913),
.Y(n_15056)
);

AOI31xp33_ASAP7_75t_L g15057 ( 
.A1(n_14905),
.A2(n_2734),
.A3(n_2732),
.B(n_2733),
.Y(n_15057)
);

INVx1_ASAP7_75t_L g15058 ( 
.A(n_14910),
.Y(n_15058)
);

OAI32xp33_ASAP7_75t_L g15059 ( 
.A1(n_14926),
.A2(n_2735),
.A3(n_2732),
.B1(n_2734),
.B2(n_2736),
.Y(n_15059)
);

INVx2_ASAP7_75t_L g15060 ( 
.A(n_14911),
.Y(n_15060)
);

NAND3xp33_ASAP7_75t_SL g15061 ( 
.A(n_14973),
.B(n_2736),
.C(n_2737),
.Y(n_15061)
);

HB1xp67_ASAP7_75t_L g15062 ( 
.A(n_14986),
.Y(n_15062)
);

INVx1_ASAP7_75t_L g15063 ( 
.A(n_14946),
.Y(n_15063)
);

INVx1_ASAP7_75t_L g15064 ( 
.A(n_14949),
.Y(n_15064)
);

AO221x1_ASAP7_75t_L g15065 ( 
.A1(n_14937),
.A2(n_2739),
.B1(n_2737),
.B2(n_2738),
.C(n_2740),
.Y(n_15065)
);

AOI222xp33_ASAP7_75t_L g15066 ( 
.A1(n_14967),
.A2(n_2741),
.B1(n_2743),
.B2(n_2739),
.C1(n_2740),
.C2(n_2742),
.Y(n_15066)
);

AND2x2_ASAP7_75t_L g15067 ( 
.A(n_14904),
.B(n_2741),
.Y(n_15067)
);

INVx1_ASAP7_75t_L g15068 ( 
.A(n_14930),
.Y(n_15068)
);

OAI22xp5_ASAP7_75t_L g15069 ( 
.A1(n_14947),
.A2(n_2744),
.B1(n_2742),
.B2(n_2743),
.Y(n_15069)
);

NAND2xp5_ASAP7_75t_L g15070 ( 
.A(n_14924),
.B(n_2745),
.Y(n_15070)
);

AND2x4_ASAP7_75t_SL g15071 ( 
.A(n_14984),
.B(n_2745),
.Y(n_15071)
);

NAND2xp5_ASAP7_75t_L g15072 ( 
.A(n_14953),
.B(n_2746),
.Y(n_15072)
);

AND2x2_ASAP7_75t_L g15073 ( 
.A(n_14906),
.B(n_14907),
.Y(n_15073)
);

INVx1_ASAP7_75t_SL g15074 ( 
.A(n_15008),
.Y(n_15074)
);

INVx2_ASAP7_75t_L g15075 ( 
.A(n_14970),
.Y(n_15075)
);

INVx2_ASAP7_75t_L g15076 ( 
.A(n_14936),
.Y(n_15076)
);

AND2x2_ASAP7_75t_L g15077 ( 
.A(n_14917),
.B(n_2746),
.Y(n_15077)
);

INVx2_ASAP7_75t_L g15078 ( 
.A(n_14901),
.Y(n_15078)
);

NAND2xp5_ASAP7_75t_L g15079 ( 
.A(n_14919),
.B(n_2747),
.Y(n_15079)
);

OAI21xp33_ASAP7_75t_L g15080 ( 
.A1(n_14897),
.A2(n_14908),
.B(n_14942),
.Y(n_15080)
);

INVx1_ASAP7_75t_L g15081 ( 
.A(n_14960),
.Y(n_15081)
);

AND2x2_ASAP7_75t_L g15082 ( 
.A(n_14921),
.B(n_2747),
.Y(n_15082)
);

OAI22xp5_ASAP7_75t_L g15083 ( 
.A1(n_15003),
.A2(n_2752),
.B1(n_2749),
.B2(n_2750),
.Y(n_15083)
);

NAND2xp33_ASAP7_75t_SL g15084 ( 
.A(n_14916),
.B(n_2749),
.Y(n_15084)
);

AND2x2_ASAP7_75t_L g15085 ( 
.A(n_14922),
.B(n_2752),
.Y(n_15085)
);

INVx1_ASAP7_75t_L g15086 ( 
.A(n_14889),
.Y(n_15086)
);

INVx1_ASAP7_75t_L g15087 ( 
.A(n_14964),
.Y(n_15087)
);

INVx2_ASAP7_75t_L g15088 ( 
.A(n_14900),
.Y(n_15088)
);

INVx1_ASAP7_75t_L g15089 ( 
.A(n_14912),
.Y(n_15089)
);

INVx1_ASAP7_75t_L g15090 ( 
.A(n_14996),
.Y(n_15090)
);

INVx1_ASAP7_75t_L g15091 ( 
.A(n_14991),
.Y(n_15091)
);

INVx1_ASAP7_75t_L g15092 ( 
.A(n_15014),
.Y(n_15092)
);

OR2x2_ASAP7_75t_L g15093 ( 
.A(n_14891),
.B(n_2753),
.Y(n_15093)
);

INVx1_ASAP7_75t_L g15094 ( 
.A(n_14893),
.Y(n_15094)
);

OAI21xp33_ASAP7_75t_L g15095 ( 
.A1(n_15012),
.A2(n_2754),
.B(n_2755),
.Y(n_15095)
);

NOR2xp67_ASAP7_75t_SL g15096 ( 
.A(n_14888),
.B(n_2754),
.Y(n_15096)
);

INVx1_ASAP7_75t_SL g15097 ( 
.A(n_15004),
.Y(n_15097)
);

INVx1_ASAP7_75t_L g15098 ( 
.A(n_14896),
.Y(n_15098)
);

BUFx2_ASAP7_75t_L g15099 ( 
.A(n_14929),
.Y(n_15099)
);

NAND3xp33_ASAP7_75t_L g15100 ( 
.A(n_15015),
.B(n_15002),
.C(n_14977),
.Y(n_15100)
);

OR2x2_ASAP7_75t_L g15101 ( 
.A(n_14902),
.B(n_2755),
.Y(n_15101)
);

NAND2xp5_ASAP7_75t_L g15102 ( 
.A(n_14999),
.B(n_14962),
.Y(n_15102)
);

INVx3_ASAP7_75t_L g15103 ( 
.A(n_14938),
.Y(n_15103)
);

NAND2xp5_ASAP7_75t_L g15104 ( 
.A(n_14932),
.B(n_2756),
.Y(n_15104)
);

INVx1_ASAP7_75t_L g15105 ( 
.A(n_15017),
.Y(n_15105)
);

INVx2_ASAP7_75t_L g15106 ( 
.A(n_14948),
.Y(n_15106)
);

AOI32xp33_ASAP7_75t_L g15107 ( 
.A1(n_14934),
.A2(n_2758),
.A3(n_2756),
.B1(n_2757),
.B2(n_2759),
.Y(n_15107)
);

AND2x2_ASAP7_75t_L g15108 ( 
.A(n_14939),
.B(n_2757),
.Y(n_15108)
);

INVx1_ASAP7_75t_SL g15109 ( 
.A(n_14920),
.Y(n_15109)
);

INVx1_ASAP7_75t_L g15110 ( 
.A(n_14969),
.Y(n_15110)
);

AOI22xp5_ASAP7_75t_L g15111 ( 
.A1(n_14952),
.A2(n_2761),
.B1(n_2758),
.B2(n_2759),
.Y(n_15111)
);

OR2x2_ASAP7_75t_L g15112 ( 
.A(n_14951),
.B(n_2761),
.Y(n_15112)
);

NAND2xp5_ASAP7_75t_L g15113 ( 
.A(n_14971),
.B(n_2762),
.Y(n_15113)
);

OAI32xp33_ASAP7_75t_L g15114 ( 
.A1(n_14898),
.A2(n_2764),
.A3(n_2762),
.B1(n_2763),
.B2(n_2765),
.Y(n_15114)
);

INVxp67_ASAP7_75t_L g15115 ( 
.A(n_14899),
.Y(n_15115)
);

INVx1_ASAP7_75t_L g15116 ( 
.A(n_14965),
.Y(n_15116)
);

INVx1_ASAP7_75t_L g15117 ( 
.A(n_14955),
.Y(n_15117)
);

NAND2xp5_ASAP7_75t_L g15118 ( 
.A(n_14958),
.B(n_2764),
.Y(n_15118)
);

INVx1_ASAP7_75t_SL g15119 ( 
.A(n_14968),
.Y(n_15119)
);

INVx2_ASAP7_75t_SL g15120 ( 
.A(n_14928),
.Y(n_15120)
);

AOI22xp5_ASAP7_75t_L g15121 ( 
.A1(n_14954),
.A2(n_2767),
.B1(n_2765),
.B2(n_2766),
.Y(n_15121)
);

AOI22xp33_ASAP7_75t_L g15122 ( 
.A1(n_14931),
.A2(n_2768),
.B1(n_2766),
.B2(n_2767),
.Y(n_15122)
);

INVx2_ASAP7_75t_L g15123 ( 
.A(n_14975),
.Y(n_15123)
);

HB1xp67_ASAP7_75t_L g15124 ( 
.A(n_14927),
.Y(n_15124)
);

AND2x2_ASAP7_75t_L g15125 ( 
.A(n_14956),
.B(n_2768),
.Y(n_15125)
);

AOI22xp5_ASAP7_75t_L g15126 ( 
.A1(n_15001),
.A2(n_2771),
.B1(n_2769),
.B2(n_2770),
.Y(n_15126)
);

OR2x2_ASAP7_75t_L g15127 ( 
.A(n_14981),
.B(n_2769),
.Y(n_15127)
);

NOR2x1_ASAP7_75t_L g15128 ( 
.A(n_14959),
.B(n_2770),
.Y(n_15128)
);

INVx1_ASAP7_75t_L g15129 ( 
.A(n_14982),
.Y(n_15129)
);

NAND2xp5_ASAP7_75t_L g15130 ( 
.A(n_14892),
.B(n_2771),
.Y(n_15130)
);

INVx2_ASAP7_75t_L g15131 ( 
.A(n_14978),
.Y(n_15131)
);

NOR4xp25_ASAP7_75t_L g15132 ( 
.A(n_14997),
.B(n_2775),
.C(n_2772),
.D(n_2774),
.Y(n_15132)
);

A2O1A1Ixp33_ASAP7_75t_L g15133 ( 
.A1(n_14966),
.A2(n_2777),
.B(n_2772),
.C(n_2776),
.Y(n_15133)
);

INVxp67_ASAP7_75t_L g15134 ( 
.A(n_14983),
.Y(n_15134)
);

AND2x2_ASAP7_75t_L g15135 ( 
.A(n_14894),
.B(n_2776),
.Y(n_15135)
);

INVx1_ASAP7_75t_L g15136 ( 
.A(n_15006),
.Y(n_15136)
);

AOI33xp33_ASAP7_75t_L g15137 ( 
.A1(n_15019),
.A2(n_2779),
.A3(n_2781),
.B1(n_2777),
.B2(n_2778),
.B3(n_2780),
.Y(n_15137)
);

INVx2_ASAP7_75t_L g15138 ( 
.A(n_15011),
.Y(n_15138)
);

INVx1_ASAP7_75t_SL g15139 ( 
.A(n_14979),
.Y(n_15139)
);

NAND2x2_ASAP7_75t_L g15140 ( 
.A(n_15021),
.B(n_2778),
.Y(n_15140)
);

INVx1_ASAP7_75t_L g15141 ( 
.A(n_15018),
.Y(n_15141)
);

OAI31xp33_ASAP7_75t_L g15142 ( 
.A1(n_14940),
.A2(n_2781),
.A3(n_2779),
.B(n_2780),
.Y(n_15142)
);

AOI22xp33_ASAP7_75t_SL g15143 ( 
.A1(n_14944),
.A2(n_2784),
.B1(n_2782),
.B2(n_2783),
.Y(n_15143)
);

INVx1_ASAP7_75t_L g15144 ( 
.A(n_15000),
.Y(n_15144)
);

INVx2_ASAP7_75t_SL g15145 ( 
.A(n_14980),
.Y(n_15145)
);

OAI21xp5_ASAP7_75t_L g15146 ( 
.A1(n_14974),
.A2(n_2783),
.B(n_2785),
.Y(n_15146)
);

INVx2_ASAP7_75t_L g15147 ( 
.A(n_14994),
.Y(n_15147)
);

INVx2_ASAP7_75t_L g15148 ( 
.A(n_14976),
.Y(n_15148)
);

AOI21xp5_ASAP7_75t_L g15149 ( 
.A1(n_15020),
.A2(n_2787),
.B(n_2788),
.Y(n_15149)
);

INVxp67_ASAP7_75t_L g15150 ( 
.A(n_15022),
.Y(n_15150)
);

NAND2xp5_ASAP7_75t_L g15151 ( 
.A(n_14972),
.B(n_2787),
.Y(n_15151)
);

INVx2_ASAP7_75t_L g15152 ( 
.A(n_14985),
.Y(n_15152)
);

INVx1_ASAP7_75t_L g15153 ( 
.A(n_14989),
.Y(n_15153)
);

OAI22xp5_ASAP7_75t_L g15154 ( 
.A1(n_14993),
.A2(n_2790),
.B1(n_2788),
.B2(n_2789),
.Y(n_15154)
);

INVx1_ASAP7_75t_L g15155 ( 
.A(n_14995),
.Y(n_15155)
);

INVx1_ASAP7_75t_L g15156 ( 
.A(n_14998),
.Y(n_15156)
);

INVx1_ASAP7_75t_L g15157 ( 
.A(n_14992),
.Y(n_15157)
);

NAND2xp5_ASAP7_75t_SL g15158 ( 
.A(n_15005),
.B(n_2789),
.Y(n_15158)
);

OAI31xp33_ASAP7_75t_L g15159 ( 
.A1(n_15007),
.A2(n_2792),
.A3(n_2790),
.B(n_2791),
.Y(n_15159)
);

NAND2xp5_ASAP7_75t_L g15160 ( 
.A(n_15025),
.B(n_15013),
.Y(n_15160)
);

INVxp67_ASAP7_75t_L g15161 ( 
.A(n_15041),
.Y(n_15161)
);

AOI22xp33_ASAP7_75t_L g15162 ( 
.A1(n_15099),
.A2(n_15028),
.B1(n_15048),
.B2(n_15056),
.Y(n_15162)
);

INVx1_ASAP7_75t_L g15163 ( 
.A(n_15071),
.Y(n_15163)
);

OAI21xp33_ASAP7_75t_SL g15164 ( 
.A1(n_15097),
.A2(n_15010),
.B(n_2791),
.Y(n_15164)
);

NAND2xp5_ASAP7_75t_L g15165 ( 
.A(n_15065),
.B(n_2792),
.Y(n_15165)
);

AND2x2_ASAP7_75t_L g15166 ( 
.A(n_15073),
.B(n_2793),
.Y(n_15166)
);

OAI22xp5_ASAP7_75t_L g15167 ( 
.A1(n_15046),
.A2(n_2796),
.B1(n_2793),
.B2(n_2794),
.Y(n_15167)
);

INVx1_ASAP7_75t_L g15168 ( 
.A(n_15026),
.Y(n_15168)
);

AOI21xp5_ASAP7_75t_L g15169 ( 
.A1(n_15124),
.A2(n_2794),
.B(n_2796),
.Y(n_15169)
);

AND2x2_ASAP7_75t_L g15170 ( 
.A(n_15038),
.B(n_2797),
.Y(n_15170)
);

INVx1_ASAP7_75t_L g15171 ( 
.A(n_15067),
.Y(n_15171)
);

OR2x2_ASAP7_75t_L g15172 ( 
.A(n_15132),
.B(n_2798),
.Y(n_15172)
);

OR2x2_ASAP7_75t_L g15173 ( 
.A(n_15061),
.B(n_15103),
.Y(n_15173)
);

OAI21xp5_ASAP7_75t_L g15174 ( 
.A1(n_15100),
.A2(n_2798),
.B(n_2799),
.Y(n_15174)
);

AND2x2_ASAP7_75t_L g15175 ( 
.A(n_15036),
.B(n_2799),
.Y(n_15175)
);

AOI222xp33_ASAP7_75t_L g15176 ( 
.A1(n_15080),
.A2(n_2802),
.B1(n_2804),
.B2(n_2800),
.C1(n_2801),
.C2(n_2803),
.Y(n_15176)
);

OAI21xp5_ASAP7_75t_L g15177 ( 
.A1(n_15150),
.A2(n_2800),
.B(n_2801),
.Y(n_15177)
);

AND2x2_ASAP7_75t_L g15178 ( 
.A(n_15040),
.B(n_2802),
.Y(n_15178)
);

AOI32xp33_ASAP7_75t_L g15179 ( 
.A1(n_15103),
.A2(n_2807),
.A3(n_2805),
.B1(n_2806),
.B2(n_2808),
.Y(n_15179)
);

NAND2xp5_ASAP7_75t_L g15180 ( 
.A(n_15077),
.B(n_2805),
.Y(n_15180)
);

OR2x2_ASAP7_75t_L g15181 ( 
.A(n_15042),
.B(n_2806),
.Y(n_15181)
);

AOI22xp5_ASAP7_75t_L g15182 ( 
.A1(n_15120),
.A2(n_2810),
.B1(n_2808),
.B2(n_2809),
.Y(n_15182)
);

AND2x2_ASAP7_75t_L g15183 ( 
.A(n_15047),
.B(n_2809),
.Y(n_15183)
);

NAND3xp33_ASAP7_75t_SL g15184 ( 
.A(n_15037),
.B(n_2810),
.C(n_2811),
.Y(n_15184)
);

INVx2_ASAP7_75t_SL g15185 ( 
.A(n_15034),
.Y(n_15185)
);

OAI22xp5_ASAP7_75t_L g15186 ( 
.A1(n_15027),
.A2(n_2813),
.B1(n_2811),
.B2(n_2812),
.Y(n_15186)
);

INVx1_ASAP7_75t_L g15187 ( 
.A(n_15082),
.Y(n_15187)
);

OR2x2_ASAP7_75t_L g15188 ( 
.A(n_15070),
.B(n_2812),
.Y(n_15188)
);

NAND2xp5_ASAP7_75t_L g15189 ( 
.A(n_15085),
.B(n_2813),
.Y(n_15189)
);

INVx3_ASAP7_75t_L g15190 ( 
.A(n_15039),
.Y(n_15190)
);

NAND2xp5_ASAP7_75t_L g15191 ( 
.A(n_15096),
.B(n_15051),
.Y(n_15191)
);

OR2x2_ASAP7_75t_L g15192 ( 
.A(n_15043),
.B(n_2814),
.Y(n_15192)
);

INVx1_ASAP7_75t_L g15193 ( 
.A(n_15093),
.Y(n_15193)
);

AOI32xp33_ASAP7_75t_L g15194 ( 
.A1(n_15029),
.A2(n_2816),
.A3(n_2814),
.B1(n_2815),
.B2(n_2817),
.Y(n_15194)
);

NAND2x1p5_ASAP7_75t_L g15195 ( 
.A(n_15032),
.B(n_2815),
.Y(n_15195)
);

AOI32xp33_ASAP7_75t_L g15196 ( 
.A1(n_15084),
.A2(n_2819),
.A3(n_2816),
.B1(n_2818),
.B2(n_2821),
.Y(n_15196)
);

AOI21xp5_ASAP7_75t_L g15197 ( 
.A1(n_15102),
.A2(n_15158),
.B(n_15072),
.Y(n_15197)
);

NAND2xp5_ASAP7_75t_L g15198 ( 
.A(n_15108),
.B(n_15143),
.Y(n_15198)
);

OAI21xp33_ASAP7_75t_L g15199 ( 
.A1(n_15145),
.A2(n_2822),
.B(n_2823),
.Y(n_15199)
);

OAI22xp5_ASAP7_75t_L g15200 ( 
.A1(n_15140),
.A2(n_15045),
.B1(n_15035),
.B2(n_15074),
.Y(n_15200)
);

OAI22xp5_ASAP7_75t_L g15201 ( 
.A1(n_15147),
.A2(n_2825),
.B1(n_2823),
.B2(n_2824),
.Y(n_15201)
);

INVx2_ASAP7_75t_L g15202 ( 
.A(n_15101),
.Y(n_15202)
);

INVxp67_ASAP7_75t_L g15203 ( 
.A(n_15062),
.Y(n_15203)
);

INVx1_ASAP7_75t_L g15204 ( 
.A(n_15137),
.Y(n_15204)
);

AOI32xp33_ASAP7_75t_L g15205 ( 
.A1(n_15128),
.A2(n_2826),
.A3(n_2824),
.B1(n_2825),
.B2(n_2827),
.Y(n_15205)
);

NAND2xp5_ASAP7_75t_L g15206 ( 
.A(n_15135),
.B(n_2827),
.Y(n_15206)
);

AOI222xp33_ASAP7_75t_L g15207 ( 
.A1(n_15144),
.A2(n_2830),
.B1(n_2832),
.B2(n_2828),
.C1(n_2829),
.C2(n_2831),
.Y(n_15207)
);

INVx2_ASAP7_75t_L g15208 ( 
.A(n_15050),
.Y(n_15208)
);

NAND4xp25_ASAP7_75t_L g15209 ( 
.A(n_15139),
.B(n_2830),
.C(n_2828),
.D(n_2829),
.Y(n_15209)
);

AOI221xp5_ASAP7_75t_L g15210 ( 
.A1(n_15092),
.A2(n_2834),
.B1(n_2831),
.B2(n_2833),
.C(n_2836),
.Y(n_15210)
);

NAND2xp5_ASAP7_75t_SL g15211 ( 
.A(n_15066),
.B(n_2833),
.Y(n_15211)
);

AOI32xp33_ASAP7_75t_L g15212 ( 
.A1(n_15148),
.A2(n_2837),
.A3(n_2834),
.B1(n_2836),
.B2(n_2838),
.Y(n_15212)
);

OAI22xp5_ASAP7_75t_L g15213 ( 
.A1(n_15058),
.A2(n_2839),
.B1(n_2837),
.B2(n_2838),
.Y(n_15213)
);

NAND2xp5_ASAP7_75t_L g15214 ( 
.A(n_15125),
.B(n_2839),
.Y(n_15214)
);

AOI22xp5_ASAP7_75t_L g15215 ( 
.A1(n_15068),
.A2(n_2842),
.B1(n_2840),
.B2(n_2841),
.Y(n_15215)
);

OR2x2_ASAP7_75t_L g15216 ( 
.A(n_15079),
.B(n_2840),
.Y(n_15216)
);

AOI32xp33_ASAP7_75t_L g15217 ( 
.A1(n_15054),
.A2(n_2843),
.A3(n_2841),
.B1(n_2842),
.B2(n_2844),
.Y(n_15217)
);

NAND3xp33_ASAP7_75t_L g15218 ( 
.A(n_15142),
.B(n_2843),
.C(n_2844),
.Y(n_15218)
);

NOR2xp33_ASAP7_75t_SL g15219 ( 
.A(n_15159),
.B(n_2845),
.Y(n_15219)
);

INVx1_ASAP7_75t_L g15220 ( 
.A(n_15057),
.Y(n_15220)
);

INVxp67_ASAP7_75t_L g15221 ( 
.A(n_15044),
.Y(n_15221)
);

AND2x2_ASAP7_75t_L g15222 ( 
.A(n_15055),
.B(n_2845),
.Y(n_15222)
);

OAI22xp5_ASAP7_75t_L g15223 ( 
.A1(n_15053),
.A2(n_2848),
.B1(n_2846),
.B2(n_2847),
.Y(n_15223)
);

INVx1_ASAP7_75t_L g15224 ( 
.A(n_15033),
.Y(n_15224)
);

OAI32xp33_ASAP7_75t_L g15225 ( 
.A1(n_15104),
.A2(n_2849),
.A3(n_2846),
.B1(n_2848),
.B2(n_2850),
.Y(n_15225)
);

OAI21xp5_ASAP7_75t_L g15226 ( 
.A1(n_15133),
.A2(n_2849),
.B(n_2850),
.Y(n_15226)
);

NOR2xp67_ASAP7_75t_L g15227 ( 
.A(n_15149),
.B(n_2851),
.Y(n_15227)
);

INVx2_ASAP7_75t_L g15228 ( 
.A(n_15112),
.Y(n_15228)
);

INVx1_ASAP7_75t_L g15229 ( 
.A(n_15031),
.Y(n_15229)
);

AND2x2_ASAP7_75t_L g15230 ( 
.A(n_15063),
.B(n_2851),
.Y(n_15230)
);

AOI21xp33_ASAP7_75t_L g15231 ( 
.A1(n_15064),
.A2(n_2852),
.B(n_2853),
.Y(n_15231)
);

INVx1_ASAP7_75t_L g15232 ( 
.A(n_15113),
.Y(n_15232)
);

INVx2_ASAP7_75t_L g15233 ( 
.A(n_15127),
.Y(n_15233)
);

INVx2_ASAP7_75t_L g15234 ( 
.A(n_15049),
.Y(n_15234)
);

INVxp33_ASAP7_75t_L g15235 ( 
.A(n_15118),
.Y(n_15235)
);

INVx1_ASAP7_75t_L g15236 ( 
.A(n_15130),
.Y(n_15236)
);

NAND4xp25_ASAP7_75t_L g15237 ( 
.A(n_15089),
.B(n_2854),
.C(n_2852),
.D(n_2853),
.Y(n_15237)
);

AND2x2_ASAP7_75t_L g15238 ( 
.A(n_15075),
.B(n_15081),
.Y(n_15238)
);

OAI21xp33_ASAP7_75t_L g15239 ( 
.A1(n_15087),
.A2(n_2854),
.B(n_2855),
.Y(n_15239)
);

INVx2_ASAP7_75t_L g15240 ( 
.A(n_15060),
.Y(n_15240)
);

AO22x1_ASAP7_75t_L g15241 ( 
.A1(n_15146),
.A2(n_2858),
.B1(n_2856),
.B2(n_2857),
.Y(n_15241)
);

OAI22xp5_ASAP7_75t_L g15242 ( 
.A1(n_15090),
.A2(n_2860),
.B1(n_2856),
.B2(n_2859),
.Y(n_15242)
);

INVx2_ASAP7_75t_L g15243 ( 
.A(n_15078),
.Y(n_15243)
);

OR2x2_ASAP7_75t_L g15244 ( 
.A(n_15076),
.B(n_15091),
.Y(n_15244)
);

INVx1_ASAP7_75t_L g15245 ( 
.A(n_15151),
.Y(n_15245)
);

NAND2xp5_ASAP7_75t_L g15246 ( 
.A(n_15052),
.B(n_2859),
.Y(n_15246)
);

OAI31xp33_ASAP7_75t_L g15247 ( 
.A1(n_15109),
.A2(n_2862),
.A3(n_2860),
.B(n_2861),
.Y(n_15247)
);

INVx1_ASAP7_75t_L g15248 ( 
.A(n_15030),
.Y(n_15248)
);

AOI22xp33_ASAP7_75t_L g15249 ( 
.A1(n_15086),
.A2(n_2863),
.B1(n_2861),
.B2(n_2862),
.Y(n_15249)
);

INVx1_ASAP7_75t_L g15250 ( 
.A(n_15095),
.Y(n_15250)
);

INVx1_ASAP7_75t_L g15251 ( 
.A(n_15105),
.Y(n_15251)
);

NAND2xp5_ASAP7_75t_L g15252 ( 
.A(n_15107),
.B(n_2863),
.Y(n_15252)
);

INVx1_ASAP7_75t_L g15253 ( 
.A(n_15088),
.Y(n_15253)
);

AOI32xp33_ASAP7_75t_L g15254 ( 
.A1(n_15119),
.A2(n_2866),
.A3(n_2864),
.B1(n_2865),
.B2(n_2867),
.Y(n_15254)
);

AOI211xp5_ASAP7_75t_L g15255 ( 
.A1(n_15155),
.A2(n_2866),
.B(n_2864),
.C(n_2865),
.Y(n_15255)
);

HB1xp67_ASAP7_75t_L g15256 ( 
.A(n_15083),
.Y(n_15256)
);

OAI21xp5_ASAP7_75t_L g15257 ( 
.A1(n_15134),
.A2(n_2867),
.B(n_2869),
.Y(n_15257)
);

INVx2_ASAP7_75t_L g15258 ( 
.A(n_15106),
.Y(n_15258)
);

NAND2xp5_ASAP7_75t_L g15259 ( 
.A(n_15122),
.B(n_2869),
.Y(n_15259)
);

NAND2xp5_ASAP7_75t_L g15260 ( 
.A(n_15126),
.B(n_2871),
.Y(n_15260)
);

INVx1_ASAP7_75t_SL g15261 ( 
.A(n_15138),
.Y(n_15261)
);

O2A1O1Ixp33_ASAP7_75t_L g15262 ( 
.A1(n_15059),
.A2(n_2874),
.B(n_2871),
.C(n_2872),
.Y(n_15262)
);

NAND2xp5_ASAP7_75t_L g15263 ( 
.A(n_15111),
.B(n_2872),
.Y(n_15263)
);

INVx2_ASAP7_75t_SL g15264 ( 
.A(n_15123),
.Y(n_15264)
);

INVx1_ASAP7_75t_L g15265 ( 
.A(n_15114),
.Y(n_15265)
);

AOI22xp33_ASAP7_75t_L g15266 ( 
.A1(n_15152),
.A2(n_2877),
.B1(n_2875),
.B2(n_2876),
.Y(n_15266)
);

AND2x2_ASAP7_75t_L g15267 ( 
.A(n_15131),
.B(n_15116),
.Y(n_15267)
);

O2A1O1Ixp33_ASAP7_75t_L g15268 ( 
.A1(n_15156),
.A2(n_2878),
.B(n_2875),
.C(n_2876),
.Y(n_15268)
);

OAI21xp33_ASAP7_75t_L g15269 ( 
.A1(n_15110),
.A2(n_2878),
.B(n_2879),
.Y(n_15269)
);

OR2x2_ASAP7_75t_L g15270 ( 
.A(n_15153),
.B(n_2879),
.Y(n_15270)
);

AOI22xp5_ASAP7_75t_L g15271 ( 
.A1(n_15157),
.A2(n_2882),
.B1(n_2880),
.B2(n_2881),
.Y(n_15271)
);

OA222x2_ASAP7_75t_L g15272 ( 
.A1(n_15115),
.A2(n_2882),
.B1(n_2884),
.B2(n_2880),
.C1(n_2881),
.C2(n_2883),
.Y(n_15272)
);

AND2x2_ASAP7_75t_L g15273 ( 
.A(n_15094),
.B(n_2883),
.Y(n_15273)
);

OR2x2_ASAP7_75t_L g15274 ( 
.A(n_15098),
.B(n_2885),
.Y(n_15274)
);

AND2x2_ASAP7_75t_L g15275 ( 
.A(n_15117),
.B(n_2886),
.Y(n_15275)
);

INVx2_ASAP7_75t_L g15276 ( 
.A(n_15129),
.Y(n_15276)
);

INVx1_ASAP7_75t_L g15277 ( 
.A(n_15121),
.Y(n_15277)
);

INVx2_ASAP7_75t_L g15278 ( 
.A(n_15136),
.Y(n_15278)
);

AOI211x1_ASAP7_75t_SL g15279 ( 
.A1(n_15069),
.A2(n_2888),
.B(n_2886),
.C(n_2887),
.Y(n_15279)
);

NAND2xp5_ASAP7_75t_L g15280 ( 
.A(n_15141),
.B(n_2888),
.Y(n_15280)
);

INVx1_ASAP7_75t_SL g15281 ( 
.A(n_15154),
.Y(n_15281)
);

NOR2xp33_ASAP7_75t_SL g15282 ( 
.A(n_15025),
.B(n_2889),
.Y(n_15282)
);

OR2x2_ASAP7_75t_L g15283 ( 
.A(n_15025),
.B(n_2889),
.Y(n_15283)
);

OAI211xp5_ASAP7_75t_L g15284 ( 
.A1(n_15080),
.A2(n_2892),
.B(n_2890),
.C(n_2891),
.Y(n_15284)
);

OAI31xp33_ASAP7_75t_L g15285 ( 
.A1(n_15025),
.A2(n_2892),
.A3(n_2890),
.B(n_2891),
.Y(n_15285)
);

NOR3xp33_ASAP7_75t_L g15286 ( 
.A(n_15190),
.B(n_2893),
.C(n_2894),
.Y(n_15286)
);

INVx1_ASAP7_75t_L g15287 ( 
.A(n_15283),
.Y(n_15287)
);

OAI22xp5_ASAP7_75t_L g15288 ( 
.A1(n_15162),
.A2(n_15161),
.B1(n_15203),
.B2(n_15173),
.Y(n_15288)
);

OAI221xp5_ASAP7_75t_L g15289 ( 
.A1(n_15247),
.A2(n_2895),
.B1(n_2893),
.B2(n_2894),
.C(n_2896),
.Y(n_15289)
);

NAND2xp5_ASAP7_75t_L g15290 ( 
.A(n_15166),
.B(n_2895),
.Y(n_15290)
);

AOI211xp5_ASAP7_75t_L g15291 ( 
.A1(n_15200),
.A2(n_2898),
.B(n_2896),
.C(n_2897),
.Y(n_15291)
);

INVxp67_ASAP7_75t_L g15292 ( 
.A(n_15282),
.Y(n_15292)
);

AOI322xp5_ASAP7_75t_L g15293 ( 
.A1(n_15261),
.A2(n_15185),
.A3(n_15281),
.B1(n_15265),
.B2(n_15220),
.C1(n_15264),
.C2(n_15253),
.Y(n_15293)
);

INVx2_ASAP7_75t_L g15294 ( 
.A(n_15195),
.Y(n_15294)
);

AOI21xp33_ASAP7_75t_SL g15295 ( 
.A1(n_15172),
.A2(n_2898),
.B(n_2899),
.Y(n_15295)
);

INVx1_ASAP7_75t_L g15296 ( 
.A(n_15178),
.Y(n_15296)
);

AOI221xp5_ASAP7_75t_L g15297 ( 
.A1(n_15262),
.A2(n_2901),
.B1(n_2899),
.B2(n_2900),
.C(n_2902),
.Y(n_15297)
);

O2A1O1Ixp33_ASAP7_75t_L g15298 ( 
.A1(n_15164),
.A2(n_2903),
.B(n_2901),
.C(n_2902),
.Y(n_15298)
);

OAI22xp5_ASAP7_75t_L g15299 ( 
.A1(n_15218),
.A2(n_2905),
.B1(n_2903),
.B2(n_2904),
.Y(n_15299)
);

INVxp67_ASAP7_75t_L g15300 ( 
.A(n_15170),
.Y(n_15300)
);

AOI321xp33_ASAP7_75t_L g15301 ( 
.A1(n_15211),
.A2(n_2907),
.A3(n_2909),
.B1(n_2905),
.B2(n_2906),
.C(n_2908),
.Y(n_15301)
);

INVx2_ASAP7_75t_L g15302 ( 
.A(n_15270),
.Y(n_15302)
);

AND2x2_ASAP7_75t_L g15303 ( 
.A(n_15238),
.B(n_15190),
.Y(n_15303)
);

AOI21xp5_ASAP7_75t_SL g15304 ( 
.A1(n_15268),
.A2(n_2906),
.B(n_2908),
.Y(n_15304)
);

INVx3_ASAP7_75t_L g15305 ( 
.A(n_15234),
.Y(n_15305)
);

OAI321xp33_ASAP7_75t_L g15306 ( 
.A1(n_15191),
.A2(n_2911),
.A3(n_2913),
.B1(n_2909),
.B2(n_2910),
.C(n_2912),
.Y(n_15306)
);

INVx1_ASAP7_75t_L g15307 ( 
.A(n_15183),
.Y(n_15307)
);

OR2x2_ASAP7_75t_L g15308 ( 
.A(n_15165),
.B(n_2910),
.Y(n_15308)
);

NAND2xp5_ASAP7_75t_L g15309 ( 
.A(n_15222),
.B(n_2911),
.Y(n_15309)
);

OAI22xp33_ASAP7_75t_L g15310 ( 
.A1(n_15219),
.A2(n_15192),
.B1(n_15240),
.B2(n_15259),
.Y(n_15310)
);

INVx1_ASAP7_75t_L g15311 ( 
.A(n_15230),
.Y(n_15311)
);

AOI221xp5_ASAP7_75t_L g15312 ( 
.A1(n_15174),
.A2(n_2916),
.B1(n_2914),
.B2(n_2915),
.C(n_2917),
.Y(n_15312)
);

OAI21xp5_ASAP7_75t_L g15313 ( 
.A1(n_15197),
.A2(n_2915),
.B(n_2918),
.Y(n_15313)
);

AOI21xp5_ASAP7_75t_L g15314 ( 
.A1(n_15160),
.A2(n_15214),
.B(n_15206),
.Y(n_15314)
);

NOR2xp33_ASAP7_75t_L g15315 ( 
.A(n_15237),
.B(n_2919),
.Y(n_15315)
);

OA22x2_ASAP7_75t_L g15316 ( 
.A1(n_15226),
.A2(n_2922),
.B1(n_2920),
.B2(n_2921),
.Y(n_15316)
);

NOR2xp33_ASAP7_75t_L g15317 ( 
.A(n_15199),
.B(n_2920),
.Y(n_15317)
);

AOI31xp33_ASAP7_75t_L g15318 ( 
.A1(n_15163),
.A2(n_2923),
.A3(n_2921),
.B(n_2922),
.Y(n_15318)
);

INVx1_ASAP7_75t_L g15319 ( 
.A(n_15175),
.Y(n_15319)
);

AND2x2_ASAP7_75t_L g15320 ( 
.A(n_15243),
.B(n_2924),
.Y(n_15320)
);

AOI22xp5_ASAP7_75t_L g15321 ( 
.A1(n_15258),
.A2(n_2926),
.B1(n_2924),
.B2(n_2925),
.Y(n_15321)
);

AOI22xp5_ASAP7_75t_L g15322 ( 
.A1(n_15251),
.A2(n_15204),
.B1(n_15248),
.B2(n_15267),
.Y(n_15322)
);

INVx1_ASAP7_75t_L g15323 ( 
.A(n_15274),
.Y(n_15323)
);

AOI22xp5_ASAP7_75t_L g15324 ( 
.A1(n_15250),
.A2(n_2927),
.B1(n_2925),
.B2(n_2926),
.Y(n_15324)
);

OAI211xp5_ASAP7_75t_SL g15325 ( 
.A1(n_15221),
.A2(n_2930),
.B(n_2928),
.C(n_2929),
.Y(n_15325)
);

INVx1_ASAP7_75t_L g15326 ( 
.A(n_15273),
.Y(n_15326)
);

AOI22xp33_ASAP7_75t_SL g15327 ( 
.A1(n_15256),
.A2(n_2932),
.B1(n_2930),
.B2(n_2931),
.Y(n_15327)
);

OAI22xp5_ASAP7_75t_L g15328 ( 
.A1(n_15244),
.A2(n_2935),
.B1(n_2933),
.B2(n_2934),
.Y(n_15328)
);

OAI22x1_ASAP7_75t_L g15329 ( 
.A1(n_15202),
.A2(n_2935),
.B1(n_2933),
.B2(n_2934),
.Y(n_15329)
);

O2A1O1Ixp33_ASAP7_75t_L g15330 ( 
.A1(n_15246),
.A2(n_2938),
.B(n_2936),
.C(n_2937),
.Y(n_15330)
);

INVx1_ASAP7_75t_L g15331 ( 
.A(n_15275),
.Y(n_15331)
);

INVx1_ASAP7_75t_SL g15332 ( 
.A(n_15181),
.Y(n_15332)
);

OR2x2_ASAP7_75t_L g15333 ( 
.A(n_15180),
.B(n_2936),
.Y(n_15333)
);

NOR2xp33_ASAP7_75t_L g15334 ( 
.A(n_15209),
.B(n_2938),
.Y(n_15334)
);

OAI21xp5_ASAP7_75t_L g15335 ( 
.A1(n_15227),
.A2(n_2939),
.B(n_2940),
.Y(n_15335)
);

OAI21xp5_ASAP7_75t_SL g15336 ( 
.A1(n_15279),
.A2(n_2939),
.B(n_2940),
.Y(n_15336)
);

OAI21xp5_ASAP7_75t_L g15337 ( 
.A1(n_15252),
.A2(n_2941),
.B(n_2942),
.Y(n_15337)
);

XOR2x2_ASAP7_75t_L g15338 ( 
.A(n_15184),
.B(n_2941),
.Y(n_15338)
);

AND2x2_ASAP7_75t_L g15339 ( 
.A(n_15171),
.B(n_2942),
.Y(n_15339)
);

AOI22xp33_ASAP7_75t_L g15340 ( 
.A1(n_15208),
.A2(n_2945),
.B1(n_2943),
.B2(n_2944),
.Y(n_15340)
);

AOI21xp33_ASAP7_75t_L g15341 ( 
.A1(n_15235),
.A2(n_2943),
.B(n_2945),
.Y(n_15341)
);

AOI22xp5_ASAP7_75t_L g15342 ( 
.A1(n_15187),
.A2(n_2948),
.B1(n_2946),
.B2(n_2947),
.Y(n_15342)
);

AOI21xp5_ASAP7_75t_L g15343 ( 
.A1(n_15198),
.A2(n_2948),
.B(n_2949),
.Y(n_15343)
);

AOI211xp5_ASAP7_75t_L g15344 ( 
.A1(n_15241),
.A2(n_2951),
.B(n_2949),
.C(n_2950),
.Y(n_15344)
);

INVx2_ASAP7_75t_L g15345 ( 
.A(n_15188),
.Y(n_15345)
);

OAI221xp5_ASAP7_75t_L g15346 ( 
.A1(n_15205),
.A2(n_2953),
.B1(n_2950),
.B2(n_2952),
.C(n_2954),
.Y(n_15346)
);

OAI221xp5_ASAP7_75t_L g15347 ( 
.A1(n_15285),
.A2(n_2955),
.B1(n_2953),
.B2(n_2954),
.C(n_2956),
.Y(n_15347)
);

AOI22xp5_ASAP7_75t_L g15348 ( 
.A1(n_15277),
.A2(n_2957),
.B1(n_2955),
.B2(n_2956),
.Y(n_15348)
);

INVx2_ASAP7_75t_L g15349 ( 
.A(n_15216),
.Y(n_15349)
);

INVx2_ASAP7_75t_L g15350 ( 
.A(n_15193),
.Y(n_15350)
);

INVx2_ASAP7_75t_L g15351 ( 
.A(n_15189),
.Y(n_15351)
);

XOR2x2_ASAP7_75t_L g15352 ( 
.A(n_15255),
.B(n_2957),
.Y(n_15352)
);

O2A1O1Ixp33_ASAP7_75t_SL g15353 ( 
.A1(n_15284),
.A2(n_2960),
.B(n_2958),
.C(n_2959),
.Y(n_15353)
);

INVxp67_ASAP7_75t_L g15354 ( 
.A(n_15207),
.Y(n_15354)
);

INVx1_ASAP7_75t_L g15355 ( 
.A(n_15263),
.Y(n_15355)
);

OAI221xp5_ASAP7_75t_L g15356 ( 
.A1(n_15196),
.A2(n_2962),
.B1(n_2958),
.B2(n_2961),
.C(n_2963),
.Y(n_15356)
);

OAI21xp5_ASAP7_75t_L g15357 ( 
.A1(n_15280),
.A2(n_2961),
.B(n_2962),
.Y(n_15357)
);

OAI22xp5_ASAP7_75t_L g15358 ( 
.A1(n_15168),
.A2(n_2965),
.B1(n_2963),
.B2(n_2964),
.Y(n_15358)
);

INVx1_ASAP7_75t_L g15359 ( 
.A(n_15260),
.Y(n_15359)
);

NAND3xp33_ASAP7_75t_L g15360 ( 
.A(n_15176),
.B(n_2964),
.C(n_2965),
.Y(n_15360)
);

INVx1_ASAP7_75t_L g15361 ( 
.A(n_15239),
.Y(n_15361)
);

AOI222xp33_ASAP7_75t_L g15362 ( 
.A1(n_15229),
.A2(n_2969),
.B1(n_2971),
.B2(n_2966),
.C1(n_2968),
.C2(n_2970),
.Y(n_15362)
);

INVx1_ASAP7_75t_L g15363 ( 
.A(n_15269),
.Y(n_15363)
);

AOI21xp33_ASAP7_75t_SL g15364 ( 
.A1(n_15186),
.A2(n_2968),
.B(n_2969),
.Y(n_15364)
);

OAI22x1_ASAP7_75t_L g15365 ( 
.A1(n_15182),
.A2(n_2972),
.B1(n_2970),
.B2(n_2971),
.Y(n_15365)
);

AOI222xp33_ASAP7_75t_L g15366 ( 
.A1(n_15276),
.A2(n_2974),
.B1(n_2977),
.B2(n_2972),
.C1(n_2973),
.C2(n_2976),
.Y(n_15366)
);

AOI322xp5_ASAP7_75t_L g15367 ( 
.A1(n_15278),
.A2(n_2980),
.A3(n_2979),
.B1(n_2976),
.B2(n_2973),
.C1(n_2974),
.C2(n_2978),
.Y(n_15367)
);

AOI211xp5_ASAP7_75t_L g15368 ( 
.A1(n_15223),
.A2(n_2980),
.B(n_2978),
.C(n_2979),
.Y(n_15368)
);

AOI22xp5_ASAP7_75t_L g15369 ( 
.A1(n_15224),
.A2(n_2983),
.B1(n_2981),
.B2(n_2982),
.Y(n_15369)
);

INVx1_ASAP7_75t_L g15370 ( 
.A(n_15177),
.Y(n_15370)
);

OA21x2_ASAP7_75t_L g15371 ( 
.A1(n_15232),
.A2(n_2981),
.B(n_2982),
.Y(n_15371)
);

INVx1_ASAP7_75t_L g15372 ( 
.A(n_15257),
.Y(n_15372)
);

OR2x2_ASAP7_75t_L g15373 ( 
.A(n_15228),
.B(n_2985),
.Y(n_15373)
);

NOR3xp33_ASAP7_75t_L g15374 ( 
.A(n_15236),
.B(n_2985),
.C(n_2986),
.Y(n_15374)
);

AOI221xp5_ASAP7_75t_L g15375 ( 
.A1(n_15245),
.A2(n_2988),
.B1(n_2986),
.B2(n_2987),
.C(n_2989),
.Y(n_15375)
);

AOI21xp33_ASAP7_75t_SL g15376 ( 
.A1(n_15254),
.A2(n_2987),
.B(n_2988),
.Y(n_15376)
);

O2A1O1Ixp5_ASAP7_75t_L g15377 ( 
.A1(n_15233),
.A2(n_2992),
.B(n_2990),
.C(n_2991),
.Y(n_15377)
);

NAND3xp33_ASAP7_75t_L g15378 ( 
.A(n_15169),
.B(n_2990),
.C(n_2991),
.Y(n_15378)
);

AOI22xp5_ASAP7_75t_L g15379 ( 
.A1(n_15210),
.A2(n_2994),
.B1(n_2992),
.B2(n_2993),
.Y(n_15379)
);

AOI22xp5_ASAP7_75t_L g15380 ( 
.A1(n_15167),
.A2(n_2995),
.B1(n_2993),
.B2(n_2994),
.Y(n_15380)
);

A2O1A1Ixp33_ASAP7_75t_L g15381 ( 
.A1(n_15212),
.A2(n_15179),
.B(n_15194),
.C(n_15217),
.Y(n_15381)
);

OAI21xp33_ASAP7_75t_L g15382 ( 
.A1(n_15266),
.A2(n_2996),
.B(n_2997),
.Y(n_15382)
);

OAI22xp5_ASAP7_75t_L g15383 ( 
.A1(n_15249),
.A2(n_2999),
.B1(n_2996),
.B2(n_2998),
.Y(n_15383)
);

OAI31xp33_ASAP7_75t_L g15384 ( 
.A1(n_15231),
.A2(n_3000),
.A3(n_2998),
.B(n_2999),
.Y(n_15384)
);

INVx2_ASAP7_75t_SL g15385 ( 
.A(n_15201),
.Y(n_15385)
);

OAI32xp33_ASAP7_75t_L g15386 ( 
.A1(n_15213),
.A2(n_3003),
.A3(n_3001),
.B1(n_3002),
.B2(n_3004),
.Y(n_15386)
);

AOI221xp5_ASAP7_75t_L g15387 ( 
.A1(n_15225),
.A2(n_3003),
.B1(n_3001),
.B2(n_3002),
.C(n_3006),
.Y(n_15387)
);

OAI211xp5_ASAP7_75t_SL g15388 ( 
.A1(n_15215),
.A2(n_15271),
.B(n_15242),
.C(n_15272),
.Y(n_15388)
);

INVx2_ASAP7_75t_L g15389 ( 
.A(n_15283),
.Y(n_15389)
);

INVxp33_ASAP7_75t_L g15390 ( 
.A(n_15170),
.Y(n_15390)
);

INVx1_ASAP7_75t_SL g15391 ( 
.A(n_15173),
.Y(n_15391)
);

INVx1_ASAP7_75t_L g15392 ( 
.A(n_15283),
.Y(n_15392)
);

AOI21xp33_ASAP7_75t_L g15393 ( 
.A1(n_15173),
.A2(n_3006),
.B(n_3007),
.Y(n_15393)
);

INVx1_ASAP7_75t_SL g15394 ( 
.A(n_15173),
.Y(n_15394)
);

NAND3xp33_ASAP7_75t_L g15395 ( 
.A(n_15162),
.B(n_3007),
.C(n_3008),
.Y(n_15395)
);

NAND2xp5_ASAP7_75t_L g15396 ( 
.A(n_15166),
.B(n_3008),
.Y(n_15396)
);

INVx1_ASAP7_75t_L g15397 ( 
.A(n_15283),
.Y(n_15397)
);

OAI21xp5_ASAP7_75t_L g15398 ( 
.A1(n_15161),
.A2(n_3009),
.B(n_3010),
.Y(n_15398)
);

OAI22xp5_ASAP7_75t_L g15399 ( 
.A1(n_15162),
.A2(n_3012),
.B1(n_3010),
.B2(n_3011),
.Y(n_15399)
);

OA33x2_ASAP7_75t_L g15400 ( 
.A1(n_15191),
.A2(n_3013),
.A3(n_3015),
.B1(n_3011),
.B2(n_3012),
.B3(n_3014),
.Y(n_15400)
);

AOI31xp33_ASAP7_75t_L g15401 ( 
.A1(n_15172),
.A2(n_3015),
.A3(n_3013),
.B(n_3014),
.Y(n_15401)
);

AOI22xp5_ASAP7_75t_L g15402 ( 
.A1(n_15185),
.A2(n_3018),
.B1(n_3016),
.B2(n_3017),
.Y(n_15402)
);

INVx1_ASAP7_75t_L g15403 ( 
.A(n_15283),
.Y(n_15403)
);

INVx1_ASAP7_75t_L g15404 ( 
.A(n_15283),
.Y(n_15404)
);

NAND2xp33_ASAP7_75t_L g15405 ( 
.A(n_15254),
.B(n_3016),
.Y(n_15405)
);

INVxp33_ASAP7_75t_L g15406 ( 
.A(n_15170),
.Y(n_15406)
);

AOI221xp5_ASAP7_75t_L g15407 ( 
.A1(n_15200),
.A2(n_3020),
.B1(n_3017),
.B2(n_3019),
.C(n_3021),
.Y(n_15407)
);

OR2x2_ASAP7_75t_L g15408 ( 
.A(n_15172),
.B(n_3019),
.Y(n_15408)
);

AOI22xp5_ASAP7_75t_L g15409 ( 
.A1(n_15185),
.A2(n_3022),
.B1(n_3020),
.B2(n_3021),
.Y(n_15409)
);

AOI21xp5_ASAP7_75t_L g15410 ( 
.A1(n_15191),
.A2(n_3023),
.B(n_3024),
.Y(n_15410)
);

INVx1_ASAP7_75t_L g15411 ( 
.A(n_15283),
.Y(n_15411)
);

INVx1_ASAP7_75t_L g15412 ( 
.A(n_15283),
.Y(n_15412)
);

AOI221xp5_ASAP7_75t_L g15413 ( 
.A1(n_15200),
.A2(n_3026),
.B1(n_3024),
.B2(n_3025),
.C(n_3027),
.Y(n_15413)
);

OAI332xp33_ASAP7_75t_L g15414 ( 
.A1(n_15261),
.A2(n_3030),
.A3(n_3029),
.B1(n_3027),
.B2(n_3031),
.B3(n_3025),
.C1(n_3026),
.C2(n_3028),
.Y(n_15414)
);

AOI22xp5_ASAP7_75t_L g15415 ( 
.A1(n_15185),
.A2(n_3030),
.B1(n_3028),
.B2(n_3029),
.Y(n_15415)
);

AOI22xp5_ASAP7_75t_L g15416 ( 
.A1(n_15185),
.A2(n_3033),
.B1(n_3031),
.B2(n_3032),
.Y(n_15416)
);

INVx3_ASAP7_75t_L g15417 ( 
.A(n_15305),
.Y(n_15417)
);

INVx1_ASAP7_75t_L g15418 ( 
.A(n_15303),
.Y(n_15418)
);

NAND2xp5_ASAP7_75t_L g15419 ( 
.A(n_15339),
.B(n_3033),
.Y(n_15419)
);

AND2x4_ASAP7_75t_L g15420 ( 
.A(n_15294),
.B(n_3034),
.Y(n_15420)
);

AND2x2_ASAP7_75t_L g15421 ( 
.A(n_15319),
.B(n_3034),
.Y(n_15421)
);

NOR2xp33_ASAP7_75t_L g15422 ( 
.A(n_15390),
.B(n_3035),
.Y(n_15422)
);

OR2x2_ASAP7_75t_L g15423 ( 
.A(n_15408),
.B(n_15290),
.Y(n_15423)
);

INVx1_ASAP7_75t_L g15424 ( 
.A(n_15320),
.Y(n_15424)
);

INVx2_ASAP7_75t_L g15425 ( 
.A(n_15371),
.Y(n_15425)
);

INVx1_ASAP7_75t_SL g15426 ( 
.A(n_15371),
.Y(n_15426)
);

NOR2xp33_ASAP7_75t_L g15427 ( 
.A(n_15406),
.B(n_15401),
.Y(n_15427)
);

OAI22xp5_ASAP7_75t_SL g15428 ( 
.A1(n_15327),
.A2(n_3038),
.B1(n_3036),
.B2(n_3037),
.Y(n_15428)
);

OAI21xp33_ASAP7_75t_SL g15429 ( 
.A1(n_15293),
.A2(n_3036),
.B(n_3037),
.Y(n_15429)
);

NAND2xp5_ASAP7_75t_L g15430 ( 
.A(n_15318),
.B(n_3038),
.Y(n_15430)
);

AO22x1_ASAP7_75t_L g15431 ( 
.A1(n_15335),
.A2(n_3041),
.B1(n_3039),
.B2(n_3040),
.Y(n_15431)
);

OAI32xp33_ASAP7_75t_L g15432 ( 
.A1(n_15391),
.A2(n_3043),
.A3(n_3041),
.B1(n_3042),
.B2(n_3044),
.Y(n_15432)
);

NAND2xp5_ASAP7_75t_L g15433 ( 
.A(n_15305),
.B(n_15286),
.Y(n_15433)
);

OR2x2_ASAP7_75t_L g15434 ( 
.A(n_15396),
.B(n_3042),
.Y(n_15434)
);

OR2x2_ASAP7_75t_L g15435 ( 
.A(n_15308),
.B(n_3043),
.Y(n_15435)
);

NAND2xp33_ASAP7_75t_L g15436 ( 
.A(n_15374),
.B(n_15329),
.Y(n_15436)
);

OAI31xp33_ASAP7_75t_L g15437 ( 
.A1(n_15336),
.A2(n_3047),
.A3(n_3045),
.B(n_3046),
.Y(n_15437)
);

OAI221xp5_ASAP7_75t_L g15438 ( 
.A1(n_15301),
.A2(n_3048),
.B1(n_3045),
.B2(n_3047),
.C(n_3049),
.Y(n_15438)
);

OR2x2_ASAP7_75t_L g15439 ( 
.A(n_15309),
.B(n_3048),
.Y(n_15439)
);

HB1xp67_ASAP7_75t_L g15440 ( 
.A(n_15365),
.Y(n_15440)
);

OAI22xp5_ASAP7_75t_L g15441 ( 
.A1(n_15322),
.A2(n_3051),
.B1(n_3049),
.B2(n_3050),
.Y(n_15441)
);

NAND4xp25_ASAP7_75t_L g15442 ( 
.A(n_15288),
.B(n_15394),
.C(n_15381),
.D(n_15297),
.Y(n_15442)
);

BUFx3_ASAP7_75t_L g15443 ( 
.A(n_15296),
.Y(n_15443)
);

INVx1_ASAP7_75t_SL g15444 ( 
.A(n_15373),
.Y(n_15444)
);

INVx1_ASAP7_75t_L g15445 ( 
.A(n_15316),
.Y(n_15445)
);

NAND2xp5_ASAP7_75t_L g15446 ( 
.A(n_15295),
.B(n_15344),
.Y(n_15446)
);

AND2x2_ASAP7_75t_L g15447 ( 
.A(n_15350),
.B(n_3050),
.Y(n_15447)
);

NOR2xp33_ASAP7_75t_L g15448 ( 
.A(n_15325),
.B(n_3051),
.Y(n_15448)
);

INVx2_ASAP7_75t_L g15449 ( 
.A(n_15333),
.Y(n_15449)
);

INVx1_ASAP7_75t_SL g15450 ( 
.A(n_15338),
.Y(n_15450)
);

AOI22xp33_ASAP7_75t_L g15451 ( 
.A1(n_15388),
.A2(n_3054),
.B1(n_3052),
.B2(n_3053),
.Y(n_15451)
);

INVx1_ASAP7_75t_L g15452 ( 
.A(n_15353),
.Y(n_15452)
);

INVx2_ASAP7_75t_L g15453 ( 
.A(n_15377),
.Y(n_15453)
);

OAI222xp33_ASAP7_75t_L g15454 ( 
.A1(n_15354),
.A2(n_3054),
.B1(n_3056),
.B2(n_3052),
.C1(n_3053),
.C2(n_3055),
.Y(n_15454)
);

OAI21xp33_ASAP7_75t_SL g15455 ( 
.A1(n_15384),
.A2(n_3055),
.B(n_3057),
.Y(n_15455)
);

OR2x2_ASAP7_75t_L g15456 ( 
.A(n_15395),
.B(n_3058),
.Y(n_15456)
);

OAI22xp33_ASAP7_75t_L g15457 ( 
.A1(n_15379),
.A2(n_3061),
.B1(n_3059),
.B2(n_3060),
.Y(n_15457)
);

OAI22xp5_ASAP7_75t_L g15458 ( 
.A1(n_15380),
.A2(n_15360),
.B1(n_15292),
.B2(n_15289),
.Y(n_15458)
);

NAND2xp5_ASAP7_75t_L g15459 ( 
.A(n_15414),
.B(n_3059),
.Y(n_15459)
);

AOI21xp5_ASAP7_75t_L g15460 ( 
.A1(n_15304),
.A2(n_3060),
.B(n_3061),
.Y(n_15460)
);

AND2x2_ASAP7_75t_L g15461 ( 
.A(n_15300),
.B(n_3063),
.Y(n_15461)
);

INVx1_ASAP7_75t_L g15462 ( 
.A(n_15298),
.Y(n_15462)
);

INVxp67_ASAP7_75t_L g15463 ( 
.A(n_15400),
.Y(n_15463)
);

INVx1_ASAP7_75t_L g15464 ( 
.A(n_15352),
.Y(n_15464)
);

OAI32xp33_ASAP7_75t_L g15465 ( 
.A1(n_15361),
.A2(n_3066),
.A3(n_3063),
.B1(n_3065),
.B2(n_3067),
.Y(n_15465)
);

OR2x2_ASAP7_75t_L g15466 ( 
.A(n_15399),
.B(n_3065),
.Y(n_15466)
);

OAI21xp33_ASAP7_75t_L g15467 ( 
.A1(n_15363),
.A2(n_3066),
.B(n_3067),
.Y(n_15467)
);

NAND2xp5_ASAP7_75t_L g15468 ( 
.A(n_15291),
.B(n_3068),
.Y(n_15468)
);

OAI221xp5_ASAP7_75t_L g15469 ( 
.A1(n_15382),
.A2(n_3071),
.B1(n_3069),
.B2(n_3070),
.C(n_3072),
.Y(n_15469)
);

INVx2_ASAP7_75t_L g15470 ( 
.A(n_15389),
.Y(n_15470)
);

INVx2_ASAP7_75t_L g15471 ( 
.A(n_15302),
.Y(n_15471)
);

AND2x4_ASAP7_75t_L g15472 ( 
.A(n_15307),
.B(n_3071),
.Y(n_15472)
);

AND2x2_ASAP7_75t_L g15473 ( 
.A(n_15311),
.B(n_3072),
.Y(n_15473)
);

INVx1_ASAP7_75t_L g15474 ( 
.A(n_15378),
.Y(n_15474)
);

INVx2_ASAP7_75t_L g15475 ( 
.A(n_15326),
.Y(n_15475)
);

AOI222xp33_ASAP7_75t_L g15476 ( 
.A1(n_15405),
.A2(n_3075),
.B1(n_3077),
.B2(n_3073),
.C1(n_3074),
.C2(n_3076),
.Y(n_15476)
);

INVxp67_ASAP7_75t_L g15477 ( 
.A(n_15315),
.Y(n_15477)
);

INVx2_ASAP7_75t_L g15478 ( 
.A(n_15331),
.Y(n_15478)
);

AOI22xp33_ASAP7_75t_L g15479 ( 
.A1(n_15385),
.A2(n_15392),
.B1(n_15397),
.B2(n_15287),
.Y(n_15479)
);

AOI22xp5_ASAP7_75t_L g15480 ( 
.A1(n_15334),
.A2(n_3076),
.B1(n_3073),
.B2(n_3074),
.Y(n_15480)
);

INVx1_ASAP7_75t_L g15481 ( 
.A(n_15317),
.Y(n_15481)
);

NAND2xp5_ASAP7_75t_L g15482 ( 
.A(n_15410),
.B(n_3077),
.Y(n_15482)
);

NAND2xp5_ASAP7_75t_L g15483 ( 
.A(n_15348),
.B(n_15387),
.Y(n_15483)
);

OAI221xp5_ASAP7_75t_L g15484 ( 
.A1(n_15313),
.A2(n_3080),
.B1(n_3078),
.B2(n_3079),
.C(n_3081),
.Y(n_15484)
);

OAI21xp5_ASAP7_75t_L g15485 ( 
.A1(n_15330),
.A2(n_3078),
.B(n_3080),
.Y(n_15485)
);

INVx1_ASAP7_75t_L g15486 ( 
.A(n_15398),
.Y(n_15486)
);

XOR2xp5_ASAP7_75t_L g15487 ( 
.A(n_15299),
.B(n_3083),
.Y(n_15487)
);

INVx1_ASAP7_75t_L g15488 ( 
.A(n_15403),
.Y(n_15488)
);

INVx1_ASAP7_75t_SL g15489 ( 
.A(n_15332),
.Y(n_15489)
);

AOI22xp33_ASAP7_75t_L g15490 ( 
.A1(n_15404),
.A2(n_3085),
.B1(n_3083),
.B2(n_3084),
.Y(n_15490)
);

INVx1_ASAP7_75t_L g15491 ( 
.A(n_15411),
.Y(n_15491)
);

INVx1_ASAP7_75t_L g15492 ( 
.A(n_15412),
.Y(n_15492)
);

AOI221xp5_ASAP7_75t_L g15493 ( 
.A1(n_15376),
.A2(n_3087),
.B1(n_3084),
.B2(n_3086),
.C(n_3088),
.Y(n_15493)
);

INVx2_ASAP7_75t_SL g15494 ( 
.A(n_15323),
.Y(n_15494)
);

OAI31xp33_ASAP7_75t_L g15495 ( 
.A1(n_15346),
.A2(n_3090),
.A3(n_3086),
.B(n_3089),
.Y(n_15495)
);

INVx1_ASAP7_75t_L g15496 ( 
.A(n_15356),
.Y(n_15496)
);

INVxp33_ASAP7_75t_L g15497 ( 
.A(n_15347),
.Y(n_15497)
);

O2A1O1Ixp33_ASAP7_75t_SL g15498 ( 
.A1(n_15310),
.A2(n_3092),
.B(n_3089),
.C(n_3091),
.Y(n_15498)
);

NAND2xp5_ASAP7_75t_SL g15499 ( 
.A(n_15306),
.B(n_3091),
.Y(n_15499)
);

OR3x2_ASAP7_75t_L g15500 ( 
.A(n_15370),
.B(n_3093),
.C(n_3094),
.Y(n_15500)
);

OAI22xp33_ASAP7_75t_SL g15501 ( 
.A1(n_15372),
.A2(n_3097),
.B1(n_3095),
.B2(n_3096),
.Y(n_15501)
);

AOI22xp5_ASAP7_75t_L g15502 ( 
.A1(n_15383),
.A2(n_3099),
.B1(n_3095),
.B2(n_3098),
.Y(n_15502)
);

INVx1_ASAP7_75t_L g15503 ( 
.A(n_15357),
.Y(n_15503)
);

NOR2xp67_ASAP7_75t_L g15504 ( 
.A(n_15364),
.B(n_3098),
.Y(n_15504)
);

INVx1_ASAP7_75t_L g15505 ( 
.A(n_15337),
.Y(n_15505)
);

AND2x2_ASAP7_75t_L g15506 ( 
.A(n_15345),
.B(n_3099),
.Y(n_15506)
);

OAI22xp5_ASAP7_75t_L g15507 ( 
.A1(n_15368),
.A2(n_3103),
.B1(n_3100),
.B2(n_3101),
.Y(n_15507)
);

NOR2x1_ASAP7_75t_L g15508 ( 
.A(n_15328),
.B(n_3100),
.Y(n_15508)
);

NAND2xp5_ASAP7_75t_L g15509 ( 
.A(n_15343),
.B(n_3103),
.Y(n_15509)
);

INVx1_ASAP7_75t_L g15510 ( 
.A(n_15402),
.Y(n_15510)
);

OAI22xp5_ASAP7_75t_L g15511 ( 
.A1(n_15324),
.A2(n_3106),
.B1(n_3104),
.B2(n_3105),
.Y(n_15511)
);

INVx2_ASAP7_75t_L g15512 ( 
.A(n_15349),
.Y(n_15512)
);

INVx2_ASAP7_75t_L g15513 ( 
.A(n_15351),
.Y(n_15513)
);

OAI221xp5_ASAP7_75t_L g15514 ( 
.A1(n_15407),
.A2(n_3107),
.B1(n_3104),
.B2(n_3106),
.C(n_3108),
.Y(n_15514)
);

AND2x2_ASAP7_75t_L g15515 ( 
.A(n_15355),
.B(n_3108),
.Y(n_15515)
);

INVx1_ASAP7_75t_L g15516 ( 
.A(n_15409),
.Y(n_15516)
);

AOI322xp5_ASAP7_75t_L g15517 ( 
.A1(n_15359),
.A2(n_3114),
.A3(n_3113),
.B1(n_3111),
.B2(n_3109),
.C1(n_3110),
.C2(n_3112),
.Y(n_15517)
);

A2O1A1Ixp33_ASAP7_75t_L g15518 ( 
.A1(n_15393),
.A2(n_3112),
.B(n_3110),
.C(n_3111),
.Y(n_15518)
);

NAND2xp5_ASAP7_75t_L g15519 ( 
.A(n_15415),
.B(n_3113),
.Y(n_15519)
);

AND2x2_ASAP7_75t_L g15520 ( 
.A(n_15312),
.B(n_3115),
.Y(n_15520)
);

OA21x2_ASAP7_75t_L g15521 ( 
.A1(n_15314),
.A2(n_3115),
.B(n_3116),
.Y(n_15521)
);

INVx2_ASAP7_75t_L g15522 ( 
.A(n_15416),
.Y(n_15522)
);

AND2x4_ASAP7_75t_L g15523 ( 
.A(n_15321),
.B(n_3116),
.Y(n_15523)
);

AOI22xp5_ASAP7_75t_L g15524 ( 
.A1(n_15413),
.A2(n_3119),
.B1(n_3117),
.B2(n_3118),
.Y(n_15524)
);

INVxp67_ASAP7_75t_L g15525 ( 
.A(n_15366),
.Y(n_15525)
);

AND2x4_ASAP7_75t_L g15526 ( 
.A(n_15342),
.B(n_3117),
.Y(n_15526)
);

OAI211xp5_ASAP7_75t_L g15527 ( 
.A1(n_15386),
.A2(n_3120),
.B(n_3118),
.C(n_3119),
.Y(n_15527)
);

AOI221xp5_ASAP7_75t_L g15528 ( 
.A1(n_15341),
.A2(n_3122),
.B1(n_3120),
.B2(n_3121),
.C(n_3124),
.Y(n_15528)
);

INVx1_ASAP7_75t_L g15529 ( 
.A(n_15358),
.Y(n_15529)
);

OAI21xp5_ASAP7_75t_L g15530 ( 
.A1(n_15340),
.A2(n_3121),
.B(n_3122),
.Y(n_15530)
);

OAI32xp33_ASAP7_75t_L g15531 ( 
.A1(n_15362),
.A2(n_3126),
.A3(n_3124),
.B1(n_3125),
.B2(n_3127),
.Y(n_15531)
);

NAND2xp5_ASAP7_75t_L g15532 ( 
.A(n_15369),
.B(n_3125),
.Y(n_15532)
);

INVx1_ASAP7_75t_SL g15533 ( 
.A(n_15367),
.Y(n_15533)
);

NAND2xp5_ASAP7_75t_L g15534 ( 
.A(n_15375),
.B(n_3126),
.Y(n_15534)
);

NAND4xp25_ASAP7_75t_L g15535 ( 
.A(n_15451),
.B(n_3130),
.C(n_3128),
.D(n_3129),
.Y(n_15535)
);

INVx1_ASAP7_75t_L g15536 ( 
.A(n_15425),
.Y(n_15536)
);

OAI211xp5_ASAP7_75t_L g15537 ( 
.A1(n_15429),
.A2(n_3130),
.B(n_3128),
.C(n_3129),
.Y(n_15537)
);

AOI22xp33_ASAP7_75t_L g15538 ( 
.A1(n_15418),
.A2(n_3133),
.B1(n_3131),
.B2(n_3132),
.Y(n_15538)
);

NAND2xp5_ASAP7_75t_L g15539 ( 
.A(n_15421),
.B(n_15447),
.Y(n_15539)
);

OAI21xp5_ASAP7_75t_L g15540 ( 
.A1(n_15455),
.A2(n_3131),
.B(n_3132),
.Y(n_15540)
);

OAI22xp5_ASAP7_75t_L g15541 ( 
.A1(n_15500),
.A2(n_15479),
.B1(n_15480),
.B2(n_15463),
.Y(n_15541)
);

OAI321xp33_ASAP7_75t_L g15542 ( 
.A1(n_15442),
.A2(n_3135),
.A3(n_3137),
.B1(n_3133),
.B2(n_3134),
.C(n_3136),
.Y(n_15542)
);

NAND4xp25_ASAP7_75t_L g15543 ( 
.A(n_15437),
.B(n_3138),
.C(n_3136),
.D(n_3137),
.Y(n_15543)
);

NAND4xp25_ASAP7_75t_L g15544 ( 
.A(n_15427),
.B(n_3140),
.C(n_3138),
.D(n_3139),
.Y(n_15544)
);

AOI221xp5_ASAP7_75t_L g15545 ( 
.A1(n_15531),
.A2(n_15498),
.B1(n_15438),
.B2(n_15458),
.C(n_15533),
.Y(n_15545)
);

NAND3xp33_ASAP7_75t_SL g15546 ( 
.A(n_15426),
.B(n_3139),
.C(n_3140),
.Y(n_15546)
);

NAND2xp5_ASAP7_75t_L g15547 ( 
.A(n_15473),
.B(n_3141),
.Y(n_15547)
);

NAND2xp5_ASAP7_75t_SL g15548 ( 
.A(n_15417),
.B(n_3142),
.Y(n_15548)
);

NAND2xp5_ASAP7_75t_SL g15549 ( 
.A(n_15504),
.B(n_3142),
.Y(n_15549)
);

NAND2xp5_ASAP7_75t_L g15550 ( 
.A(n_15506),
.B(n_3143),
.Y(n_15550)
);

O2A1O1Ixp33_ASAP7_75t_L g15551 ( 
.A1(n_15454),
.A2(n_3146),
.B(n_3144),
.C(n_3145),
.Y(n_15551)
);

AO22x2_ASAP7_75t_L g15552 ( 
.A1(n_15452),
.A2(n_3146),
.B1(n_3144),
.B2(n_3145),
.Y(n_15552)
);

NAND4xp25_ASAP7_75t_L g15553 ( 
.A(n_15495),
.B(n_3149),
.C(n_3147),
.D(n_3148),
.Y(n_15553)
);

INVx1_ASAP7_75t_L g15554 ( 
.A(n_15521),
.Y(n_15554)
);

AOI222xp33_ASAP7_75t_L g15555 ( 
.A1(n_15436),
.A2(n_3150),
.B1(n_3152),
.B2(n_3147),
.C1(n_3149),
.C2(n_3151),
.Y(n_15555)
);

OAI211xp5_ASAP7_75t_L g15556 ( 
.A1(n_15476),
.A2(n_3154),
.B(n_3150),
.C(n_3153),
.Y(n_15556)
);

INVx1_ASAP7_75t_L g15557 ( 
.A(n_15521),
.Y(n_15557)
);

AOI221xp5_ASAP7_75t_L g15558 ( 
.A1(n_15445),
.A2(n_3155),
.B1(n_3153),
.B2(n_3154),
.C(n_3156),
.Y(n_15558)
);

AOI211xp5_ASAP7_75t_L g15559 ( 
.A1(n_15457),
.A2(n_3159),
.B(n_3156),
.C(n_3158),
.Y(n_15559)
);

NOR2xp33_ASAP7_75t_L g15560 ( 
.A(n_15467),
.B(n_3158),
.Y(n_15560)
);

OAI211xp5_ASAP7_75t_SL g15561 ( 
.A1(n_15525),
.A2(n_3161),
.B(n_3159),
.C(n_3160),
.Y(n_15561)
);

NAND2xp5_ASAP7_75t_L g15562 ( 
.A(n_15515),
.B(n_3160),
.Y(n_15562)
);

NAND2xp5_ASAP7_75t_L g15563 ( 
.A(n_15431),
.B(n_15420),
.Y(n_15563)
);

AOI22xp33_ASAP7_75t_SL g15564 ( 
.A1(n_15443),
.A2(n_3163),
.B1(n_3161),
.B2(n_3162),
.Y(n_15564)
);

AOI322xp5_ASAP7_75t_L g15565 ( 
.A1(n_15489),
.A2(n_15440),
.A3(n_15450),
.B1(n_15494),
.B2(n_15492),
.C1(n_15491),
.C2(n_15488),
.Y(n_15565)
);

NAND2xp5_ASAP7_75t_SL g15566 ( 
.A(n_15493),
.B(n_3162),
.Y(n_15566)
);

NAND2xp5_ASAP7_75t_L g15567 ( 
.A(n_15461),
.B(n_3164),
.Y(n_15567)
);

INVx1_ASAP7_75t_L g15568 ( 
.A(n_15430),
.Y(n_15568)
);

NAND2xp5_ASAP7_75t_SL g15569 ( 
.A(n_15460),
.B(n_3164),
.Y(n_15569)
);

OAI21xp33_ASAP7_75t_L g15570 ( 
.A1(n_15497),
.A2(n_3165),
.B(n_3166),
.Y(n_15570)
);

NAND2xp5_ASAP7_75t_SL g15571 ( 
.A(n_15501),
.B(n_3166),
.Y(n_15571)
);

A2O1A1Ixp33_ASAP7_75t_L g15572 ( 
.A1(n_15448),
.A2(n_3169),
.B(n_3167),
.C(n_3168),
.Y(n_15572)
);

NOR3xp33_ASAP7_75t_L g15573 ( 
.A(n_15433),
.B(n_3168),
.C(n_3169),
.Y(n_15573)
);

INVx1_ASAP7_75t_L g15574 ( 
.A(n_15472),
.Y(n_15574)
);

OA21x2_ASAP7_75t_L g15575 ( 
.A1(n_15475),
.A2(n_3170),
.B(n_3171),
.Y(n_15575)
);

OAI21xp5_ASAP7_75t_SL g15576 ( 
.A1(n_15524),
.A2(n_3170),
.B(n_3171),
.Y(n_15576)
);

NAND4xp25_ASAP7_75t_SL g15577 ( 
.A(n_15527),
.B(n_3174),
.C(n_3172),
.D(n_3173),
.Y(n_15577)
);

AOI322xp5_ASAP7_75t_L g15578 ( 
.A1(n_15499),
.A2(n_3178),
.A3(n_3177),
.B1(n_3175),
.B2(n_3172),
.C1(n_3174),
.C2(n_3176),
.Y(n_15578)
);

NAND2xp5_ASAP7_75t_L g15579 ( 
.A(n_15422),
.B(n_3176),
.Y(n_15579)
);

NOR2x1_ASAP7_75t_L g15580 ( 
.A(n_15435),
.B(n_3177),
.Y(n_15580)
);

INVxp67_ASAP7_75t_SL g15581 ( 
.A(n_15428),
.Y(n_15581)
);

NAND4xp25_ASAP7_75t_L g15582 ( 
.A(n_15459),
.B(n_3180),
.C(n_3178),
.D(n_3179),
.Y(n_15582)
);

NAND2xp5_ASAP7_75t_L g15583 ( 
.A(n_15518),
.B(n_3180),
.Y(n_15583)
);

OAI21xp33_ASAP7_75t_SL g15584 ( 
.A1(n_15508),
.A2(n_3181),
.B(n_3182),
.Y(n_15584)
);

AOI222xp33_ASAP7_75t_L g15585 ( 
.A1(n_15462),
.A2(n_15529),
.B1(n_15485),
.B2(n_15496),
.C1(n_15474),
.C2(n_15516),
.Y(n_15585)
);

OAI211xp5_ASAP7_75t_L g15586 ( 
.A1(n_15530),
.A2(n_3184),
.B(n_3182),
.C(n_3183),
.Y(n_15586)
);

AOI22xp5_ASAP7_75t_L g15587 ( 
.A1(n_15470),
.A2(n_3186),
.B1(n_3184),
.B2(n_3185),
.Y(n_15587)
);

NAND2xp5_ASAP7_75t_SL g15588 ( 
.A(n_15453),
.B(n_3185),
.Y(n_15588)
);

OAI32xp33_ASAP7_75t_L g15589 ( 
.A1(n_15456),
.A2(n_3188),
.A3(n_3186),
.B1(n_3187),
.B2(n_3189),
.Y(n_15589)
);

AOI211xp5_ASAP7_75t_SL g15590 ( 
.A1(n_15482),
.A2(n_3191),
.B(n_3188),
.C(n_3190),
.Y(n_15590)
);

OAI21xp33_ASAP7_75t_L g15591 ( 
.A1(n_15471),
.A2(n_15512),
.B(n_15478),
.Y(n_15591)
);

NAND3xp33_ASAP7_75t_L g15592 ( 
.A(n_15528),
.B(n_3190),
.C(n_3192),
.Y(n_15592)
);

OAI322xp33_ASAP7_75t_L g15593 ( 
.A1(n_15446),
.A2(n_3197),
.A3(n_3196),
.B1(n_3194),
.B2(n_3192),
.C1(n_3193),
.C2(n_3195),
.Y(n_15593)
);

OAI221xp5_ASAP7_75t_SL g15594 ( 
.A1(n_15466),
.A2(n_3196),
.B1(n_3193),
.B2(n_3195),
.C(n_3197),
.Y(n_15594)
);

NAND2xp5_ASAP7_75t_SL g15595 ( 
.A(n_15502),
.B(n_3198),
.Y(n_15595)
);

O2A1O1Ixp33_ASAP7_75t_L g15596 ( 
.A1(n_15468),
.A2(n_3200),
.B(n_3198),
.C(n_3199),
.Y(n_15596)
);

OAI21xp33_ASAP7_75t_SL g15597 ( 
.A1(n_15534),
.A2(n_3199),
.B(n_3200),
.Y(n_15597)
);

AOI221xp5_ASAP7_75t_L g15598 ( 
.A1(n_15514),
.A2(n_3203),
.B1(n_3201),
.B2(n_3202),
.C(n_3204),
.Y(n_15598)
);

AOI21xp33_ASAP7_75t_L g15599 ( 
.A1(n_15487),
.A2(n_3201),
.B(n_3202),
.Y(n_15599)
);

OAI22xp5_ASAP7_75t_L g15600 ( 
.A1(n_15469),
.A2(n_3205),
.B1(n_3203),
.B2(n_3204),
.Y(n_15600)
);

O2A1O1Ixp33_ASAP7_75t_L g15601 ( 
.A1(n_15507),
.A2(n_3207),
.B(n_3205),
.C(n_3206),
.Y(n_15601)
);

OAI21xp5_ASAP7_75t_SL g15602 ( 
.A1(n_15444),
.A2(n_3207),
.B(n_3208),
.Y(n_15602)
);

AOI21xp33_ASAP7_75t_SL g15603 ( 
.A1(n_15441),
.A2(n_3208),
.B(n_3209),
.Y(n_15603)
);

NAND2xp5_ASAP7_75t_L g15604 ( 
.A(n_15424),
.B(n_15526),
.Y(n_15604)
);

AOI211xp5_ASAP7_75t_L g15605 ( 
.A1(n_15484),
.A2(n_3211),
.B(n_3209),
.C(n_3210),
.Y(n_15605)
);

AO22x1_ASAP7_75t_L g15606 ( 
.A1(n_15523),
.A2(n_15509),
.B1(n_15486),
.B2(n_15505),
.Y(n_15606)
);

NOR2xp33_ASAP7_75t_L g15607 ( 
.A(n_15419),
.B(n_3210),
.Y(n_15607)
);

OAI221xp5_ASAP7_75t_SL g15608 ( 
.A1(n_15483),
.A2(n_3213),
.B1(n_3211),
.B2(n_3212),
.C(n_3214),
.Y(n_15608)
);

NAND2xp5_ASAP7_75t_L g15609 ( 
.A(n_15490),
.B(n_3212),
.Y(n_15609)
);

OAI21xp5_ASAP7_75t_L g15610 ( 
.A1(n_15519),
.A2(n_3213),
.B(n_3214),
.Y(n_15610)
);

AOI21xp5_ASAP7_75t_L g15611 ( 
.A1(n_15532),
.A2(n_3215),
.B(n_3216),
.Y(n_15611)
);

INVx2_ASAP7_75t_L g15612 ( 
.A(n_15434),
.Y(n_15612)
);

OAI22xp5_ASAP7_75t_L g15613 ( 
.A1(n_15439),
.A2(n_3217),
.B1(n_3215),
.B2(n_3216),
.Y(n_15613)
);

AOI21xp5_ASAP7_75t_L g15614 ( 
.A1(n_15511),
.A2(n_3217),
.B(n_3218),
.Y(n_15614)
);

OAI21xp5_ASAP7_75t_SL g15615 ( 
.A1(n_15520),
.A2(n_15510),
.B(n_15477),
.Y(n_15615)
);

NOR3xp33_ASAP7_75t_L g15616 ( 
.A(n_15513),
.B(n_3218),
.C(n_3219),
.Y(n_15616)
);

AOI211xp5_ASAP7_75t_SL g15617 ( 
.A1(n_15464),
.A2(n_3221),
.B(n_3219),
.C(n_3220),
.Y(n_15617)
);

NOR2xp33_ASAP7_75t_L g15618 ( 
.A(n_15522),
.B(n_3220),
.Y(n_15618)
);

OAI221xp5_ASAP7_75t_L g15619 ( 
.A1(n_15503),
.A2(n_3223),
.B1(n_3221),
.B2(n_3222),
.C(n_3224),
.Y(n_15619)
);

OAI221xp5_ASAP7_75t_L g15620 ( 
.A1(n_15481),
.A2(n_3227),
.B1(n_3222),
.B2(n_3226),
.C(n_3228),
.Y(n_15620)
);

OAI21xp33_ASAP7_75t_SL g15621 ( 
.A1(n_15423),
.A2(n_3228),
.B(n_3229),
.Y(n_15621)
);

AOI32xp33_ASAP7_75t_L g15622 ( 
.A1(n_15449),
.A2(n_3231),
.A3(n_3229),
.B1(n_3230),
.B2(n_3232),
.Y(n_15622)
);

OAI21xp33_ASAP7_75t_L g15623 ( 
.A1(n_15432),
.A2(n_3230),
.B(n_3231),
.Y(n_15623)
);

INVxp67_ASAP7_75t_L g15624 ( 
.A(n_15465),
.Y(n_15624)
);

INVx1_ASAP7_75t_L g15625 ( 
.A(n_15517),
.Y(n_15625)
);

AOI21xp5_ASAP7_75t_L g15626 ( 
.A1(n_15436),
.A2(n_3233),
.B(n_3234),
.Y(n_15626)
);

OA22x2_ASAP7_75t_L g15627 ( 
.A1(n_15524),
.A2(n_3235),
.B1(n_3233),
.B2(n_3234),
.Y(n_15627)
);

OR2x2_ASAP7_75t_L g15628 ( 
.A(n_15430),
.B(n_3235),
.Y(n_15628)
);

A2O1A1Ixp33_ASAP7_75t_L g15629 ( 
.A1(n_15448),
.A2(n_3239),
.B(n_3237),
.C(n_3238),
.Y(n_15629)
);

AOI221xp5_ASAP7_75t_L g15630 ( 
.A1(n_15531),
.A2(n_3239),
.B1(n_3237),
.B2(n_3238),
.C(n_3240),
.Y(n_15630)
);

NAND3xp33_ASAP7_75t_L g15631 ( 
.A(n_15451),
.B(n_3241),
.C(n_3242),
.Y(n_15631)
);

OAI221xp5_ASAP7_75t_L g15632 ( 
.A1(n_15451),
.A2(n_3243),
.B1(n_3241),
.B2(n_3242),
.C(n_3244),
.Y(n_15632)
);

OAI222xp33_ASAP7_75t_L g15633 ( 
.A1(n_15533),
.A2(n_3245),
.B1(n_3247),
.B2(n_3243),
.C1(n_3244),
.C2(n_3246),
.Y(n_15633)
);

AOI211x1_ASAP7_75t_L g15634 ( 
.A1(n_15485),
.A2(n_3247),
.B(n_3245),
.C(n_3246),
.Y(n_15634)
);

AOI21xp5_ASAP7_75t_L g15635 ( 
.A1(n_15436),
.A2(n_3248),
.B(n_3249),
.Y(n_15635)
);

AO22x1_ASAP7_75t_L g15636 ( 
.A1(n_15425),
.A2(n_3250),
.B1(n_3248),
.B2(n_3249),
.Y(n_15636)
);

OAI22xp5_ASAP7_75t_L g15637 ( 
.A1(n_15451),
.A2(n_3252),
.B1(n_3250),
.B2(n_3251),
.Y(n_15637)
);

OA22x2_ASAP7_75t_L g15638 ( 
.A1(n_15524),
.A2(n_3255),
.B1(n_3253),
.B2(n_3254),
.Y(n_15638)
);

NAND2xp5_ASAP7_75t_L g15639 ( 
.A(n_15421),
.B(n_3253),
.Y(n_15639)
);

OA22x2_ASAP7_75t_L g15640 ( 
.A1(n_15524),
.A2(n_3256),
.B1(n_3254),
.B2(n_3255),
.Y(n_15640)
);

NAND2xp5_ASAP7_75t_SL g15641 ( 
.A(n_15542),
.B(n_3257),
.Y(n_15641)
);

NOR2xp33_ASAP7_75t_L g15642 ( 
.A(n_15544),
.B(n_3257),
.Y(n_15642)
);

NOR2xp67_ASAP7_75t_L g15643 ( 
.A(n_15554),
.B(n_3258),
.Y(n_15643)
);

NAND3xp33_ASAP7_75t_SL g15644 ( 
.A(n_15565),
.B(n_3258),
.C(n_3260),
.Y(n_15644)
);

NOR2xp33_ASAP7_75t_SL g15645 ( 
.A(n_15633),
.B(n_3261),
.Y(n_15645)
);

OAI211xp5_ASAP7_75t_L g15646 ( 
.A1(n_15621),
.A2(n_3263),
.B(n_3261),
.C(n_3262),
.Y(n_15646)
);

NAND2xp5_ASAP7_75t_SL g15647 ( 
.A(n_15584),
.B(n_3263),
.Y(n_15647)
);

NAND3xp33_ASAP7_75t_L g15648 ( 
.A(n_15578),
.B(n_3264),
.C(n_3265),
.Y(n_15648)
);

NOR3xp33_ASAP7_75t_L g15649 ( 
.A(n_15591),
.B(n_3264),
.C(n_3266),
.Y(n_15649)
);

OAI221xp5_ASAP7_75t_L g15650 ( 
.A1(n_15602),
.A2(n_15630),
.B1(n_15623),
.B2(n_15576),
.C(n_15535),
.Y(n_15650)
);

AOI21xp5_ASAP7_75t_L g15651 ( 
.A1(n_15549),
.A2(n_3266),
.B(n_3267),
.Y(n_15651)
);

NOR2xp33_ASAP7_75t_L g15652 ( 
.A(n_15561),
.B(n_3267),
.Y(n_15652)
);

AOI21xp33_ASAP7_75t_L g15653 ( 
.A1(n_15601),
.A2(n_3269),
.B(n_3270),
.Y(n_15653)
);

AOI222xp33_ASAP7_75t_L g15654 ( 
.A1(n_15557),
.A2(n_3271),
.B1(n_3273),
.B2(n_3269),
.C1(n_3270),
.C2(n_3272),
.Y(n_15654)
);

NOR2xp33_ASAP7_75t_L g15655 ( 
.A(n_15570),
.B(n_3271),
.Y(n_15655)
);

AOI21xp5_ASAP7_75t_L g15656 ( 
.A1(n_15569),
.A2(n_3273),
.B(n_3274),
.Y(n_15656)
);

OAI22xp5_ASAP7_75t_L g15657 ( 
.A1(n_15624),
.A2(n_3276),
.B1(n_3274),
.B2(n_3275),
.Y(n_15657)
);

INVx1_ASAP7_75t_L g15658 ( 
.A(n_15580),
.Y(n_15658)
);

AOI211x1_ASAP7_75t_L g15659 ( 
.A1(n_15537),
.A2(n_3277),
.B(n_3275),
.C(n_3276),
.Y(n_15659)
);

AOI211xp5_ASAP7_75t_L g15660 ( 
.A1(n_15603),
.A2(n_3279),
.B(n_3277),
.C(n_3278),
.Y(n_15660)
);

INVx1_ASAP7_75t_SL g15661 ( 
.A(n_15575),
.Y(n_15661)
);

O2A1O1Ixp33_ASAP7_75t_L g15662 ( 
.A1(n_15546),
.A2(n_3280),
.B(n_3278),
.C(n_3279),
.Y(n_15662)
);

NAND2xp5_ASAP7_75t_L g15663 ( 
.A(n_15617),
.B(n_3280),
.Y(n_15663)
);

AOI221xp5_ASAP7_75t_SL g15664 ( 
.A1(n_15541),
.A2(n_3283),
.B1(n_3281),
.B2(n_3282),
.C(n_3284),
.Y(n_15664)
);

NOR4xp25_ASAP7_75t_L g15665 ( 
.A(n_15597),
.B(n_3283),
.C(n_3281),
.D(n_3282),
.Y(n_15665)
);

AOI221xp5_ASAP7_75t_SL g15666 ( 
.A1(n_15551),
.A2(n_3286),
.B1(n_3284),
.B2(n_3285),
.C(n_3287),
.Y(n_15666)
);

NOR4xp25_ASAP7_75t_L g15667 ( 
.A(n_15536),
.B(n_3287),
.C(n_3285),
.D(n_3286),
.Y(n_15667)
);

NAND4xp25_ASAP7_75t_L g15668 ( 
.A(n_15545),
.B(n_15585),
.C(n_15634),
.D(n_15631),
.Y(n_15668)
);

OAI221xp5_ASAP7_75t_L g15669 ( 
.A1(n_15540),
.A2(n_3290),
.B1(n_3288),
.B2(n_3289),
.C(n_3291),
.Y(n_15669)
);

NAND4xp25_ASAP7_75t_L g15670 ( 
.A(n_15605),
.B(n_3292),
.C(n_3290),
.D(n_3291),
.Y(n_15670)
);

NOR2xp33_ASAP7_75t_SL g15671 ( 
.A(n_15608),
.B(n_3292),
.Y(n_15671)
);

AOI221x1_ASAP7_75t_L g15672 ( 
.A1(n_15582),
.A2(n_3295),
.B1(n_3293),
.B2(n_3294),
.C(n_3296),
.Y(n_15672)
);

NAND2xp5_ASAP7_75t_L g15673 ( 
.A(n_15590),
.B(n_3293),
.Y(n_15673)
);

OAI221xp5_ASAP7_75t_SL g15674 ( 
.A1(n_15615),
.A2(n_15556),
.B1(n_15625),
.B2(n_15609),
.C(n_15581),
.Y(n_15674)
);

AOI22xp5_ASAP7_75t_L g15675 ( 
.A1(n_15577),
.A2(n_3296),
.B1(n_3294),
.B2(n_3295),
.Y(n_15675)
);

NOR3xp33_ASAP7_75t_L g15676 ( 
.A(n_15606),
.B(n_15599),
.C(n_15579),
.Y(n_15676)
);

NOR2x1_ASAP7_75t_L g15677 ( 
.A(n_15575),
.B(n_3297),
.Y(n_15677)
);

NAND2xp5_ASAP7_75t_SL g15678 ( 
.A(n_15598),
.B(n_3298),
.Y(n_15678)
);

NAND2xp5_ASAP7_75t_L g15679 ( 
.A(n_15618),
.B(n_3298),
.Y(n_15679)
);

AOI21xp5_ASAP7_75t_L g15680 ( 
.A1(n_15588),
.A2(n_3299),
.B(n_3300),
.Y(n_15680)
);

AOI21xp5_ASAP7_75t_L g15681 ( 
.A1(n_15563),
.A2(n_3299),
.B(n_3300),
.Y(n_15681)
);

INVx1_ASAP7_75t_L g15682 ( 
.A(n_15627),
.Y(n_15682)
);

AOI211xp5_ASAP7_75t_L g15683 ( 
.A1(n_15637),
.A2(n_3303),
.B(n_3301),
.C(n_3302),
.Y(n_15683)
);

AOI21xp5_ASAP7_75t_L g15684 ( 
.A1(n_15571),
.A2(n_3301),
.B(n_3302),
.Y(n_15684)
);

AOI211xp5_ASAP7_75t_SL g15685 ( 
.A1(n_15586),
.A2(n_3305),
.B(n_3303),
.C(n_3304),
.Y(n_15685)
);

AOI31xp33_ASAP7_75t_L g15686 ( 
.A1(n_15559),
.A2(n_3306),
.A3(n_3304),
.B(n_3305),
.Y(n_15686)
);

BUFx3_ASAP7_75t_L g15687 ( 
.A(n_15574),
.Y(n_15687)
);

OAI21xp33_ASAP7_75t_SL g15688 ( 
.A1(n_15553),
.A2(n_3307),
.B(n_3308),
.Y(n_15688)
);

NOR3xp33_ASAP7_75t_L g15689 ( 
.A(n_15604),
.B(n_3307),
.C(n_3308),
.Y(n_15689)
);

NOR4xp25_ASAP7_75t_SL g15690 ( 
.A(n_15594),
.B(n_3311),
.C(n_3309),
.D(n_3310),
.Y(n_15690)
);

NOR4xp25_ASAP7_75t_SL g15691 ( 
.A(n_15595),
.B(n_3312),
.C(n_3309),
.D(n_3311),
.Y(n_15691)
);

OAI21xp33_ASAP7_75t_L g15692 ( 
.A1(n_15543),
.A2(n_15539),
.B(n_15560),
.Y(n_15692)
);

NOR2xp33_ASAP7_75t_SL g15693 ( 
.A(n_15593),
.B(n_3312),
.Y(n_15693)
);

AOI22xp5_ASAP7_75t_L g15694 ( 
.A1(n_15573),
.A2(n_3315),
.B1(n_3313),
.B2(n_3314),
.Y(n_15694)
);

OAI21xp5_ASAP7_75t_L g15695 ( 
.A1(n_15592),
.A2(n_3315),
.B(n_3316),
.Y(n_15695)
);

OAI21xp5_ASAP7_75t_L g15696 ( 
.A1(n_15614),
.A2(n_3316),
.B(n_3317),
.Y(n_15696)
);

AOI21xp5_ASAP7_75t_L g15697 ( 
.A1(n_15566),
.A2(n_3317),
.B(n_3318),
.Y(n_15697)
);

INVx3_ASAP7_75t_L g15698 ( 
.A(n_15552),
.Y(n_15698)
);

AOI21xp33_ASAP7_75t_L g15699 ( 
.A1(n_15596),
.A2(n_3318),
.B(n_3319),
.Y(n_15699)
);

NAND2xp5_ASAP7_75t_L g15700 ( 
.A(n_15636),
.B(n_15622),
.Y(n_15700)
);

NOR2x1_ASAP7_75t_L g15701 ( 
.A(n_15548),
.B(n_3322),
.Y(n_15701)
);

NOR4xp25_ASAP7_75t_L g15702 ( 
.A(n_15568),
.B(n_4271),
.C(n_4263),
.D(n_3323),
.Y(n_15702)
);

OAI22xp5_ASAP7_75t_L g15703 ( 
.A1(n_15632),
.A2(n_3329),
.B1(n_3338),
.B2(n_3321),
.Y(n_15703)
);

A2O1A1Ixp33_ASAP7_75t_L g15704 ( 
.A1(n_15626),
.A2(n_3323),
.B(n_3321),
.C(n_3322),
.Y(n_15704)
);

OAI22xp33_ASAP7_75t_L g15705 ( 
.A1(n_15547),
.A2(n_3326),
.B1(n_3324),
.B2(n_3325),
.Y(n_15705)
);

NAND3xp33_ASAP7_75t_L g15706 ( 
.A(n_15572),
.B(n_15629),
.C(n_15555),
.Y(n_15706)
);

INVx1_ASAP7_75t_L g15707 ( 
.A(n_15638),
.Y(n_15707)
);

NOR3xp33_ASAP7_75t_L g15708 ( 
.A(n_15550),
.B(n_3324),
.C(n_3327),
.Y(n_15708)
);

AOI211xp5_ASAP7_75t_SL g15709 ( 
.A1(n_15628),
.A2(n_3329),
.B(n_3327),
.C(n_3328),
.Y(n_15709)
);

NOR4xp25_ASAP7_75t_L g15710 ( 
.A(n_15583),
.B(n_4271),
.C(n_3331),
.D(n_3328),
.Y(n_15710)
);

AOI221xp5_ASAP7_75t_L g15711 ( 
.A1(n_15600),
.A2(n_3332),
.B1(n_3330),
.B2(n_3331),
.C(n_3333),
.Y(n_15711)
);

OAI221xp5_ASAP7_75t_L g15712 ( 
.A1(n_15635),
.A2(n_4276),
.B1(n_4277),
.B2(n_4275),
.C(n_4274),
.Y(n_15712)
);

INVx1_ASAP7_75t_L g15713 ( 
.A(n_15640),
.Y(n_15713)
);

O2A1O1Ixp33_ASAP7_75t_SL g15714 ( 
.A1(n_15567),
.A2(n_4276),
.B(n_4274),
.C(n_3333),
.Y(n_15714)
);

NAND2xp5_ASAP7_75t_L g15715 ( 
.A(n_15616),
.B(n_3330),
.Y(n_15715)
);

NAND2xp5_ASAP7_75t_L g15716 ( 
.A(n_15607),
.B(n_3332),
.Y(n_15716)
);

OAI322xp33_ASAP7_75t_L g15717 ( 
.A1(n_15612),
.A2(n_3340),
.A3(n_3339),
.B1(n_3337),
.B2(n_3334),
.C1(n_3335),
.C2(n_3338),
.Y(n_15717)
);

AOI221x1_ASAP7_75t_L g15718 ( 
.A1(n_15611),
.A2(n_3337),
.B1(n_3334),
.B2(n_3335),
.C(n_3339),
.Y(n_15718)
);

INVx1_ASAP7_75t_L g15719 ( 
.A(n_15639),
.Y(n_15719)
);

NAND2xp5_ASAP7_75t_L g15720 ( 
.A(n_15564),
.B(n_3340),
.Y(n_15720)
);

NAND3xp33_ASAP7_75t_SL g15721 ( 
.A(n_15610),
.B(n_3341),
.C(n_3342),
.Y(n_15721)
);

AOI21xp33_ASAP7_75t_L g15722 ( 
.A1(n_15562),
.A2(n_3341),
.B(n_3343),
.Y(n_15722)
);

AOI322xp5_ASAP7_75t_L g15723 ( 
.A1(n_15558),
.A2(n_3348),
.A3(n_3347),
.B1(n_3345),
.B2(n_3343),
.C1(n_3344),
.C2(n_3346),
.Y(n_15723)
);

NAND4xp25_ASAP7_75t_L g15724 ( 
.A(n_15589),
.B(n_3346),
.C(n_3344),
.D(n_3345),
.Y(n_15724)
);

NOR2xp33_ASAP7_75t_L g15725 ( 
.A(n_15613),
.B(n_3347),
.Y(n_15725)
);

OAI22xp33_ASAP7_75t_SL g15726 ( 
.A1(n_15620),
.A2(n_15619),
.B1(n_15587),
.B2(n_15552),
.Y(n_15726)
);

NOR2xp33_ASAP7_75t_L g15727 ( 
.A(n_15538),
.B(n_3348),
.Y(n_15727)
);

AOI221xp5_ASAP7_75t_L g15728 ( 
.A1(n_15541),
.A2(n_3351),
.B1(n_3349),
.B2(n_3350),
.C(n_3353),
.Y(n_15728)
);

NOR3xp33_ASAP7_75t_L g15729 ( 
.A(n_15591),
.B(n_3349),
.C(n_3354),
.Y(n_15729)
);

OAI211xp5_ASAP7_75t_SL g15730 ( 
.A1(n_15565),
.A2(n_3362),
.B(n_3370),
.C(n_3354),
.Y(n_15730)
);

OAI221xp5_ASAP7_75t_L g15731 ( 
.A1(n_15591),
.A2(n_4266),
.B1(n_4267),
.B2(n_4265),
.C(n_4264),
.Y(n_15731)
);

INVx1_ASAP7_75t_L g15732 ( 
.A(n_15554),
.Y(n_15732)
);

AOI221xp5_ASAP7_75t_L g15733 ( 
.A1(n_15541),
.A2(n_3357),
.B1(n_3355),
.B2(n_3356),
.C(n_3358),
.Y(n_15733)
);

AOI211xp5_ASAP7_75t_L g15734 ( 
.A1(n_15561),
.A2(n_3359),
.B(n_3357),
.C(n_3358),
.Y(n_15734)
);

NAND4xp25_ASAP7_75t_SL g15735 ( 
.A(n_15565),
.B(n_3362),
.C(n_3360),
.D(n_3361),
.Y(n_15735)
);

AOI22xp5_ASAP7_75t_L g15736 ( 
.A1(n_15591),
.A2(n_3363),
.B1(n_3360),
.B2(n_3361),
.Y(n_15736)
);

AO22x1_ASAP7_75t_L g15737 ( 
.A1(n_15554),
.A2(n_3372),
.B1(n_3380),
.B2(n_3363),
.Y(n_15737)
);

OAI22xp5_ASAP7_75t_SL g15738 ( 
.A1(n_15554),
.A2(n_3366),
.B1(n_3364),
.B2(n_3365),
.Y(n_15738)
);

AOI21xp5_ASAP7_75t_L g15739 ( 
.A1(n_15549),
.A2(n_3365),
.B(n_3367),
.Y(n_15739)
);

AOI322xp5_ASAP7_75t_L g15740 ( 
.A1(n_15591),
.A2(n_3373),
.A3(n_3372),
.B1(n_3369),
.B2(n_3367),
.C1(n_3368),
.C2(n_3371),
.Y(n_15740)
);

OAI21xp33_ASAP7_75t_L g15741 ( 
.A1(n_15565),
.A2(n_3368),
.B(n_3371),
.Y(n_15741)
);

NAND2xp5_ASAP7_75t_L g15742 ( 
.A(n_15617),
.B(n_3373),
.Y(n_15742)
);

INVx1_ASAP7_75t_SL g15743 ( 
.A(n_15575),
.Y(n_15743)
);

OAI21xp33_ASAP7_75t_L g15744 ( 
.A1(n_15565),
.A2(n_3374),
.B(n_3375),
.Y(n_15744)
);

NOR2xp33_ASAP7_75t_SL g15745 ( 
.A(n_15633),
.B(n_3374),
.Y(n_15745)
);

OAI21xp5_ASAP7_75t_L g15746 ( 
.A1(n_15631),
.A2(n_3375),
.B(n_3376),
.Y(n_15746)
);

INVx1_ASAP7_75t_L g15747 ( 
.A(n_15677),
.Y(n_15747)
);

NOR4xp25_ASAP7_75t_L g15748 ( 
.A(n_15741),
.B(n_3378),
.C(n_3376),
.D(n_3377),
.Y(n_15748)
);

NOR2xp33_ASAP7_75t_L g15749 ( 
.A(n_15744),
.B(n_3377),
.Y(n_15749)
);

NOR2xp67_ASAP7_75t_L g15750 ( 
.A(n_15698),
.B(n_3379),
.Y(n_15750)
);

OAI322xp33_ASAP7_75t_L g15751 ( 
.A1(n_15645),
.A2(n_3383),
.A3(n_3382),
.B1(n_3380),
.B2(n_3378),
.C1(n_3379),
.C2(n_3381),
.Y(n_15751)
);

NOR3xp33_ASAP7_75t_L g15752 ( 
.A(n_15674),
.B(n_4259),
.C(n_4258),
.Y(n_15752)
);

OAI221xp5_ASAP7_75t_L g15753 ( 
.A1(n_15675),
.A2(n_3383),
.B1(n_3381),
.B2(n_3382),
.C(n_3384),
.Y(n_15753)
);

INVx1_ASAP7_75t_L g15754 ( 
.A(n_15698),
.Y(n_15754)
);

NOR2xp33_ASAP7_75t_L g15755 ( 
.A(n_15730),
.B(n_3384),
.Y(n_15755)
);

NAND2xp5_ASAP7_75t_L g15756 ( 
.A(n_15709),
.B(n_3385),
.Y(n_15756)
);

OAI21xp5_ASAP7_75t_SL g15757 ( 
.A1(n_15685),
.A2(n_4263),
.B(n_4262),
.Y(n_15757)
);

NAND2xp5_ASAP7_75t_L g15758 ( 
.A(n_15643),
.B(n_3385),
.Y(n_15758)
);

NOR2xp33_ASAP7_75t_L g15759 ( 
.A(n_15644),
.B(n_3386),
.Y(n_15759)
);

OAI211xp5_ASAP7_75t_L g15760 ( 
.A1(n_15710),
.A2(n_4268),
.B(n_4269),
.C(n_4267),
.Y(n_15760)
);

HB1xp67_ASAP7_75t_L g15761 ( 
.A(n_15661),
.Y(n_15761)
);

NAND2xp5_ASAP7_75t_L g15762 ( 
.A(n_15743),
.B(n_3386),
.Y(n_15762)
);

OAI22xp5_ASAP7_75t_L g15763 ( 
.A1(n_15694),
.A2(n_3389),
.B1(n_3387),
.B2(n_3388),
.Y(n_15763)
);

INVx2_ASAP7_75t_L g15764 ( 
.A(n_15687),
.Y(n_15764)
);

NOR3xp33_ASAP7_75t_SL g15765 ( 
.A(n_15735),
.B(n_3387),
.C(n_3388),
.Y(n_15765)
);

AO21x1_ASAP7_75t_L g15766 ( 
.A1(n_15647),
.A2(n_3389),
.B(n_3390),
.Y(n_15766)
);

INVx1_ASAP7_75t_L g15767 ( 
.A(n_15663),
.Y(n_15767)
);

NAND5xp2_ASAP7_75t_L g15768 ( 
.A(n_15745),
.B(n_3407),
.C(n_3415),
.D(n_3399),
.E(n_3390),
.Y(n_15768)
);

AOI322xp5_ASAP7_75t_L g15769 ( 
.A1(n_15688),
.A2(n_3396),
.A3(n_3395),
.B1(n_3393),
.B2(n_3391),
.C1(n_3392),
.C2(n_3394),
.Y(n_15769)
);

NOR2xp67_ASAP7_75t_L g15770 ( 
.A(n_15646),
.B(n_3393),
.Y(n_15770)
);

INVx1_ASAP7_75t_L g15771 ( 
.A(n_15742),
.Y(n_15771)
);

INVxp67_ASAP7_75t_SL g15772 ( 
.A(n_15738),
.Y(n_15772)
);

INVxp67_ASAP7_75t_L g15773 ( 
.A(n_15652),
.Y(n_15773)
);

NAND4xp25_ASAP7_75t_L g15774 ( 
.A(n_15734),
.B(n_3395),
.C(n_3392),
.D(n_3394),
.Y(n_15774)
);

AOI211xp5_ASAP7_75t_L g15775 ( 
.A1(n_15653),
.A2(n_3399),
.B(n_3396),
.C(n_3397),
.Y(n_15775)
);

AND2x2_ASAP7_75t_L g15776 ( 
.A(n_15690),
.B(n_3397),
.Y(n_15776)
);

NOR2xp33_ASAP7_75t_L g15777 ( 
.A(n_15670),
.B(n_3400),
.Y(n_15777)
);

NAND3xp33_ASAP7_75t_SL g15778 ( 
.A(n_15691),
.B(n_3400),
.C(n_3401),
.Y(n_15778)
);

NOR3xp33_ASAP7_75t_L g15779 ( 
.A(n_15668),
.B(n_4268),
.C(n_4266),
.Y(n_15779)
);

INVx1_ASAP7_75t_L g15780 ( 
.A(n_15673),
.Y(n_15780)
);

NOR2xp33_ASAP7_75t_L g15781 ( 
.A(n_15686),
.B(n_3401),
.Y(n_15781)
);

NAND2xp5_ASAP7_75t_L g15782 ( 
.A(n_15667),
.B(n_3402),
.Y(n_15782)
);

INVx2_ASAP7_75t_L g15783 ( 
.A(n_15737),
.Y(n_15783)
);

INVx1_ASAP7_75t_L g15784 ( 
.A(n_15714),
.Y(n_15784)
);

NOR2xp33_ASAP7_75t_L g15785 ( 
.A(n_15669),
.B(n_3403),
.Y(n_15785)
);

NOR3xp33_ASAP7_75t_SL g15786 ( 
.A(n_15692),
.B(n_3403),
.C(n_3404),
.Y(n_15786)
);

NOR3x1_ASAP7_75t_L g15787 ( 
.A(n_15648),
.B(n_3404),
.C(n_3405),
.Y(n_15787)
);

AOI221xp5_ASAP7_75t_SL g15788 ( 
.A1(n_15697),
.A2(n_3422),
.B1(n_3430),
.B2(n_3414),
.C(n_3405),
.Y(n_15788)
);

AOI21xp5_ASAP7_75t_L g15789 ( 
.A1(n_15658),
.A2(n_3406),
.B(n_3408),
.Y(n_15789)
);

INVx2_ASAP7_75t_L g15790 ( 
.A(n_15659),
.Y(n_15790)
);

INVx2_ASAP7_75t_L g15791 ( 
.A(n_15732),
.Y(n_15791)
);

OAI221xp5_ASAP7_75t_L g15792 ( 
.A1(n_15666),
.A2(n_3409),
.B1(n_3406),
.B2(n_3408),
.C(n_3410),
.Y(n_15792)
);

OAI21xp33_ASAP7_75t_SL g15793 ( 
.A1(n_15641),
.A2(n_15724),
.B(n_15701),
.Y(n_15793)
);

OAI22xp33_ASAP7_75t_L g15794 ( 
.A1(n_15693),
.A2(n_3412),
.B1(n_3410),
.B2(n_3411),
.Y(n_15794)
);

AOI211xp5_ASAP7_75t_L g15795 ( 
.A1(n_15699),
.A2(n_3414),
.B(n_3412),
.C(n_3413),
.Y(n_15795)
);

NAND4xp25_ASAP7_75t_L g15796 ( 
.A(n_15676),
.B(n_3416),
.C(n_3413),
.D(n_3415),
.Y(n_15796)
);

NOR2x1_ASAP7_75t_L g15797 ( 
.A(n_15657),
.B(n_3416),
.Y(n_15797)
);

AOI211x1_ASAP7_75t_L g15798 ( 
.A1(n_15650),
.A2(n_3419),
.B(n_3417),
.C(n_3418),
.Y(n_15798)
);

NAND4xp25_ASAP7_75t_L g15799 ( 
.A(n_15642),
.B(n_3419),
.C(n_3417),
.D(n_3418),
.Y(n_15799)
);

NAND2xp33_ASAP7_75t_L g15800 ( 
.A(n_15649),
.B(n_3420),
.Y(n_15800)
);

NAND4xp25_ASAP7_75t_SL g15801 ( 
.A(n_15664),
.B(n_3422),
.C(n_3420),
.D(n_3421),
.Y(n_15801)
);

NOR2xp33_ASAP7_75t_L g15802 ( 
.A(n_15721),
.B(n_3421),
.Y(n_15802)
);

NAND3xp33_ASAP7_75t_L g15803 ( 
.A(n_15729),
.B(n_3423),
.C(n_3424),
.Y(n_15803)
);

INVx1_ASAP7_75t_L g15804 ( 
.A(n_15720),
.Y(n_15804)
);

OAI211xp5_ASAP7_75t_L g15805 ( 
.A1(n_15672),
.A2(n_4253),
.B(n_4254),
.C(n_4252),
.Y(n_15805)
);

NAND4xp25_ASAP7_75t_L g15806 ( 
.A(n_15671),
.B(n_3426),
.C(n_3424),
.D(n_3425),
.Y(n_15806)
);

NAND2xp5_ASAP7_75t_L g15807 ( 
.A(n_15702),
.B(n_15665),
.Y(n_15807)
);

HB1xp67_ASAP7_75t_L g15808 ( 
.A(n_15718),
.Y(n_15808)
);

AOI22xp33_ASAP7_75t_L g15809 ( 
.A1(n_15682),
.A2(n_3427),
.B1(n_3425),
.B2(n_3426),
.Y(n_15809)
);

AOI21xp5_ASAP7_75t_L g15810 ( 
.A1(n_15684),
.A2(n_3427),
.B(n_3428),
.Y(n_15810)
);

NOR3x1_ASAP7_75t_L g15811 ( 
.A(n_15712),
.B(n_3429),
.C(n_3430),
.Y(n_15811)
);

NOR4xp75_ASAP7_75t_L g15812 ( 
.A(n_15695),
.B(n_3432),
.C(n_3429),
.D(n_3431),
.Y(n_15812)
);

NAND3xp33_ASAP7_75t_L g15813 ( 
.A(n_15711),
.B(n_3431),
.C(n_3432),
.Y(n_15813)
);

NOR2xp33_ASAP7_75t_L g15814 ( 
.A(n_15707),
.B(n_3433),
.Y(n_15814)
);

NAND3xp33_ASAP7_75t_L g15815 ( 
.A(n_15660),
.B(n_3434),
.C(n_3435),
.Y(n_15815)
);

NOR2x1_ASAP7_75t_L g15816 ( 
.A(n_15717),
.B(n_3434),
.Y(n_15816)
);

AND4x1_ASAP7_75t_L g15817 ( 
.A(n_15683),
.B(n_3443),
.C(n_3451),
.D(n_3435),
.Y(n_15817)
);

NOR2xp33_ASAP7_75t_L g15818 ( 
.A(n_15713),
.B(n_3436),
.Y(n_15818)
);

AND4x1_ASAP7_75t_L g15819 ( 
.A(n_15681),
.B(n_3445),
.C(n_3454),
.D(n_3436),
.Y(n_15819)
);

NAND3xp33_ASAP7_75t_L g15820 ( 
.A(n_15689),
.B(n_3437),
.C(n_3438),
.Y(n_15820)
);

NOR2xp67_ASAP7_75t_L g15821 ( 
.A(n_15731),
.B(n_3438),
.Y(n_15821)
);

NAND2xp5_ASAP7_75t_L g15822 ( 
.A(n_15708),
.B(n_3437),
.Y(n_15822)
);

NAND4xp25_ASAP7_75t_L g15823 ( 
.A(n_15662),
.B(n_3441),
.C(n_3439),
.D(n_3440),
.Y(n_15823)
);

AND3x2_ASAP7_75t_L g15824 ( 
.A(n_15728),
.B(n_4256),
.C(n_4255),
.Y(n_15824)
);

NAND2xp5_ASAP7_75t_SL g15825 ( 
.A(n_15726),
.B(n_3441),
.Y(n_15825)
);

AOI21xp5_ASAP7_75t_L g15826 ( 
.A1(n_15700),
.A2(n_3442),
.B(n_3444),
.Y(n_15826)
);

AOI211xp5_ASAP7_75t_L g15827 ( 
.A1(n_15703),
.A2(n_3445),
.B(n_3442),
.C(n_3444),
.Y(n_15827)
);

OAI21xp5_ASAP7_75t_SL g15828 ( 
.A1(n_15655),
.A2(n_4261),
.B(n_4260),
.Y(n_15828)
);

NAND2xp5_ASAP7_75t_L g15829 ( 
.A(n_15705),
.B(n_3446),
.Y(n_15829)
);

NOR4xp25_ASAP7_75t_SL g15830 ( 
.A(n_15678),
.B(n_4260),
.C(n_3448),
.D(n_3446),
.Y(n_15830)
);

NOR3xp33_ASAP7_75t_L g15831 ( 
.A(n_15716),
.B(n_4270),
.C(n_4269),
.Y(n_15831)
);

NAND2xp5_ASAP7_75t_SL g15832 ( 
.A(n_15723),
.B(n_3447),
.Y(n_15832)
);

INVx1_ASAP7_75t_L g15833 ( 
.A(n_15715),
.Y(n_15833)
);

OAI21xp5_ASAP7_75t_L g15834 ( 
.A1(n_15651),
.A2(n_3448),
.B(n_3449),
.Y(n_15834)
);

INVxp67_ASAP7_75t_SL g15835 ( 
.A(n_15736),
.Y(n_15835)
);

NAND2xp5_ASAP7_75t_L g15836 ( 
.A(n_15704),
.B(n_3449),
.Y(n_15836)
);

AOI222xp33_ASAP7_75t_L g15837 ( 
.A1(n_15727),
.A2(n_3453),
.B1(n_3456),
.B2(n_3457),
.C1(n_3452),
.C2(n_3455),
.Y(n_15837)
);

NOR3x1_ASAP7_75t_L g15838 ( 
.A(n_15746),
.B(n_3450),
.C(n_3452),
.Y(n_15838)
);

NAND3xp33_ASAP7_75t_L g15839 ( 
.A(n_15733),
.B(n_3450),
.C(n_3453),
.Y(n_15839)
);

INVx1_ASAP7_75t_L g15840 ( 
.A(n_15679),
.Y(n_15840)
);

INVx1_ASAP7_75t_L g15841 ( 
.A(n_15725),
.Y(n_15841)
);

NAND2xp5_ASAP7_75t_L g15842 ( 
.A(n_15680),
.B(n_3456),
.Y(n_15842)
);

INVx2_ASAP7_75t_L g15843 ( 
.A(n_15719),
.Y(n_15843)
);

AND2x2_ASAP7_75t_L g15844 ( 
.A(n_15696),
.B(n_3457),
.Y(n_15844)
);

NOR3x1_ASAP7_75t_L g15845 ( 
.A(n_15706),
.B(n_3458),
.C(n_3459),
.Y(n_15845)
);

INVx1_ASAP7_75t_L g15846 ( 
.A(n_15739),
.Y(n_15846)
);

AOI21xp5_ASAP7_75t_L g15847 ( 
.A1(n_15656),
.A2(n_15722),
.B(n_15654),
.Y(n_15847)
);

AOI21xp33_ASAP7_75t_L g15848 ( 
.A1(n_15740),
.A2(n_3458),
.B(n_3459),
.Y(n_15848)
);

A2O1A1Ixp33_ASAP7_75t_L g15849 ( 
.A1(n_15643),
.A2(n_3462),
.B(n_3460),
.C(n_3461),
.Y(n_15849)
);

OAI21xp5_ASAP7_75t_L g15850 ( 
.A1(n_15688),
.A2(n_3460),
.B(n_3461),
.Y(n_15850)
);

NAND2xp5_ASAP7_75t_L g15851 ( 
.A(n_15709),
.B(n_3462),
.Y(n_15851)
);

AOI221xp5_ASAP7_75t_L g15852 ( 
.A1(n_15748),
.A2(n_3465),
.B1(n_3463),
.B2(n_3464),
.C(n_3466),
.Y(n_15852)
);

NOR2xp33_ASAP7_75t_SL g15853 ( 
.A(n_15750),
.B(n_3463),
.Y(n_15853)
);

NAND3xp33_ASAP7_75t_L g15854 ( 
.A(n_15779),
.B(n_3465),
.C(n_3466),
.Y(n_15854)
);

NOR2x1_ASAP7_75t_L g15855 ( 
.A(n_15747),
.B(n_3468),
.Y(n_15855)
);

INVx1_ASAP7_75t_L g15856 ( 
.A(n_15776),
.Y(n_15856)
);

NOR3xp33_ASAP7_75t_SL g15857 ( 
.A(n_15794),
.B(n_3468),
.C(n_3469),
.Y(n_15857)
);

NOR3xp33_ASAP7_75t_SL g15858 ( 
.A(n_15825),
.B(n_3469),
.C(n_3470),
.Y(n_15858)
);

NAND4xp25_ASAP7_75t_L g15859 ( 
.A(n_15768),
.B(n_15752),
.C(n_15838),
.D(n_15755),
.Y(n_15859)
);

NAND2xp5_ASAP7_75t_L g15860 ( 
.A(n_15814),
.B(n_15818),
.Y(n_15860)
);

AND2x2_ASAP7_75t_L g15861 ( 
.A(n_15765),
.B(n_3470),
.Y(n_15861)
);

INVx1_ASAP7_75t_L g15862 ( 
.A(n_15762),
.Y(n_15862)
);

AND2x2_ASAP7_75t_L g15863 ( 
.A(n_15786),
.B(n_3471),
.Y(n_15863)
);

AOI21x1_ASAP7_75t_L g15864 ( 
.A1(n_15808),
.A2(n_15784),
.B(n_15761),
.Y(n_15864)
);

OR2x2_ASAP7_75t_L g15865 ( 
.A(n_15778),
.B(n_4250),
.Y(n_15865)
);

NAND2xp5_ASAP7_75t_SL g15866 ( 
.A(n_15837),
.B(n_3472),
.Y(n_15866)
);

NAND4xp75_ASAP7_75t_L g15867 ( 
.A(n_15845),
.B(n_3474),
.C(n_3472),
.D(n_3473),
.Y(n_15867)
);

NOR2xp33_ASAP7_75t_L g15868 ( 
.A(n_15799),
.B(n_3473),
.Y(n_15868)
);

INVx1_ASAP7_75t_L g15869 ( 
.A(n_15758),
.Y(n_15869)
);

AND2x2_ASAP7_75t_L g15870 ( 
.A(n_15790),
.B(n_3475),
.Y(n_15870)
);

OR2x2_ASAP7_75t_L g15871 ( 
.A(n_15782),
.B(n_4253),
.Y(n_15871)
);

NAND2xp5_ASAP7_75t_L g15872 ( 
.A(n_15769),
.B(n_3475),
.Y(n_15872)
);

NOR3xp33_ASAP7_75t_L g15873 ( 
.A(n_15754),
.B(n_3476),
.C(n_3477),
.Y(n_15873)
);

INVx1_ASAP7_75t_L g15874 ( 
.A(n_15756),
.Y(n_15874)
);

NOR3xp33_ASAP7_75t_SL g15875 ( 
.A(n_15793),
.B(n_15806),
.C(n_15760),
.Y(n_15875)
);

NAND2xp5_ASAP7_75t_L g15876 ( 
.A(n_15849),
.B(n_3476),
.Y(n_15876)
);

NAND2xp5_ASAP7_75t_L g15877 ( 
.A(n_15789),
.B(n_3477),
.Y(n_15877)
);

OR2x2_ASAP7_75t_L g15878 ( 
.A(n_15851),
.B(n_4257),
.Y(n_15878)
);

HB1xp67_ASAP7_75t_L g15879 ( 
.A(n_15812),
.Y(n_15879)
);

INVx1_ASAP7_75t_L g15880 ( 
.A(n_15766),
.Y(n_15880)
);

NOR2xp33_ASAP7_75t_L g15881 ( 
.A(n_15823),
.B(n_15792),
.Y(n_15881)
);

NOR3xp33_ASAP7_75t_L g15882 ( 
.A(n_15791),
.B(n_3478),
.C(n_3479),
.Y(n_15882)
);

INVx2_ASAP7_75t_L g15883 ( 
.A(n_15798),
.Y(n_15883)
);

NAND3xp33_ASAP7_75t_L g15884 ( 
.A(n_15775),
.B(n_3478),
.C(n_3480),
.Y(n_15884)
);

NAND2xp5_ASAP7_75t_L g15885 ( 
.A(n_15770),
.B(n_3481),
.Y(n_15885)
);

OR2x2_ASAP7_75t_L g15886 ( 
.A(n_15774),
.B(n_15796),
.Y(n_15886)
);

INVx1_ASAP7_75t_L g15887 ( 
.A(n_15819),
.Y(n_15887)
);

NOR3xp33_ASAP7_75t_L g15888 ( 
.A(n_15764),
.B(n_15772),
.C(n_15843),
.Y(n_15888)
);

NAND2xp33_ASAP7_75t_SL g15889 ( 
.A(n_15830),
.B(n_3481),
.Y(n_15889)
);

NOR2xp33_ASAP7_75t_L g15890 ( 
.A(n_15757),
.B(n_3482),
.Y(n_15890)
);

INVx1_ASAP7_75t_L g15891 ( 
.A(n_15807),
.Y(n_15891)
);

NAND2xp33_ASAP7_75t_L g15892 ( 
.A(n_15831),
.B(n_3482),
.Y(n_15892)
);

AOI21xp5_ASAP7_75t_L g15893 ( 
.A1(n_15800),
.A2(n_3484),
.B(n_3485),
.Y(n_15893)
);

INVx2_ASAP7_75t_L g15894 ( 
.A(n_15824),
.Y(n_15894)
);

INVx1_ASAP7_75t_L g15895 ( 
.A(n_15817),
.Y(n_15895)
);

INVx1_ASAP7_75t_L g15896 ( 
.A(n_15781),
.Y(n_15896)
);

AOI221x1_ASAP7_75t_L g15897 ( 
.A1(n_15783),
.A2(n_3486),
.B1(n_3484),
.B2(n_3485),
.C(n_3487),
.Y(n_15897)
);

NAND2xp5_ASAP7_75t_SL g15898 ( 
.A(n_15795),
.B(n_3486),
.Y(n_15898)
);

INVx1_ASAP7_75t_L g15899 ( 
.A(n_15805),
.Y(n_15899)
);

AND2x2_ASAP7_75t_L g15900 ( 
.A(n_15816),
.B(n_3487),
.Y(n_15900)
);

AND2x2_ASAP7_75t_L g15901 ( 
.A(n_15844),
.B(n_3488),
.Y(n_15901)
);

AND2x2_ASAP7_75t_L g15902 ( 
.A(n_15850),
.B(n_3488),
.Y(n_15902)
);

INVx1_ASAP7_75t_L g15903 ( 
.A(n_15759),
.Y(n_15903)
);

NOR3xp33_ASAP7_75t_L g15904 ( 
.A(n_15773),
.B(n_3489),
.C(n_3490),
.Y(n_15904)
);

INVx2_ASAP7_75t_SL g15905 ( 
.A(n_15797),
.Y(n_15905)
);

NOR3xp33_ASAP7_75t_L g15906 ( 
.A(n_15841),
.B(n_3489),
.C(n_3490),
.Y(n_15906)
);

NOR3xp33_ASAP7_75t_L g15907 ( 
.A(n_15846),
.B(n_3491),
.C(n_3492),
.Y(n_15907)
);

INVx1_ASAP7_75t_L g15908 ( 
.A(n_15822),
.Y(n_15908)
);

OAI211xp5_ASAP7_75t_L g15909 ( 
.A1(n_15828),
.A2(n_15826),
.B(n_15848),
.C(n_15827),
.Y(n_15909)
);

NOR2x1_ASAP7_75t_L g15910 ( 
.A(n_15751),
.B(n_15820),
.Y(n_15910)
);

AND2x2_ASAP7_75t_L g15911 ( 
.A(n_15777),
.B(n_15787),
.Y(n_15911)
);

OAI21xp33_ASAP7_75t_SL g15912 ( 
.A1(n_15801),
.A2(n_3491),
.B(n_3492),
.Y(n_15912)
);

AOI221xp5_ASAP7_75t_L g15913 ( 
.A1(n_15749),
.A2(n_3495),
.B1(n_3493),
.B2(n_3494),
.C(n_3496),
.Y(n_15913)
);

NOR2xp33_ASAP7_75t_L g15914 ( 
.A(n_15803),
.B(n_3493),
.Y(n_15914)
);

AOI22xp33_ASAP7_75t_SL g15915 ( 
.A1(n_15802),
.A2(n_3496),
.B1(n_3494),
.B2(n_3495),
.Y(n_15915)
);

NAND4xp25_ASAP7_75t_L g15916 ( 
.A(n_15811),
.B(n_3499),
.C(n_3497),
.D(n_3498),
.Y(n_15916)
);

OAI22xp5_ASAP7_75t_L g15917 ( 
.A1(n_15815),
.A2(n_3500),
.B1(n_3497),
.B2(n_3498),
.Y(n_15917)
);

CKINVDCx20_ASAP7_75t_L g15918 ( 
.A(n_15788),
.Y(n_15918)
);

NAND3xp33_ASAP7_75t_L g15919 ( 
.A(n_15829),
.B(n_3500),
.C(n_3501),
.Y(n_15919)
);

AOI22xp5_ASAP7_75t_L g15920 ( 
.A1(n_15835),
.A2(n_3503),
.B1(n_3501),
.B2(n_3502),
.Y(n_15920)
);

NOR2xp33_ASAP7_75t_L g15921 ( 
.A(n_15753),
.B(n_3502),
.Y(n_15921)
);

NOR2xp33_ASAP7_75t_L g15922 ( 
.A(n_15842),
.B(n_3504),
.Y(n_15922)
);

INVx1_ASAP7_75t_L g15923 ( 
.A(n_15836),
.Y(n_15923)
);

INVx1_ASAP7_75t_L g15924 ( 
.A(n_15839),
.Y(n_15924)
);

AOI221x1_ASAP7_75t_L g15925 ( 
.A1(n_15767),
.A2(n_3507),
.B1(n_3505),
.B2(n_3506),
.C(n_3508),
.Y(n_15925)
);

NOR3xp33_ASAP7_75t_L g15926 ( 
.A(n_15780),
.B(n_3505),
.C(n_3506),
.Y(n_15926)
);

INVx1_ASAP7_75t_SL g15927 ( 
.A(n_15810),
.Y(n_15927)
);

A2O1A1Ixp33_ASAP7_75t_L g15928 ( 
.A1(n_15785),
.A2(n_3509),
.B(n_3507),
.C(n_3508),
.Y(n_15928)
);

NOR4xp25_ASAP7_75t_L g15929 ( 
.A(n_15832),
.B(n_3511),
.C(n_3509),
.D(n_3510),
.Y(n_15929)
);

NOR3x1_ASAP7_75t_L g15930 ( 
.A(n_15834),
.B(n_3512),
.C(n_3513),
.Y(n_15930)
);

NAND3xp33_ASAP7_75t_L g15931 ( 
.A(n_15813),
.B(n_3512),
.C(n_3514),
.Y(n_15931)
);

AOI221x1_ASAP7_75t_L g15932 ( 
.A1(n_15771),
.A2(n_3516),
.B1(n_3514),
.B2(n_3515),
.C(n_3517),
.Y(n_15932)
);

NAND2xp5_ASAP7_75t_L g15933 ( 
.A(n_15809),
.B(n_3515),
.Y(n_15933)
);

NAND4xp25_ASAP7_75t_L g15934 ( 
.A(n_15821),
.B(n_3518),
.C(n_3516),
.D(n_3517),
.Y(n_15934)
);

NAND2xp5_ASAP7_75t_SL g15935 ( 
.A(n_15763),
.B(n_3519),
.Y(n_15935)
);

NOR4xp25_ASAP7_75t_L g15936 ( 
.A(n_15804),
.B(n_3521),
.C(n_3519),
.D(n_3520),
.Y(n_15936)
);

NOR3xp33_ASAP7_75t_L g15937 ( 
.A(n_15840),
.B(n_3520),
.C(n_3521),
.Y(n_15937)
);

NAND2xp5_ASAP7_75t_L g15938 ( 
.A(n_15847),
.B(n_3522),
.Y(n_15938)
);

NOR3xp33_ASAP7_75t_SL g15939 ( 
.A(n_15833),
.B(n_3522),
.C(n_3523),
.Y(n_15939)
);

NAND3xp33_ASAP7_75t_L g15940 ( 
.A(n_15779),
.B(n_3524),
.C(n_3525),
.Y(n_15940)
);

AND2x2_ASAP7_75t_L g15941 ( 
.A(n_15779),
.B(n_3525),
.Y(n_15941)
);

AOI21xp5_ASAP7_75t_L g15942 ( 
.A1(n_15825),
.A2(n_3526),
.B(n_3527),
.Y(n_15942)
);

NOR2x1_ASAP7_75t_L g15943 ( 
.A(n_15750),
.B(n_3528),
.Y(n_15943)
);

INVx1_ASAP7_75t_L g15944 ( 
.A(n_15776),
.Y(n_15944)
);

NAND2xp5_ASAP7_75t_L g15945 ( 
.A(n_15750),
.B(n_3528),
.Y(n_15945)
);

OAI21xp5_ASAP7_75t_L g15946 ( 
.A1(n_15912),
.A2(n_3529),
.B(n_3530),
.Y(n_15946)
);

INVx1_ASAP7_75t_L g15947 ( 
.A(n_15855),
.Y(n_15947)
);

OA22x2_ASAP7_75t_L g15948 ( 
.A1(n_15870),
.A2(n_3533),
.B1(n_3531),
.B2(n_3532),
.Y(n_15948)
);

NOR2xp33_ASAP7_75t_L g15949 ( 
.A(n_15916),
.B(n_3531),
.Y(n_15949)
);

NAND2xp5_ASAP7_75t_L g15950 ( 
.A(n_15943),
.B(n_4273),
.Y(n_15950)
);

NAND2xp5_ASAP7_75t_SL g15951 ( 
.A(n_15936),
.B(n_3532),
.Y(n_15951)
);

NOR2xp67_ASAP7_75t_L g15952 ( 
.A(n_15934),
.B(n_3534),
.Y(n_15952)
);

OAI211xp5_ASAP7_75t_SL g15953 ( 
.A1(n_15875),
.A2(n_3536),
.B(n_3534),
.C(n_3535),
.Y(n_15953)
);

AOI211xp5_ASAP7_75t_L g15954 ( 
.A1(n_15917),
.A2(n_3537),
.B(n_3535),
.C(n_3536),
.Y(n_15954)
);

NAND3xp33_ASAP7_75t_SL g15955 ( 
.A(n_15853),
.B(n_3546),
.C(n_3538),
.Y(n_15955)
);

INVx1_ASAP7_75t_L g15956 ( 
.A(n_15945),
.Y(n_15956)
);

INVx1_ASAP7_75t_SL g15957 ( 
.A(n_15889),
.Y(n_15957)
);

INVx1_ASAP7_75t_SL g15958 ( 
.A(n_15865),
.Y(n_15958)
);

NAND2xp5_ASAP7_75t_L g15959 ( 
.A(n_15907),
.B(n_4252),
.Y(n_15959)
);

NOR2xp33_ASAP7_75t_SL g15960 ( 
.A(n_15879),
.B(n_15856),
.Y(n_15960)
);

INVx1_ASAP7_75t_L g15961 ( 
.A(n_15901),
.Y(n_15961)
);

INVx1_ASAP7_75t_L g15962 ( 
.A(n_15861),
.Y(n_15962)
);

NOR3x1_ASAP7_75t_L g15963 ( 
.A(n_15867),
.B(n_3538),
.C(n_3539),
.Y(n_15963)
);

NAND2xp5_ASAP7_75t_L g15964 ( 
.A(n_15873),
.B(n_4255),
.Y(n_15964)
);

AND2x2_ASAP7_75t_L g15965 ( 
.A(n_15863),
.B(n_3539),
.Y(n_15965)
);

NOR2x1_ASAP7_75t_L g15966 ( 
.A(n_15880),
.B(n_3540),
.Y(n_15966)
);

NOR2xp33_ASAP7_75t_L g15967 ( 
.A(n_15854),
.B(n_3540),
.Y(n_15967)
);

INVx1_ASAP7_75t_L g15968 ( 
.A(n_15885),
.Y(n_15968)
);

NOR3xp33_ASAP7_75t_L g15969 ( 
.A(n_15938),
.B(n_3541),
.C(n_3542),
.Y(n_15969)
);

HB1xp67_ASAP7_75t_L g15970 ( 
.A(n_15897),
.Y(n_15970)
);

NOR2x1p5_ASAP7_75t_L g15971 ( 
.A(n_15859),
.B(n_3541),
.Y(n_15971)
);

NOR3xp33_ASAP7_75t_L g15972 ( 
.A(n_15864),
.B(n_15888),
.C(n_15944),
.Y(n_15972)
);

INVx1_ASAP7_75t_L g15973 ( 
.A(n_15941),
.Y(n_15973)
);

INVx1_ASAP7_75t_L g15974 ( 
.A(n_15871),
.Y(n_15974)
);

NAND2xp5_ASAP7_75t_L g15975 ( 
.A(n_15915),
.B(n_15882),
.Y(n_15975)
);

AND2x2_ASAP7_75t_L g15976 ( 
.A(n_15939),
.B(n_15900),
.Y(n_15976)
);

NAND2x1p5_ASAP7_75t_L g15977 ( 
.A(n_15887),
.B(n_3544),
.Y(n_15977)
);

NAND3xp33_ASAP7_75t_L g15978 ( 
.A(n_15919),
.B(n_3543),
.C(n_3544),
.Y(n_15978)
);

NAND2xp5_ASAP7_75t_L g15979 ( 
.A(n_15926),
.B(n_4270),
.Y(n_15979)
);

INVx1_ASAP7_75t_L g15980 ( 
.A(n_15878),
.Y(n_15980)
);

AND2x2_ASAP7_75t_L g15981 ( 
.A(n_15858),
.B(n_3543),
.Y(n_15981)
);

NOR3xp33_ASAP7_75t_L g15982 ( 
.A(n_15891),
.B(n_3545),
.C(n_3547),
.Y(n_15982)
);

OAI322xp33_ASAP7_75t_L g15983 ( 
.A1(n_15890),
.A2(n_3552),
.A3(n_3551),
.B1(n_3549),
.B2(n_3547),
.C1(n_3548),
.C2(n_3550),
.Y(n_15983)
);

INVx1_ASAP7_75t_L g15984 ( 
.A(n_15872),
.Y(n_15984)
);

AOI211xp5_ASAP7_75t_L g15985 ( 
.A1(n_15929),
.A2(n_3550),
.B(n_3548),
.C(n_3549),
.Y(n_15985)
);

OR2x2_ASAP7_75t_L g15986 ( 
.A(n_15940),
.B(n_3551),
.Y(n_15986)
);

AND3x4_ASAP7_75t_L g15987 ( 
.A(n_15857),
.B(n_3552),
.C(n_3553),
.Y(n_15987)
);

NAND3xp33_ASAP7_75t_L g15988 ( 
.A(n_15928),
.B(n_3553),
.C(n_3554),
.Y(n_15988)
);

NAND2xp5_ASAP7_75t_L g15989 ( 
.A(n_15906),
.B(n_4251),
.Y(n_15989)
);

XOR2x1_ASAP7_75t_L g15990 ( 
.A(n_15905),
.B(n_3554),
.Y(n_15990)
);

NAND2xp5_ASAP7_75t_L g15991 ( 
.A(n_15937),
.B(n_4254),
.Y(n_15991)
);

BUFx12f_ASAP7_75t_L g15992 ( 
.A(n_15918),
.Y(n_15992)
);

HB1xp67_ASAP7_75t_L g15993 ( 
.A(n_15925),
.Y(n_15993)
);

AO22x2_ASAP7_75t_L g15994 ( 
.A1(n_15899),
.A2(n_4256),
.B1(n_3557),
.B2(n_3555),
.Y(n_15994)
);

OAI211xp5_ASAP7_75t_SL g15995 ( 
.A1(n_15892),
.A2(n_3558),
.B(n_3555),
.C(n_3556),
.Y(n_15995)
);

OA22x2_ASAP7_75t_L g15996 ( 
.A1(n_15895),
.A2(n_3560),
.B1(n_3556),
.B2(n_3559),
.Y(n_15996)
);

NAND4xp75_ASAP7_75t_L g15997 ( 
.A(n_15930),
.B(n_3561),
.C(n_3559),
.D(n_3560),
.Y(n_15997)
);

NAND3xp33_ASAP7_75t_L g15998 ( 
.A(n_15922),
.B(n_15868),
.C(n_15913),
.Y(n_15998)
);

AND2x2_ASAP7_75t_L g15999 ( 
.A(n_15902),
.B(n_3561),
.Y(n_15999)
);

NOR3xp33_ASAP7_75t_L g16000 ( 
.A(n_15860),
.B(n_15894),
.C(n_15924),
.Y(n_16000)
);

OAI211xp5_ASAP7_75t_SL g16001 ( 
.A1(n_15910),
.A2(n_3564),
.B(n_3562),
.C(n_3563),
.Y(n_16001)
);

NAND4xp75_ASAP7_75t_L g16002 ( 
.A(n_15911),
.B(n_3564),
.C(n_3562),
.D(n_3563),
.Y(n_16002)
);

INVx1_ASAP7_75t_L g16003 ( 
.A(n_15877),
.Y(n_16003)
);

INVx2_ASAP7_75t_L g16004 ( 
.A(n_15886),
.Y(n_16004)
);

NAND2xp5_ASAP7_75t_SL g16005 ( 
.A(n_15852),
.B(n_3566),
.Y(n_16005)
);

NAND2x1p5_ASAP7_75t_L g16006 ( 
.A(n_15927),
.B(n_3567),
.Y(n_16006)
);

HB1xp67_ASAP7_75t_L g16007 ( 
.A(n_15932),
.Y(n_16007)
);

HB1xp67_ASAP7_75t_L g16008 ( 
.A(n_15904),
.Y(n_16008)
);

NOR2xp33_ASAP7_75t_L g16009 ( 
.A(n_15884),
.B(n_3566),
.Y(n_16009)
);

AOI21xp5_ASAP7_75t_L g16010 ( 
.A1(n_15866),
.A2(n_3567),
.B(n_3568),
.Y(n_16010)
);

NAND2xp5_ASAP7_75t_L g16011 ( 
.A(n_15942),
.B(n_4248),
.Y(n_16011)
);

INVx2_ASAP7_75t_L g16012 ( 
.A(n_15883),
.Y(n_16012)
);

AOI21xp5_ASAP7_75t_L g16013 ( 
.A1(n_15898),
.A2(n_3568),
.B(n_3569),
.Y(n_16013)
);

CKINVDCx6p67_ASAP7_75t_R g16014 ( 
.A(n_15874),
.Y(n_16014)
);

NAND2xp5_ASAP7_75t_L g16015 ( 
.A(n_15893),
.B(n_4250),
.Y(n_16015)
);

NAND2xp5_ASAP7_75t_L g16016 ( 
.A(n_15914),
.B(n_4251),
.Y(n_16016)
);

NAND2xp5_ASAP7_75t_L g16017 ( 
.A(n_15920),
.B(n_4257),
.Y(n_16017)
);

INVx2_ASAP7_75t_L g16018 ( 
.A(n_15876),
.Y(n_16018)
);

NAND4xp75_ASAP7_75t_L g16019 ( 
.A(n_15903),
.B(n_3572),
.C(n_3570),
.D(n_3571),
.Y(n_16019)
);

NOR2xp33_ASAP7_75t_L g16020 ( 
.A(n_15931),
.B(n_3572),
.Y(n_16020)
);

NOR2xp67_ASAP7_75t_L g16021 ( 
.A(n_15909),
.B(n_15933),
.Y(n_16021)
);

NAND4xp25_ASAP7_75t_SL g16022 ( 
.A(n_15862),
.B(n_3575),
.C(n_3573),
.D(n_3574),
.Y(n_16022)
);

NOR2xp67_ASAP7_75t_L g16023 ( 
.A(n_15921),
.B(n_3573),
.Y(n_16023)
);

INVx3_ASAP7_75t_L g16024 ( 
.A(n_15896),
.Y(n_16024)
);

NAND3xp33_ASAP7_75t_L g16025 ( 
.A(n_15881),
.B(n_3574),
.C(n_3575),
.Y(n_16025)
);

INVx1_ASAP7_75t_L g16026 ( 
.A(n_15935),
.Y(n_16026)
);

NAND2xp5_ASAP7_75t_L g16027 ( 
.A(n_15869),
.B(n_4240),
.Y(n_16027)
);

INVx1_ASAP7_75t_SL g16028 ( 
.A(n_15923),
.Y(n_16028)
);

NOR3xp33_ASAP7_75t_L g16029 ( 
.A(n_15908),
.B(n_3576),
.C(n_3577),
.Y(n_16029)
);

INVx1_ASAP7_75t_L g16030 ( 
.A(n_15855),
.Y(n_16030)
);

NOR3xp33_ASAP7_75t_L g16031 ( 
.A(n_15938),
.B(n_3577),
.C(n_3578),
.Y(n_16031)
);

NOR3x1_ASAP7_75t_L g16032 ( 
.A(n_15934),
.B(n_3578),
.C(n_3579),
.Y(n_16032)
);

INVx1_ASAP7_75t_L g16033 ( 
.A(n_15855),
.Y(n_16033)
);

AOI211xp5_ASAP7_75t_SL g16034 ( 
.A1(n_15938),
.A2(n_3582),
.B(n_3580),
.C(n_3581),
.Y(n_16034)
);

NAND4xp25_ASAP7_75t_SL g16035 ( 
.A(n_15852),
.B(n_3583),
.C(n_3581),
.D(n_3582),
.Y(n_16035)
);

NOR2x1_ASAP7_75t_L g16036 ( 
.A(n_15855),
.B(n_3584),
.Y(n_16036)
);

AND4x1_ASAP7_75t_L g16037 ( 
.A(n_15875),
.B(n_3587),
.C(n_3585),
.D(n_3586),
.Y(n_16037)
);

NAND3xp33_ASAP7_75t_SL g16038 ( 
.A(n_15853),
.B(n_3595),
.C(n_3585),
.Y(n_16038)
);

INVx1_ASAP7_75t_L g16039 ( 
.A(n_15855),
.Y(n_16039)
);

AND5x1_ASAP7_75t_L g16040 ( 
.A(n_15921),
.B(n_3589),
.C(n_3587),
.D(n_3588),
.E(n_3590),
.Y(n_16040)
);

NOR3xp33_ASAP7_75t_L g16041 ( 
.A(n_15938),
.B(n_3588),
.C(n_3589),
.Y(n_16041)
);

NAND2xp5_ASAP7_75t_L g16042 ( 
.A(n_15870),
.B(n_3591),
.Y(n_16042)
);

NAND2xp5_ASAP7_75t_SL g16043 ( 
.A(n_15972),
.B(n_3591),
.Y(n_16043)
);

AOI211xp5_ASAP7_75t_L g16044 ( 
.A1(n_15995),
.A2(n_3595),
.B(n_3593),
.C(n_3594),
.Y(n_16044)
);

NOR2x1_ASAP7_75t_L g16045 ( 
.A(n_15966),
.B(n_3596),
.Y(n_16045)
);

OAI211xp5_ASAP7_75t_SL g16046 ( 
.A1(n_15957),
.A2(n_3597),
.B(n_3594),
.C(n_3596),
.Y(n_16046)
);

INVx1_ASAP7_75t_L g16047 ( 
.A(n_15990),
.Y(n_16047)
);

AO22x2_ASAP7_75t_L g16048 ( 
.A1(n_15947),
.A2(n_3599),
.B1(n_3600),
.B2(n_3598),
.Y(n_16048)
);

NOR3xp33_ASAP7_75t_L g16049 ( 
.A(n_16024),
.B(n_3597),
.C(n_3598),
.Y(n_16049)
);

NAND3x1_ASAP7_75t_SL g16050 ( 
.A(n_16036),
.B(n_3601),
.C(n_3600),
.Y(n_16050)
);

INVxp33_ASAP7_75t_SL g16051 ( 
.A(n_15960),
.Y(n_16051)
);

NAND2xp5_ASAP7_75t_L g16052 ( 
.A(n_16034),
.B(n_3601),
.Y(n_16052)
);

NOR2x1_ASAP7_75t_L g16053 ( 
.A(n_16030),
.B(n_3602),
.Y(n_16053)
);

NOR4xp25_ASAP7_75t_L g16054 ( 
.A(n_16028),
.B(n_4248),
.C(n_3603),
.D(n_3599),
.Y(n_16054)
);

AND4x1_ASAP7_75t_L g16055 ( 
.A(n_16000),
.B(n_3605),
.C(n_3602),
.D(n_3604),
.Y(n_16055)
);

NOR3xp33_ASAP7_75t_L g16056 ( 
.A(n_16024),
.B(n_16012),
.C(n_16039),
.Y(n_16056)
);

NAND4xp75_ASAP7_75t_L g16057 ( 
.A(n_16021),
.B(n_3606),
.C(n_3604),
.D(n_3605),
.Y(n_16057)
);

NOR3x1_ASAP7_75t_L g16058 ( 
.A(n_15997),
.B(n_3606),
.C(n_3607),
.Y(n_16058)
);

NOR3xp33_ASAP7_75t_L g16059 ( 
.A(n_16033),
.B(n_3608),
.C(n_3609),
.Y(n_16059)
);

INVx1_ASAP7_75t_L g16060 ( 
.A(n_16042),
.Y(n_16060)
);

INVxp33_ASAP7_75t_L g16061 ( 
.A(n_15987),
.Y(n_16061)
);

NOR3xp33_ASAP7_75t_SL g16062 ( 
.A(n_15955),
.B(n_3608),
.C(n_3609),
.Y(n_16062)
);

INVx2_ASAP7_75t_L g16063 ( 
.A(n_15994),
.Y(n_16063)
);

NOR3xp33_ASAP7_75t_L g16064 ( 
.A(n_15961),
.B(n_3610),
.C(n_3611),
.Y(n_16064)
);

NAND4xp25_ASAP7_75t_L g16065 ( 
.A(n_16032),
.B(n_15963),
.C(n_15949),
.D(n_15985),
.Y(n_16065)
);

AOI211xp5_ASAP7_75t_L g16066 ( 
.A1(n_16035),
.A2(n_16038),
.B(n_16001),
.C(n_15953),
.Y(n_16066)
);

NOR3xp33_ASAP7_75t_L g16067 ( 
.A(n_16004),
.B(n_3610),
.C(n_3611),
.Y(n_16067)
);

NAND4xp25_ASAP7_75t_L g16068 ( 
.A(n_15954),
.B(n_3614),
.C(n_3612),
.D(n_3613),
.Y(n_16068)
);

AOI211xp5_ASAP7_75t_L g16069 ( 
.A1(n_15978),
.A2(n_15988),
.B(n_15946),
.C(n_16009),
.Y(n_16069)
);

NOR2x1_ASAP7_75t_L g16070 ( 
.A(n_16002),
.B(n_3614),
.Y(n_16070)
);

HB1xp67_ASAP7_75t_L g16071 ( 
.A(n_16037),
.Y(n_16071)
);

NOR2x1_ASAP7_75t_L g16072 ( 
.A(n_16019),
.B(n_3615),
.Y(n_16072)
);

NAND4xp75_ASAP7_75t_L g16073 ( 
.A(n_16023),
.B(n_3617),
.C(n_3612),
.D(n_3616),
.Y(n_16073)
);

AND2x2_ASAP7_75t_L g16074 ( 
.A(n_15965),
.B(n_3616),
.Y(n_16074)
);

NAND4xp25_ASAP7_75t_L g16075 ( 
.A(n_15952),
.B(n_3620),
.C(n_3618),
.D(n_3619),
.Y(n_16075)
);

NAND4xp75_ASAP7_75t_L g16076 ( 
.A(n_15976),
.B(n_3621),
.C(n_3618),
.D(n_3619),
.Y(n_16076)
);

NOR3xp33_ASAP7_75t_L g16077 ( 
.A(n_15962),
.B(n_3621),
.C(n_3622),
.Y(n_16077)
);

NOR2x1_ASAP7_75t_L g16078 ( 
.A(n_16022),
.B(n_3623),
.Y(n_16078)
);

AND2x4_ASAP7_75t_L g16079 ( 
.A(n_16040),
.B(n_3622),
.Y(n_16079)
);

INVx1_ASAP7_75t_L g16080 ( 
.A(n_16006),
.Y(n_16080)
);

OAI211xp5_ASAP7_75t_L g16081 ( 
.A1(n_15950),
.A2(n_3626),
.B(n_3627),
.C(n_3625),
.Y(n_16081)
);

NOR2x1_ASAP7_75t_L g16082 ( 
.A(n_15971),
.B(n_3625),
.Y(n_16082)
);

NOR2x1_ASAP7_75t_L g16083 ( 
.A(n_16025),
.B(n_15983),
.Y(n_16083)
);

AND2x2_ASAP7_75t_L g16084 ( 
.A(n_15999),
.B(n_3624),
.Y(n_16084)
);

OAI211xp5_ASAP7_75t_L g16085 ( 
.A1(n_16010),
.A2(n_3627),
.B(n_3628),
.C(n_3626),
.Y(n_16085)
);

NAND2xp33_ASAP7_75t_SL g16086 ( 
.A(n_15970),
.B(n_3624),
.Y(n_16086)
);

NOR3xp33_ASAP7_75t_L g16087 ( 
.A(n_15984),
.B(n_3629),
.C(n_3630),
.Y(n_16087)
);

NAND4xp75_ASAP7_75t_L g16088 ( 
.A(n_16026),
.B(n_3632),
.C(n_3630),
.D(n_3631),
.Y(n_16088)
);

XNOR2x1_ASAP7_75t_L g16089 ( 
.A(n_15986),
.B(n_4245),
.Y(n_16089)
);

OR2x2_ASAP7_75t_L g16090 ( 
.A(n_16015),
.B(n_3631),
.Y(n_16090)
);

AOI21xp5_ASAP7_75t_L g16091 ( 
.A1(n_15951),
.A2(n_3632),
.B(n_3633),
.Y(n_16091)
);

NOR3xp33_ASAP7_75t_L g16092 ( 
.A(n_15998),
.B(n_3633),
.C(n_3634),
.Y(n_16092)
);

NOR2xp33_ASAP7_75t_L g16093 ( 
.A(n_15992),
.B(n_4259),
.Y(n_16093)
);

INVx1_ASAP7_75t_L g16094 ( 
.A(n_15977),
.Y(n_16094)
);

NOR3xp33_ASAP7_75t_L g16095 ( 
.A(n_15958),
.B(n_3634),
.C(n_3635),
.Y(n_16095)
);

INVx2_ASAP7_75t_SL g16096 ( 
.A(n_15948),
.Y(n_16096)
);

NOR2xp33_ASAP7_75t_SL g16097 ( 
.A(n_15993),
.B(n_3635),
.Y(n_16097)
);

AOI21xp5_ASAP7_75t_SL g16098 ( 
.A1(n_16007),
.A2(n_3638),
.B(n_3637),
.Y(n_16098)
);

AND4x1_ASAP7_75t_L g16099 ( 
.A(n_15969),
.B(n_3640),
.C(n_3636),
.D(n_3639),
.Y(n_16099)
);

NAND2xp5_ASAP7_75t_SL g16100 ( 
.A(n_16031),
.B(n_3639),
.Y(n_16100)
);

NOR3x1_ASAP7_75t_L g16101 ( 
.A(n_16016),
.B(n_3641),
.C(n_3642),
.Y(n_16101)
);

NAND4xp75_ASAP7_75t_L g16102 ( 
.A(n_16013),
.B(n_3644),
.C(n_3641),
.D(n_3643),
.Y(n_16102)
);

NAND4xp25_ASAP7_75t_L g16103 ( 
.A(n_15967),
.B(n_3645),
.C(n_3643),
.D(n_3644),
.Y(n_16103)
);

NOR2x1_ASAP7_75t_L g16104 ( 
.A(n_15974),
.B(n_3646),
.Y(n_16104)
);

NAND3xp33_ASAP7_75t_L g16105 ( 
.A(n_16041),
.B(n_3645),
.C(n_3646),
.Y(n_16105)
);

NAND3xp33_ASAP7_75t_L g16106 ( 
.A(n_15982),
.B(n_3647),
.C(n_3648),
.Y(n_16106)
);

NAND3xp33_ASAP7_75t_L g16107 ( 
.A(n_16020),
.B(n_3647),
.C(n_3648),
.Y(n_16107)
);

NOR3xp33_ASAP7_75t_L g16108 ( 
.A(n_15973),
.B(n_3649),
.C(n_3651),
.Y(n_16108)
);

INVx1_ASAP7_75t_L g16109 ( 
.A(n_15996),
.Y(n_16109)
);

NAND2xp5_ASAP7_75t_L g16110 ( 
.A(n_16029),
.B(n_3652),
.Y(n_16110)
);

NOR2x1_ASAP7_75t_L g16111 ( 
.A(n_15980),
.B(n_3652),
.Y(n_16111)
);

NAND2xp5_ASAP7_75t_L g16112 ( 
.A(n_15981),
.B(n_3653),
.Y(n_16112)
);

AND2x4_ASAP7_75t_L g16113 ( 
.A(n_16011),
.B(n_15956),
.Y(n_16113)
);

NOR3xp33_ASAP7_75t_L g16114 ( 
.A(n_16008),
.B(n_3649),
.C(n_3654),
.Y(n_16114)
);

NOR2x1_ASAP7_75t_L g16115 ( 
.A(n_16027),
.B(n_3655),
.Y(n_16115)
);

NAND2x1p5_ASAP7_75t_L g16116 ( 
.A(n_15968),
.B(n_3654),
.Y(n_16116)
);

INVx1_ASAP7_75t_SL g16117 ( 
.A(n_15964),
.Y(n_16117)
);

INVx1_ASAP7_75t_L g16118 ( 
.A(n_15959),
.Y(n_16118)
);

NAND3xp33_ASAP7_75t_L g16119 ( 
.A(n_15979),
.B(n_3655),
.C(n_3656),
.Y(n_16119)
);

NAND4xp75_ASAP7_75t_L g16120 ( 
.A(n_16003),
.B(n_3658),
.C(n_3656),
.D(n_3657),
.Y(n_16120)
);

NOR3x1_ASAP7_75t_L g16121 ( 
.A(n_15991),
.B(n_3658),
.C(n_3659),
.Y(n_16121)
);

NAND3xp33_ASAP7_75t_SL g16122 ( 
.A(n_15989),
.B(n_15975),
.C(n_16017),
.Y(n_16122)
);

NOR2xp67_ASAP7_75t_L g16123 ( 
.A(n_16005),
.B(n_3660),
.Y(n_16123)
);

NOR2x1_ASAP7_75t_L g16124 ( 
.A(n_16018),
.B(n_3660),
.Y(n_16124)
);

NOR3xp33_ASAP7_75t_L g16125 ( 
.A(n_16014),
.B(n_3659),
.C(n_3661),
.Y(n_16125)
);

NAND4xp25_ASAP7_75t_L g16126 ( 
.A(n_15994),
.B(n_3663),
.C(n_3661),
.D(n_3662),
.Y(n_16126)
);

NAND3xp33_ASAP7_75t_L g16127 ( 
.A(n_15972),
.B(n_3662),
.C(n_3663),
.Y(n_16127)
);

NAND4xp25_ASAP7_75t_L g16128 ( 
.A(n_15960),
.B(n_3666),
.C(n_3664),
.D(n_3665),
.Y(n_16128)
);

AOI22xp5_ASAP7_75t_L g16129 ( 
.A1(n_15960),
.A2(n_3666),
.B1(n_3664),
.B2(n_3665),
.Y(n_16129)
);

NOR2xp33_ASAP7_75t_L g16130 ( 
.A(n_15995),
.B(n_4261),
.Y(n_16130)
);

NAND4xp25_ASAP7_75t_L g16131 ( 
.A(n_15960),
.B(n_3669),
.C(n_3667),
.D(n_3668),
.Y(n_16131)
);

OAI211xp5_ASAP7_75t_L g16132 ( 
.A1(n_16042),
.A2(n_3670),
.B(n_3671),
.C(n_3668),
.Y(n_16132)
);

NAND2xp5_ASAP7_75t_L g16133 ( 
.A(n_16034),
.B(n_3670),
.Y(n_16133)
);

NOR2xp33_ASAP7_75t_L g16134 ( 
.A(n_15995),
.B(n_3667),
.Y(n_16134)
);

NAND3xp33_ASAP7_75t_L g16135 ( 
.A(n_15972),
.B(n_3671),
.C(n_3672),
.Y(n_16135)
);

AND4x1_ASAP7_75t_L g16136 ( 
.A(n_15960),
.B(n_3675),
.C(n_3673),
.D(n_3674),
.Y(n_16136)
);

NAND3xp33_ASAP7_75t_L g16137 ( 
.A(n_15972),
.B(n_3673),
.C(n_3674),
.Y(n_16137)
);

INVx2_ASAP7_75t_L g16138 ( 
.A(n_15994),
.Y(n_16138)
);

NOR2x1_ASAP7_75t_L g16139 ( 
.A(n_15966),
.B(n_3676),
.Y(n_16139)
);

INVx1_ASAP7_75t_L g16140 ( 
.A(n_15990),
.Y(n_16140)
);

NOR4xp25_ASAP7_75t_L g16141 ( 
.A(n_15957),
.B(n_4265),
.C(n_4241),
.D(n_3677),
.Y(n_16141)
);

INVx1_ASAP7_75t_L g16142 ( 
.A(n_15990),
.Y(n_16142)
);

NOR2xp33_ASAP7_75t_L g16143 ( 
.A(n_15995),
.B(n_4242),
.Y(n_16143)
);

OAI211xp5_ASAP7_75t_L g16144 ( 
.A1(n_16042),
.A2(n_3677),
.B(n_3678),
.C(n_3676),
.Y(n_16144)
);

NAND4xp25_ASAP7_75t_L g16145 ( 
.A(n_15960),
.B(n_3679),
.C(n_3675),
.D(n_3678),
.Y(n_16145)
);

NAND2xp5_ASAP7_75t_SL g16146 ( 
.A(n_15972),
.B(n_3679),
.Y(n_16146)
);

NAND2xp5_ASAP7_75t_L g16147 ( 
.A(n_16034),
.B(n_3681),
.Y(n_16147)
);

NAND3x1_ASAP7_75t_L g16148 ( 
.A(n_16036),
.B(n_3680),
.C(n_3682),
.Y(n_16148)
);

NOR2x1_ASAP7_75t_L g16149 ( 
.A(n_15966),
.B(n_3682),
.Y(n_16149)
);

NOR2x1_ASAP7_75t_L g16150 ( 
.A(n_15966),
.B(n_3683),
.Y(n_16150)
);

NAND3xp33_ASAP7_75t_L g16151 ( 
.A(n_15972),
.B(n_3680),
.C(n_3683),
.Y(n_16151)
);

NOR3xp33_ASAP7_75t_L g16152 ( 
.A(n_15972),
.B(n_3684),
.C(n_3685),
.Y(n_16152)
);

NAND4xp75_ASAP7_75t_L g16153 ( 
.A(n_15966),
.B(n_3686),
.C(n_3684),
.D(n_3685),
.Y(n_16153)
);

NAND2xp5_ASAP7_75t_L g16154 ( 
.A(n_16034),
.B(n_3688),
.Y(n_16154)
);

AND2x2_ASAP7_75t_L g16155 ( 
.A(n_15965),
.B(n_3687),
.Y(n_16155)
);

NOR2x1_ASAP7_75t_SL g16156 ( 
.A(n_15955),
.B(n_3688),
.Y(n_16156)
);

NAND2xp5_ASAP7_75t_L g16157 ( 
.A(n_16034),
.B(n_3689),
.Y(n_16157)
);

NOR2x1_ASAP7_75t_L g16158 ( 
.A(n_15966),
.B(n_3689),
.Y(n_16158)
);

INVx1_ASAP7_75t_L g16159 ( 
.A(n_15990),
.Y(n_16159)
);

NAND3xp33_ASAP7_75t_L g16160 ( 
.A(n_15972),
.B(n_3687),
.C(n_3691),
.Y(n_16160)
);

NAND2xp5_ASAP7_75t_L g16161 ( 
.A(n_16034),
.B(n_3693),
.Y(n_16161)
);

NOR2xp33_ASAP7_75t_L g16162 ( 
.A(n_15995),
.B(n_4242),
.Y(n_16162)
);

NAND3xp33_ASAP7_75t_L g16163 ( 
.A(n_16097),
.B(n_3692),
.C(n_3693),
.Y(n_16163)
);

OAI211xp5_ASAP7_75t_L g16164 ( 
.A1(n_16043),
.A2(n_3695),
.B(n_3696),
.C(n_3694),
.Y(n_16164)
);

OAI211xp5_ASAP7_75t_L g16165 ( 
.A1(n_16146),
.A2(n_3696),
.B(n_3697),
.C(n_3694),
.Y(n_16165)
);

AOI221x1_ASAP7_75t_L g16166 ( 
.A1(n_16056),
.A2(n_3699),
.B1(n_3692),
.B2(n_3698),
.C(n_3700),
.Y(n_16166)
);

OAI21x1_ASAP7_75t_L g16167 ( 
.A1(n_16148),
.A2(n_4273),
.B(n_4272),
.Y(n_16167)
);

AOI22xp5_ASAP7_75t_L g16168 ( 
.A1(n_16051),
.A2(n_3700),
.B1(n_3698),
.B2(n_3699),
.Y(n_16168)
);

AOI221xp5_ASAP7_75t_L g16169 ( 
.A1(n_16086),
.A2(n_16134),
.B1(n_16162),
.B2(n_16143),
.C(n_16130),
.Y(n_16169)
);

AOI211xp5_ASAP7_75t_L g16170 ( 
.A1(n_16127),
.A2(n_3703),
.B(n_3701),
.C(n_3702),
.Y(n_16170)
);

AOI21xp5_ASAP7_75t_L g16171 ( 
.A1(n_16052),
.A2(n_3702),
.B(n_3703),
.Y(n_16171)
);

AOI22xp33_ASAP7_75t_L g16172 ( 
.A1(n_16079),
.A2(n_3706),
.B1(n_3704),
.B2(n_3705),
.Y(n_16172)
);

OAI211xp5_ASAP7_75t_L g16173 ( 
.A1(n_16098),
.A2(n_3708),
.B(n_3709),
.C(n_3705),
.Y(n_16173)
);

XOR2xp5_ASAP7_75t_L g16174 ( 
.A(n_16089),
.B(n_3704),
.Y(n_16174)
);

OAI21xp5_ASAP7_75t_L g16175 ( 
.A1(n_16091),
.A2(n_3708),
.B(n_3709),
.Y(n_16175)
);

NAND3xp33_ASAP7_75t_L g16176 ( 
.A(n_16152),
.B(n_3710),
.C(n_3712),
.Y(n_16176)
);

XNOR2x1_ASAP7_75t_L g16177 ( 
.A(n_16073),
.B(n_4244),
.Y(n_16177)
);

AOI22xp5_ASAP7_75t_L g16178 ( 
.A1(n_16079),
.A2(n_3713),
.B1(n_3710),
.B2(n_3712),
.Y(n_16178)
);

NAND2xp5_ASAP7_75t_L g16179 ( 
.A(n_16093),
.B(n_16155),
.Y(n_16179)
);

AOI321xp33_ASAP7_75t_L g16180 ( 
.A1(n_16066),
.A2(n_3716),
.A3(n_3718),
.B1(n_3714),
.B2(n_3715),
.C(n_3717),
.Y(n_16180)
);

OAI222xp33_ASAP7_75t_L g16181 ( 
.A1(n_16082),
.A2(n_3717),
.B1(n_3720),
.B2(n_3714),
.C1(n_3715),
.C2(n_3719),
.Y(n_16181)
);

NAND2xp5_ASAP7_75t_SL g16182 ( 
.A(n_16141),
.B(n_16054),
.Y(n_16182)
);

INVx2_ASAP7_75t_SL g16183 ( 
.A(n_16045),
.Y(n_16183)
);

A2O1A1Ixp33_ASAP7_75t_SL g16184 ( 
.A1(n_16047),
.A2(n_4238),
.B(n_4239),
.C(n_4237),
.Y(n_16184)
);

NAND2xp5_ASAP7_75t_L g16185 ( 
.A(n_16074),
.B(n_3721),
.Y(n_16185)
);

CKINVDCx20_ASAP7_75t_R g16186 ( 
.A(n_16071),
.Y(n_16186)
);

AO22x1_ASAP7_75t_L g16187 ( 
.A1(n_16139),
.A2(n_3723),
.B1(n_3721),
.B2(n_3722),
.Y(n_16187)
);

OAI31xp33_ASAP7_75t_L g16188 ( 
.A1(n_16085),
.A2(n_16046),
.A3(n_16105),
.B(n_16106),
.Y(n_16188)
);

OAI31xp33_ASAP7_75t_L g16189 ( 
.A1(n_16135),
.A2(n_3724),
.A3(n_3722),
.B(n_3723),
.Y(n_16189)
);

NAND4xp25_ASAP7_75t_L g16190 ( 
.A(n_16058),
.B(n_4272),
.C(n_4239),
.D(n_3726),
.Y(n_16190)
);

INVx1_ASAP7_75t_SL g16191 ( 
.A(n_16084),
.Y(n_16191)
);

OAI22xp5_ASAP7_75t_L g16192 ( 
.A1(n_16137),
.A2(n_3726),
.B1(n_3724),
.B2(n_3725),
.Y(n_16192)
);

INVx1_ASAP7_75t_L g16193 ( 
.A(n_16053),
.Y(n_16193)
);

AOI22xp5_ASAP7_75t_L g16194 ( 
.A1(n_16096),
.A2(n_16095),
.B1(n_16109),
.B2(n_16092),
.Y(n_16194)
);

NOR3xp33_ASAP7_75t_L g16195 ( 
.A(n_16122),
.B(n_3725),
.C(n_3727),
.Y(n_16195)
);

AOI22xp5_ASAP7_75t_L g16196 ( 
.A1(n_16151),
.A2(n_3729),
.B1(n_3727),
.B2(n_3728),
.Y(n_16196)
);

OAI21xp5_ASAP7_75t_L g16197 ( 
.A1(n_16133),
.A2(n_3728),
.B(n_3729),
.Y(n_16197)
);

OAI31xp33_ASAP7_75t_L g16198 ( 
.A1(n_16160),
.A2(n_3732),
.A3(n_3730),
.B(n_3731),
.Y(n_16198)
);

OAI21xp5_ASAP7_75t_SL g16199 ( 
.A1(n_16107),
.A2(n_3730),
.B(n_3731),
.Y(n_16199)
);

NAND3xp33_ASAP7_75t_SL g16200 ( 
.A(n_16112),
.B(n_3732),
.C(n_3733),
.Y(n_16200)
);

INVx1_ASAP7_75t_L g16201 ( 
.A(n_16104),
.Y(n_16201)
);

INVx2_ASAP7_75t_L g16202 ( 
.A(n_16048),
.Y(n_16202)
);

O2A1O1Ixp33_ASAP7_75t_L g16203 ( 
.A1(n_16063),
.A2(n_3742),
.B(n_3750),
.C(n_3733),
.Y(n_16203)
);

OAI211xp5_ASAP7_75t_SL g16204 ( 
.A1(n_16069),
.A2(n_3736),
.B(n_3734),
.C(n_3735),
.Y(n_16204)
);

AOI21xp33_ASAP7_75t_SL g16205 ( 
.A1(n_16116),
.A2(n_3734),
.B(n_3735),
.Y(n_16205)
);

AOI221xp5_ASAP7_75t_L g16206 ( 
.A1(n_16140),
.A2(n_3739),
.B1(n_3736),
.B2(n_3738),
.C(n_3740),
.Y(n_16206)
);

HB1xp67_ASAP7_75t_L g16207 ( 
.A(n_16136),
.Y(n_16207)
);

OAI22xp5_ASAP7_75t_L g16208 ( 
.A1(n_16119),
.A2(n_3743),
.B1(n_3740),
.B2(n_3741),
.Y(n_16208)
);

AOI211x1_ASAP7_75t_SL g16209 ( 
.A1(n_16123),
.A2(n_3745),
.B(n_3743),
.C(n_3744),
.Y(n_16209)
);

NOR3xp33_ASAP7_75t_L g16210 ( 
.A(n_16142),
.B(n_3744),
.C(n_3745),
.Y(n_16210)
);

AOI21xp5_ASAP7_75t_L g16211 ( 
.A1(n_16147),
.A2(n_3746),
.B(n_3747),
.Y(n_16211)
);

AOI22xp5_ASAP7_75t_L g16212 ( 
.A1(n_16068),
.A2(n_3748),
.B1(n_3746),
.B2(n_3747),
.Y(n_16212)
);

OAI211xp5_ASAP7_75t_SL g16213 ( 
.A1(n_16159),
.A2(n_3750),
.B(n_3748),
.C(n_3749),
.Y(n_16213)
);

AOI222xp33_ASAP7_75t_L g16214 ( 
.A1(n_16100),
.A2(n_3752),
.B1(n_3754),
.B2(n_3749),
.C1(n_3751),
.C2(n_3753),
.Y(n_16214)
);

NOR2xp33_ASAP7_75t_R g16215 ( 
.A(n_16080),
.B(n_3752),
.Y(n_16215)
);

AOI221xp5_ASAP7_75t_L g16216 ( 
.A1(n_16154),
.A2(n_3754),
.B1(n_3751),
.B2(n_3753),
.C(n_3755),
.Y(n_16216)
);

AOI211xp5_ASAP7_75t_L g16217 ( 
.A1(n_16081),
.A2(n_3757),
.B(n_3755),
.C(n_3756),
.Y(n_16217)
);

HB1xp67_ASAP7_75t_L g16218 ( 
.A(n_16111),
.Y(n_16218)
);

AOI221xp5_ASAP7_75t_L g16219 ( 
.A1(n_16157),
.A2(n_3759),
.B1(n_3757),
.B2(n_3758),
.C(n_3760),
.Y(n_16219)
);

NAND3x1_ASAP7_75t_SL g16220 ( 
.A(n_16149),
.B(n_16158),
.C(n_16150),
.Y(n_16220)
);

NAND3xp33_ASAP7_75t_SL g16221 ( 
.A(n_16099),
.B(n_3758),
.C(n_3759),
.Y(n_16221)
);

OAI321xp33_ASAP7_75t_L g16222 ( 
.A1(n_16161),
.A2(n_3763),
.A3(n_3765),
.B1(n_3760),
.B2(n_3762),
.C(n_3764),
.Y(n_16222)
);

AOI221xp5_ASAP7_75t_L g16223 ( 
.A1(n_16044),
.A2(n_3767),
.B1(n_3763),
.B2(n_3766),
.C(n_3768),
.Y(n_16223)
);

NOR2xp33_ASAP7_75t_SL g16224 ( 
.A(n_16065),
.B(n_3766),
.Y(n_16224)
);

AOI21xp33_ASAP7_75t_L g16225 ( 
.A1(n_16061),
.A2(n_16110),
.B(n_16094),
.Y(n_16225)
);

AOI221xp5_ASAP7_75t_L g16226 ( 
.A1(n_16138),
.A2(n_3770),
.B1(n_3768),
.B2(n_3769),
.C(n_3771),
.Y(n_16226)
);

BUFx6f_ASAP7_75t_L g16227 ( 
.A(n_16113),
.Y(n_16227)
);

OAI311xp33_ASAP7_75t_L g16228 ( 
.A1(n_16118),
.A2(n_3771),
.A3(n_3769),
.B1(n_3770),
.C1(n_3772),
.Y(n_16228)
);

NAND2xp5_ASAP7_75t_L g16229 ( 
.A(n_16125),
.B(n_3772),
.Y(n_16229)
);

AOI211xp5_ASAP7_75t_L g16230 ( 
.A1(n_16126),
.A2(n_3775),
.B(n_3773),
.C(n_3774),
.Y(n_16230)
);

INVx1_ASAP7_75t_L g16231 ( 
.A(n_16124),
.Y(n_16231)
);

AOI21xp5_ASAP7_75t_L g16232 ( 
.A1(n_16156),
.A2(n_3774),
.B(n_3776),
.Y(n_16232)
);

AND2x2_ASAP7_75t_L g16233 ( 
.A(n_16062),
.B(n_3776),
.Y(n_16233)
);

NOR4xp25_ASAP7_75t_L g16234 ( 
.A(n_16117),
.B(n_3779),
.C(n_3777),
.D(n_3778),
.Y(n_16234)
);

AOI22xp5_ASAP7_75t_L g16235 ( 
.A1(n_16102),
.A2(n_3779),
.B1(n_3777),
.B2(n_3778),
.Y(n_16235)
);

NOR2xp67_ASAP7_75t_L g16236 ( 
.A(n_16075),
.B(n_3781),
.Y(n_16236)
);

OAI22xp5_ASAP7_75t_L g16237 ( 
.A1(n_16090),
.A2(n_3782),
.B1(n_3780),
.B2(n_3781),
.Y(n_16237)
);

OAI221xp5_ASAP7_75t_SL g16238 ( 
.A1(n_16060),
.A2(n_3783),
.B1(n_3780),
.B2(n_3782),
.C(n_3784),
.Y(n_16238)
);

AOI321xp33_ASAP7_75t_L g16239 ( 
.A1(n_16078),
.A2(n_3785),
.A3(n_3787),
.B1(n_3783),
.B2(n_3784),
.C(n_3786),
.Y(n_16239)
);

NOR2x1_ASAP7_75t_L g16240 ( 
.A(n_16153),
.B(n_16057),
.Y(n_16240)
);

OA22x2_ASAP7_75t_L g16241 ( 
.A1(n_16132),
.A2(n_3787),
.B1(n_3785),
.B2(n_3786),
.Y(n_16241)
);

OAI21xp5_ASAP7_75t_L g16242 ( 
.A1(n_16070),
.A2(n_3788),
.B(n_3789),
.Y(n_16242)
);

NOR4xp25_ASAP7_75t_L g16243 ( 
.A(n_16103),
.B(n_3791),
.C(n_3789),
.D(n_3790),
.Y(n_16243)
);

NOR2x1_ASAP7_75t_L g16244 ( 
.A(n_16076),
.B(n_4244),
.Y(n_16244)
);

AOI21xp33_ASAP7_75t_L g16245 ( 
.A1(n_16083),
.A2(n_3790),
.B(n_3792),
.Y(n_16245)
);

AOI221xp5_ASAP7_75t_L g16246 ( 
.A1(n_16113),
.A2(n_3794),
.B1(n_3792),
.B2(n_3793),
.C(n_3795),
.Y(n_16246)
);

AOI222xp33_ASAP7_75t_L g16247 ( 
.A1(n_16072),
.A2(n_3795),
.B1(n_3798),
.B2(n_3793),
.C1(n_3794),
.C2(n_3797),
.Y(n_16247)
);

NOR3xp33_ASAP7_75t_L g16248 ( 
.A(n_16220),
.B(n_16050),
.C(n_16115),
.Y(n_16248)
);

INVx1_ASAP7_75t_L g16249 ( 
.A(n_16167),
.Y(n_16249)
);

NAND3xp33_ASAP7_75t_SL g16250 ( 
.A(n_16186),
.B(n_16055),
.C(n_16067),
.Y(n_16250)
);

INVxp67_ASAP7_75t_L g16251 ( 
.A(n_16224),
.Y(n_16251)
);

NOR2xp33_ASAP7_75t_SL g16252 ( 
.A(n_16191),
.B(n_16120),
.Y(n_16252)
);

INVx1_ASAP7_75t_L g16253 ( 
.A(n_16241),
.Y(n_16253)
);

OAI21xp5_ASAP7_75t_SL g16254 ( 
.A1(n_16209),
.A2(n_16144),
.B(n_16087),
.Y(n_16254)
);

NAND3xp33_ASAP7_75t_L g16255 ( 
.A(n_16247),
.B(n_16077),
.C(n_16114),
.Y(n_16255)
);

NOR3x2_ASAP7_75t_L g16256 ( 
.A(n_16183),
.B(n_16088),
.C(n_16218),
.Y(n_16256)
);

NAND3x2_ASAP7_75t_L g16257 ( 
.A(n_16233),
.B(n_16121),
.C(n_16101),
.Y(n_16257)
);

NOR2x1_ASAP7_75t_L g16258 ( 
.A(n_16202),
.B(n_16128),
.Y(n_16258)
);

INVx2_ASAP7_75t_SL g16259 ( 
.A(n_16177),
.Y(n_16259)
);

AND2x4_ASAP7_75t_L g16260 ( 
.A(n_16240),
.B(n_16064),
.Y(n_16260)
);

AOI21xp5_ASAP7_75t_SL g16261 ( 
.A1(n_16182),
.A2(n_16129),
.B(n_16131),
.Y(n_16261)
);

NOR2xp67_ASAP7_75t_L g16262 ( 
.A(n_16190),
.B(n_16145),
.Y(n_16262)
);

AND2x4_ASAP7_75t_L g16263 ( 
.A(n_16244),
.B(n_16108),
.Y(n_16263)
);

NAND2xp5_ASAP7_75t_SL g16264 ( 
.A(n_16239),
.B(n_16059),
.Y(n_16264)
);

NOR3x2_ASAP7_75t_L g16265 ( 
.A(n_16187),
.B(n_16049),
.C(n_16048),
.Y(n_16265)
);

NOR2x1_ASAP7_75t_L g16266 ( 
.A(n_16201),
.B(n_3797),
.Y(n_16266)
);

NOR2x1p5_ASAP7_75t_L g16267 ( 
.A(n_16221),
.B(n_3798),
.Y(n_16267)
);

OAI22xp5_ASAP7_75t_L g16268 ( 
.A1(n_16172),
.A2(n_3801),
.B1(n_3799),
.B2(n_3800),
.Y(n_16268)
);

NOR3xp33_ASAP7_75t_L g16269 ( 
.A(n_16225),
.B(n_3799),
.C(n_3800),
.Y(n_16269)
);

NOR3xp33_ASAP7_75t_L g16270 ( 
.A(n_16231),
.B(n_3801),
.C(n_3802),
.Y(n_16270)
);

NOR3xp33_ASAP7_75t_L g16271 ( 
.A(n_16193),
.B(n_3802),
.C(n_3803),
.Y(n_16271)
);

INVx1_ASAP7_75t_L g16272 ( 
.A(n_16174),
.Y(n_16272)
);

NAND2xp5_ASAP7_75t_L g16273 ( 
.A(n_16178),
.B(n_3803),
.Y(n_16273)
);

NOR2x1p5_ASAP7_75t_L g16274 ( 
.A(n_16229),
.B(n_3804),
.Y(n_16274)
);

INVxp33_ASAP7_75t_L g16275 ( 
.A(n_16215),
.Y(n_16275)
);

INVx2_ASAP7_75t_SL g16276 ( 
.A(n_16185),
.Y(n_16276)
);

NOR3xp33_ASAP7_75t_L g16277 ( 
.A(n_16179),
.B(n_3804),
.C(n_3805),
.Y(n_16277)
);

NOR2x1p5_ASAP7_75t_L g16278 ( 
.A(n_16200),
.B(n_3805),
.Y(n_16278)
);

NOR2x1_ASAP7_75t_SL g16279 ( 
.A(n_16173),
.B(n_3806),
.Y(n_16279)
);

NAND2x1p5_ASAP7_75t_L g16280 ( 
.A(n_16227),
.B(n_16194),
.Y(n_16280)
);

NOR2x1_ASAP7_75t_L g16281 ( 
.A(n_16163),
.B(n_16181),
.Y(n_16281)
);

NAND3x2_ASAP7_75t_L g16282 ( 
.A(n_16189),
.B(n_4240),
.C(n_3807),
.Y(n_16282)
);

NOR2x1_ASAP7_75t_L g16283 ( 
.A(n_16242),
.B(n_3808),
.Y(n_16283)
);

XNOR2xp5_ASAP7_75t_L g16284 ( 
.A(n_16243),
.B(n_3809),
.Y(n_16284)
);

OR2x2_ASAP7_75t_L g16285 ( 
.A(n_16234),
.B(n_3809),
.Y(n_16285)
);

NAND2x1p5_ASAP7_75t_L g16286 ( 
.A(n_16227),
.B(n_3810),
.Y(n_16286)
);

NAND2xp5_ASAP7_75t_L g16287 ( 
.A(n_16205),
.B(n_16230),
.Y(n_16287)
);

NOR2x1_ASAP7_75t_L g16288 ( 
.A(n_16213),
.B(n_3810),
.Y(n_16288)
);

INVx1_ASAP7_75t_L g16289 ( 
.A(n_16235),
.Y(n_16289)
);

AND3x4_ASAP7_75t_L g16290 ( 
.A(n_16236),
.B(n_3819),
.C(n_3811),
.Y(n_16290)
);

NOR2x1_ASAP7_75t_L g16291 ( 
.A(n_16197),
.B(n_3811),
.Y(n_16291)
);

NOR2x1_ASAP7_75t_L g16292 ( 
.A(n_16176),
.B(n_3812),
.Y(n_16292)
);

NAND2xp5_ASAP7_75t_L g16293 ( 
.A(n_16195),
.B(n_3813),
.Y(n_16293)
);

NOR3x1_ASAP7_75t_L g16294 ( 
.A(n_16184),
.B(n_4231),
.C(n_4230),
.Y(n_16294)
);

NOR2x1_ASAP7_75t_L g16295 ( 
.A(n_16164),
.B(n_3813),
.Y(n_16295)
);

INVx1_ASAP7_75t_L g16296 ( 
.A(n_16212),
.Y(n_16296)
);

AND2x2_ASAP7_75t_L g16297 ( 
.A(n_16175),
.B(n_3814),
.Y(n_16297)
);

NAND3xp33_ASAP7_75t_L g16298 ( 
.A(n_16169),
.B(n_3822),
.C(n_3814),
.Y(n_16298)
);

INVx1_ASAP7_75t_L g16299 ( 
.A(n_16207),
.Y(n_16299)
);

NAND2xp5_ASAP7_75t_L g16300 ( 
.A(n_16232),
.B(n_3815),
.Y(n_16300)
);

NOR2x1_ASAP7_75t_L g16301 ( 
.A(n_16165),
.B(n_3816),
.Y(n_16301)
);

NOR3x1_ASAP7_75t_L g16302 ( 
.A(n_16199),
.B(n_4234),
.C(n_4233),
.Y(n_16302)
);

NOR2x1p5_ASAP7_75t_L g16303 ( 
.A(n_16227),
.B(n_3816),
.Y(n_16303)
);

NAND2xp5_ASAP7_75t_L g16304 ( 
.A(n_16217),
.B(n_3817),
.Y(n_16304)
);

NOR2x1p5_ASAP7_75t_L g16305 ( 
.A(n_16188),
.B(n_3817),
.Y(n_16305)
);

NOR2x1p5_ASAP7_75t_L g16306 ( 
.A(n_16198),
.B(n_3818),
.Y(n_16306)
);

OAI32xp33_ASAP7_75t_L g16307 ( 
.A1(n_16204),
.A2(n_3820),
.A3(n_3818),
.B1(n_3819),
.B2(n_3821),
.Y(n_16307)
);

INVxp67_ASAP7_75t_L g16308 ( 
.A(n_16171),
.Y(n_16308)
);

AND3x4_ASAP7_75t_L g16309 ( 
.A(n_16210),
.B(n_3829),
.C(n_3820),
.Y(n_16309)
);

INVx1_ASAP7_75t_L g16310 ( 
.A(n_16208),
.Y(n_16310)
);

NAND4xp75_ASAP7_75t_L g16311 ( 
.A(n_16211),
.B(n_3824),
.C(n_3822),
.D(n_3823),
.Y(n_16311)
);

NAND2xp5_ASAP7_75t_SL g16312 ( 
.A(n_16223),
.B(n_3824),
.Y(n_16312)
);

NAND4xp75_ASAP7_75t_L g16313 ( 
.A(n_16258),
.B(n_16166),
.C(n_16219),
.D(n_16216),
.Y(n_16313)
);

INVx1_ASAP7_75t_L g16314 ( 
.A(n_16303),
.Y(n_16314)
);

NOR2x1_ASAP7_75t_L g16315 ( 
.A(n_16266),
.B(n_16203),
.Y(n_16315)
);

INVxp67_ASAP7_75t_L g16316 ( 
.A(n_16300),
.Y(n_16316)
);

AND2x2_ASAP7_75t_L g16317 ( 
.A(n_16305),
.B(n_16170),
.Y(n_16317)
);

NAND3xp33_ASAP7_75t_L g16318 ( 
.A(n_16248),
.B(n_16214),
.C(n_16196),
.Y(n_16318)
);

AND2x2_ASAP7_75t_L g16319 ( 
.A(n_16288),
.B(n_16192),
.Y(n_16319)
);

INVx1_ASAP7_75t_L g16320 ( 
.A(n_16290),
.Y(n_16320)
);

NAND4xp75_ASAP7_75t_L g16321 ( 
.A(n_16299),
.B(n_16245),
.C(n_16206),
.D(n_16226),
.Y(n_16321)
);

INVx1_ASAP7_75t_L g16322 ( 
.A(n_16284),
.Y(n_16322)
);

INVx1_ASAP7_75t_L g16323 ( 
.A(n_16274),
.Y(n_16323)
);

INVxp67_ASAP7_75t_L g16324 ( 
.A(n_16283),
.Y(n_16324)
);

XOR2xp5_ASAP7_75t_L g16325 ( 
.A(n_16280),
.B(n_16237),
.Y(n_16325)
);

INVx1_ASAP7_75t_L g16326 ( 
.A(n_16309),
.Y(n_16326)
);

AND2x4_ASAP7_75t_L g16327 ( 
.A(n_16262),
.B(n_16168),
.Y(n_16327)
);

INVx1_ASAP7_75t_L g16328 ( 
.A(n_16285),
.Y(n_16328)
);

AOI22xp5_ASAP7_75t_L g16329 ( 
.A1(n_16252),
.A2(n_16246),
.B1(n_16228),
.B2(n_16222),
.Y(n_16329)
);

INVx1_ASAP7_75t_L g16330 ( 
.A(n_16279),
.Y(n_16330)
);

XOR2xp5_ASAP7_75t_L g16331 ( 
.A(n_16250),
.B(n_16180),
.Y(n_16331)
);

XNOR2x1_ASAP7_75t_L g16332 ( 
.A(n_16257),
.B(n_16238),
.Y(n_16332)
);

INVx1_ASAP7_75t_L g16333 ( 
.A(n_16294),
.Y(n_16333)
);

AND2x2_ASAP7_75t_L g16334 ( 
.A(n_16297),
.B(n_3825),
.Y(n_16334)
);

HB1xp67_ASAP7_75t_L g16335 ( 
.A(n_16286),
.Y(n_16335)
);

OAI22xp5_ASAP7_75t_L g16336 ( 
.A1(n_16282),
.A2(n_16293),
.B1(n_16298),
.B2(n_16304),
.Y(n_16336)
);

AND2x4_ASAP7_75t_L g16337 ( 
.A(n_16278),
.B(n_3825),
.Y(n_16337)
);

INVx1_ASAP7_75t_L g16338 ( 
.A(n_16311),
.Y(n_16338)
);

AND2x2_ASAP7_75t_L g16339 ( 
.A(n_16302),
.B(n_3826),
.Y(n_16339)
);

NAND4xp75_ASAP7_75t_L g16340 ( 
.A(n_16253),
.B(n_16281),
.C(n_16289),
.D(n_16249),
.Y(n_16340)
);

NAND2xp5_ASAP7_75t_L g16341 ( 
.A(n_16269),
.B(n_16270),
.Y(n_16341)
);

INVx1_ASAP7_75t_L g16342 ( 
.A(n_16273),
.Y(n_16342)
);

INVx1_ASAP7_75t_L g16343 ( 
.A(n_16291),
.Y(n_16343)
);

NOR2x1_ASAP7_75t_L g16344 ( 
.A(n_16267),
.B(n_3827),
.Y(n_16344)
);

NAND2xp5_ASAP7_75t_L g16345 ( 
.A(n_16271),
.B(n_3827),
.Y(n_16345)
);

INVx1_ASAP7_75t_L g16346 ( 
.A(n_16265),
.Y(n_16346)
);

INVx1_ASAP7_75t_L g16347 ( 
.A(n_16292),
.Y(n_16347)
);

INVx1_ASAP7_75t_L g16348 ( 
.A(n_16295),
.Y(n_16348)
);

INVx1_ASAP7_75t_L g16349 ( 
.A(n_16301),
.Y(n_16349)
);

XOR2xp5_ASAP7_75t_L g16350 ( 
.A(n_16272),
.B(n_3829),
.Y(n_16350)
);

INVx1_ASAP7_75t_L g16351 ( 
.A(n_16306),
.Y(n_16351)
);

INVx1_ASAP7_75t_L g16352 ( 
.A(n_16307),
.Y(n_16352)
);

NAND3xp33_ASAP7_75t_L g16353 ( 
.A(n_16251),
.B(n_3828),
.C(n_3830),
.Y(n_16353)
);

OR2x2_ASAP7_75t_L g16354 ( 
.A(n_16268),
.B(n_3828),
.Y(n_16354)
);

NAND2x1p5_ASAP7_75t_L g16355 ( 
.A(n_16263),
.B(n_3830),
.Y(n_16355)
);

AND2x4_ASAP7_75t_L g16356 ( 
.A(n_16260),
.B(n_3831),
.Y(n_16356)
);

OAI22xp5_ASAP7_75t_L g16357 ( 
.A1(n_16255),
.A2(n_3833),
.B1(n_3831),
.B2(n_3832),
.Y(n_16357)
);

INVx1_ASAP7_75t_L g16358 ( 
.A(n_16287),
.Y(n_16358)
);

NAND2xp5_ASAP7_75t_L g16359 ( 
.A(n_16277),
.B(n_3833),
.Y(n_16359)
);

NOR3xp33_ASAP7_75t_L g16360 ( 
.A(n_16259),
.B(n_16308),
.C(n_16276),
.Y(n_16360)
);

OR2x2_ASAP7_75t_L g16361 ( 
.A(n_16264),
.B(n_3834),
.Y(n_16361)
);

NAND2xp5_ASAP7_75t_L g16362 ( 
.A(n_16263),
.B(n_3834),
.Y(n_16362)
);

INVx1_ASAP7_75t_L g16363 ( 
.A(n_16256),
.Y(n_16363)
);

XOR2xp5_ASAP7_75t_L g16364 ( 
.A(n_16275),
.B(n_16260),
.Y(n_16364)
);

NOR3xp33_ASAP7_75t_L g16365 ( 
.A(n_16310),
.B(n_3836),
.C(n_3837),
.Y(n_16365)
);

AND2x4_ASAP7_75t_L g16366 ( 
.A(n_16296),
.B(n_3836),
.Y(n_16366)
);

XNOR2xp5_ASAP7_75t_L g16367 ( 
.A(n_16312),
.B(n_3837),
.Y(n_16367)
);

AND2x2_ASAP7_75t_SL g16368 ( 
.A(n_16261),
.B(n_3838),
.Y(n_16368)
);

NAND2x1_ASAP7_75t_L g16369 ( 
.A(n_16254),
.B(n_3838),
.Y(n_16369)
);

INVx1_ASAP7_75t_L g16370 ( 
.A(n_16368),
.Y(n_16370)
);

INVx1_ASAP7_75t_L g16371 ( 
.A(n_16334),
.Y(n_16371)
);

INVx1_ASAP7_75t_L g16372 ( 
.A(n_16369),
.Y(n_16372)
);

NAND4xp75_ASAP7_75t_L g16373 ( 
.A(n_16346),
.B(n_3841),
.C(n_3839),
.D(n_3840),
.Y(n_16373)
);

AND2x4_ASAP7_75t_L g16374 ( 
.A(n_16337),
.B(n_3840),
.Y(n_16374)
);

AND2x2_ASAP7_75t_L g16375 ( 
.A(n_16339),
.B(n_3841),
.Y(n_16375)
);

NOR2xp33_ASAP7_75t_L g16376 ( 
.A(n_16354),
.B(n_3842),
.Y(n_16376)
);

NOR2x1_ASAP7_75t_L g16377 ( 
.A(n_16340),
.B(n_3843),
.Y(n_16377)
);

INVx2_ASAP7_75t_SL g16378 ( 
.A(n_16361),
.Y(n_16378)
);

INVx2_ASAP7_75t_SL g16379 ( 
.A(n_16355),
.Y(n_16379)
);

XNOR2x1_ASAP7_75t_L g16380 ( 
.A(n_16332),
.B(n_3844),
.Y(n_16380)
);

INVx1_ASAP7_75t_L g16381 ( 
.A(n_16344),
.Y(n_16381)
);

AOI22xp5_ASAP7_75t_L g16382 ( 
.A1(n_16363),
.A2(n_3853),
.B1(n_3861),
.B2(n_3845),
.Y(n_16382)
);

XNOR2xp5_ASAP7_75t_L g16383 ( 
.A(n_16364),
.B(n_3845),
.Y(n_16383)
);

OAI21xp33_ASAP7_75t_L g16384 ( 
.A1(n_16329),
.A2(n_3846),
.B(n_3847),
.Y(n_16384)
);

NOR3xp33_ASAP7_75t_L g16385 ( 
.A(n_16324),
.B(n_3846),
.C(n_3847),
.Y(n_16385)
);

XNOR2x1_ASAP7_75t_L g16386 ( 
.A(n_16331),
.B(n_3848),
.Y(n_16386)
);

AND2x2_ASAP7_75t_L g16387 ( 
.A(n_16317),
.B(n_3848),
.Y(n_16387)
);

NOR3xp33_ASAP7_75t_L g16388 ( 
.A(n_16343),
.B(n_3849),
.C(n_3850),
.Y(n_16388)
);

NOR3xp33_ASAP7_75t_L g16389 ( 
.A(n_16335),
.B(n_16330),
.C(n_16360),
.Y(n_16389)
);

NAND4xp75_ASAP7_75t_L g16390 ( 
.A(n_16333),
.B(n_3851),
.C(n_3849),
.D(n_3850),
.Y(n_16390)
);

NOR2xp67_ASAP7_75t_L g16391 ( 
.A(n_16318),
.B(n_3852),
.Y(n_16391)
);

INVx1_ASAP7_75t_L g16392 ( 
.A(n_16345),
.Y(n_16392)
);

XNOR2xp5_ASAP7_75t_L g16393 ( 
.A(n_16325),
.B(n_3852),
.Y(n_16393)
);

OR3x2_ASAP7_75t_L g16394 ( 
.A(n_16338),
.B(n_3855),
.C(n_3854),
.Y(n_16394)
);

INVx3_ASAP7_75t_SL g16395 ( 
.A(n_16327),
.Y(n_16395)
);

OR2x2_ASAP7_75t_L g16396 ( 
.A(n_16359),
.B(n_3853),
.Y(n_16396)
);

XNOR2xp5_ASAP7_75t_L g16397 ( 
.A(n_16367),
.B(n_16358),
.Y(n_16397)
);

NOR2xp67_ASAP7_75t_L g16398 ( 
.A(n_16314),
.B(n_3854),
.Y(n_16398)
);

AND2x4_ASAP7_75t_L g16399 ( 
.A(n_16320),
.B(n_3855),
.Y(n_16399)
);

NOR2x1_ASAP7_75t_L g16400 ( 
.A(n_16348),
.B(n_3856),
.Y(n_16400)
);

AOI22xp5_ASAP7_75t_L g16401 ( 
.A1(n_16322),
.A2(n_3865),
.B1(n_3873),
.B2(n_3856),
.Y(n_16401)
);

INVx3_ASAP7_75t_L g16402 ( 
.A(n_16321),
.Y(n_16402)
);

AND2x2_ASAP7_75t_L g16403 ( 
.A(n_16319),
.B(n_16315),
.Y(n_16403)
);

INVx2_ASAP7_75t_L g16404 ( 
.A(n_16350),
.Y(n_16404)
);

INVx3_ASAP7_75t_L g16405 ( 
.A(n_16313),
.Y(n_16405)
);

INVx1_ASAP7_75t_L g16406 ( 
.A(n_16353),
.Y(n_16406)
);

XNOR2xp5_ASAP7_75t_L g16407 ( 
.A(n_16336),
.B(n_3857),
.Y(n_16407)
);

NAND4xp75_ASAP7_75t_L g16408 ( 
.A(n_16349),
.B(n_3860),
.C(n_3858),
.D(n_3859),
.Y(n_16408)
);

NOR2xp67_ASAP7_75t_L g16409 ( 
.A(n_16352),
.B(n_3859),
.Y(n_16409)
);

INVx2_ASAP7_75t_L g16410 ( 
.A(n_16356),
.Y(n_16410)
);

NOR2x1_ASAP7_75t_L g16411 ( 
.A(n_16347),
.B(n_16323),
.Y(n_16411)
);

NAND4xp75_ASAP7_75t_L g16412 ( 
.A(n_16328),
.B(n_16351),
.C(n_16326),
.D(n_16342),
.Y(n_16412)
);

AOI22xp5_ASAP7_75t_L g16413 ( 
.A1(n_16316),
.A2(n_3870),
.B1(n_3878),
.B2(n_3861),
.Y(n_16413)
);

XNOR2xp5_ASAP7_75t_L g16414 ( 
.A(n_16341),
.B(n_3862),
.Y(n_16414)
);

XOR2xp5_ASAP7_75t_SL g16415 ( 
.A(n_16365),
.B(n_3863),
.Y(n_16415)
);

INVx1_ASAP7_75t_L g16416 ( 
.A(n_16357),
.Y(n_16416)
);

AND2x4_ASAP7_75t_L g16417 ( 
.A(n_16366),
.B(n_3865),
.Y(n_16417)
);

AND2x4_ASAP7_75t_L g16418 ( 
.A(n_16362),
.B(n_3866),
.Y(n_16418)
);

AND2x4_ASAP7_75t_L g16419 ( 
.A(n_16334),
.B(n_3867),
.Y(n_16419)
);

XOR2x2_ASAP7_75t_L g16420 ( 
.A(n_16344),
.B(n_3867),
.Y(n_16420)
);

INVx1_ASAP7_75t_L g16421 ( 
.A(n_16368),
.Y(n_16421)
);

AOI21xp5_ASAP7_75t_L g16422 ( 
.A1(n_16364),
.A2(n_3868),
.B(n_3869),
.Y(n_16422)
);

NOR3xp33_ASAP7_75t_L g16423 ( 
.A(n_16340),
.B(n_3868),
.C(n_3869),
.Y(n_16423)
);

INVx2_ASAP7_75t_L g16424 ( 
.A(n_16355),
.Y(n_16424)
);

INVx1_ASAP7_75t_L g16425 ( 
.A(n_16368),
.Y(n_16425)
);

INVx2_ASAP7_75t_SL g16426 ( 
.A(n_16368),
.Y(n_16426)
);

OAI21xp5_ASAP7_75t_SL g16427 ( 
.A1(n_16367),
.A2(n_3870),
.B(n_3871),
.Y(n_16427)
);

INVx2_ASAP7_75t_L g16428 ( 
.A(n_16355),
.Y(n_16428)
);

NAND4xp75_ASAP7_75t_L g16429 ( 
.A(n_16346),
.B(n_3874),
.C(n_3872),
.D(n_3873),
.Y(n_16429)
);

NAND2xp5_ASAP7_75t_L g16430 ( 
.A(n_16368),
.B(n_3874),
.Y(n_16430)
);

NOR3xp33_ASAP7_75t_L g16431 ( 
.A(n_16340),
.B(n_3872),
.C(n_3875),
.Y(n_16431)
);

XOR2x1_ASAP7_75t_L g16432 ( 
.A(n_16335),
.B(n_3876),
.Y(n_16432)
);

INVx1_ASAP7_75t_L g16433 ( 
.A(n_16368),
.Y(n_16433)
);

XNOR2x1_ASAP7_75t_L g16434 ( 
.A(n_16340),
.B(n_3876),
.Y(n_16434)
);

INVx1_ASAP7_75t_L g16435 ( 
.A(n_16375),
.Y(n_16435)
);

OAI222xp33_ASAP7_75t_L g16436 ( 
.A1(n_16377),
.A2(n_3881),
.B1(n_3883),
.B2(n_3877),
.C1(n_3879),
.C2(n_3882),
.Y(n_16436)
);

AOI311xp33_ASAP7_75t_L g16437 ( 
.A1(n_16389),
.A2(n_3883),
.A3(n_3879),
.B(n_3881),
.C(n_3884),
.Y(n_16437)
);

OAI22xp5_ASAP7_75t_L g16438 ( 
.A1(n_16394),
.A2(n_3887),
.B1(n_3885),
.B2(n_3886),
.Y(n_16438)
);

INVx1_ASAP7_75t_L g16439 ( 
.A(n_16432),
.Y(n_16439)
);

NAND2xp5_ASAP7_75t_L g16440 ( 
.A(n_16409),
.B(n_3885),
.Y(n_16440)
);

INVx1_ASAP7_75t_L g16441 ( 
.A(n_16430),
.Y(n_16441)
);

NAND4xp25_ASAP7_75t_L g16442 ( 
.A(n_16423),
.B(n_3888),
.C(n_3886),
.D(n_3887),
.Y(n_16442)
);

NOR3xp33_ASAP7_75t_L g16443 ( 
.A(n_16405),
.B(n_3888),
.C(n_3889),
.Y(n_16443)
);

AOI22xp5_ASAP7_75t_L g16444 ( 
.A1(n_16431),
.A2(n_3891),
.B1(n_3889),
.B2(n_3890),
.Y(n_16444)
);

NAND3xp33_ASAP7_75t_SL g16445 ( 
.A(n_16370),
.B(n_3892),
.C(n_3893),
.Y(n_16445)
);

NAND5xp2_ASAP7_75t_L g16446 ( 
.A(n_16403),
.B(n_3895),
.C(n_3897),
.D(n_3894),
.E(n_3896),
.Y(n_16446)
);

NOR2xp33_ASAP7_75t_L g16447 ( 
.A(n_16395),
.B(n_3893),
.Y(n_16447)
);

NOR2x1p5_ASAP7_75t_L g16448 ( 
.A(n_16412),
.B(n_3894),
.Y(n_16448)
);

NOR3x2_ASAP7_75t_L g16449 ( 
.A(n_16396),
.B(n_3895),
.C(n_3896),
.Y(n_16449)
);

AOI22xp33_ASAP7_75t_SL g16450 ( 
.A1(n_16402),
.A2(n_3899),
.B1(n_3897),
.B2(n_3898),
.Y(n_16450)
);

AO22x2_ASAP7_75t_L g16451 ( 
.A1(n_16434),
.A2(n_3906),
.B1(n_3914),
.B2(n_3898),
.Y(n_16451)
);

INVx2_ASAP7_75t_L g16452 ( 
.A(n_16386),
.Y(n_16452)
);

OAI211xp5_ASAP7_75t_L g16453 ( 
.A1(n_16411),
.A2(n_16391),
.B(n_16372),
.C(n_16427),
.Y(n_16453)
);

AND2x2_ASAP7_75t_L g16454 ( 
.A(n_16426),
.B(n_3899),
.Y(n_16454)
);

NAND5xp2_ASAP7_75t_L g16455 ( 
.A(n_16421),
.B(n_3902),
.C(n_3904),
.D(n_3901),
.E(n_3903),
.Y(n_16455)
);

AO22x2_ASAP7_75t_L g16456 ( 
.A1(n_16425),
.A2(n_3910),
.B1(n_3919),
.B2(n_3900),
.Y(n_16456)
);

OAI22xp5_ASAP7_75t_L g16457 ( 
.A1(n_16380),
.A2(n_3904),
.B1(n_3900),
.B2(n_3902),
.Y(n_16457)
);

NOR3xp33_ASAP7_75t_L g16458 ( 
.A(n_16433),
.B(n_3905),
.C(n_3906),
.Y(n_16458)
);

NOR2xp33_ASAP7_75t_L g16459 ( 
.A(n_16379),
.B(n_3907),
.Y(n_16459)
);

INVx1_ASAP7_75t_L g16460 ( 
.A(n_16374),
.Y(n_16460)
);

INVx1_ASAP7_75t_L g16461 ( 
.A(n_16420),
.Y(n_16461)
);

NOR2x1p5_ASAP7_75t_L g16462 ( 
.A(n_16410),
.B(n_3907),
.Y(n_16462)
);

AOI22xp5_ASAP7_75t_L g16463 ( 
.A1(n_16376),
.A2(n_3911),
.B1(n_3908),
.B2(n_3909),
.Y(n_16463)
);

INVxp67_ASAP7_75t_L g16464 ( 
.A(n_16400),
.Y(n_16464)
);

NAND2xp5_ASAP7_75t_L g16465 ( 
.A(n_16398),
.B(n_3908),
.Y(n_16465)
);

AOI211xp5_ASAP7_75t_L g16466 ( 
.A1(n_16381),
.A2(n_3912),
.B(n_3909),
.C(n_3911),
.Y(n_16466)
);

NOR3xp33_ASAP7_75t_L g16467 ( 
.A(n_16378),
.B(n_3912),
.C(n_3913),
.Y(n_16467)
);

NAND4xp25_ASAP7_75t_L g16468 ( 
.A(n_16371),
.B(n_3916),
.C(n_3913),
.D(n_3915),
.Y(n_16468)
);

INVx1_ASAP7_75t_L g16469 ( 
.A(n_16407),
.Y(n_16469)
);

OAI22xp5_ASAP7_75t_L g16470 ( 
.A1(n_16424),
.A2(n_3917),
.B1(n_3915),
.B2(n_3916),
.Y(n_16470)
);

NAND3xp33_ASAP7_75t_SL g16471 ( 
.A(n_16428),
.B(n_3917),
.C(n_3918),
.Y(n_16471)
);

INVx1_ASAP7_75t_L g16472 ( 
.A(n_16417),
.Y(n_16472)
);

AND2x4_ASAP7_75t_L g16473 ( 
.A(n_16416),
.B(n_3918),
.Y(n_16473)
);

NAND3xp33_ASAP7_75t_L g16474 ( 
.A(n_16397),
.B(n_3919),
.C(n_3920),
.Y(n_16474)
);

XNOR2xp5_ASAP7_75t_SL g16475 ( 
.A(n_16406),
.B(n_3922),
.Y(n_16475)
);

INVx2_ASAP7_75t_L g16476 ( 
.A(n_16373),
.Y(n_16476)
);

AND3x2_ASAP7_75t_L g16477 ( 
.A(n_16388),
.B(n_3921),
.C(n_3922),
.Y(n_16477)
);

NAND3xp33_ASAP7_75t_L g16478 ( 
.A(n_16392),
.B(n_3921),
.C(n_3923),
.Y(n_16478)
);

INVx1_ASAP7_75t_L g16479 ( 
.A(n_16419),
.Y(n_16479)
);

AOI211xp5_ASAP7_75t_L g16480 ( 
.A1(n_16404),
.A2(n_3925),
.B(n_3923),
.C(n_3924),
.Y(n_16480)
);

OAI22xp5_ASAP7_75t_L g16481 ( 
.A1(n_16422),
.A2(n_3927),
.B1(n_3924),
.B2(n_3926),
.Y(n_16481)
);

O2A1O1Ixp33_ASAP7_75t_L g16482 ( 
.A1(n_16384),
.A2(n_3928),
.B(n_3926),
.C(n_3927),
.Y(n_16482)
);

AOI211xp5_ASAP7_75t_L g16483 ( 
.A1(n_16385),
.A2(n_3930),
.B(n_3928),
.C(n_3929),
.Y(n_16483)
);

NOR2x1p5_ASAP7_75t_L g16484 ( 
.A(n_16415),
.B(n_3929),
.Y(n_16484)
);

INVx1_ASAP7_75t_L g16485 ( 
.A(n_16418),
.Y(n_16485)
);

NOR3xp33_ASAP7_75t_L g16486 ( 
.A(n_16429),
.B(n_3930),
.C(n_3931),
.Y(n_16486)
);

NAND2x1p5_ASAP7_75t_L g16487 ( 
.A(n_16382),
.B(n_16401),
.Y(n_16487)
);

INVx1_ASAP7_75t_L g16488 ( 
.A(n_16383),
.Y(n_16488)
);

AOI21xp5_ASAP7_75t_L g16489 ( 
.A1(n_16393),
.A2(n_16414),
.B(n_16413),
.Y(n_16489)
);

AOI22xp5_ASAP7_75t_L g16490 ( 
.A1(n_16390),
.A2(n_16408),
.B1(n_16387),
.B2(n_16399),
.Y(n_16490)
);

AND2x4_ASAP7_75t_L g16491 ( 
.A(n_16374),
.B(n_3931),
.Y(n_16491)
);

OAI222xp33_ASAP7_75t_L g16492 ( 
.A1(n_16377),
.A2(n_3934),
.B1(n_3936),
.B2(n_3932),
.C1(n_3933),
.C2(n_3935),
.Y(n_16492)
);

OAI22xp5_ASAP7_75t_L g16493 ( 
.A1(n_16394),
.A2(n_3934),
.B1(n_3932),
.B2(n_3933),
.Y(n_16493)
);

CKINVDCx20_ASAP7_75t_R g16494 ( 
.A(n_16395),
.Y(n_16494)
);

NAND4xp25_ASAP7_75t_L g16495 ( 
.A(n_16389),
.B(n_3937),
.C(n_3935),
.D(n_3936),
.Y(n_16495)
);

NAND3xp33_ASAP7_75t_SL g16496 ( 
.A(n_16389),
.B(n_3937),
.C(n_3938),
.Y(n_16496)
);

NAND3xp33_ASAP7_75t_L g16497 ( 
.A(n_16434),
.B(n_3938),
.C(n_3939),
.Y(n_16497)
);

NAND4xp25_ASAP7_75t_L g16498 ( 
.A(n_16389),
.B(n_3941),
.C(n_3939),
.D(n_3940),
.Y(n_16498)
);

OAI211xp5_ASAP7_75t_SL g16499 ( 
.A1(n_16411),
.A2(n_3943),
.B(n_3941),
.C(n_3942),
.Y(n_16499)
);

AOI21xp5_ASAP7_75t_L g16500 ( 
.A1(n_16426),
.A2(n_3944),
.B(n_3945),
.Y(n_16500)
);

NAND4xp25_ASAP7_75t_SL g16501 ( 
.A(n_16423),
.B(n_3947),
.C(n_3944),
.D(n_3946),
.Y(n_16501)
);

AOI22xp5_ASAP7_75t_L g16502 ( 
.A1(n_16423),
.A2(n_3949),
.B1(n_3946),
.B2(n_3948),
.Y(n_16502)
);

AO22x2_ASAP7_75t_L g16503 ( 
.A1(n_16434),
.A2(n_3956),
.B1(n_3964),
.B2(n_3948),
.Y(n_16503)
);

NOR3xp33_ASAP7_75t_L g16504 ( 
.A(n_16405),
.B(n_3949),
.C(n_3950),
.Y(n_16504)
);

NAND2xp5_ASAP7_75t_L g16505 ( 
.A(n_16432),
.B(n_3951),
.Y(n_16505)
);

NOR2x1p5_ASAP7_75t_L g16506 ( 
.A(n_16432),
.B(n_3951),
.Y(n_16506)
);

NOR3xp33_ASAP7_75t_L g16507 ( 
.A(n_16405),
.B(n_3952),
.C(n_3953),
.Y(n_16507)
);

NAND2xp5_ASAP7_75t_SL g16508 ( 
.A(n_16423),
.B(n_3952),
.Y(n_16508)
);

NAND3xp33_ASAP7_75t_L g16509 ( 
.A(n_16434),
.B(n_3953),
.C(n_3954),
.Y(n_16509)
);

OAI211xp5_ASAP7_75t_SL g16510 ( 
.A1(n_16411),
.A2(n_3956),
.B(n_3954),
.C(n_3955),
.Y(n_16510)
);

NOR2x1_ASAP7_75t_L g16511 ( 
.A(n_16506),
.B(n_16439),
.Y(n_16511)
);

NAND2xp5_ASAP7_75t_L g16512 ( 
.A(n_16477),
.B(n_4245),
.Y(n_16512)
);

HB1xp67_ASAP7_75t_L g16513 ( 
.A(n_16448),
.Y(n_16513)
);

NOR2x1p5_ASAP7_75t_L g16514 ( 
.A(n_16476),
.B(n_3955),
.Y(n_16514)
);

NAND2xp5_ASAP7_75t_L g16515 ( 
.A(n_16486),
.B(n_4249),
.Y(n_16515)
);

AND2x2_ASAP7_75t_L g16516 ( 
.A(n_16484),
.B(n_3957),
.Y(n_16516)
);

AOI221xp5_ASAP7_75t_L g16517 ( 
.A1(n_16482),
.A2(n_3960),
.B1(n_3958),
.B2(n_3959),
.C(n_3961),
.Y(n_16517)
);

AND2x4_ASAP7_75t_L g16518 ( 
.A(n_16494),
.B(n_3960),
.Y(n_16518)
);

HB1xp67_ASAP7_75t_L g16519 ( 
.A(n_16462),
.Y(n_16519)
);

NOR3xp33_ASAP7_75t_SL g16520 ( 
.A(n_16453),
.B(n_3969),
.C(n_3961),
.Y(n_16520)
);

AOI22xp33_ASAP7_75t_SL g16521 ( 
.A1(n_16497),
.A2(n_3964),
.B1(n_3962),
.B2(n_3963),
.Y(n_16521)
);

NAND2x1p5_ASAP7_75t_L g16522 ( 
.A(n_16479),
.B(n_3962),
.Y(n_16522)
);

INVx2_ASAP7_75t_SL g16523 ( 
.A(n_16491),
.Y(n_16523)
);

BUFx6f_ASAP7_75t_L g16524 ( 
.A(n_16435),
.Y(n_16524)
);

INVx1_ASAP7_75t_L g16525 ( 
.A(n_16465),
.Y(n_16525)
);

NOR2xp33_ASAP7_75t_L g16526 ( 
.A(n_16464),
.B(n_4235),
.Y(n_16526)
);

INVx3_ASAP7_75t_L g16527 ( 
.A(n_16449),
.Y(n_16527)
);

NAND2xp5_ASAP7_75t_L g16528 ( 
.A(n_16438),
.B(n_16493),
.Y(n_16528)
);

OAI221xp5_ASAP7_75t_L g16529 ( 
.A1(n_16509),
.A2(n_3966),
.B1(n_3963),
.B2(n_3965),
.C(n_3967),
.Y(n_16529)
);

BUFx2_ASAP7_75t_L g16530 ( 
.A(n_16475),
.Y(n_16530)
);

INVxp67_ASAP7_75t_L g16531 ( 
.A(n_16505),
.Y(n_16531)
);

OAI22x1_ASAP7_75t_L g16532 ( 
.A1(n_16490),
.A2(n_3967),
.B1(n_3965),
.B2(n_3966),
.Y(n_16532)
);

AND3x4_ASAP7_75t_L g16533 ( 
.A(n_16452),
.B(n_16504),
.C(n_16443),
.Y(n_16533)
);

AO22x2_ASAP7_75t_L g16534 ( 
.A1(n_16472),
.A2(n_3976),
.B1(n_3984),
.B2(n_3968),
.Y(n_16534)
);

AOI22xp5_ASAP7_75t_L g16535 ( 
.A1(n_16501),
.A2(n_3970),
.B1(n_3968),
.B2(n_3969),
.Y(n_16535)
);

NAND4xp75_ASAP7_75t_L g16536 ( 
.A(n_16460),
.B(n_3972),
.C(n_3970),
.D(n_3971),
.Y(n_16536)
);

INVx3_ASAP7_75t_L g16537 ( 
.A(n_16487),
.Y(n_16537)
);

AND2x2_ASAP7_75t_L g16538 ( 
.A(n_16485),
.B(n_3971),
.Y(n_16538)
);

NAND2xp5_ASAP7_75t_L g16539 ( 
.A(n_16440),
.B(n_16483),
.Y(n_16539)
);

OAI22xp5_ASAP7_75t_L g16540 ( 
.A1(n_16444),
.A2(n_3974),
.B1(n_3975),
.B2(n_3973),
.Y(n_16540)
);

AND2x4_ASAP7_75t_L g16541 ( 
.A(n_16508),
.B(n_16488),
.Y(n_16541)
);

OAI22xp5_ASAP7_75t_SL g16542 ( 
.A1(n_16469),
.A2(n_16461),
.B1(n_16441),
.B2(n_16502),
.Y(n_16542)
);

XNOR2xp5_ASAP7_75t_L g16543 ( 
.A(n_16451),
.B(n_3972),
.Y(n_16543)
);

NOR2x1_ASAP7_75t_L g16544 ( 
.A(n_16496),
.B(n_3974),
.Y(n_16544)
);

NAND5xp2_ASAP7_75t_L g16545 ( 
.A(n_16489),
.B(n_3976),
.C(n_3973),
.D(n_3975),
.E(n_3977),
.Y(n_16545)
);

NAND2x1_ASAP7_75t_SL g16546 ( 
.A(n_16463),
.B(n_3977),
.Y(n_16546)
);

XNOR2xp5_ASAP7_75t_L g16547 ( 
.A(n_16451),
.B(n_3978),
.Y(n_16547)
);

INVx1_ASAP7_75t_L g16548 ( 
.A(n_16503),
.Y(n_16548)
);

AOI32xp33_ASAP7_75t_L g16549 ( 
.A1(n_16499),
.A2(n_3980),
.A3(n_3978),
.B1(n_3979),
.B2(n_3981),
.Y(n_16549)
);

INVx2_ASAP7_75t_L g16550 ( 
.A(n_16503),
.Y(n_16550)
);

INVx1_ASAP7_75t_L g16551 ( 
.A(n_16442),
.Y(n_16551)
);

NAND4xp25_ASAP7_75t_L g16552 ( 
.A(n_16437),
.B(n_3981),
.C(n_3979),
.D(n_3980),
.Y(n_16552)
);

OR3x1_ASAP7_75t_L g16553 ( 
.A(n_16510),
.B(n_3982),
.C(n_3983),
.Y(n_16553)
);

INVx2_ASAP7_75t_L g16554 ( 
.A(n_16456),
.Y(n_16554)
);

AOI222xp33_ASAP7_75t_L g16555 ( 
.A1(n_16481),
.A2(n_3986),
.B1(n_3988),
.B2(n_3984),
.C1(n_3985),
.C2(n_3987),
.Y(n_16555)
);

NOR2xp33_ASAP7_75t_L g16556 ( 
.A(n_16471),
.B(n_4246),
.Y(n_16556)
);

AND2x4_ASAP7_75t_L g16557 ( 
.A(n_16507),
.B(n_3985),
.Y(n_16557)
);

AOI22xp5_ASAP7_75t_L g16558 ( 
.A1(n_16445),
.A2(n_3989),
.B1(n_3986),
.B2(n_3987),
.Y(n_16558)
);

OAI22xp5_ASAP7_75t_L g16559 ( 
.A1(n_16500),
.A2(n_3991),
.B1(n_3992),
.B2(n_3990),
.Y(n_16559)
);

NAND2xp5_ASAP7_75t_L g16560 ( 
.A(n_16467),
.B(n_4229),
.Y(n_16560)
);

OAI22xp5_ASAP7_75t_L g16561 ( 
.A1(n_16457),
.A2(n_3991),
.B1(n_3993),
.B2(n_3990),
.Y(n_16561)
);

CKINVDCx5p33_ASAP7_75t_R g16562 ( 
.A(n_16524),
.Y(n_16562)
);

NAND4xp75_ASAP7_75t_L g16563 ( 
.A(n_16511),
.B(n_16447),
.C(n_16459),
.D(n_16454),
.Y(n_16563)
);

INVx2_ASAP7_75t_L g16564 ( 
.A(n_16522),
.Y(n_16564)
);

AOI22xp5_ASAP7_75t_L g16565 ( 
.A1(n_16516),
.A2(n_16537),
.B1(n_16561),
.B2(n_16540),
.Y(n_16565)
);

AOI22xp33_ASAP7_75t_L g16566 ( 
.A1(n_16524),
.A2(n_16458),
.B1(n_16446),
.B2(n_16455),
.Y(n_16566)
);

NAND2xp5_ASAP7_75t_L g16567 ( 
.A(n_16549),
.B(n_16480),
.Y(n_16567)
);

NOR2x1_ASAP7_75t_L g16568 ( 
.A(n_16548),
.B(n_16436),
.Y(n_16568)
);

AND2x4_ASAP7_75t_L g16569 ( 
.A(n_16523),
.B(n_16474),
.Y(n_16569)
);

INVx3_ASAP7_75t_L g16570 ( 
.A(n_16557),
.Y(n_16570)
);

AND2x2_ASAP7_75t_L g16571 ( 
.A(n_16519),
.B(n_16450),
.Y(n_16571)
);

INVx2_ASAP7_75t_L g16572 ( 
.A(n_16514),
.Y(n_16572)
);

INVx2_ASAP7_75t_L g16573 ( 
.A(n_16536),
.Y(n_16573)
);

INVx1_ASAP7_75t_SL g16574 ( 
.A(n_16515),
.Y(n_16574)
);

XNOR2xp5_ASAP7_75t_L g16575 ( 
.A(n_16543),
.B(n_16547),
.Y(n_16575)
);

AND2x4_ASAP7_75t_L g16576 ( 
.A(n_16544),
.B(n_16520),
.Y(n_16576)
);

INVx1_ASAP7_75t_L g16577 ( 
.A(n_16512),
.Y(n_16577)
);

AND2x4_ASAP7_75t_L g16578 ( 
.A(n_16551),
.B(n_16478),
.Y(n_16578)
);

HB1xp67_ASAP7_75t_L g16579 ( 
.A(n_16554),
.Y(n_16579)
);

NAND2xp5_ASAP7_75t_L g16580 ( 
.A(n_16556),
.B(n_16466),
.Y(n_16580)
);

XNOR2x1_ASAP7_75t_L g16581 ( 
.A(n_16533),
.B(n_16541),
.Y(n_16581)
);

AND2x2_ASAP7_75t_L g16582 ( 
.A(n_16513),
.B(n_16470),
.Y(n_16582)
);

INVx1_ASAP7_75t_L g16583 ( 
.A(n_16560),
.Y(n_16583)
);

INVx3_ASAP7_75t_L g16584 ( 
.A(n_16550),
.Y(n_16584)
);

NAND2xp5_ASAP7_75t_L g16585 ( 
.A(n_16535),
.B(n_16495),
.Y(n_16585)
);

INVx1_ASAP7_75t_L g16586 ( 
.A(n_16546),
.Y(n_16586)
);

INVx4_ASAP7_75t_L g16587 ( 
.A(n_16527),
.Y(n_16587)
);

NAND4xp75_ASAP7_75t_L g16588 ( 
.A(n_16525),
.B(n_16492),
.C(n_16498),
.D(n_16468),
.Y(n_16588)
);

INVx1_ASAP7_75t_L g16589 ( 
.A(n_16553),
.Y(n_16589)
);

INVx2_ASAP7_75t_L g16590 ( 
.A(n_16532),
.Y(n_16590)
);

AND2x2_ASAP7_75t_SL g16591 ( 
.A(n_16530),
.B(n_16473),
.Y(n_16591)
);

INVx1_ASAP7_75t_L g16592 ( 
.A(n_16552),
.Y(n_16592)
);

INVx1_ASAP7_75t_L g16593 ( 
.A(n_16558),
.Y(n_16593)
);

INVx1_ASAP7_75t_L g16594 ( 
.A(n_16539),
.Y(n_16594)
);

NAND3x1_ASAP7_75t_L g16595 ( 
.A(n_16528),
.B(n_16456),
.C(n_3989),
.Y(n_16595)
);

INVx2_ASAP7_75t_L g16596 ( 
.A(n_16518),
.Y(n_16596)
);

OR4x1_ASAP7_75t_L g16597 ( 
.A(n_16592),
.B(n_16542),
.C(n_16531),
.D(n_16517),
.Y(n_16597)
);

INVxp67_ASAP7_75t_SL g16598 ( 
.A(n_16579),
.Y(n_16598)
);

XOR2xp5_ASAP7_75t_L g16599 ( 
.A(n_16581),
.B(n_16521),
.Y(n_16599)
);

OAI21xp5_ASAP7_75t_L g16600 ( 
.A1(n_16568),
.A2(n_16559),
.B(n_16529),
.Y(n_16600)
);

NAND3xp33_ASAP7_75t_L g16601 ( 
.A(n_16562),
.B(n_16555),
.C(n_16526),
.Y(n_16601)
);

INVx1_ASAP7_75t_L g16602 ( 
.A(n_16595),
.Y(n_16602)
);

AND3x2_ASAP7_75t_L g16603 ( 
.A(n_16586),
.B(n_16538),
.C(n_16545),
.Y(n_16603)
);

INVx2_ASAP7_75t_L g16604 ( 
.A(n_16576),
.Y(n_16604)
);

INVx1_ASAP7_75t_L g16605 ( 
.A(n_16585),
.Y(n_16605)
);

XNOR2x1_ASAP7_75t_L g16606 ( 
.A(n_16575),
.B(n_16534),
.Y(n_16606)
);

NAND2x1p5_ASAP7_75t_L g16607 ( 
.A(n_16564),
.B(n_16534),
.Y(n_16607)
);

AOI22xp5_ASAP7_75t_L g16608 ( 
.A1(n_16584),
.A2(n_4001),
.B1(n_4009),
.B2(n_3993),
.Y(n_16608)
);

INVx1_ASAP7_75t_L g16609 ( 
.A(n_16572),
.Y(n_16609)
);

HB1xp67_ASAP7_75t_L g16610 ( 
.A(n_16588),
.Y(n_16610)
);

NAND2xp5_ASAP7_75t_L g16611 ( 
.A(n_16566),
.B(n_3994),
.Y(n_16611)
);

OAI22xp33_ASAP7_75t_L g16612 ( 
.A1(n_16587),
.A2(n_16590),
.B1(n_16565),
.B2(n_16573),
.Y(n_16612)
);

NAND4xp75_ASAP7_75t_L g16613 ( 
.A(n_16591),
.B(n_3996),
.C(n_3994),
.D(n_3995),
.Y(n_16613)
);

OAI22xp5_ASAP7_75t_L g16614 ( 
.A1(n_16589),
.A2(n_3999),
.B1(n_3997),
.B2(n_3998),
.Y(n_16614)
);

AOI22x1_ASAP7_75t_L g16615 ( 
.A1(n_16596),
.A2(n_3999),
.B1(n_3997),
.B2(n_3998),
.Y(n_16615)
);

XOR2xp5_ASAP7_75t_L g16616 ( 
.A(n_16563),
.B(n_4000),
.Y(n_16616)
);

OAI22xp5_ASAP7_75t_L g16617 ( 
.A1(n_16594),
.A2(n_4002),
.B1(n_4000),
.B2(n_4001),
.Y(n_16617)
);

NAND2xp5_ASAP7_75t_L g16618 ( 
.A(n_16570),
.B(n_4002),
.Y(n_16618)
);

INVx2_ASAP7_75t_L g16619 ( 
.A(n_16569),
.Y(n_16619)
);

OAI22xp5_ASAP7_75t_L g16620 ( 
.A1(n_16567),
.A2(n_4005),
.B1(n_4003),
.B2(n_4004),
.Y(n_16620)
);

OAI21x1_ASAP7_75t_L g16621 ( 
.A1(n_16580),
.A2(n_4003),
.B(n_4004),
.Y(n_16621)
);

AOI22x1_ASAP7_75t_L g16622 ( 
.A1(n_16571),
.A2(n_4008),
.B1(n_4006),
.B2(n_4007),
.Y(n_16622)
);

INVx1_ASAP7_75t_L g16623 ( 
.A(n_16616),
.Y(n_16623)
);

BUFx2_ASAP7_75t_L g16624 ( 
.A(n_16611),
.Y(n_16624)
);

BUFx2_ASAP7_75t_L g16625 ( 
.A(n_16598),
.Y(n_16625)
);

INVx1_ASAP7_75t_L g16626 ( 
.A(n_16607),
.Y(n_16626)
);

OAI31xp33_ASAP7_75t_L g16627 ( 
.A1(n_16612),
.A2(n_16582),
.A3(n_16593),
.B(n_16574),
.Y(n_16627)
);

INVx1_ASAP7_75t_L g16628 ( 
.A(n_16610),
.Y(n_16628)
);

INVx1_ASAP7_75t_L g16629 ( 
.A(n_16606),
.Y(n_16629)
);

INVx2_ASAP7_75t_SL g16630 ( 
.A(n_16603),
.Y(n_16630)
);

OAI22xp33_ASAP7_75t_L g16631 ( 
.A1(n_16604),
.A2(n_16577),
.B1(n_16583),
.B2(n_16578),
.Y(n_16631)
);

INVx1_ASAP7_75t_L g16632 ( 
.A(n_16599),
.Y(n_16632)
);

OAI22xp5_ASAP7_75t_L g16633 ( 
.A1(n_16619),
.A2(n_4008),
.B1(n_4006),
.B2(n_4007),
.Y(n_16633)
);

OAI31xp33_ASAP7_75t_L g16634 ( 
.A1(n_16609),
.A2(n_4011),
.A3(n_4009),
.B(n_4010),
.Y(n_16634)
);

NAND2xp5_ASAP7_75t_L g16635 ( 
.A(n_16602),
.B(n_4012),
.Y(n_16635)
);

AOI22xp33_ASAP7_75t_SL g16636 ( 
.A1(n_16605),
.A2(n_4013),
.B1(n_4014),
.B2(n_4012),
.Y(n_16636)
);

NAND2xp5_ASAP7_75t_L g16637 ( 
.A(n_16600),
.B(n_4013),
.Y(n_16637)
);

AND2x2_ASAP7_75t_L g16638 ( 
.A(n_16601),
.B(n_4010),
.Y(n_16638)
);

NAND2xp5_ASAP7_75t_L g16639 ( 
.A(n_16621),
.B(n_4016),
.Y(n_16639)
);

INVx1_ASAP7_75t_L g16640 ( 
.A(n_16597),
.Y(n_16640)
);

AO22x2_ASAP7_75t_L g16641 ( 
.A1(n_16613),
.A2(n_16614),
.B1(n_16617),
.B2(n_16620),
.Y(n_16641)
);

A2O1A1Ixp33_ASAP7_75t_SL g16642 ( 
.A1(n_16608),
.A2(n_4018),
.B(n_4015),
.C(n_4017),
.Y(n_16642)
);

INVx1_ASAP7_75t_L g16643 ( 
.A(n_16622),
.Y(n_16643)
);

INVx1_ASAP7_75t_L g16644 ( 
.A(n_16615),
.Y(n_16644)
);

CKINVDCx20_ASAP7_75t_R g16645 ( 
.A(n_16632),
.Y(n_16645)
);

OAI22xp5_ASAP7_75t_L g16646 ( 
.A1(n_16639),
.A2(n_16618),
.B1(n_4020),
.B2(n_4017),
.Y(n_16646)
);

AOI22xp5_ASAP7_75t_L g16647 ( 
.A1(n_16625),
.A2(n_4021),
.B1(n_4019),
.B2(n_4020),
.Y(n_16647)
);

OAI22xp5_ASAP7_75t_L g16648 ( 
.A1(n_16628),
.A2(n_4023),
.B1(n_4021),
.B2(n_4022),
.Y(n_16648)
);

NAND3xp33_ASAP7_75t_L g16649 ( 
.A(n_16627),
.B(n_4022),
.C(n_4024),
.Y(n_16649)
);

NAND2xp5_ASAP7_75t_L g16650 ( 
.A(n_16626),
.B(n_16630),
.Y(n_16650)
);

INVx2_ASAP7_75t_L g16651 ( 
.A(n_16638),
.Y(n_16651)
);

INVx2_ASAP7_75t_L g16652 ( 
.A(n_16637),
.Y(n_16652)
);

OAI21xp5_ASAP7_75t_L g16653 ( 
.A1(n_16640),
.A2(n_4024),
.B(n_4025),
.Y(n_16653)
);

INVx1_ASAP7_75t_L g16654 ( 
.A(n_16641),
.Y(n_16654)
);

INVx2_ASAP7_75t_SL g16655 ( 
.A(n_16641),
.Y(n_16655)
);

OAI21xp33_ASAP7_75t_L g16656 ( 
.A1(n_16629),
.A2(n_4025),
.B(n_4026),
.Y(n_16656)
);

XOR2x1_ASAP7_75t_L g16657 ( 
.A(n_16644),
.B(n_4027),
.Y(n_16657)
);

OAI21xp5_ASAP7_75t_SL g16658 ( 
.A1(n_16623),
.A2(n_4026),
.B(n_4027),
.Y(n_16658)
);

NAND3xp33_ASAP7_75t_L g16659 ( 
.A(n_16624),
.B(n_4028),
.C(n_4029),
.Y(n_16659)
);

CKINVDCx20_ASAP7_75t_R g16660 ( 
.A(n_16645),
.Y(n_16660)
);

BUFx4f_ASAP7_75t_SL g16661 ( 
.A(n_16655),
.Y(n_16661)
);

OAI22xp5_ASAP7_75t_L g16662 ( 
.A1(n_16650),
.A2(n_16643),
.B1(n_16631),
.B2(n_16642),
.Y(n_16662)
);

INVx1_ASAP7_75t_L g16663 ( 
.A(n_16654),
.Y(n_16663)
);

AOI22xp5_ASAP7_75t_L g16664 ( 
.A1(n_16651),
.A2(n_16633),
.B1(n_16636),
.B2(n_16634),
.Y(n_16664)
);

HB1xp67_ASAP7_75t_L g16665 ( 
.A(n_16652),
.Y(n_16665)
);

OAI22xp33_ASAP7_75t_SL g16666 ( 
.A1(n_16646),
.A2(n_16635),
.B1(n_4030),
.B2(n_4028),
.Y(n_16666)
);

AOI22x1_ASAP7_75t_L g16667 ( 
.A1(n_16657),
.A2(n_4031),
.B1(n_4029),
.B2(n_4030),
.Y(n_16667)
);

OAI22x1_ASAP7_75t_L g16668 ( 
.A1(n_16649),
.A2(n_4033),
.B1(n_4031),
.B2(n_4032),
.Y(n_16668)
);

OAI21xp5_ASAP7_75t_L g16669 ( 
.A1(n_16663),
.A2(n_16658),
.B(n_16653),
.Y(n_16669)
);

OA21x2_ASAP7_75t_L g16670 ( 
.A1(n_16662),
.A2(n_16659),
.B(n_16656),
.Y(n_16670)
);

OR2x2_ASAP7_75t_L g16671 ( 
.A(n_16665),
.B(n_16648),
.Y(n_16671)
);

OR2x2_ASAP7_75t_L g16672 ( 
.A(n_16664),
.B(n_16647),
.Y(n_16672)
);

INVx1_ASAP7_75t_L g16673 ( 
.A(n_16661),
.Y(n_16673)
);

AND2x2_ASAP7_75t_L g16674 ( 
.A(n_16660),
.B(n_4032),
.Y(n_16674)
);

AO21x2_ASAP7_75t_L g16675 ( 
.A1(n_16666),
.A2(n_4042),
.B(n_4033),
.Y(n_16675)
);

OAI21xp5_ASAP7_75t_SL g16676 ( 
.A1(n_16673),
.A2(n_16668),
.B(n_16667),
.Y(n_16676)
);

XNOR2x1_ASAP7_75t_L g16677 ( 
.A(n_16672),
.B(n_4034),
.Y(n_16677)
);

AOI22xp5_ASAP7_75t_L g16678 ( 
.A1(n_16675),
.A2(n_4037),
.B1(n_4034),
.B2(n_4035),
.Y(n_16678)
);

NAND2xp5_ASAP7_75t_L g16679 ( 
.A(n_16669),
.B(n_4035),
.Y(n_16679)
);

AOI21xp5_ASAP7_75t_L g16680 ( 
.A1(n_16676),
.A2(n_16671),
.B(n_16670),
.Y(n_16680)
);

OAI21xp5_ASAP7_75t_SL g16681 ( 
.A1(n_16678),
.A2(n_16674),
.B(n_4037),
.Y(n_16681)
);

AOI22xp33_ASAP7_75t_L g16682 ( 
.A1(n_16680),
.A2(n_16677),
.B1(n_16679),
.B2(n_4040),
.Y(n_16682)
);

OR2x6_ASAP7_75t_L g16683 ( 
.A(n_16682),
.B(n_16681),
.Y(n_16683)
);

AOI322xp5_ASAP7_75t_L g16684 ( 
.A1(n_16683),
.A2(n_4043),
.A3(n_4042),
.B1(n_4040),
.B2(n_4038),
.C1(n_4039),
.C2(n_4041),
.Y(n_16684)
);

INVx2_ASAP7_75t_L g16685 ( 
.A(n_16684),
.Y(n_16685)
);

OAI22xp5_ASAP7_75t_SL g16686 ( 
.A1(n_16685),
.A2(n_4041),
.B1(n_4038),
.B2(n_4039),
.Y(n_16686)
);

AOI22xp5_ASAP7_75t_L g16687 ( 
.A1(n_16686),
.A2(n_4045),
.B1(n_4043),
.B2(n_4044),
.Y(n_16687)
);

AOI211xp5_ASAP7_75t_L g16688 ( 
.A1(n_16687),
.A2(n_4047),
.B(n_4045),
.C(n_4046),
.Y(n_16688)
);


endmodule