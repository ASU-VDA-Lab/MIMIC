module fake_jpeg_594_n_533 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_533);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_533;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_18),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_51),
.Y(n_157)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_23),
.B(n_17),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_54),
.B(n_67),
.Y(n_115)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_60),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_17),
.B1(n_16),
.B2(n_2),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_61),
.A2(n_50),
.B1(n_26),
.B2(n_47),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_66),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_21),
.B(n_16),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_30),
.B(n_16),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_68),
.B(n_70),
.Y(n_124)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_21),
.B(n_0),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_37),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_72),
.B(n_38),
.Y(n_129)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_75),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_77),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_80),
.Y(n_150)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g121 ( 
.A(n_83),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_84),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_24),
.B(n_0),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_38),
.Y(n_128)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_94),
.Y(n_154)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_97),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_38),
.Y(n_135)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_32),
.Y(n_100)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

AND2x4_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_68),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_104),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_88),
.A2(n_33),
.B1(n_32),
.B2(n_42),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_110),
.A2(n_83),
.B1(n_77),
.B2(n_75),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_91),
.A2(n_33),
.B1(n_32),
.B2(n_44),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_122),
.A2(n_153),
.B1(n_28),
.B2(n_26),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_128),
.B(n_129),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_67),
.B(n_70),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_134),
.B(n_138),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_135),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_54),
.B(n_45),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

AO22x2_ASAP7_75t_L g140 ( 
.A1(n_76),
.A2(n_89),
.B1(n_97),
.B2(n_78),
.Y(n_140)
);

AND2x4_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_86),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_76),
.B(n_50),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_145),
.B(n_159),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_89),
.A2(n_33),
.B1(n_38),
.B2(n_39),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_148),
.A2(n_39),
.B1(n_85),
.B2(n_79),
.Y(n_201)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_78),
.B(n_36),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_85),
.B(n_28),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_117),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_164),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_165),
.B(n_180),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_166),
.A2(n_179),
.B1(n_187),
.B2(n_201),
.Y(n_236)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_167),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_118),
.Y(n_171)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_171),
.Y(n_264)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_109),
.Y(n_173)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_173),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_124),
.A2(n_115),
.B1(n_122),
.B2(n_128),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_175),
.A2(n_218),
.B1(n_142),
.B2(n_141),
.Y(n_229)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_109),
.Y(n_176)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_176),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_177),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_106),
.Y(n_178)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_178),
.Y(n_275)
);

INVx11_ASAP7_75t_L g179 ( 
.A(n_117),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_159),
.Y(n_180)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_181),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_183),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_184),
.Y(n_243)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_116),
.Y(n_185)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_185),
.Y(n_248)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_125),
.Y(n_186)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_186),
.Y(n_250)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_127),
.Y(n_188)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_188),
.Y(n_252)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_103),
.Y(n_189)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_189),
.Y(n_256)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_120),
.Y(n_190)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_190),
.Y(n_257)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_191),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_106),
.Y(n_192)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_192),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_126),
.Y(n_193)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_193),
.Y(n_274)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_157),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_197),
.Y(n_234)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_124),
.A2(n_31),
.B(n_34),
.C(n_47),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_196),
.A2(n_0),
.B(n_1),
.Y(n_253)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_157),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_155),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_198),
.B(n_199),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_145),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_133),
.Y(n_200)
);

INVx13_ASAP7_75t_L g266 ( 
.A(n_200),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_135),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_208),
.Y(n_227)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_119),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_203),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_204),
.A2(n_217),
.B1(n_223),
.B2(n_3),
.Y(n_261)
);

BUFx8_ASAP7_75t_L g205 ( 
.A(n_140),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_131),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_154),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_102),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_115),
.B(n_114),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_211),
.Y(n_228)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_161),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_136),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_213),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_144),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_107),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_214),
.B(n_216),
.Y(n_255)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_130),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_147),
.A2(n_110),
.B1(n_112),
.B2(n_42),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_104),
.A2(n_64),
.B1(n_62),
.B2(n_60),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_121),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_219),
.B(n_220),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_126),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_104),
.B(n_39),
.Y(n_221)
);

MAJx2_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_27),
.C(n_39),
.Y(n_249)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_132),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_222),
.A2(n_219),
.B1(n_174),
.B2(n_182),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_111),
.A2(n_59),
.B1(n_42),
.B2(n_45),
.Y(n_223)
);

AOI32xp33_ASAP7_75t_L g224 ( 
.A1(n_184),
.A2(n_108),
.A3(n_158),
.B1(n_149),
.B2(n_148),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_224),
.B(n_181),
.Y(n_283)
);

OA21x2_ASAP7_75t_L g226 ( 
.A1(n_187),
.A2(n_121),
.B(n_48),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_226),
.B(n_259),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_229),
.A2(n_233),
.B1(n_247),
.B2(n_273),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_164),
.A2(n_123),
.B1(n_162),
.B2(n_163),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_205),
.A2(n_142),
.B1(n_141),
.B2(n_113),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_235),
.A2(n_245),
.B1(n_267),
.B2(n_269),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_48),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_238),
.B(n_239),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_168),
.B(n_36),
.C(n_31),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_168),
.B(n_163),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_240),
.B(n_249),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_205),
.A2(n_113),
.B1(n_162),
.B2(n_34),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_217),
.A2(n_39),
.B1(n_27),
.B2(n_2),
.Y(n_247)
);

INVxp67_ASAP7_75t_SL g282 ( 
.A(n_251),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_253),
.B(n_12),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_187),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_254),
.A2(n_265),
.B1(n_14),
.B2(n_267),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_221),
.B(n_3),
.C(n_4),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_215),
.B(n_3),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_260),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_261),
.A2(n_186),
.B1(n_189),
.B2(n_179),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_187),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_174),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_209),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_269)
);

OAI32xp33_ASAP7_75t_L g270 ( 
.A1(n_194),
.A2(n_8),
.A3(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_10),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_201),
.A2(n_196),
.B1(n_172),
.B2(n_220),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_276),
.B(n_279),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_234),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_277),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_253),
.A2(n_169),
.B(n_208),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_278),
.A2(n_283),
.B(n_290),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_255),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_228),
.B(n_198),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_281),
.B(n_288),
.Y(n_331)
);

OA21x2_ASAP7_75t_L g284 ( 
.A1(n_245),
.A2(n_197),
.B(n_195),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_284),
.Y(n_362)
);

CKINVDCx14_ASAP7_75t_R g357 ( 
.A(n_285),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_246),
.A2(n_178),
.B1(n_193),
.B2(n_192),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_287),
.A2(n_289),
.B1(n_314),
.B2(n_274),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_228),
.B(n_213),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_246),
.A2(n_176),
.B1(n_212),
.B2(n_173),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_237),
.A2(n_177),
.B(n_171),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_255),
.Y(n_292)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_292),
.Y(n_324)
);

OAI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_293),
.A2(n_225),
.B1(n_266),
.B2(n_282),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_242),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_294),
.B(n_295),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_243),
.B(n_12),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_242),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_296),
.B(n_312),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_248),
.B(n_13),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_298),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_227),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_300),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_244),
.A2(n_15),
.B(n_13),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_301),
.A2(n_272),
.B(n_263),
.Y(n_338)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_268),
.Y(n_302)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_302),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_236),
.A2(n_14),
.B1(n_229),
.B2(n_235),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_304),
.A2(n_286),
.B1(n_284),
.B2(n_301),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_257),
.B(n_14),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_305),
.Y(n_334)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_275),
.Y(n_306)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_306),
.Y(n_340)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_268),
.Y(n_307)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_307),
.Y(n_348)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_275),
.Y(n_308)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_308),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_234),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_309),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_241),
.A2(n_273),
.B(n_244),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_310),
.A2(n_264),
.B(n_262),
.Y(n_342)
);

INVxp33_ASAP7_75t_L g311 ( 
.A(n_244),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_311),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_240),
.B(n_14),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_313),
.B(n_276),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_233),
.A2(n_226),
.B1(n_227),
.B2(n_247),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_239),
.B(n_238),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_315),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_234),
.Y(n_316)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_316),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_260),
.B(n_270),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_317),
.B(n_318),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_249),
.B(n_259),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_269),
.B(n_226),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_319),
.B(n_320),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_272),
.B(n_263),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_252),
.Y(n_321)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_321),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_230),
.B(n_232),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_322),
.Y(n_345)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_271),
.Y(n_323)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_323),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_299),
.B(n_258),
.C(n_250),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_326),
.B(n_353),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_299),
.B(n_256),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_327),
.B(n_336),
.Y(n_374)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_332),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_318),
.B(n_231),
.Y(n_336)
);

CKINVDCx14_ASAP7_75t_R g391 ( 
.A(n_338),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_320),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_341),
.B(n_355),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_342),
.A2(n_343),
.B(n_346),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_310),
.A2(n_264),
.B(n_262),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_344),
.A2(n_347),
.B1(n_284),
.B2(n_292),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_294),
.A2(n_225),
.B(n_266),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_280),
.A2(n_314),
.B1(n_279),
.B2(n_319),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_351),
.A2(n_354),
.B1(n_359),
.B2(n_284),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_291),
.B(n_297),
.C(n_312),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_281),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_304),
.A2(n_280),
.B1(n_296),
.B2(n_286),
.Y(n_359)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_321),
.Y(n_365)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_365),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_362),
.A2(n_277),
.B1(n_316),
.B2(n_309),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_366),
.A2(n_379),
.B1(n_383),
.B2(n_384),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_346),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_368),
.B(n_376),
.Y(n_409)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_356),
.Y(n_370)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_370),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_359),
.A2(n_307),
.B1(n_302),
.B2(n_317),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_371),
.A2(n_335),
.B1(n_324),
.B2(n_348),
.Y(n_405)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_356),
.Y(n_372)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_372),
.Y(n_413)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_365),
.Y(n_375)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_375),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_331),
.Y(n_376)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_364),
.Y(n_378)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_378),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_330),
.A2(n_278),
.B(n_290),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_380),
.A2(n_352),
.B(n_335),
.Y(n_429)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_364),
.Y(n_381)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_381),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_331),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_382),
.B(n_388),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_347),
.A2(n_303),
.B1(n_288),
.B2(n_291),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_345),
.B(n_297),
.Y(n_385)
);

CKINVDCx14_ASAP7_75t_R g404 ( 
.A(n_385),
.Y(n_404)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_339),
.Y(n_386)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_386),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_351),
.A2(n_303),
.B1(n_287),
.B2(n_293),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_387),
.A2(n_394),
.B1(n_397),
.B2(n_400),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_358),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_360),
.Y(n_389)
);

CKINVDCx14_ASAP7_75t_R g430 ( 
.A(n_389),
.Y(n_430)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_339),
.Y(n_390)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_390),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_345),
.B(n_328),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_393),
.Y(n_406)
);

AOI22x1_ASAP7_75t_L g394 ( 
.A1(n_362),
.A2(n_303),
.B1(n_323),
.B2(n_306),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_361),
.Y(n_395)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_395),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_360),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_396),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_362),
.A2(n_289),
.B1(n_308),
.B2(n_355),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_348),
.Y(n_398)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_398),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_334),
.B(n_329),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_399),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_329),
.B(n_333),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_373),
.B(n_327),
.C(n_353),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_401),
.B(n_363),
.C(n_376),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_405),
.A2(n_420),
.B1(n_424),
.B2(n_426),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_373),
.B(n_374),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_410),
.B(n_412),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_389),
.A2(n_341),
.B1(n_324),
.B2(n_337),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_411),
.B(n_416),
.Y(n_441)
);

XNOR2x1_ASAP7_75t_SL g412 ( 
.A(n_384),
.B(n_337),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_396),
.A2(n_325),
.B1(n_342),
.B2(n_333),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_374),
.B(n_336),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_417),
.B(n_378),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_371),
.B(n_326),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_419),
.B(n_369),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_391),
.A2(n_330),
.B1(n_361),
.B2(n_325),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_379),
.A2(n_357),
.B1(n_354),
.B2(n_343),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_377),
.A2(n_338),
.B(n_349),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_425),
.A2(n_377),
.B(n_380),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_392),
.A2(n_332),
.B1(n_354),
.B2(n_352),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_429),
.A2(n_372),
.B(n_375),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_418),
.B(n_388),
.Y(n_432)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_432),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_406),
.B(n_401),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_433),
.B(n_440),
.Y(n_464)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_431),
.Y(n_434)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_434),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_435),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_425),
.A2(n_368),
.B(n_394),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_437),
.Y(n_466)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_421),
.Y(n_438)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_438),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_439),
.B(n_417),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_404),
.B(n_357),
.Y(n_440)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_421),
.Y(n_442)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_442),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_410),
.B(n_395),
.C(n_367),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_443),
.B(n_447),
.C(n_439),
.Y(n_462)
);

NAND3xp33_ASAP7_75t_L g444 ( 
.A(n_408),
.B(n_382),
.C(n_367),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_444),
.A2(n_452),
.B1(n_453),
.B2(n_454),
.Y(n_460)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_403),
.Y(n_445)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_445),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_405),
.A2(n_392),
.B1(n_387),
.B2(n_397),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_446),
.A2(n_422),
.B1(n_416),
.B2(n_423),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_419),
.B(n_394),
.C(n_398),
.Y(n_447)
);

A2O1A1Ixp33_ASAP7_75t_SL g448 ( 
.A1(n_409),
.A2(n_392),
.B(n_390),
.C(n_386),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_448),
.A2(n_450),
.B(n_436),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_451),
.B(n_455),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_429),
.B(n_369),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_431),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g454 ( 
.A(n_402),
.Y(n_454)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_403),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_456),
.A2(n_457),
.B1(n_454),
.B2(n_423),
.Y(n_468)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_402),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_458),
.B(n_461),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_441),
.A2(n_430),
.B1(n_426),
.B2(n_420),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_459),
.A2(n_473),
.B1(n_466),
.B2(n_463),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_443),
.B(n_412),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_462),
.B(n_465),
.C(n_471),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_447),
.B(n_414),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_468),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_449),
.B(n_409),
.C(n_411),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_473),
.A2(n_450),
.B1(n_448),
.B2(n_453),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_449),
.B(n_415),
.C(n_381),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_475),
.B(n_457),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_441),
.A2(n_407),
.B1(n_428),
.B2(n_427),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_476),
.B(n_477),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_477),
.A2(n_448),
.B(n_407),
.Y(n_489)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_469),
.Y(n_480)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_480),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_459),
.A2(n_446),
.B1(n_435),
.B2(n_437),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_481),
.B(n_489),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_464),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_482),
.B(n_483),
.Y(n_504)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_484),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_463),
.A2(n_448),
.B(n_434),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_486),
.B(n_490),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_488),
.B(n_493),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_470),
.A2(n_428),
.B1(n_427),
.B2(n_451),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_474),
.A2(n_413),
.B1(n_415),
.B2(n_370),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_491),
.B(n_492),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_465),
.A2(n_455),
.B1(n_340),
.B2(n_350),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_460),
.A2(n_340),
.B1(n_350),
.B2(n_466),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_467),
.B(n_471),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_494),
.B(n_495),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_494),
.B(n_462),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_498),
.B(n_500),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_487),
.B(n_458),
.C(n_475),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_487),
.B(n_461),
.C(n_472),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_503),
.B(n_485),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_480),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_506),
.B(n_495),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_482),
.B(n_478),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_507),
.B(n_485),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_500),
.B(n_483),
.Y(n_509)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_509),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_503),
.B(n_479),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_510),
.A2(n_511),
.B(n_513),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_504),
.A2(n_496),
.B(n_505),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_514),
.A2(n_515),
.B(n_516),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_501),
.B(n_492),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_506),
.B(n_484),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_517),
.A2(n_502),
.B1(n_488),
.B2(n_493),
.Y(n_518)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_518),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_512),
.B(n_499),
.C(n_508),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_521),
.A2(n_522),
.B(n_517),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_516),
.B(n_499),
.C(n_501),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_524),
.B(n_525),
.Y(n_527)
);

OAI31xp33_ASAP7_75t_SL g525 ( 
.A1(n_520),
.A2(n_489),
.A3(n_490),
.B(n_486),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_526),
.B(n_521),
.Y(n_528)
);

A2O1A1O1Ixp25_ASAP7_75t_L g529 ( 
.A1(n_528),
.A2(n_523),
.B(n_522),
.C(n_519),
.D(n_497),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_529),
.B(n_527),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_530),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_531),
.B(n_481),
.C(n_491),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_472),
.Y(n_533)
);


endmodule