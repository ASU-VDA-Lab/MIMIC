module fake_jpeg_13552_n_61 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_61);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_61;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

OR2x2_ASAP7_75t_L g8 ( 
.A(n_7),
.B(n_0),
.Y(n_8)
);

INVx8_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_3),
.A2(n_7),
.B1(n_1),
.B2(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_21),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g19 ( 
.A1(n_17),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_19),
.A2(n_16),
.B1(n_20),
.B2(n_23),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVxp33_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_12),
.B(n_15),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_12),
.B(n_5),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_25),
.Y(n_28)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_8),
.B(n_14),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

AO22x2_ASAP7_75t_L g30 ( 
.A1(n_22),
.A2(n_10),
.B1(n_11),
.B2(n_17),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_30),
.A2(n_22),
.B1(n_34),
.B2(n_36),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_8),
.C(n_15),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_27),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_25),
.A2(n_24),
.B(n_11),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_36),
.B(n_30),
.Y(n_43)
);

AO22x1_ASAP7_75t_L g36 ( 
.A1(n_19),
.A2(n_10),
.B1(n_16),
.B2(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_33),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_18),
.B1(n_34),
.B2(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_41),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_47),
.B1(n_31),
.B2(n_42),
.Y(n_51)
);

FAx1_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_28),
.CI(n_30),
.CON(n_41),
.SN(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_29),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_42),
.B(n_45),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_40),
.B1(n_41),
.B2(n_44),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_29),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_50),
.B(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_53),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_50),
.B1(n_51),
.B2(n_48),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_56),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

FAx1_ASAP7_75t_SL g60 ( 
.A(n_59),
.B(n_54),
.CI(n_56),
.CON(n_60),
.SN(n_60)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_49),
.B(n_58),
.Y(n_61)
);


endmodule