module real_jpeg_21818_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_49;
wire n_10;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_9;
wire n_72;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_0),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_1),
.A2(n_4),
.B1(n_17),
.B2(n_18),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_1),
.Y(n_18)
);

OAI22xp33_ASAP7_75t_L g31 ( 
.A1(n_1),
.A2(n_6),
.B1(n_18),
.B2(n_29),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_1),
.A2(n_7),
.B1(n_18),
.B2(n_23),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_1),
.A2(n_23),
.B(n_29),
.C(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_2),
.A2(n_6),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_2),
.A2(n_7),
.B1(n_23),
.B2(n_28),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_2),
.B(n_39),
.Y(n_40)
);

AOI21xp33_ASAP7_75t_L g66 ( 
.A1(n_2),
.A2(n_6),
.B(n_7),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_3),
.A2(n_4),
.B1(n_17),
.B2(n_21),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_3),
.A2(n_7),
.B1(n_21),
.B2(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_3),
.A2(n_5),
.B1(n_21),
.B2(n_55),
.Y(n_54)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

O2A1O1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_4),
.A2(n_7),
.B(n_21),
.C(n_42),
.Y(n_41)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_7),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_7),
.B(n_16),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_61),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_10),
.B(n_60),
.Y(n_9)
);

INVxp67_ASAP7_75t_L g10 ( 
.A(n_11),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_46),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_12),
.B(n_46),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_24),
.B(n_33),
.C(n_44),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_13),
.B(n_24),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_13),
.A2(n_14),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_13),
.A2(n_14),
.B1(n_24),
.B2(n_25),
.Y(n_88)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_22),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_19),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_20),
.Y(n_19)
);

OAI21xp33_ASAP7_75t_L g42 ( 
.A1(n_17),
.A2(n_18),
.B(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_23),
.B(n_27),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_23),
.B(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_24),
.A2(n_25),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_24),
.B(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_24),
.A2(n_25),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_24),
.A2(n_25),
.B1(n_65),
.B2(n_82),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_25),
.B(n_36),
.C(n_69),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_27),
.B(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_28),
.B(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_33),
.A2(n_34),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_41),
.B2(n_43),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_36),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_35),
.A2(n_36),
.B1(n_68),
.B2(n_71),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_35),
.B(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2x1_ASAP7_75t_SL g59 ( 
.A(n_36),
.B(n_41),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_36),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_36),
.B(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_41),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_56),
.B2(n_57),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_84),
.B(n_89),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_72),
.B(n_83),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_67),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_65),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_68),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_80),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_76),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_86),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);


endmodule