module fake_ariane_3201_n_1488 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_332, n_294, n_197, n_176, n_34, n_172, n_347, n_183, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_349, n_346, n_214, n_348, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_327, n_77, n_372, n_15, n_23, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_267, n_335, n_350, n_291, n_344, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_333, n_221, n_321, n_86, n_361, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_118, n_121, n_353, n_22, n_241, n_29, n_357, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_351, n_39, n_359, n_155, n_127, n_1488);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_347;
input n_183;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_327;
input n_77;
input n_372;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_333;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_118;
input n_121;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_351;
input n_39;
input n_359;
input n_155;
input n_127;

output n_1488;

wire n_913;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_559;
wire n_495;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1314;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_611;
wire n_1295;
wire n_1013;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1396;
wire n_1230;
wire n_612;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1432;
wire n_1108;
wire n_851;
wire n_444;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_436;
wire n_669;
wire n_931;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1455;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_706;
wire n_1401;
wire n_1419;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1456;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_529;
wire n_502;
wire n_1467;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1371;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1218;
wire n_861;
wire n_1431;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1478;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_1466;
wire n_608;
wire n_1037;
wire n_1329;
wire n_1257;
wire n_1480;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_1352;
wire n_643;
wire n_1441;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_1450;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1438;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_467;
wire n_1422;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1440;
wire n_1370;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1444;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_1482;
wire n_1361;
wire n_1057;
wire n_978;
wire n_1011;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1458;
wire n_679;
wire n_663;
wire n_443;
wire n_1412;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_1452;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_1470;
wire n_671;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_1479;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1474;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_1434;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_363),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_247),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_140),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_56),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_34),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_192),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_46),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_74),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_327),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_158),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_48),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_238),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_26),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_182),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_345),
.Y(n_389)
);

CKINVDCx14_ASAP7_75t_R g390 ( 
.A(n_355),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_183),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_152),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_97),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_75),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_258),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_256),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_262),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_126),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_233),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_239),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_347),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_311),
.Y(n_402)
);

BUFx10_ASAP7_75t_L g403 ( 
.A(n_81),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_255),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_241),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_31),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_341),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_181),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_44),
.Y(n_409)
);

BUFx10_ASAP7_75t_L g410 ( 
.A(n_112),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_185),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_157),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_127),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_20),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_354),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_69),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_36),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_43),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_122),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_312),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_215),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_147),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_28),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_68),
.Y(n_424)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_42),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_100),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_362),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_359),
.Y(n_428)
);

BUFx10_ASAP7_75t_L g429 ( 
.A(n_320),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_344),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_252),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_33),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_95),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_149),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_213),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_348),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_370),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_304),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_3),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_361),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_10),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_191),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_136),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_356),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_23),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_138),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_186),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_336),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_260),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_87),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_220),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_334),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_236),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_67),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_318),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_174),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_364),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_130),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_107),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_176),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_42),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_177),
.Y(n_462)
);

CKINVDCx14_ASAP7_75t_R g463 ( 
.A(n_209),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_62),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_353),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_123),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_3),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_224),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_214),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_120),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_226),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_110),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_234),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_240),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_367),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_199),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_50),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_321),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_144),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_35),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_373),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_45),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_263),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_230),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_281),
.Y(n_485)
);

BUFx5_ASAP7_75t_L g486 ( 
.A(n_141),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g487 ( 
.A(n_246),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_268),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_43),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_78),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_61),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_328),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_124),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_13),
.Y(n_494)
);

HB1xp67_ASAP7_75t_SL g495 ( 
.A(n_128),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_47),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_205),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_227),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_235),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_194),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_217),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_88),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_131),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_48),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_64),
.Y(n_505)
);

CKINVDCx16_ASAP7_75t_R g506 ( 
.A(n_374),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_219),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_71),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_305),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_231),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_58),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_352),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_108),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_27),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_70),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_207),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_245),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_23),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_360),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_34),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_310),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_8),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_49),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_73),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_294),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_190),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_326),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_98),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_27),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_16),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_121),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_366),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_161),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_72),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_357),
.Y(n_535)
);

CKINVDCx16_ASAP7_75t_R g536 ( 
.A(n_365),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_317),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_6),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_165),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_175),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_119),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_270),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_31),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_115),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_1),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_349),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_346),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_358),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_18),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_83),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_153),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_52),
.Y(n_552)
);

BUFx10_ASAP7_75t_L g553 ( 
.A(n_168),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_267),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_278),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_342),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_21),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_164),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_193),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_295),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_271),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_111),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_313),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_116),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_7),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_173),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_11),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_28),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_376),
.Y(n_569)
);

BUFx2_ASAP7_75t_L g570 ( 
.A(n_417),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_440),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_520),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_448),
.Y(n_573)
);

BUFx8_ASAP7_75t_L g574 ( 
.A(n_544),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_425),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_403),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_482),
.A2(n_4),
.B1(n_0),
.B2(n_2),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_385),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_440),
.B(n_4),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_520),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_376),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_432),
.B(n_5),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_376),
.Y(n_583)
);

INVx5_ASAP7_75t_L g584 ( 
.A(n_403),
.Y(n_584)
);

INVx5_ASAP7_75t_L g585 ( 
.A(n_410),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_460),
.Y(n_586)
);

BUFx12f_ASAP7_75t_L g587 ( 
.A(n_410),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_460),
.Y(n_588)
);

BUFx12f_ASAP7_75t_L g589 ( 
.A(n_429),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_379),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_520),
.Y(n_591)
);

OAI22x1_ASAP7_75t_R g592 ( 
.A1(n_406),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_592)
);

OAI21x1_ASAP7_75t_L g593 ( 
.A1(n_411),
.A2(n_53),
.B(n_51),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_467),
.B(n_8),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_530),
.Y(n_595)
);

OAI21x1_ASAP7_75t_L g596 ( 
.A1(n_442),
.A2(n_55),
.B(n_54),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_409),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_472),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_530),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_429),
.Y(n_600)
);

OAI21x1_ASAP7_75t_L g601 ( 
.A1(n_469),
.A2(n_59),
.B(n_57),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_375),
.Y(n_602)
);

OAI22x1_ASAP7_75t_SL g603 ( 
.A1(n_518),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_470),
.B(n_9),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_553),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_418),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_414),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_439),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_447),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_530),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_423),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_441),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_472),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_445),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_377),
.B(n_12),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_472),
.Y(n_616)
);

BUFx8_ASAP7_75t_SL g617 ( 
.A(n_473),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_480),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_490),
.Y(n_619)
);

BUFx12f_ASAP7_75t_L g620 ( 
.A(n_553),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_461),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_489),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_381),
.B(n_12),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_387),
.B(n_13),
.Y(n_624)
);

CKINVDCx16_ASAP7_75t_R g625 ( 
.A(n_438),
.Y(n_625)
);

INVxp67_ASAP7_75t_L g626 ( 
.A(n_565),
.Y(n_626)
);

OAI22x1_ASAP7_75t_SL g627 ( 
.A1(n_494),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_504),
.Y(n_628)
);

BUFx12f_ASAP7_75t_L g629 ( 
.A(n_496),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_490),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_522),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_490),
.Y(n_632)
);

OAI22x1_ASAP7_75t_R g633 ( 
.A1(n_529),
.A2(n_17),
.B1(n_14),
.B2(n_15),
.Y(n_633)
);

INVx5_ASAP7_75t_L g634 ( 
.A(n_550),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_514),
.B(n_17),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_476),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_636)
);

BUFx12f_ASAP7_75t_L g637 ( 
.A(n_557),
.Y(n_637)
);

CKINVDCx16_ASAP7_75t_R g638 ( 
.A(n_487),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_538),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_550),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_477),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_550),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_543),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_545),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_380),
.B(n_19),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_567),
.Y(n_646)
);

BUFx8_ASAP7_75t_SL g647 ( 
.A(n_491),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_383),
.B(n_21),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_390),
.B(n_22),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_L g650 ( 
.A1(n_495),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_650)
);

AOI22x1_ASAP7_75t_SL g651 ( 
.A1(n_532),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_533),
.A2(n_32),
.B1(n_29),
.B2(n_30),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_386),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_549),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_568),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_384),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_398),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_388),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_506),
.A2(n_32),
.B1(n_29),
.B2(n_30),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_408),
.B(n_33),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_536),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_412),
.B(n_35),
.Y(n_662)
);

BUFx12f_ASAP7_75t_L g663 ( 
.A(n_561),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_465),
.Y(n_664)
);

BUFx12f_ASAP7_75t_L g665 ( 
.A(n_378),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_382),
.Y(n_666)
);

BUFx2_ASAP7_75t_L g667 ( 
.A(n_463),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_466),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_495),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_617),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_647),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_R g672 ( 
.A(n_602),
.B(n_391),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_569),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_609),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_R g675 ( 
.A(n_641),
.B(n_625),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_667),
.B(n_393),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_665),
.Y(n_677)
);

NAND2xp33_ASAP7_75t_R g678 ( 
.A(n_606),
.B(n_392),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_638),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_629),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_R g681 ( 
.A(n_667),
.B(n_395),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_584),
.B(n_389),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_569),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_637),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_569),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_587),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_589),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_581),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_590),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_620),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_574),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_661),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_574),
.Y(n_693)
);

OA21x2_ASAP7_75t_L g694 ( 
.A1(n_615),
.A2(n_407),
.B(n_394),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_653),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_669),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_607),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_666),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_R g699 ( 
.A(n_606),
.B(n_396),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_573),
.B(n_466),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_666),
.Y(n_701)
);

CKINVDCx20_ASAP7_75t_R g702 ( 
.A(n_576),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_611),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_663),
.Y(n_704)
);

INVx4_ASAP7_75t_L g705 ( 
.A(n_634),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_584),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_584),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_585),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_585),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_585),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_612),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_581),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_605),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_597),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_605),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_605),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_608),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_621),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_646),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_R g720 ( 
.A(n_631),
.B(n_399),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_581),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_664),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_649),
.A2(n_579),
.B1(n_570),
.B2(n_668),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_R g724 ( 
.A(n_600),
.B(n_400),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_616),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_664),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_614),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_570),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_583),
.Y(n_729)
);

BUFx2_ASAP7_75t_L g730 ( 
.A(n_668),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_583),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_616),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_657),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_578),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_632),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_632),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_660),
.B(n_662),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_571),
.B(n_548),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_619),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_618),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_654),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_583),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_619),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_622),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_630),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_630),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_640),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_586),
.Y(n_748)
);

CKINVDCx20_ASAP7_75t_R g749 ( 
.A(n_588),
.Y(n_749)
);

BUFx2_ASAP7_75t_L g750 ( 
.A(n_626),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_628),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_640),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_642),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_651),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_598),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_639),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_725),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_689),
.Y(n_758)
);

AO221x1_ASAP7_75t_L g759 ( 
.A1(n_714),
.A2(n_575),
.B1(n_650),
.B2(n_592),
.C(n_633),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_725),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_698),
.B(n_701),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_673),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_697),
.Y(n_763)
);

NOR3xp33_ASAP7_75t_L g764 ( 
.A(n_714),
.B(n_604),
.C(n_645),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_683),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_725),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_685),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_688),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_681),
.B(n_660),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_737),
.B(n_662),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_676),
.B(n_656),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_730),
.B(n_635),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_703),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_700),
.B(n_582),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_712),
.Y(n_775)
);

BUFx6f_ASAP7_75t_SL g776 ( 
.A(n_700),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_735),
.B(n_658),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_741),
.B(n_750),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_736),
.B(n_634),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_711),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_727),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_748),
.B(n_634),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_696),
.B(n_582),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_748),
.B(n_642),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_738),
.B(n_635),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_721),
.Y(n_786)
);

OR2x6_ASAP7_75t_L g787 ( 
.A(n_695),
.B(n_594),
.Y(n_787)
);

NOR2xp67_ASAP7_75t_L g788 ( 
.A(n_686),
.B(n_643),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_740),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_694),
.B(n_594),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_729),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_682),
.B(n_648),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_744),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_751),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_694),
.B(n_756),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_672),
.B(n_659),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_728),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_734),
.B(n_623),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_733),
.B(n_624),
.Y(n_799)
);

INVxp33_ASAP7_75t_L g800 ( 
.A(n_692),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_670),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_731),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_705),
.B(n_419),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_720),
.B(n_724),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_742),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_706),
.B(n_655),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_755),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_707),
.B(n_644),
.Y(n_808)
);

BUFx2_ASAP7_75t_L g809 ( 
.A(n_717),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_753),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_708),
.B(n_598),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_709),
.B(n_548),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_692),
.B(n_572),
.Y(n_813)
);

NOR2xp67_ASAP7_75t_L g814 ( 
.A(n_687),
.B(n_401),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_SL g815 ( 
.A(n_677),
.B(n_397),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_710),
.B(n_598),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_753),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_743),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_718),
.B(n_636),
.Y(n_819)
);

NOR3xp33_ASAP7_75t_L g820 ( 
.A(n_719),
.B(n_652),
.C(n_424),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_745),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_746),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_713),
.B(n_613),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_715),
.B(n_577),
.Y(n_824)
);

AOI221xp5_ASAP7_75t_L g825 ( 
.A1(n_723),
.A2(n_603),
.B1(n_627),
.B2(n_428),
.C(n_435),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_716),
.B(n_599),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_747),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_SL g828 ( 
.A(n_679),
.B(n_421),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_752),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_705),
.B(n_613),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_722),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_732),
.B(n_613),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_732),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_726),
.B(n_675),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_732),
.B(n_580),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_739),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_739),
.B(n_591),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_739),
.B(n_595),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_704),
.B(n_599),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_690),
.B(n_610),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_702),
.B(n_610),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_749),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_680),
.B(n_402),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_684),
.B(n_422),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_691),
.B(n_431),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_674),
.B(n_436),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_678),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_699),
.B(n_404),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_693),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_671),
.B(n_484),
.Y(n_850)
);

BUFx2_ASAP7_75t_L g851 ( 
.A(n_797),
.Y(n_851)
);

AND2x6_ASAP7_75t_SL g852 ( 
.A(n_846),
.B(n_778),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_761),
.B(n_507),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_758),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_757),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_820),
.A2(n_509),
.B1(n_451),
.B2(n_453),
.Y(n_856)
);

NAND3xp33_ASAP7_75t_L g857 ( 
.A(n_783),
.B(n_455),
.C(n_450),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_763),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_792),
.B(n_405),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_785),
.B(n_413),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_762),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_809),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_790),
.A2(n_459),
.B1(n_471),
.B2(n_456),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_765),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_790),
.A2(n_481),
.B1(n_483),
.B2(n_479),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_757),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_801),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_800),
.B(n_754),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_787),
.B(n_488),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_773),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_847),
.B(n_799),
.Y(n_871)
);

O2A1O1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_770),
.A2(n_501),
.B(n_510),
.C(n_493),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_SL g873 ( 
.A1(n_828),
.A2(n_515),
.B1(n_521),
.B2(n_511),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_780),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_777),
.A2(n_596),
.B(n_593),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_781),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_767),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_776),
.Y(n_878)
);

INVx1_ASAP7_75t_SL g879 ( 
.A(n_842),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_789),
.Y(n_880)
);

BUFx6f_ASAP7_75t_SL g881 ( 
.A(n_849),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_799),
.B(n_415),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_L g883 ( 
.A1(n_764),
.A2(n_537),
.B1(n_542),
.B2(n_534),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_793),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_834),
.B(n_36),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_794),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_804),
.B(n_416),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_771),
.B(n_420),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_828),
.B(n_426),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_796),
.A2(n_547),
.B1(n_554),
.B2(n_546),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_806),
.B(n_427),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_768),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_787),
.B(n_556),
.Y(n_893)
);

OAI21xp33_ASAP7_75t_L g894 ( 
.A1(n_812),
.A2(n_566),
.B(n_562),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_795),
.B(n_430),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_775),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_776),
.Y(n_897)
);

OR2x6_ASAP7_75t_L g898 ( 
.A(n_831),
.B(n_516),
.Y(n_898)
);

BUFx4f_ASAP7_75t_L g899 ( 
.A(n_818),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_772),
.A2(n_528),
.B1(n_519),
.B2(n_434),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_795),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_769),
.B(n_433),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_810),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_817),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_807),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_786),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_R g907 ( 
.A(n_815),
.B(n_437),
.Y(n_907)
);

INVx5_ASAP7_75t_L g908 ( 
.A(n_787),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_819),
.A2(n_486),
.B1(n_444),
.B2(n_446),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_791),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_813),
.B(n_37),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_774),
.B(n_808),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_848),
.B(n_443),
.Y(n_913)
);

OR2x6_ASAP7_75t_L g914 ( 
.A(n_788),
.B(n_601),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_798),
.B(n_449),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_784),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_757),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_782),
.B(n_452),
.Y(n_918)
);

INVx5_ASAP7_75t_L g919 ( 
.A(n_760),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_802),
.Y(n_920)
);

CKINVDCx20_ASAP7_75t_R g921 ( 
.A(n_841),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_844),
.B(n_454),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_844),
.B(n_457),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_805),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_837),
.Y(n_925)
);

NOR2x2_ASAP7_75t_L g926 ( 
.A(n_759),
.B(n_37),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_L g927 ( 
.A1(n_825),
.A2(n_486),
.B1(n_462),
.B2(n_464),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_838),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_833),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_760),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_760),
.Y(n_931)
);

CKINVDCx20_ASAP7_75t_R g932 ( 
.A(n_850),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_803),
.A2(n_468),
.B(n_458),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_779),
.A2(n_475),
.B(n_474),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_840),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_815),
.B(n_38),
.Y(n_936)
);

NAND2x1p5_ASAP7_75t_L g937 ( 
.A(n_821),
.B(n_38),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_803),
.B(n_478),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_845),
.B(n_39),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_845),
.B(n_485),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_830),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_814),
.B(n_492),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_766),
.Y(n_943)
);

INVx5_ASAP7_75t_L g944 ( 
.A(n_766),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_836),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_822),
.B(n_497),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_839),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_836),
.B(n_498),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_827),
.Y(n_949)
);

INVxp67_ASAP7_75t_L g950 ( 
.A(n_829),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_811),
.B(n_816),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_853),
.B(n_824),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_871),
.B(n_843),
.Y(n_953)
);

INVx3_ASAP7_75t_L g954 ( 
.A(n_855),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_933),
.A2(n_835),
.B(n_823),
.C(n_826),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_950),
.B(n_832),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_859),
.B(n_499),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_854),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_879),
.B(n_500),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_939),
.B(n_502),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_891),
.A2(n_505),
.B1(n_508),
.B2(n_503),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_875),
.A2(n_513),
.B(n_512),
.Y(n_962)
);

OAI21xp33_ASAP7_75t_SL g963 ( 
.A1(n_883),
.A2(n_39),
.B(n_40),
.Y(n_963)
);

A2O1A1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_894),
.A2(n_523),
.B(n_524),
.C(n_517),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_860),
.A2(n_870),
.B(n_874),
.C(n_858),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_R g966 ( 
.A(n_867),
.B(n_525),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_935),
.B(n_526),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_899),
.B(n_527),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_855),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_861),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_SL g971 ( 
.A1(n_927),
.A2(n_932),
.B1(n_873),
.B2(n_856),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_949),
.B(n_531),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_901),
.A2(n_539),
.B(n_535),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_951),
.A2(n_541),
.B(n_540),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_895),
.A2(n_552),
.B(n_551),
.Y(n_975)
);

OA22x2_ASAP7_75t_L g976 ( 
.A1(n_868),
.A2(n_558),
.B1(n_559),
.B2(n_555),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_882),
.A2(n_563),
.B(n_560),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_R g978 ( 
.A(n_878),
.B(n_564),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_881),
.Y(n_979)
);

CKINVDCx20_ASAP7_75t_R g980 ( 
.A(n_921),
.Y(n_980)
);

INVx4_ASAP7_75t_L g981 ( 
.A(n_908),
.Y(n_981)
);

NAND2xp33_ASAP7_75t_L g982 ( 
.A(n_876),
.B(n_486),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_912),
.B(n_40),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_940),
.B(n_41),
.Y(n_984)
);

BUFx12f_ASAP7_75t_L g985 ( 
.A(n_851),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_922),
.A2(n_486),
.B(n_63),
.Y(n_986)
);

NOR2xp67_ASAP7_75t_L g987 ( 
.A(n_908),
.B(n_60),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_880),
.B(n_884),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_923),
.A2(n_938),
.B(n_918),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_R g990 ( 
.A(n_881),
.B(n_65),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_862),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_888),
.A2(n_941),
.B(n_948),
.Y(n_992)
);

OR2x6_ASAP7_75t_L g993 ( 
.A(n_897),
.B(n_41),
.Y(n_993)
);

BUFx8_ASAP7_75t_L g994 ( 
.A(n_936),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_886),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_863),
.A2(n_47),
.B1(n_486),
.B2(n_76),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_908),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_905),
.Y(n_998)
);

AOI21x1_ASAP7_75t_L g999 ( 
.A1(n_914),
.A2(n_486),
.B(n_66),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_945),
.A2(n_77),
.B(n_79),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_916),
.B(n_80),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_920),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_924),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_925),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_864),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_R g1006 ( 
.A(n_852),
.B(n_82),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_887),
.A2(n_84),
.B(n_85),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_877),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_902),
.A2(n_86),
.B(n_89),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_890),
.B(n_90),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_885),
.B(n_928),
.Y(n_1011)
);

A2O1A1Ixp33_ASAP7_75t_SL g1012 ( 
.A1(n_934),
.A2(n_91),
.B(n_92),
.C(n_93),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_892),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_865),
.B(n_94),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_866),
.A2(n_96),
.B(n_99),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_R g1016 ( 
.A(n_919),
.B(n_101),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_946),
.A2(n_102),
.B(n_103),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_942),
.A2(n_914),
.B(n_913),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_949),
.B(n_372),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_855),
.Y(n_1020)
);

A2O1A1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_915),
.A2(n_104),
.B(n_105),
.C(n_106),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_947),
.B(n_109),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_911),
.B(n_113),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_872),
.A2(n_114),
.B(n_117),
.C(n_118),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_898),
.B(n_125),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_896),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_906),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_889),
.A2(n_129),
.B1(n_132),
.B2(n_133),
.Y(n_1028)
);

INVx8_ASAP7_75t_L g1029 ( 
.A(n_985),
.Y(n_1029)
);

INVx2_ASAP7_75t_SL g1030 ( 
.A(n_980),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_981),
.B(n_919),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_969),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_991),
.Y(n_1033)
);

AOI22x1_ASAP7_75t_L g1034 ( 
.A1(n_989),
.A2(n_937),
.B1(n_929),
.B2(n_866),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_958),
.Y(n_1035)
);

INVx6_ASAP7_75t_L g1036 ( 
.A(n_994),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_969),
.Y(n_1037)
);

AO21x2_ASAP7_75t_L g1038 ( 
.A1(n_1018),
.A2(n_904),
.B(n_903),
.Y(n_1038)
);

AO21x2_ASAP7_75t_L g1039 ( 
.A1(n_992),
.A2(n_857),
.B(n_910),
.Y(n_1039)
);

INVx4_ASAP7_75t_L g1040 ( 
.A(n_981),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_982),
.A2(n_917),
.B(n_943),
.Y(n_1041)
);

BUFx10_ASAP7_75t_L g1042 ( 
.A(n_979),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_983),
.A2(n_909),
.B(n_917),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_997),
.B(n_919),
.Y(n_1044)
);

BUFx8_ASAP7_75t_SL g1045 ( 
.A(n_993),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_1002),
.Y(n_1046)
);

INVxp67_ASAP7_75t_SL g1047 ( 
.A(n_969),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_952),
.B(n_907),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_966),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_998),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_1015),
.A2(n_900),
.B(n_944),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_999),
.A2(n_944),
.B(n_943),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_994),
.Y(n_1053)
);

BUFx12f_ASAP7_75t_L g1054 ( 
.A(n_993),
.Y(n_1054)
);

AO21x2_ASAP7_75t_L g1055 ( 
.A1(n_1001),
.A2(n_893),
.B(n_869),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_1020),
.Y(n_1056)
);

NAND2x1p5_ASAP7_75t_L g1057 ( 
.A(n_1020),
.B(n_930),
.Y(n_1057)
);

CKINVDCx12_ASAP7_75t_R g1058 ( 
.A(n_971),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_1020),
.Y(n_1059)
);

OA21x2_ASAP7_75t_L g1060 ( 
.A1(n_1009),
.A2(n_893),
.B(n_869),
.Y(n_1060)
);

CKINVDCx20_ASAP7_75t_R g1061 ( 
.A(n_978),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_1016),
.Y(n_1062)
);

BUFx12f_ASAP7_75t_L g1063 ( 
.A(n_990),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_1004),
.B(n_931),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_954),
.Y(n_1065)
);

OAI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_1011),
.A2(n_898),
.B1(n_944),
.B2(n_943),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_988),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_986),
.A2(n_134),
.B(n_135),
.Y(n_1068)
);

INVxp33_ASAP7_75t_L g1069 ( 
.A(n_959),
.Y(n_1069)
);

AO21x2_ASAP7_75t_L g1070 ( 
.A1(n_1023),
.A2(n_926),
.B(n_137),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1003),
.Y(n_1071)
);

INVx5_ASAP7_75t_L g1072 ( 
.A(n_954),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_967),
.B(n_139),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_970),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1013),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_953),
.B(n_142),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1026),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_1005),
.Y(n_1078)
);

NAND2x1p5_ASAP7_75t_L g1079 ( 
.A(n_987),
.B(n_143),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1027),
.Y(n_1080)
);

INVx5_ASAP7_75t_L g1081 ( 
.A(n_1008),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_965),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_1022),
.Y(n_1083)
);

OA21x2_ASAP7_75t_L g1084 ( 
.A1(n_962),
.A2(n_145),
.B(n_146),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_1000),
.A2(n_148),
.B(n_150),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_976),
.Y(n_1086)
);

AO21x2_ASAP7_75t_L g1087 ( 
.A1(n_955),
.A2(n_1014),
.B(n_975),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_1007),
.A2(n_151),
.B(n_154),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1010),
.Y(n_1089)
);

NAND2x1p5_ASAP7_75t_L g1090 ( 
.A(n_968),
.B(n_155),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_957),
.A2(n_156),
.B(n_159),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_996),
.Y(n_1092)
);

CKINVDCx6p67_ASAP7_75t_R g1093 ( 
.A(n_972),
.Y(n_1093)
);

BUFx12f_ASAP7_75t_L g1094 ( 
.A(n_1006),
.Y(n_1094)
);

CKINVDCx16_ASAP7_75t_R g1095 ( 
.A(n_1025),
.Y(n_1095)
);

AOI21x1_ASAP7_75t_L g1096 ( 
.A1(n_1082),
.A2(n_974),
.B(n_977),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1046),
.Y(n_1097)
);

INVx1_ASAP7_75t_SL g1098 ( 
.A(n_1033),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1069),
.B(n_956),
.Y(n_1099)
);

BUFx8_ASAP7_75t_SL g1100 ( 
.A(n_1045),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1075),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1048),
.A2(n_984),
.B1(n_960),
.B2(n_1019),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1075),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_1052),
.A2(n_1017),
.B(n_1028),
.Y(n_1104)
);

AOI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1058),
.A2(n_963),
.B1(n_961),
.B2(n_995),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_SL g1106 ( 
.A1(n_1095),
.A2(n_973),
.B1(n_1024),
.B2(n_1021),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_1029),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1035),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1077),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1035),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1092),
.A2(n_1070),
.B1(n_1067),
.B2(n_1086),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_1061),
.Y(n_1112)
);

NAND2xp33_ASAP7_75t_L g1113 ( 
.A(n_1073),
.B(n_964),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_1051),
.A2(n_1012),
.B(n_160),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1050),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1067),
.B(n_1062),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1050),
.Y(n_1117)
);

BUFx4f_ASAP7_75t_SL g1118 ( 
.A(n_1063),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1071),
.Y(n_1119)
);

AOI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1049),
.A2(n_162),
.B1(n_163),
.B2(n_166),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1077),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1080),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1068),
.A2(n_1088),
.B(n_1085),
.Y(n_1123)
);

OR2x6_ASAP7_75t_L g1124 ( 
.A(n_1029),
.B(n_167),
.Y(n_1124)
);

INVx2_ASAP7_75t_SL g1125 ( 
.A(n_1036),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_1036),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1034),
.A2(n_169),
.B(n_170),
.Y(n_1127)
);

AOI22xp33_ASAP7_75t_SL g1128 ( 
.A1(n_1070),
.A2(n_171),
.B1(n_172),
.B2(n_178),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_1056),
.Y(n_1129)
);

CKINVDCx11_ASAP7_75t_R g1130 ( 
.A(n_1042),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_SL g1131 ( 
.A1(n_1092),
.A2(n_179),
.B1(n_180),
.B2(n_184),
.Y(n_1131)
);

AO21x2_ASAP7_75t_L g1132 ( 
.A1(n_1038),
.A2(n_187),
.B(n_188),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1071),
.B(n_189),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1064),
.B(n_371),
.Y(n_1134)
);

NAND2x1p5_ASAP7_75t_L g1135 ( 
.A(n_1072),
.B(n_195),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1080),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1074),
.Y(n_1137)
);

INVx3_ASAP7_75t_L g1138 ( 
.A(n_1056),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1074),
.Y(n_1139)
);

AO21x1_ASAP7_75t_SL g1140 ( 
.A1(n_1082),
.A2(n_196),
.B(n_197),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_1030),
.Y(n_1141)
);

OA21x2_ASAP7_75t_L g1142 ( 
.A1(n_1089),
.A2(n_198),
.B(n_200),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1064),
.B(n_369),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_1056),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1078),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_1031),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1039),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_SL g1148 ( 
.A1(n_1054),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_1044),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1078),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1078),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_1044),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1055),
.A2(n_204),
.B1(n_206),
.B2(n_208),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1039),
.Y(n_1154)
);

NOR3xp33_ASAP7_75t_SL g1155 ( 
.A(n_1112),
.B(n_1102),
.C(n_1130),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_1100),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_1149),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_1118),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1099),
.B(n_1093),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1097),
.Y(n_1160)
);

AO31x2_ASAP7_75t_L g1161 ( 
.A1(n_1147),
.A2(n_1089),
.A3(n_1083),
.B(n_1076),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_1116),
.B(n_1066),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1101),
.Y(n_1163)
);

NAND3xp33_ASAP7_75t_SL g1164 ( 
.A(n_1105),
.B(n_1090),
.C(n_1043),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1149),
.B(n_1053),
.Y(n_1165)
);

BUFx10_ASAP7_75t_L g1166 ( 
.A(n_1124),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_SL g1167 ( 
.A(n_1107),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1103),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1098),
.B(n_1081),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1108),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1109),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_1152),
.B(n_1081),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1110),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1109),
.B(n_1081),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1152),
.B(n_1031),
.Y(n_1175)
);

NOR3xp33_ASAP7_75t_SL g1176 ( 
.A(n_1130),
.B(n_1091),
.C(n_1042),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1121),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1115),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1111),
.A2(n_1055),
.B1(n_1094),
.B2(n_1087),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_SL g1180 ( 
.A1(n_1133),
.A2(n_1041),
.B(n_1047),
.C(n_1037),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1121),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1122),
.Y(n_1182)
);

AOI21xp33_ASAP7_75t_L g1183 ( 
.A1(n_1113),
.A2(n_1087),
.B(n_1034),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_1146),
.B(n_1059),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1111),
.A2(n_1040),
.B1(n_1065),
.B2(n_1072),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1141),
.B(n_1032),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1146),
.B(n_1072),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_1117),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1143),
.B(n_1032),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_1119),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1122),
.B(n_1037),
.Y(n_1191)
);

AO31x2_ASAP7_75t_L g1192 ( 
.A1(n_1147),
.A2(n_1084),
.A3(n_1060),
.B(n_1079),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1124),
.B(n_1057),
.Y(n_1193)
);

OR2x2_ASAP7_75t_L g1194 ( 
.A(n_1136),
.B(n_1040),
.Y(n_1194)
);

OR2x2_ASAP7_75t_L g1195 ( 
.A(n_1136),
.B(n_1060),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1139),
.Y(n_1196)
);

NAND2xp33_ASAP7_75t_SL g1197 ( 
.A(n_1107),
.B(n_1084),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1137),
.Y(n_1198)
);

NAND2xp33_ASAP7_75t_SL g1199 ( 
.A(n_1125),
.B(n_210),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_1100),
.Y(n_1200)
);

INVx4_ASAP7_75t_L g1201 ( 
.A(n_1118),
.Y(n_1201)
);

NAND2xp33_ASAP7_75t_R g1202 ( 
.A(n_1124),
.B(n_211),
.Y(n_1202)
);

NOR3xp33_ASAP7_75t_SL g1203 ( 
.A(n_1134),
.B(n_212),
.C(n_216),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1139),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_1126),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1145),
.Y(n_1206)
);

NOR3xp33_ASAP7_75t_SL g1207 ( 
.A(n_1150),
.B(n_218),
.C(n_221),
.Y(n_1207)
);

NAND2xp33_ASAP7_75t_R g1208 ( 
.A(n_1142),
.B(n_222),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1138),
.B(n_223),
.Y(n_1209)
);

OR2x2_ASAP7_75t_L g1210 ( 
.A(n_1151),
.B(n_225),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1129),
.Y(n_1211)
);

BUFx10_ASAP7_75t_L g1212 ( 
.A(n_1129),
.Y(n_1212)
);

O2A1O1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_1113),
.A2(n_228),
.B(n_229),
.C(n_232),
.Y(n_1213)
);

NOR3xp33_ASAP7_75t_SL g1214 ( 
.A(n_1140),
.B(n_237),
.C(n_242),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1138),
.B(n_243),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1129),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1129),
.Y(n_1217)
);

NAND2xp33_ASAP7_75t_R g1218 ( 
.A(n_1142),
.B(n_244),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1106),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_1219)
);

AO31x2_ASAP7_75t_L g1220 ( 
.A1(n_1154),
.A2(n_251),
.A3(n_253),
.B(n_254),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1144),
.Y(n_1221)
);

INVxp67_ASAP7_75t_L g1222 ( 
.A(n_1144),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1135),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_1153),
.B(n_257),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1128),
.B(n_1106),
.Y(n_1225)
);

INVx4_ASAP7_75t_L g1226 ( 
.A(n_1166),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1188),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1170),
.B(n_1128),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1195),
.Y(n_1229)
);

AND2x4_ASAP7_75t_SL g1230 ( 
.A(n_1166),
.B(n_1153),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_1190),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_1212),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1173),
.B(n_1131),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1178),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1171),
.Y(n_1235)
);

INVxp67_ASAP7_75t_L g1236 ( 
.A(n_1159),
.Y(n_1236)
);

OR2x2_ASAP7_75t_L g1237 ( 
.A(n_1225),
.B(n_1132),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1177),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1163),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1181),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1157),
.B(n_1148),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1221),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1198),
.B(n_1131),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1224),
.A2(n_1148),
.B1(n_1142),
.B2(n_1132),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1191),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_1211),
.Y(n_1246)
);

INVx2_ASAP7_75t_SL g1247 ( 
.A(n_1212),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1182),
.B(n_1135),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1161),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1168),
.B(n_1096),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1196),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_1223),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1216),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1186),
.B(n_1120),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1162),
.B(n_1127),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_1217),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1160),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1206),
.B(n_1104),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1204),
.Y(n_1259)
);

INVxp67_ASAP7_75t_L g1260 ( 
.A(n_1169),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1161),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1194),
.B(n_1123),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1174),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1224),
.B(n_1189),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1161),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1222),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_1165),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1155),
.B(n_1114),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1220),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1179),
.B(n_259),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1209),
.B(n_261),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1215),
.B(n_1219),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1192),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1192),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1192),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1220),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1220),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1187),
.Y(n_1278)
);

OR2x2_ASAP7_75t_L g1279 ( 
.A(n_1164),
.B(n_264),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1210),
.Y(n_1280)
);

NOR2x1_ASAP7_75t_L g1281 ( 
.A(n_1205),
.B(n_265),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1180),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1193),
.B(n_266),
.Y(n_1283)
);

NAND2xp33_ASAP7_75t_SL g1284 ( 
.A(n_1202),
.B(n_269),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1185),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1214),
.B(n_272),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1172),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1172),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1184),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1183),
.B(n_273),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1267),
.B(n_1175),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1231),
.B(n_1176),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1231),
.B(n_1201),
.Y(n_1293)
);

BUFx3_ASAP7_75t_L g1294 ( 
.A(n_1267),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1227),
.Y(n_1295)
);

HB1xp67_ASAP7_75t_L g1296 ( 
.A(n_1250),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1264),
.B(n_1175),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1263),
.B(n_1184),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1284),
.A2(n_1199),
.B1(n_1197),
.B2(n_1187),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1264),
.B(n_1158),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1234),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1253),
.B(n_1201),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1242),
.B(n_1203),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1246),
.B(n_1156),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1253),
.B(n_1200),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1235),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1256),
.B(n_1207),
.Y(n_1307)
);

OR2x2_ASAP7_75t_L g1308 ( 
.A(n_1245),
.B(n_274),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1235),
.Y(n_1309)
);

OR2x2_ASAP7_75t_L g1310 ( 
.A(n_1257),
.B(n_275),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1256),
.B(n_1213),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1239),
.Y(n_1312)
);

OAI21xp33_ASAP7_75t_L g1313 ( 
.A1(n_1233),
.A2(n_1218),
.B(n_1208),
.Y(n_1313)
);

OR2x2_ASAP7_75t_L g1314 ( 
.A(n_1229),
.B(n_276),
.Y(n_1314)
);

INVx4_ASAP7_75t_L g1315 ( 
.A(n_1232),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1238),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1226),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1238),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_1229),
.B(n_277),
.Y(n_1319)
);

NAND3xp33_ASAP7_75t_L g1320 ( 
.A(n_1279),
.B(n_1167),
.C(n_280),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_SL g1321 ( 
.A1(n_1279),
.A2(n_279),
.B(n_282),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1250),
.Y(n_1322)
);

AND2x4_ASAP7_75t_L g1323 ( 
.A(n_1278),
.B(n_283),
.Y(n_1323)
);

NOR2x1_ASAP7_75t_L g1324 ( 
.A(n_1226),
.B(n_284),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_SL g1325 ( 
.A(n_1285),
.B(n_285),
.Y(n_1325)
);

AND2x4_ASAP7_75t_SL g1326 ( 
.A(n_1278),
.B(n_286),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1236),
.B(n_287),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1228),
.B(n_288),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1228),
.B(n_289),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_1260),
.B(n_290),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1289),
.B(n_291),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1266),
.B(n_292),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1233),
.B(n_293),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1289),
.B(n_1278),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1252),
.B(n_296),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1251),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1301),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1294),
.B(n_1243),
.Y(n_1338)
);

HB1xp67_ASAP7_75t_L g1339 ( 
.A(n_1296),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1296),
.B(n_1243),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1312),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1295),
.B(n_1252),
.Y(n_1342)
);

INVx1_ASAP7_75t_SL g1343 ( 
.A(n_1305),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1322),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_L g1345 ( 
.A(n_1292),
.B(n_1268),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1294),
.B(n_1262),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1334),
.B(n_1311),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1297),
.B(n_1258),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1336),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1306),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1302),
.B(n_1252),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1293),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1304),
.B(n_1226),
.Y(n_1353)
);

INVx5_ASAP7_75t_L g1354 ( 
.A(n_1335),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1325),
.A2(n_1284),
.B(n_1244),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1293),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1300),
.B(n_1302),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1291),
.B(n_1237),
.Y(n_1358)
);

OR2x2_ASAP7_75t_L g1359 ( 
.A(n_1298),
.B(n_1237),
.Y(n_1359)
);

INVx1_ASAP7_75t_SL g1360 ( 
.A(n_1327),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1303),
.B(n_1292),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1317),
.B(n_1241),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1306),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1315),
.B(n_1282),
.Y(n_1364)
);

INVxp67_ASAP7_75t_L g1365 ( 
.A(n_1332),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1315),
.B(n_1282),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1307),
.B(n_1268),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1349),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1347),
.B(n_1307),
.Y(n_1369)
);

O2A1O1Ixp5_ASAP7_75t_R g1370 ( 
.A1(n_1342),
.A2(n_1328),
.B(n_1329),
.C(n_1333),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1337),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1347),
.B(n_1232),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1365),
.A2(n_1313),
.B1(n_1328),
.B2(n_1329),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1339),
.Y(n_1374)
);

OAI33xp33_ASAP7_75t_L g1375 ( 
.A1(n_1341),
.A2(n_1333),
.A3(n_1330),
.B1(n_1320),
.B2(n_1308),
.B3(n_1314),
.Y(n_1375)
);

NAND2x2_ASAP7_75t_L g1376 ( 
.A(n_1356),
.B(n_1247),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1344),
.Y(n_1377)
);

OAI31xp67_ASAP7_75t_L g1378 ( 
.A1(n_1343),
.A2(n_1280),
.A3(n_1332),
.B(n_1321),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1340),
.B(n_1232),
.Y(n_1379)
);

INVx1_ASAP7_75t_SL g1380 ( 
.A(n_1361),
.Y(n_1380)
);

OAI33xp33_ASAP7_75t_L g1381 ( 
.A1(n_1362),
.A2(n_1319),
.A3(n_1254),
.B1(n_1325),
.B2(n_1310),
.B3(n_1255),
.Y(n_1381)
);

O2A1O1Ixp5_ASAP7_75t_R g1382 ( 
.A1(n_1345),
.A2(n_1286),
.B(n_1247),
.C(n_1324),
.Y(n_1382)
);

AOI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1355),
.A2(n_1230),
.B1(n_1272),
.B2(n_1281),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1361),
.A2(n_1270),
.B1(n_1272),
.B2(n_1230),
.Y(n_1384)
);

INVx1_ASAP7_75t_SL g1385 ( 
.A(n_1367),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1359),
.Y(n_1386)
);

NOR2xp67_ASAP7_75t_L g1387 ( 
.A(n_1354),
.B(n_1335),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1340),
.B(n_1358),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1345),
.B(n_1248),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1368),
.Y(n_1390)
);

AOI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1374),
.A2(n_1367),
.B(n_1353),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1382),
.A2(n_1360),
.B(n_1338),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1371),
.Y(n_1393)
);

XNOR2x1_ASAP7_75t_L g1394 ( 
.A(n_1373),
.B(n_1357),
.Y(n_1394)
);

INVxp67_ASAP7_75t_L g1395 ( 
.A(n_1370),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1378),
.A2(n_1354),
.B(n_1364),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1381),
.A2(n_1354),
.B(n_1364),
.Y(n_1397)
);

NOR3xp33_ASAP7_75t_L g1398 ( 
.A(n_1375),
.B(n_1366),
.C(n_1286),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1383),
.A2(n_1358),
.B1(n_1354),
.B2(n_1270),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1377),
.Y(n_1400)
);

INVxp67_ASAP7_75t_L g1401 ( 
.A(n_1369),
.Y(n_1401)
);

OAI21xp33_ASAP7_75t_L g1402 ( 
.A1(n_1380),
.A2(n_1346),
.B(n_1366),
.Y(n_1402)
);

AOI322xp5_ASAP7_75t_L g1403 ( 
.A1(n_1398),
.A2(n_1380),
.A3(n_1384),
.B1(n_1389),
.B2(n_1385),
.C1(n_1386),
.C2(n_1299),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1390),
.Y(n_1404)
);

OAI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1399),
.A2(n_1373),
.B1(n_1354),
.B2(n_1385),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1393),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1395),
.B(n_1388),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1400),
.B(n_1348),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1397),
.B(n_1348),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1396),
.A2(n_1387),
.B(n_1352),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_SL g1411 ( 
.A(n_1392),
.B(n_1356),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1394),
.B(n_1379),
.Y(n_1412)
);

INVx1_ASAP7_75t_SL g1413 ( 
.A(n_1402),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1401),
.A2(n_1280),
.B1(n_1277),
.B2(n_1248),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1391),
.B(n_1357),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1390),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_1407),
.Y(n_1417)
);

NOR3x1_ASAP7_75t_L g1418 ( 
.A(n_1411),
.B(n_1376),
.C(n_1288),
.Y(n_1418)
);

NOR3x1_ASAP7_75t_L g1419 ( 
.A(n_1409),
.B(n_1287),
.C(n_1351),
.Y(n_1419)
);

NOR2xp67_ASAP7_75t_L g1420 ( 
.A(n_1410),
.B(n_1372),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1412),
.B(n_1351),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1404),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1416),
.Y(n_1423)
);

AOI211xp5_ASAP7_75t_L g1424 ( 
.A1(n_1405),
.A2(n_1346),
.B(n_1290),
.C(n_1271),
.Y(n_1424)
);

A2O1A1Ixp33_ASAP7_75t_L g1425 ( 
.A1(n_1424),
.A2(n_1403),
.B(n_1413),
.C(n_1415),
.Y(n_1425)
);

AND4x1_ASAP7_75t_L g1426 ( 
.A(n_1418),
.B(n_1299),
.C(n_1408),
.D(n_1414),
.Y(n_1426)
);

OA22x2_ASAP7_75t_L g1427 ( 
.A1(n_1417),
.A2(n_1413),
.B1(n_1406),
.B2(n_1351),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1422),
.Y(n_1428)
);

OAI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1420),
.A2(n_1290),
.B(n_1323),
.Y(n_1429)
);

A2O1A1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1421),
.A2(n_1326),
.B(n_1271),
.C(n_1283),
.Y(n_1430)
);

AOI222xp33_ASAP7_75t_L g1431 ( 
.A1(n_1425),
.A2(n_1423),
.B1(n_1419),
.B2(n_1277),
.C1(n_1269),
.C2(n_1276),
.Y(n_1431)
);

AOI322xp5_ASAP7_75t_L g1432 ( 
.A1(n_1426),
.A2(n_1428),
.A3(n_1427),
.B1(n_1430),
.B2(n_1429),
.C1(n_1283),
.C2(n_1276),
.Y(n_1432)
);

AOI211xp5_ASAP7_75t_L g1433 ( 
.A1(n_1425),
.A2(n_1323),
.B(n_1331),
.C(n_1363),
.Y(n_1433)
);

AOI311xp33_ASAP7_75t_L g1434 ( 
.A1(n_1425),
.A2(n_1261),
.A3(n_1249),
.B(n_1265),
.C(n_1326),
.Y(n_1434)
);

AOI221x1_ASAP7_75t_L g1435 ( 
.A1(n_1425),
.A2(n_1350),
.B1(n_1249),
.B2(n_1261),
.C(n_1309),
.Y(n_1435)
);

AOI221x1_ASAP7_75t_L g1436 ( 
.A1(n_1425),
.A2(n_1350),
.B1(n_1318),
.B2(n_1309),
.C(n_1274),
.Y(n_1436)
);

NOR2x1_ASAP7_75t_L g1437 ( 
.A(n_1434),
.B(n_1273),
.Y(n_1437)
);

NOR2x1_ASAP7_75t_L g1438 ( 
.A(n_1432),
.B(n_1273),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1433),
.Y(n_1439)
);

NOR2x1_ASAP7_75t_L g1440 ( 
.A(n_1435),
.B(n_1274),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1431),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1436),
.B(n_1318),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1433),
.Y(n_1443)
);

CKINVDCx20_ASAP7_75t_R g1444 ( 
.A(n_1434),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1444),
.B(n_297),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1439),
.B(n_1316),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1443),
.B(n_1441),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1437),
.B(n_1259),
.Y(n_1448)
);

NOR2xp67_ASAP7_75t_SL g1449 ( 
.A(n_1442),
.B(n_298),
.Y(n_1449)
);

AND2x4_ASAP7_75t_SL g1450 ( 
.A(n_1438),
.B(n_1259),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1440),
.Y(n_1451)
);

INVx1_ASAP7_75t_SL g1452 ( 
.A(n_1447),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1445),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1451),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1446),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1449),
.B(n_299),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1448),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1450),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1454),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1453),
.A2(n_1251),
.B1(n_1240),
.B2(n_1275),
.Y(n_1460)
);

INVx1_ASAP7_75t_SL g1461 ( 
.A(n_1452),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1456),
.Y(n_1462)
);

OAI22xp33_ASAP7_75t_R g1463 ( 
.A1(n_1457),
.A2(n_1275),
.B1(n_1240),
.B2(n_302),
.Y(n_1463)
);

INVxp67_ASAP7_75t_SL g1464 ( 
.A(n_1455),
.Y(n_1464)
);

INVxp67_ASAP7_75t_L g1465 ( 
.A(n_1458),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1458),
.B(n_300),
.Y(n_1466)
);

INVxp67_ASAP7_75t_SL g1467 ( 
.A(n_1454),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1454),
.Y(n_1468)
);

OAI31xp33_ASAP7_75t_SL g1469 ( 
.A1(n_1461),
.A2(n_1464),
.A3(n_1459),
.B(n_1468),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1463),
.A2(n_1462),
.B1(n_1460),
.B2(n_1466),
.Y(n_1470)
);

OAI31xp33_ASAP7_75t_L g1471 ( 
.A1(n_1465),
.A2(n_368),
.A3(n_303),
.B(n_306),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_SL g1472 ( 
.A1(n_1461),
.A2(n_301),
.B1(n_307),
.B2(n_308),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1459),
.Y(n_1473)
);

AOI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1463),
.A2(n_309),
.B1(n_314),
.B2(n_315),
.Y(n_1474)
);

AOI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1463),
.A2(n_316),
.B1(n_319),
.B2(n_322),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1467),
.Y(n_1476)
);

OAI22x1_ASAP7_75t_L g1477 ( 
.A1(n_1473),
.A2(n_323),
.B1(n_324),
.B2(n_325),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1469),
.B(n_329),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1476),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1472),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1474),
.A2(n_330),
.B1(n_331),
.B2(n_332),
.Y(n_1481)
);

OAI22x1_ASAP7_75t_L g1482 ( 
.A1(n_1479),
.A2(n_1475),
.B1(n_1470),
.B2(n_1471),
.Y(n_1482)
);

XNOR2xp5_ASAP7_75t_L g1483 ( 
.A(n_1478),
.B(n_333),
.Y(n_1483)
);

AOI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1480),
.A2(n_335),
.B1(n_337),
.B2(n_338),
.Y(n_1484)
);

AOI21xp33_ASAP7_75t_L g1485 ( 
.A1(n_1483),
.A2(n_1477),
.B(n_1481),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1485),
.A2(n_1482),
.B1(n_1484),
.B2(n_340),
.Y(n_1486)
);

OR2x6_ASAP7_75t_L g1487 ( 
.A(n_1486),
.B(n_339),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1487),
.A2(n_343),
.B1(n_350),
.B2(n_351),
.Y(n_1488)
);


endmodule