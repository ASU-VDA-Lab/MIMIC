module fake_aes_3176_n_27 (n_1, n_2, n_4, n_3, n_5, n_0, n_27);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_27;
wire n_20;
wire n_23;
wire n_8;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_6;
wire n_7;
CKINVDCx20_ASAP7_75t_R g6 ( .A(n_5), .Y(n_6) );
CKINVDCx5p33_ASAP7_75t_R g7 ( .A(n_2), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_1), .Y(n_8) );
NAND2xp5_ASAP7_75t_L g9 ( .A(n_1), .B(n_0), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_2), .Y(n_10) );
NOR2x1_ASAP7_75t_L g11 ( .A(n_8), .B(n_0), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_7), .B(n_0), .Y(n_12) );
O2A1O1Ixp33_ASAP7_75t_SL g13 ( .A1(n_8), .A2(n_1), .B(n_2), .C(n_3), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_11), .Y(n_14) );
NOR2xp33_ASAP7_75t_L g15 ( .A(n_12), .B(n_7), .Y(n_15) );
NOR3xp33_ASAP7_75t_SL g16 ( .A(n_13), .B(n_10), .C(n_9), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_15), .B(n_9), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_15), .B(n_6), .Y(n_18) );
AOI21xp5_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_14), .B(n_16), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_18), .B(n_6), .Y(n_20) );
AOI21xp5_ASAP7_75t_L g21 ( .A1(n_19), .A2(n_3), .B(n_4), .Y(n_21) );
OAI221xp5_ASAP7_75t_L g22 ( .A1(n_20), .A2(n_3), .B1(n_4), .B2(n_5), .C(n_18), .Y(n_22) );
INVx1_ASAP7_75t_SL g23 ( .A(n_21), .Y(n_23) );
CKINVDCx14_ASAP7_75t_R g24 ( .A(n_22), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_24), .B(n_4), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_23), .Y(n_26) );
AOI22xp33_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_5), .B1(n_23), .B2(n_25), .Y(n_27) );
endmodule