module real_jpeg_32223_n_15 (n_123, n_8, n_116, n_0, n_2, n_114, n_10, n_9, n_12, n_6, n_121, n_11, n_14, n_120, n_7, n_117, n_3, n_119, n_5, n_4, n_115, n_122, n_1, n_118, n_13, n_113, n_15);

input n_123;
input n_8;
input n_116;
input n_0;
input n_2;
input n_114;
input n_10;
input n_9;
input n_12;
input n_6;
input n_121;
input n_11;
input n_14;
input n_120;
input n_7;
input n_117;
input n_3;
input n_119;
input n_5;
input n_4;
input n_115;
input n_122;
input n_1;
input n_118;
input n_13;
input n_113;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx1_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

AOI221xp5_ASAP7_75t_L g43 ( 
.A1(n_1),
.A2(n_8),
.B1(n_44),
.B2(n_51),
.C(n_53),
.Y(n_43)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_2),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_2),
.B(n_86),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_3),
.A2(n_17),
.B1(n_18),
.B2(n_24),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_4),
.B(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_4),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_5),
.B(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_7),
.Y(n_82)
);

AOI322xp5_ASAP7_75t_L g105 ( 
.A1(n_7),
.A2(n_78),
.A3(n_80),
.B1(n_84),
.B2(n_106),
.C1(n_108),
.C2(n_123),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_8),
.B(n_44),
.C(n_51),
.Y(n_56)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_9),
.B(n_28),
.Y(n_111)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_10),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_11),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_11),
.B(n_91),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_13),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_13),
.B(n_96),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_29),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_25),
.Y(n_15)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_20),
.Y(n_18)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_20),
.B(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_31),
.B(n_111),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI31xp33_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_72),
.A3(n_94),
.B(n_101),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_66),
.C(n_67),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_57),
.B(n_65),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_43),
.B1(n_55),
.B2(n_56),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_45),
.B(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_115),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_64),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_64),
.Y(n_65)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NOR3xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_83),
.C(n_90),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_73),
.A2(n_102),
.B(n_105),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NOR3xp33_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_90),
.C(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_119),
.Y(n_80)
);

OA21x2_ASAP7_75t_SL g102 ( 
.A1(n_83),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_89),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

NOR2x1_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_100),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_113),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_114),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_116),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_117),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_118),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_120),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_121),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_122),
.Y(n_97)
);


endmodule