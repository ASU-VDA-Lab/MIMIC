module fake_jpeg_2588_n_189 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_189);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_189;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_26),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx24_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_67),
.Y(n_70)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_73),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_66),
.A2(n_45),
.B1(n_48),
.B2(n_56),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_59),
.B1(n_67),
.B2(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_63),
.B(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_79),
.Y(n_89)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_50),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_48),
.B(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_81),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_61),
.Y(n_81)
);

CKINVDCx9p33_ASAP7_75t_R g82 ( 
.A(n_78),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_82),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_83),
.A2(n_49),
.B1(n_3),
.B2(n_4),
.Y(n_106)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_79),
.A2(n_55),
.B1(n_60),
.B2(n_54),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_85),
.A2(n_90),
.B1(n_10),
.B2(n_11),
.Y(n_118)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_55),
.B1(n_64),
.B2(n_53),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_74),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_3),
.Y(n_108)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_51),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_94),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_1),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_1),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_2),
.Y(n_99)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_107),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_70),
.B1(n_80),
.B2(n_58),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_103),
.A2(n_83),
.B1(n_86),
.B2(n_28),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_88),
.A2(n_58),
.B(n_49),
.Y(n_105)
);

NAND2x1_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_115),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_2),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_108),
.B(n_111),
.Y(n_119)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_4),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_6),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_112),
.B(n_117),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_97),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_98),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_115)
);

AND2x6_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_25),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_118),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_113),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_127),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_103),
.A2(n_109),
.B1(n_102),
.B2(n_106),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_141)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_23),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_22),
.C(n_27),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_113),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_136),
.Y(n_146)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_116),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_133),
.B(n_135),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_106),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_101),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_42),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_105),
.A2(n_10),
.B(n_11),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_19),
.B(n_20),
.Y(n_147)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_119),
.B(n_13),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_147),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_17),
.C(n_18),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_154),
.C(n_155),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_153),
.Y(n_165)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_149),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_128),
.B(n_29),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_151),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_30),
.Y(n_153)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_32),
.C(n_34),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_134),
.B(n_122),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_134),
.B(n_36),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_129),
.Y(n_166)
);

FAx1_ASAP7_75t_SL g158 ( 
.A(n_154),
.B(n_121),
.CI(n_124),
.CON(n_158),
.SN(n_158)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_166),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_146),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_159),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_151),
.B(n_139),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_163),
.A2(n_161),
.B(n_167),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_170),
.Y(n_177)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_140),
.C(n_143),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_173),
.Y(n_179)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_172),
.A2(n_157),
.B(n_165),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_160),
.A2(n_143),
.B1(n_124),
.B2(n_132),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_148),
.Y(n_175)
);

XNOR2x1_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_157),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_171),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_175),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_180),
.A2(n_181),
.B1(n_174),
.B2(n_178),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_177),
.Y(n_183)
);

INVx11_ASAP7_75t_L g184 ( 
.A(n_183),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_184),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_185),
.A2(n_184),
.B(n_179),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_168),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_39),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_40),
.Y(n_189)
);


endmodule