module real_aes_6240_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_183;
wire n_312;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_0), .B(n_105), .C(n_106), .Y(n_104) );
INVx1_ASAP7_75t_L g121 ( .A(n_0), .Y(n_121) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_1), .A2(n_148), .B(n_153), .C(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g260 ( .A(n_2), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_3), .A2(n_143), .B(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_4), .B(n_220), .Y(n_468) );
AOI21xp33_ASAP7_75t_L g221 ( .A1(n_5), .A2(n_143), .B(n_222), .Y(n_221) );
AND2x6_ASAP7_75t_L g148 ( .A(n_6), .B(n_149), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_7), .A2(n_142), .B(n_150), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_8), .B(n_40), .Y(n_110) );
INVx1_ASAP7_75t_L g557 ( .A(n_9), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_10), .B(n_192), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_11), .B(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g227 ( .A(n_12), .Y(n_227) );
INVx1_ASAP7_75t_L g140 ( .A(n_13), .Y(n_140) );
INVx1_ASAP7_75t_L g160 ( .A(n_14), .Y(n_160) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_15), .A2(n_161), .B(n_175), .C(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_16), .B(n_220), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_17), .B(n_177), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_18), .B(n_143), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_19), .B(n_481), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_20), .A2(n_208), .B(n_234), .C(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_21), .B(n_220), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_22), .B(n_192), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g156 ( .A1(n_23), .A2(n_157), .B(n_159), .C(n_161), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_24), .B(n_192), .Y(n_454) );
CKINVDCx16_ASAP7_75t_R g485 ( .A(n_25), .Y(n_485) );
INVx1_ASAP7_75t_L g453 ( .A(n_26), .Y(n_453) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_27), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_28), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_29), .B(n_192), .Y(n_261) );
INVx1_ASAP7_75t_L g478 ( .A(n_30), .Y(n_478) );
INVx1_ASAP7_75t_L g239 ( .A(n_31), .Y(n_239) );
INVx2_ASAP7_75t_L g146 ( .A(n_32), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_33), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g465 ( .A1(n_34), .A2(n_208), .B(n_228), .C(n_466), .Y(n_465) );
INVxp67_ASAP7_75t_L g479 ( .A(n_35), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_L g171 ( .A1(n_36), .A2(n_148), .B(n_153), .C(n_172), .Y(n_171) );
A2O1A1Ixp33_ASAP7_75t_L g451 ( .A1(n_37), .A2(n_153), .B(n_452), .C(n_457), .Y(n_451) );
CKINVDCx14_ASAP7_75t_R g464 ( .A(n_38), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g124 ( .A1(n_39), .A2(n_67), .B1(n_125), .B2(n_126), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_39), .Y(n_125) );
INVx1_ASAP7_75t_L g237 ( .A(n_41), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g555 ( .A1(n_42), .A2(n_179), .B(n_225), .C(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_43), .B(n_192), .Y(n_191) );
OAI22xp5_ASAP7_75t_SL g716 ( .A1(n_44), .A2(n_84), .B1(n_717), .B2(n_718), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_44), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_45), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_46), .Y(n_475) );
INVx1_ASAP7_75t_L g523 ( .A(n_47), .Y(n_523) );
CKINVDCx16_ASAP7_75t_R g240 ( .A(n_48), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_49), .B(n_143), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_50), .A2(n_153), .B1(n_234), .B2(n_236), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_51), .Y(n_183) );
CKINVDCx16_ASAP7_75t_R g257 ( .A(n_52), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_53), .A2(n_225), .B(n_226), .C(n_228), .Y(n_224) );
CKINVDCx14_ASAP7_75t_R g554 ( .A(n_54), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_55), .Y(n_196) );
INVx1_ASAP7_75t_L g223 ( .A(n_56), .Y(n_223) );
AOI222xp33_ASAP7_75t_SL g123 ( .A1(n_57), .A2(n_124), .B1(n_127), .B2(n_707), .C1(n_708), .C2(n_709), .Y(n_123) );
INVx1_ASAP7_75t_L g149 ( .A(n_58), .Y(n_149) );
INVx1_ASAP7_75t_L g139 ( .A(n_59), .Y(n_139) );
INVx1_ASAP7_75t_SL g467 ( .A(n_60), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_61), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_62), .B(n_220), .Y(n_527) );
INVx1_ASAP7_75t_L g488 ( .A(n_63), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_SL g247 ( .A1(n_64), .A2(n_177), .B(n_228), .C(n_248), .Y(n_247) );
INVxp67_ASAP7_75t_L g249 ( .A(n_65), .Y(n_249) );
INVx1_ASAP7_75t_L g108 ( .A(n_66), .Y(n_108) );
INVx1_ASAP7_75t_L g126 ( .A(n_67), .Y(n_126) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_68), .A2(n_143), .B(n_553), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_69), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_70), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_71), .A2(n_143), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g187 ( .A(n_72), .Y(n_187) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_73), .A2(n_102), .B1(n_111), .B2(n_720), .Y(n_101) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_74), .A2(n_142), .B(n_474), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g450 ( .A(n_75), .Y(n_450) );
INVx1_ASAP7_75t_L g515 ( .A(n_76), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g189 ( .A1(n_77), .A2(n_148), .B(n_153), .C(n_190), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_78), .A2(n_143), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g518 ( .A(n_79), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_80), .B(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g137 ( .A(n_81), .Y(n_137) );
INVx1_ASAP7_75t_L g507 ( .A(n_82), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_83), .B(n_177), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_84), .Y(n_717) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_85), .A2(n_148), .B(n_153), .C(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g105 ( .A(n_86), .Y(n_105) );
OR2x2_ASAP7_75t_L g118 ( .A(n_86), .B(n_119), .Y(n_118) );
OR2x2_ASAP7_75t_L g706 ( .A(n_86), .B(n_120), .Y(n_706) );
A2O1A1Ixp33_ASAP7_75t_L g486 ( .A1(n_87), .A2(n_153), .B(n_487), .C(n_491), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_88), .B(n_136), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g264 ( .A(n_89), .Y(n_264) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_90), .A2(n_148), .B(n_153), .C(n_205), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_91), .Y(n_213) );
INVx1_ASAP7_75t_L g246 ( .A(n_92), .Y(n_246) );
CKINVDCx16_ASAP7_75t_R g151 ( .A(n_93), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_94), .B(n_174), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_95), .B(n_165), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_96), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_97), .B(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_98), .A2(n_143), .B(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g526 ( .A(n_99), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_100), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_103), .Y(n_721) );
OR2x2_ASAP7_75t_SL g103 ( .A(n_104), .B(n_109), .Y(n_103) );
OR2x2_ASAP7_75t_L g439 ( .A(n_105), .B(n_120), .Y(n_439) );
NOR2x2_ASAP7_75t_L g711 ( .A(n_105), .B(n_119), .Y(n_711) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVxp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g120 ( .A(n_110), .B(n_121), .Y(n_120) );
AOI22x1_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_123), .B1(n_712), .B2(n_714), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_113), .B(n_116), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g713 ( .A(n_115), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_116), .A2(n_715), .B(n_719), .Y(n_714) );
NOR2xp33_ASAP7_75t_SL g116 ( .A(n_117), .B(n_122), .Y(n_116) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_118), .Y(n_719) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g707 ( .A(n_124), .Y(n_707) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_437), .B1(n_440), .B2(n_704), .Y(n_127) );
INVx2_ASAP7_75t_SL g128 ( .A(n_129), .Y(n_128) );
OAI22xp5_ASAP7_75t_SL g708 ( .A1(n_129), .A2(n_439), .B1(n_441), .B2(n_706), .Y(n_708) );
OR4x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_333), .C(n_392), .D(n_419), .Y(n_129) );
NAND3xp33_ASAP7_75t_SL g130 ( .A(n_131), .B(n_275), .C(n_300), .Y(n_130) );
O2A1O1Ixp33_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_198), .B(n_218), .C(n_251), .Y(n_131) );
AOI211xp5_ASAP7_75t_SL g423 ( .A1(n_132), .A2(n_424), .B(n_426), .C(n_429), .Y(n_423) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_167), .Y(n_132) );
INVx1_ASAP7_75t_L g298 ( .A(n_133), .Y(n_298) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OR2x2_ASAP7_75t_L g273 ( .A(n_134), .B(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g305 ( .A(n_134), .Y(n_305) );
AND2x2_ASAP7_75t_L g360 ( .A(n_134), .B(n_329), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_134), .B(n_216), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_134), .B(n_217), .Y(n_418) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g279 ( .A(n_135), .Y(n_279) );
AND2x2_ASAP7_75t_L g322 ( .A(n_135), .B(n_185), .Y(n_322) );
AND2x2_ASAP7_75t_L g340 ( .A(n_135), .B(n_217), .Y(n_340) );
OA21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_141), .B(n_164), .Y(n_135) );
INVx1_ASAP7_75t_L g197 ( .A(n_136), .Y(n_197) );
INVx2_ASAP7_75t_L g202 ( .A(n_136), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_L g449 ( .A1(n_136), .A2(n_188), .B(n_450), .C(n_451), .Y(n_449) );
OA21x2_ASAP7_75t_L g551 ( .A1(n_136), .A2(n_552), .B(n_558), .Y(n_551) );
AND2x2_ASAP7_75t_SL g136 ( .A(n_137), .B(n_138), .Y(n_136) );
AND2x2_ASAP7_75t_L g166 ( .A(n_137), .B(n_138), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
BUFx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_148), .Y(n_143) );
NAND2x1p5_ASAP7_75t_L g188 ( .A(n_144), .B(n_148), .Y(n_188) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
INVx1_ASAP7_75t_L g456 ( .A(n_145), .Y(n_456) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g154 ( .A(n_146), .Y(n_154) );
INVx1_ASAP7_75t_L g235 ( .A(n_146), .Y(n_235) );
INVx1_ASAP7_75t_L g155 ( .A(n_147), .Y(n_155) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_147), .Y(n_158) );
INVx3_ASAP7_75t_L g175 ( .A(n_147), .Y(n_175) );
INVx1_ASAP7_75t_L g177 ( .A(n_147), .Y(n_177) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_147), .Y(n_192) );
INVx4_ASAP7_75t_SL g163 ( .A(n_148), .Y(n_163) );
BUFx3_ASAP7_75t_L g457 ( .A(n_148), .Y(n_457) );
O2A1O1Ixp33_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_156), .C(n_163), .Y(n_150) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_152), .A2(n_163), .B(n_223), .C(n_224), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g245 ( .A1(n_152), .A2(n_163), .B(n_246), .C(n_247), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g463 ( .A1(n_152), .A2(n_163), .B(n_464), .C(n_465), .Y(n_463) );
O2A1O1Ixp33_ASAP7_75t_SL g474 ( .A1(n_152), .A2(n_163), .B(n_475), .C(n_476), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_SL g514 ( .A1(n_152), .A2(n_163), .B(n_515), .C(n_516), .Y(n_514) );
O2A1O1Ixp33_ASAP7_75t_SL g522 ( .A1(n_152), .A2(n_163), .B(n_523), .C(n_524), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_SL g553 ( .A1(n_152), .A2(n_163), .B(n_554), .C(n_555), .Y(n_553) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x6_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
BUFx3_ASAP7_75t_L g162 ( .A(n_154), .Y(n_162) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_154), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_157), .B(n_160), .Y(n_159) );
OAI22xp33_ASAP7_75t_L g477 ( .A1(n_157), .A2(n_174), .B1(n_478), .B2(n_479), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_157), .B(n_518), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_157), .B(n_526), .Y(n_525) );
INVx4_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
OAI22xp5_ASAP7_75t_SL g236 ( .A1(n_158), .A2(n_237), .B1(n_238), .B2(n_239), .Y(n_236) );
INVx2_ASAP7_75t_L g238 ( .A(n_158), .Y(n_238) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g179 ( .A(n_162), .Y(n_179) );
OAI22xp33_ASAP7_75t_L g232 ( .A1(n_163), .A2(n_188), .B1(n_233), .B2(n_240), .Y(n_232) );
INVx1_ASAP7_75t_L g491 ( .A(n_163), .Y(n_491) );
INVx4_ASAP7_75t_L g184 ( .A(n_165), .Y(n_184) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_165), .A2(n_244), .B(n_250), .Y(n_243) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_165), .Y(n_461) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g181 ( .A(n_166), .Y(n_181) );
INVx4_ASAP7_75t_L g272 ( .A(n_167), .Y(n_272) );
OAI21xp5_ASAP7_75t_L g327 ( .A1(n_167), .A2(n_328), .B(n_330), .Y(n_327) );
AND2x2_ASAP7_75t_L g408 ( .A(n_167), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_185), .Y(n_167) );
INVx1_ASAP7_75t_L g215 ( .A(n_168), .Y(n_215) );
AND2x2_ASAP7_75t_L g277 ( .A(n_168), .B(n_217), .Y(n_277) );
OR2x2_ASAP7_75t_L g306 ( .A(n_168), .B(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g320 ( .A(n_168), .Y(n_320) );
INVx3_ASAP7_75t_L g329 ( .A(n_168), .Y(n_329) );
AND2x2_ASAP7_75t_L g339 ( .A(n_168), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g372 ( .A(n_168), .B(n_278), .Y(n_372) );
AND2x2_ASAP7_75t_L g396 ( .A(n_168), .B(n_352), .Y(n_396) );
OR2x6_ASAP7_75t_L g168 ( .A(n_169), .B(n_182), .Y(n_168) );
AOI21xp5_ASAP7_75t_SL g169 ( .A1(n_170), .A2(n_171), .B(n_180), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_176), .B(n_178), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_L g259 ( .A1(n_174), .A2(n_260), .B(n_261), .C(n_262), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g452 ( .A1(n_174), .A2(n_453), .B(n_454), .C(n_455), .Y(n_452) );
INVx5_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_175), .B(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_175), .B(n_249), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_175), .B(n_557), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_178), .A2(n_191), .B(n_193), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g487 ( .A1(n_178), .A2(n_488), .B(n_489), .C(n_490), .Y(n_487) );
O2A1O1Ixp5_ASAP7_75t_L g506 ( .A1(n_178), .A2(n_489), .B(n_507), .C(n_508), .Y(n_506) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g194 ( .A(n_180), .Y(n_194) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_181), .A2(n_232), .B(n_241), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_181), .B(n_242), .Y(n_241) );
AO21x2_ASAP7_75t_L g255 ( .A1(n_181), .A2(n_256), .B(n_263), .Y(n_255) );
NOR2xp33_ASAP7_75t_SL g182 ( .A(n_183), .B(n_184), .Y(n_182) );
INVx3_ASAP7_75t_L g220 ( .A(n_184), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_184), .B(n_459), .Y(n_458) );
AO21x2_ASAP7_75t_L g483 ( .A1(n_184), .A2(n_484), .B(n_492), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_184), .B(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g217 ( .A(n_185), .Y(n_217) );
AND2x2_ASAP7_75t_L g432 ( .A(n_185), .B(n_274), .Y(n_432) );
AO21x2_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_194), .B(n_195), .Y(n_185) );
OAI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_189), .Y(n_186) );
OAI21xp5_ASAP7_75t_L g256 ( .A1(n_188), .A2(n_257), .B(n_258), .Y(n_256) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_188), .A2(n_485), .B(n_486), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g503 ( .A1(n_188), .A2(n_504), .B(n_505), .Y(n_503) );
INVx4_ASAP7_75t_L g208 ( .A(n_192), .Y(n_208) );
INVx2_ASAP7_75t_L g225 ( .A(n_192), .Y(n_225) );
INVx1_ASAP7_75t_L g472 ( .A(n_194), .Y(n_472) );
AO21x2_ASAP7_75t_L g496 ( .A1(n_194), .A2(n_497), .B(n_498), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_197), .B(n_213), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_197), .B(n_264), .Y(n_263) );
AO21x2_ASAP7_75t_L g502 ( .A1(n_197), .A2(n_503), .B(n_509), .Y(n_502) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_214), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_200), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g352 ( .A(n_200), .B(n_340), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_200), .B(n_329), .Y(n_414) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g274 ( .A(n_201), .Y(n_274) );
AND2x2_ASAP7_75t_L g278 ( .A(n_201), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g319 ( .A(n_201), .B(n_320), .Y(n_319) );
AO21x2_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B(n_212), .Y(n_201) );
INVx1_ASAP7_75t_L g481 ( .A(n_202), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_202), .B(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_204), .B(n_211), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_209), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_208), .B(n_467), .Y(n_466) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx3_ASAP7_75t_L g228 ( .A(n_210), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_214), .B(n_315), .Y(n_337) );
INVx1_ASAP7_75t_L g376 ( .A(n_214), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_214), .B(n_303), .Y(n_420) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
AND2x2_ASAP7_75t_L g283 ( .A(n_215), .B(n_278), .Y(n_283) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_217), .B(n_274), .Y(n_307) );
INVx1_ASAP7_75t_L g386 ( .A(n_217), .Y(n_386) );
AOI322xp5_ASAP7_75t_L g410 ( .A1(n_218), .A2(n_325), .A3(n_385), .B1(n_411), .B2(n_413), .C1(n_415), .C2(n_417), .Y(n_410) );
AND2x2_ASAP7_75t_SL g218 ( .A(n_219), .B(n_230), .Y(n_218) );
AND2x2_ASAP7_75t_L g265 ( .A(n_219), .B(n_243), .Y(n_265) );
INVx1_ASAP7_75t_SL g268 ( .A(n_219), .Y(n_268) );
AND2x2_ASAP7_75t_L g270 ( .A(n_219), .B(n_231), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_219), .B(n_287), .Y(n_293) );
INVx2_ASAP7_75t_L g312 ( .A(n_219), .Y(n_312) );
AND2x2_ASAP7_75t_L g325 ( .A(n_219), .B(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g363 ( .A(n_219), .B(n_287), .Y(n_363) );
BUFx2_ASAP7_75t_L g380 ( .A(n_219), .Y(n_380) );
AND2x2_ASAP7_75t_L g394 ( .A(n_219), .B(n_254), .Y(n_394) );
OA21x2_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_229), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_230), .B(n_282), .Y(n_309) );
AND2x2_ASAP7_75t_L g436 ( .A(n_230), .B(n_312), .Y(n_436) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_243), .Y(n_230) );
OR2x2_ASAP7_75t_L g281 ( .A(n_231), .B(n_282), .Y(n_281) );
INVx3_ASAP7_75t_L g287 ( .A(n_231), .Y(n_287) );
AND2x2_ASAP7_75t_L g332 ( .A(n_231), .B(n_255), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_231), .B(n_380), .Y(n_379) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_231), .Y(n_416) );
INVx2_ASAP7_75t_L g262 ( .A(n_234), .Y(n_262) );
INVx3_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g489 ( .A(n_238), .Y(n_489) );
AND2x2_ASAP7_75t_L g267 ( .A(n_243), .B(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g289 ( .A(n_243), .Y(n_289) );
BUFx2_ASAP7_75t_L g295 ( .A(n_243), .Y(n_295) );
AND2x2_ASAP7_75t_L g314 ( .A(n_243), .B(n_287), .Y(n_314) );
INVx3_ASAP7_75t_L g326 ( .A(n_243), .Y(n_326) );
OR2x2_ASAP7_75t_L g336 ( .A(n_243), .B(n_287), .Y(n_336) );
AOI31xp33_ASAP7_75t_SL g251 ( .A1(n_252), .A2(n_266), .A3(n_269), .B(n_271), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_265), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_253), .B(n_288), .Y(n_299) );
OR2x2_ASAP7_75t_L g323 ( .A(n_253), .B(n_293), .Y(n_323) );
INVx1_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_254), .B(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g344 ( .A(n_254), .B(n_336), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_254), .B(n_326), .Y(n_354) );
AND2x2_ASAP7_75t_L g361 ( .A(n_254), .B(n_362), .Y(n_361) );
NAND2x1_ASAP7_75t_L g389 ( .A(n_254), .B(n_325), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_254), .B(n_380), .Y(n_390) );
AND2x2_ASAP7_75t_L g402 ( .A(n_254), .B(n_287), .Y(n_402) );
INVx3_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx3_ASAP7_75t_L g282 ( .A(n_255), .Y(n_282) );
INVx1_ASAP7_75t_L g348 ( .A(n_265), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_265), .B(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_267), .B(n_343), .Y(n_377) );
AND2x4_ASAP7_75t_L g288 ( .A(n_268), .B(n_289), .Y(n_288) );
CKINVDCx16_ASAP7_75t_R g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx2_ASAP7_75t_L g367 ( .A(n_273), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_273), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g315 ( .A(n_274), .B(n_305), .Y(n_315) );
AND2x2_ASAP7_75t_L g409 ( .A(n_274), .B(n_279), .Y(n_409) );
INVx1_ASAP7_75t_L g434 ( .A(n_274), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_280), .B1(n_283), .B2(n_284), .C(n_290), .Y(n_275) );
CKINVDCx14_ASAP7_75t_R g296 ( .A(n_276), .Y(n_296) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_277), .B(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_280), .B(n_331), .Y(n_350) );
INVx3_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g399 ( .A(n_281), .B(n_295), .Y(n_399) );
AND2x2_ASAP7_75t_L g313 ( .A(n_282), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g343 ( .A(n_282), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_282), .B(n_326), .Y(n_371) );
NOR3xp33_ASAP7_75t_L g413 ( .A(n_282), .B(n_383), .C(n_414), .Y(n_413) );
AOI211xp5_ASAP7_75t_SL g346 ( .A1(n_283), .A2(n_347), .B(n_349), .C(n_357), .Y(n_346) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OAI22xp33_ASAP7_75t_L g335 ( .A1(n_285), .A2(n_336), .B1(n_337), .B2(n_338), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_286), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_286), .B(n_370), .Y(n_369) );
BUFx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g428 ( .A(n_288), .B(n_402), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_296), .B1(n_297), .B2(n_299), .Y(n_290) );
NOR2xp33_ASAP7_75t_SL g291 ( .A(n_292), .B(n_294), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_294), .B(n_343), .Y(n_374) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_297), .A2(n_389), .B1(n_420), .B2(n_427), .Y(n_426) );
AOI221xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_308), .B1(n_310), .B2(n_315), .C(n_316), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_306), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVxp67_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OAI221xp5_ASAP7_75t_L g316 ( .A1(n_306), .A2(n_317), .B1(n_323), .B2(n_324), .C(n_327), .Y(n_316) );
INVx1_ASAP7_75t_L g359 ( .A(n_307), .Y(n_359) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx1_ASAP7_75t_SL g331 ( .A(n_312), .Y(n_331) );
OR2x2_ASAP7_75t_L g404 ( .A(n_312), .B(n_336), .Y(n_404) );
AND2x2_ASAP7_75t_L g406 ( .A(n_312), .B(n_314), .Y(n_406) );
INVx1_ASAP7_75t_L g345 ( .A(n_315), .Y(n_345) );
OR2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_321), .Y(n_317) );
AOI21xp33_ASAP7_75t_SL g375 ( .A1(n_318), .A2(n_376), .B(n_377), .Y(n_375) );
OR2x2_ASAP7_75t_L g382 ( .A(n_318), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g356 ( .A(n_319), .B(n_340), .Y(n_356) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp33_ASAP7_75t_SL g373 ( .A(n_324), .B(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_325), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_326), .B(n_362), .Y(n_425) );
O2A1O1Ixp33_ASAP7_75t_L g341 ( .A1(n_329), .A2(n_342), .B(n_344), .C(n_345), .Y(n_341) );
NAND2x1_ASAP7_75t_SL g366 ( .A(n_329), .B(n_367), .Y(n_366) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_330), .A2(n_379), .B1(n_381), .B2(n_384), .Y(n_378) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_332), .B(n_422), .Y(n_421) );
NAND5xp2_ASAP7_75t_L g333 ( .A(n_334), .B(n_346), .C(n_364), .D(n_378), .E(n_387), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_335), .B(n_341), .Y(n_334) );
INVx1_ASAP7_75t_L g391 ( .A(n_337), .Y(n_391) );
INVx1_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_339), .A2(n_358), .B1(n_398), .B2(n_400), .C(n_403), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_340), .B(n_434), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_343), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_343), .B(n_409), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_351), .B1(n_353), .B2(n_355), .Y(n_349) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_361), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
AND2x2_ASAP7_75t_L g431 ( .A(n_360), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_368), .B1(n_372), .B2(n_373), .C(n_375), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g415 ( .A(n_370), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_SL g422 ( .A(n_380), .Y(n_422) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OAI21xp5_ASAP7_75t_SL g387 ( .A1(n_388), .A2(n_390), .B(n_391), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OAI211xp5_ASAP7_75t_SL g392 ( .A1(n_393), .A2(n_395), .B(n_397), .C(n_410), .Y(n_392) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
A2O1A1Ixp33_ASAP7_75t_L g419 ( .A1(n_395), .A2(n_420), .B(n_421), .C(n_423), .Y(n_419) );
INVx1_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_399), .B(n_401), .Y(n_400) );
AOI21xp33_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B(n_407), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AOI21xp33_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_433), .B(n_435), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
XOR2xp5_ASAP7_75t_L g715 ( .A(n_441), .B(n_716), .Y(n_715) );
OR3x1_ASAP7_75t_L g441 ( .A(n_442), .B(n_615), .C(n_662), .Y(n_441) );
NAND3xp33_ASAP7_75t_SL g442 ( .A(n_443), .B(n_561), .C(n_586), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_501), .B1(n_528), .B2(n_531), .C(n_539), .Y(n_443) );
OAI21xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_469), .B(n_494), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_446), .B(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_446), .B(n_544), .Y(n_659) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_460), .Y(n_446) );
AND2x2_ASAP7_75t_L g530 ( .A(n_447), .B(n_500), .Y(n_530) );
AND2x2_ASAP7_75t_L g579 ( .A(n_447), .B(n_499), .Y(n_579) );
AND2x2_ASAP7_75t_L g600 ( .A(n_447), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g605 ( .A(n_447), .B(n_572), .Y(n_605) );
OR2x2_ASAP7_75t_L g613 ( .A(n_447), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g685 ( .A(n_447), .B(n_482), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_447), .B(n_634), .Y(n_699) );
INVx3_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g545 ( .A(n_448), .B(n_460), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_448), .B(n_482), .Y(n_546) );
AND2x4_ASAP7_75t_L g567 ( .A(n_448), .B(n_500), .Y(n_567) );
AND2x2_ASAP7_75t_L g597 ( .A(n_448), .B(n_471), .Y(n_597) );
AND2x2_ASAP7_75t_L g606 ( .A(n_448), .B(n_596), .Y(n_606) );
AND2x2_ASAP7_75t_L g622 ( .A(n_448), .B(n_483), .Y(n_622) );
OR2x2_ASAP7_75t_L g631 ( .A(n_448), .B(n_614), .Y(n_631) );
AND2x2_ASAP7_75t_L g637 ( .A(n_448), .B(n_572), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_448), .B(n_643), .Y(n_642) );
OR2x2_ASAP7_75t_L g651 ( .A(n_448), .B(n_496), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_448), .B(n_541), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_448), .B(n_601), .Y(n_690) );
OR2x6_ASAP7_75t_L g448 ( .A(n_449), .B(n_458), .Y(n_448) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_456), .B(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g500 ( .A(n_460), .Y(n_500) );
AND2x2_ASAP7_75t_L g596 ( .A(n_460), .B(n_482), .Y(n_596) );
AND2x2_ASAP7_75t_L g601 ( .A(n_460), .B(n_483), .Y(n_601) );
INVx1_ASAP7_75t_L g657 ( .A(n_460), .Y(n_657) );
OA21x2_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_462), .B(n_468), .Y(n_460) );
OA21x2_ASAP7_75t_L g512 ( .A1(n_461), .A2(n_513), .B(n_519), .Y(n_512) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_461), .A2(n_521), .B(n_527), .Y(n_520) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g566 ( .A(n_470), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_482), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_471), .B(n_530), .Y(n_529) );
BUFx3_ASAP7_75t_L g544 ( .A(n_471), .Y(n_544) );
OR2x2_ASAP7_75t_L g614 ( .A(n_471), .B(n_482), .Y(n_614) );
OR2x2_ASAP7_75t_L g675 ( .A(n_471), .B(n_582), .Y(n_675) );
OA21x2_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B(n_480), .Y(n_471) );
INVx1_ASAP7_75t_L g497 ( .A(n_473), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_480), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_482), .B(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g634 ( .A(n_482), .B(n_496), .Y(n_634) );
INVx2_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
BUFx2_ASAP7_75t_L g573 ( .A(n_483), .Y(n_573) );
INVx1_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_495), .A2(n_679), .B1(n_683), .B2(n_686), .C(n_687), .Y(n_678) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_499), .Y(n_495) );
INVx1_ASAP7_75t_SL g542 ( .A(n_496), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_496), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g673 ( .A(n_496), .B(n_530), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_499), .B(n_544), .Y(n_665) );
AND2x2_ASAP7_75t_L g572 ( .A(n_500), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_SL g576 ( .A(n_501), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g612 ( .A(n_501), .B(n_582), .Y(n_612) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_511), .Y(n_501) );
AND2x2_ASAP7_75t_L g538 ( .A(n_502), .B(n_512), .Y(n_538) );
INVx4_ASAP7_75t_L g550 ( .A(n_502), .Y(n_550) );
BUFx3_ASAP7_75t_L g592 ( .A(n_502), .Y(n_592) );
AND3x2_ASAP7_75t_L g607 ( .A(n_502), .B(n_608), .C(n_609), .Y(n_607) );
AND2x2_ASAP7_75t_L g689 ( .A(n_511), .B(n_603), .Y(n_689) );
AND2x2_ASAP7_75t_L g697 ( .A(n_511), .B(n_582), .Y(n_697) );
INVx1_ASAP7_75t_SL g702 ( .A(n_511), .Y(n_702) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_520), .Y(n_511) );
INVx1_ASAP7_75t_SL g560 ( .A(n_512), .Y(n_560) );
AND2x2_ASAP7_75t_L g583 ( .A(n_512), .B(n_550), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_512), .B(n_534), .Y(n_585) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_512), .Y(n_625) );
OR2x2_ASAP7_75t_L g630 ( .A(n_512), .B(n_550), .Y(n_630) );
INVx2_ASAP7_75t_L g536 ( .A(n_520), .Y(n_536) );
AND2x2_ASAP7_75t_L g570 ( .A(n_520), .B(n_551), .Y(n_570) );
OR2x2_ASAP7_75t_L g590 ( .A(n_520), .B(n_551), .Y(n_590) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_520), .Y(n_610) );
INVx1_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
AOI21xp33_ASAP7_75t_L g660 ( .A1(n_529), .A2(n_569), .B(n_661), .Y(n_660) );
AOI322xp5_ASAP7_75t_L g696 ( .A1(n_531), .A2(n_541), .A3(n_567), .B1(n_697), .B2(n_698), .C1(n_700), .C2(n_703), .Y(n_696) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_537), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_533), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_534), .B(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g559 ( .A(n_535), .B(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g627 ( .A(n_536), .B(n_550), .Y(n_627) );
AND2x2_ASAP7_75t_L g694 ( .A(n_536), .B(n_551), .Y(n_694) );
INVx1_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g635 ( .A(n_538), .B(n_589), .Y(n_635) );
AOI31xp33_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_543), .A3(n_546), .B(n_547), .Y(n_539) );
AND2x2_ASAP7_75t_L g594 ( .A(n_541), .B(n_572), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_541), .B(n_564), .Y(n_676) );
AND2x2_ASAP7_75t_L g695 ( .A(n_541), .B(n_600), .Y(n_695) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_544), .B(n_572), .Y(n_584) );
NAND2x1p5_ASAP7_75t_L g618 ( .A(n_544), .B(n_601), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_544), .B(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_544), .B(n_685), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_545), .B(n_601), .Y(n_633) );
INVx1_ASAP7_75t_L g677 ( .A(n_545), .Y(n_677) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_559), .Y(n_548) );
INVxp67_ASAP7_75t_L g629 ( .A(n_549), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_550), .B(n_560), .Y(n_565) );
INVx1_ASAP7_75t_L g671 ( .A(n_550), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_550), .B(n_648), .Y(n_682) );
BUFx3_ASAP7_75t_L g582 ( .A(n_551), .Y(n_582) );
AND2x2_ASAP7_75t_L g608 ( .A(n_551), .B(n_560), .Y(n_608) );
INVx2_ASAP7_75t_L g648 ( .A(n_551), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g680 ( .A(n_559), .B(n_681), .Y(n_680) );
AOI211xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_566), .B(n_568), .C(n_577), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AOI21xp33_ASAP7_75t_L g611 ( .A1(n_563), .A2(n_612), .B(n_613), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_564), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_564), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g644 ( .A(n_565), .B(n_590), .Y(n_644) );
INVx3_ASAP7_75t_L g575 ( .A(n_567), .Y(n_575) );
OAI22xp5_ASAP7_75t_SL g568 ( .A1(n_569), .A2(n_571), .B1(n_574), .B2(n_576), .Y(n_568) );
OAI21xp5_ASAP7_75t_SL g593 ( .A1(n_570), .A2(n_594), .B(n_595), .Y(n_593) );
AND2x2_ASAP7_75t_L g619 ( .A(n_570), .B(n_583), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_570), .B(n_671), .Y(n_670) );
INVxp67_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OR2x2_ASAP7_75t_L g574 ( .A(n_573), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g643 ( .A(n_573), .Y(n_643) );
OAI21xp5_ASAP7_75t_SL g587 ( .A1(n_574), .A2(n_588), .B(n_593), .Y(n_587) );
OAI22xp33_ASAP7_75t_SL g577 ( .A1(n_578), .A2(n_580), .B1(n_584), .B2(n_585), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_579), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
INVx1_ASAP7_75t_L g603 ( .A(n_582), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_582), .B(n_625), .Y(n_624) );
NOR3xp33_ASAP7_75t_L g586 ( .A(n_587), .B(n_598), .C(n_611), .Y(n_586) );
OAI22xp5_ASAP7_75t_SL g653 ( .A1(n_588), .A2(n_654), .B1(n_658), .B2(n_659), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_589), .B(n_591), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g658 ( .A(n_590), .B(n_591), .Y(n_658) );
AND2x2_ASAP7_75t_L g666 ( .A(n_591), .B(n_647), .Y(n_666) );
CKINVDCx16_ASAP7_75t_R g591 ( .A(n_592), .Y(n_591) );
O2A1O1Ixp33_ASAP7_75t_SL g674 ( .A1(n_592), .A2(n_675), .B(n_676), .C(n_677), .Y(n_674) );
OR2x2_ASAP7_75t_L g701 ( .A(n_592), .B(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
OAI21xp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_602), .B(n_604), .Y(n_598) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
O2A1O1Ixp33_ASAP7_75t_L g636 ( .A1(n_600), .A2(n_637), .B(n_638), .C(n_641), .Y(n_636) );
OAI21xp33_ASAP7_75t_SL g604 ( .A1(n_605), .A2(n_606), .B(n_607), .Y(n_604) );
AND2x2_ASAP7_75t_L g669 ( .A(n_608), .B(n_627), .Y(n_669) );
INVxp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g647 ( .A(n_610), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g652 ( .A(n_612), .Y(n_652) );
NAND3xp33_ASAP7_75t_SL g615 ( .A(n_616), .B(n_636), .C(n_649), .Y(n_615) );
AOI211xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_619), .B(n_620), .C(n_628), .Y(n_616) );
INVx1_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .Y(n_620) );
INVx1_ASAP7_75t_L g686 ( .A(n_623), .Y(n_686) );
OR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
INVx1_ASAP7_75t_L g646 ( .A(n_625), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_625), .B(n_694), .Y(n_693) );
INVxp67_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
A2O1A1Ixp33_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_630), .B(n_631), .C(n_632), .Y(n_628) );
INVx2_ASAP7_75t_SL g640 ( .A(n_630), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_631), .A2(n_642), .B1(n_644), .B2(n_645), .Y(n_641) );
OAI21xp33_ASAP7_75t_SL g632 ( .A1(n_633), .A2(n_634), .B(n_635), .Y(n_632) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
AOI211xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_652), .B(n_653), .C(n_660), .Y(n_649) );
INVx1_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
INVxp33_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g703 ( .A(n_657), .Y(n_703) );
NAND4xp25_ASAP7_75t_L g662 ( .A(n_663), .B(n_678), .C(n_691), .D(n_696), .Y(n_662) );
AOI211xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_666), .B(n_667), .C(n_674), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_670), .B(n_672), .Y(n_667) );
AOI21xp33_ASAP7_75t_L g687 ( .A1(n_668), .A2(n_688), .B(n_690), .Y(n_687) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_675), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_695), .Y(n_691) );
INVxp67_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_721), .Y(n_720) );
endmodule