module fake_jpeg_28757_n_457 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_457);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_457;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_50),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_52),
.Y(n_130)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g96 ( 
.A(n_54),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_60),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_67),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_16),
.B(n_7),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_77),
.Y(n_119)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx5_ASAP7_75t_SL g102 ( 
.A(n_75),
.Y(n_102)
);

NAND2xp33_ASAP7_75t_SL g76 ( 
.A(n_33),
.B(n_7),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_26),
.C(n_29),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_16),
.B(n_9),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_19),
.B(n_27),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_81),
.B(n_90),
.Y(n_128)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_39),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_91),
.B(n_46),
.Y(n_113)
);

INVx6_ASAP7_75t_SL g92 ( 
.A(n_39),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_92),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_82),
.A2(n_41),
.B1(n_39),
.B2(n_44),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_100),
.A2(n_118),
.B1(n_125),
.B2(n_127),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_75),
.A2(n_41),
.B1(n_27),
.B2(n_19),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_124),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_113),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_61),
.A2(n_25),
.B1(n_23),
.B2(n_44),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_62),
.A2(n_25),
.B1(n_23),
.B2(n_46),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_56),
.A2(n_22),
.B1(n_43),
.B2(n_20),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_63),
.B(n_28),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_136),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_66),
.B(n_22),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_47),
.A2(n_29),
.B1(n_26),
.B2(n_40),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_141),
.A2(n_15),
.B1(n_21),
.B2(n_31),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_50),
.B(n_20),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_142),
.B(n_72),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_119),
.B(n_43),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_147),
.B(n_162),
.Y(n_197)
);

O2A1O1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_131),
.A2(n_40),
.B(n_28),
.C(n_15),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_148),
.A2(n_141),
.B(n_96),
.C(n_138),
.Y(n_198)
);

INVx11_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_149),
.Y(n_207)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_150),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_151),
.A2(n_159),
.B1(n_182),
.B2(n_10),
.Y(n_220)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_117),
.Y(n_152)
);

INVx4_ASAP7_75t_SL g227 ( 
.A(n_152),
.Y(n_227)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_84),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_167),
.Y(n_200)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_101),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_156),
.Y(n_196)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_107),
.Y(n_157)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_157),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_127),
.A2(n_89),
.B(n_52),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_158),
.A2(n_100),
.B(n_65),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_130),
.A2(n_69),
.B1(n_68),
.B2(n_48),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_102),
.A2(n_74),
.B1(n_86),
.B2(n_51),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_160),
.Y(n_214)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_145),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_163),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_108),
.Y(n_164)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_165),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_102),
.A2(n_60),
.B1(n_57),
.B2(n_54),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_166),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_21),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_168),
.Y(n_216)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_170),
.Y(n_217)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_97),
.Y(n_171)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_171),
.Y(n_223)
);

AND2x2_ASAP7_75t_SL g172 ( 
.A(n_116),
.B(n_0),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_172),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_98),
.Y(n_174)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_174),
.A2(n_179),
.B(n_180),
.Y(n_193)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_95),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_177),
.Y(n_202)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_176),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_126),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_178),
.Y(n_218)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_93),
.B(n_31),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_183),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_130),
.A2(n_55),
.B1(n_83),
.B2(n_80),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_144),
.B(n_71),
.Y(n_183)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_129),
.Y(n_184)
);

OA22x2_ASAP7_75t_L g201 ( 
.A1(n_184),
.A2(n_187),
.B1(n_120),
.B2(n_94),
.Y(n_201)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_L g226 ( 
.A1(n_185),
.A2(n_188),
.B1(n_18),
.B2(n_45),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_103),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_186),
.A2(n_114),
.B1(n_138),
.B2(n_133),
.Y(n_194)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_133),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_103),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_SL g219 ( 
.A1(n_189),
.A2(n_190),
.B(n_18),
.Y(n_219)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_94),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_104),
.B(n_140),
.C(n_122),
.Y(n_191)
);

AOI32xp33_ASAP7_75t_L g211 ( 
.A1(n_191),
.A2(n_96),
.A3(n_109),
.B1(n_88),
.B2(n_59),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_192),
.B(n_201),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_194),
.Y(n_261)
);

NOR3xp33_ASAP7_75t_L g237 ( 
.A(n_198),
.B(n_148),
.C(n_151),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_155),
.A2(n_105),
.B1(n_114),
.B2(n_110),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_203),
.A2(n_205),
.B1(n_209),
.B2(n_215),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_158),
.A2(n_109),
.B1(n_108),
.B2(n_110),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_169),
.A2(n_146),
.B1(n_191),
.B2(n_154),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_211),
.A2(n_222),
.B(n_167),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_146),
.A2(n_120),
.B1(n_18),
.B2(n_45),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_219),
.A2(n_224),
.B1(n_221),
.B2(n_214),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_220),
.A2(n_164),
.B1(n_152),
.B2(n_163),
.Y(n_244)
);

A2O1A1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_146),
.A2(n_10),
.B(n_14),
.C(n_13),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_154),
.A2(n_18),
.B1(n_45),
.B2(n_2),
.Y(n_224)
);

INVx3_ASAP7_75t_SL g259 ( 
.A(n_226),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_172),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_229),
.B(n_231),
.Y(n_276)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_230),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_172),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_216),
.Y(n_232)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_232),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_209),
.B(n_173),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_233),
.B(n_235),
.Y(n_267)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_234),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_167),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_236),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_237),
.A2(n_205),
.B1(n_201),
.B2(n_227),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_192),
.C(n_215),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_203),
.C(n_201),
.Y(n_274)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_195),
.Y(n_239)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_239),
.Y(n_292)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_240),
.B(n_248),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_197),
.B(n_177),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_241),
.B(n_253),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_221),
.A2(n_190),
.B1(n_180),
.B2(n_179),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_242),
.A2(n_255),
.B(n_207),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_244),
.A2(n_260),
.B1(n_227),
.B2(n_225),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_199),
.B(n_153),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_245),
.B(n_251),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_247),
.Y(n_270)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_204),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_195),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_256),
.Y(n_265)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_204),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_250),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_199),
.B(n_156),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_214),
.A2(n_157),
.B(n_175),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_252),
.A2(n_257),
.B(n_242),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_222),
.B(n_13),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_223),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_254),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_198),
.A2(n_171),
.B(n_176),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_168),
.Y(n_256)
);

NAND2xp33_ASAP7_75t_SL g257 ( 
.A(n_211),
.B(n_187),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_212),
.Y(n_258)
);

INVx11_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_220),
.A2(n_178),
.B1(n_184),
.B2(n_149),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_224),
.B(n_0),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_196),
.Y(n_286)
);

AO21x1_ASAP7_75t_L g311 ( 
.A1(n_264),
.A2(n_269),
.B(n_255),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_268),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_255),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_271),
.B(n_286),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_283),
.C(n_289),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_246),
.A2(n_193),
.B1(n_201),
.B2(n_213),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_275),
.A2(n_291),
.B(n_242),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_243),
.A2(n_213),
.B1(n_212),
.B2(n_206),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_277),
.A2(n_278),
.B1(n_280),
.B2(n_259),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_243),
.A2(n_227),
.B1(n_206),
.B2(n_202),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_259),
.A2(n_207),
.B1(n_210),
.B2(n_218),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_279),
.A2(n_285),
.B1(n_288),
.B2(n_259),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_246),
.A2(n_210),
.B1(n_196),
.B2(n_195),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_229),
.B(n_223),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_246),
.A2(n_218),
.B1(n_196),
.B2(n_217),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_244),
.A2(n_260),
.B1(n_259),
.B2(n_233),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_238),
.B(n_217),
.C(n_207),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_238),
.B(n_18),
.C(n_45),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_247),
.C(n_236),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_231),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_297),
.B(n_298),
.C(n_304),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_235),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_265),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_299),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_273),
.B(n_245),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_300),
.B(n_303),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_301),
.A2(n_302),
.B1(n_287),
.B2(n_290),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_264),
.A2(n_274),
.B1(n_271),
.B2(n_266),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_265),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_241),
.Y(n_305)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_305),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_276),
.B(n_251),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_306),
.B(n_312),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_307),
.A2(n_292),
.B1(n_249),
.B2(n_258),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_265),
.B(n_237),
.Y(n_309)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_309),
.Y(n_328)
);

NOR2xp67_ASAP7_75t_SL g310 ( 
.A(n_269),
.B(n_257),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_310),
.A2(n_311),
.B(n_315),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_252),
.C(n_232),
.Y(n_312)
);

AO22x1_ASAP7_75t_L g313 ( 
.A1(n_271),
.A2(n_291),
.B1(n_275),
.B2(n_278),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_323),
.Y(n_327)
);

OAI32xp33_ASAP7_75t_L g314 ( 
.A1(n_266),
.A2(n_262),
.A3(n_253),
.B1(n_256),
.B2(n_248),
.Y(n_314)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_314),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_294),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_316),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_284),
.B(n_250),
.Y(n_317)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_317),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_294),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_318),
.B(n_321),
.Y(n_344)
);

XOR2x1_ASAP7_75t_L g319 ( 
.A(n_267),
.B(n_286),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_319),
.B(n_293),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_270),
.A2(n_277),
.B1(n_280),
.B2(n_286),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_320),
.A2(n_285),
.B1(n_288),
.B2(n_268),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_279),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_284),
.B(n_240),
.Y(n_322)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_322),
.Y(n_346)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_263),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_267),
.B(n_254),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_324),
.B(n_282),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_325),
.A2(n_339),
.B1(n_341),
.B2(n_345),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_332),
.A2(n_295),
.B1(n_313),
.B2(n_301),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_334),
.B(n_338),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_296),
.B(n_282),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_335),
.B(n_297),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_336),
.B(n_324),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_319),
.B(n_272),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_320),
.A2(n_272),
.B1(n_263),
.B2(n_261),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_307),
.A2(n_292),
.B1(n_281),
.B2(n_234),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_309),
.Y(n_343)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_343),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_313),
.A2(n_281),
.B1(n_230),
.B2(n_258),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_347),
.A2(n_314),
.B1(n_298),
.B2(n_308),
.Y(n_370)
);

NAND3xp33_ASAP7_75t_L g348 ( 
.A(n_316),
.B(n_239),
.C(n_9),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_348),
.B(n_9),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_296),
.B(n_281),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_349),
.B(n_302),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_295),
.A2(n_321),
.B1(n_299),
.B2(n_318),
.Y(n_351)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_351),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_306),
.B(n_6),
.Y(n_352)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_352),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_355),
.B(n_366),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_356),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_349),
.B(n_312),
.C(n_304),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_357),
.B(n_373),
.C(n_330),
.Y(n_377)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_336),
.Y(n_359)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_359),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_350),
.B(n_323),
.Y(n_361)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_361),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_332),
.A2(n_295),
.B1(n_308),
.B2(n_311),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_362),
.A2(n_370),
.B1(n_337),
.B2(n_327),
.Y(n_384)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_328),
.Y(n_363)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_363),
.Y(n_392)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_328),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_364),
.Y(n_385)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_344),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_347),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_367),
.B(n_374),
.Y(n_386)
);

AOI21x1_ASAP7_75t_SL g368 ( 
.A1(n_329),
.A2(n_310),
.B(n_315),
.Y(n_368)
);

FAx1_ASAP7_75t_L g389 ( 
.A(n_368),
.B(n_333),
.CI(n_338),
.CON(n_389),
.SN(n_389)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_369),
.B(n_372),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_371),
.B(n_375),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_335),
.B(n_322),
.C(n_317),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_327),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_331),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_377),
.B(n_346),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_369),
.B(n_372),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_378),
.B(n_382),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_357),
.B(n_330),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_365),
.B(n_326),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_383),
.B(n_388),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_384),
.A2(n_325),
.B1(n_339),
.B2(n_340),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_373),
.B(n_326),
.C(n_365),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_387),
.B(n_366),
.C(n_354),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_370),
.B(n_334),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_389),
.B(n_374),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_362),
.B(n_333),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_390),
.B(n_360),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_368),
.B(n_337),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_393),
.B(n_355),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_395),
.B(n_402),
.C(n_407),
.Y(n_418)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_396),
.Y(n_414)
);

FAx1_ASAP7_75t_SL g398 ( 
.A(n_393),
.B(n_356),
.CI(n_342),
.CON(n_398),
.SN(n_398)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_398),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_399),
.B(n_405),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_394),
.B(n_361),
.Y(n_400)
);

CKINVDCx14_ASAP7_75t_R g424 ( 
.A(n_400),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_401),
.B(n_404),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_382),
.B(n_360),
.C(n_353),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_386),
.B(n_384),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_391),
.B(n_364),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_406),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_377),
.B(n_359),
.C(n_340),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_380),
.B(n_363),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_408),
.B(n_409),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_387),
.B(n_346),
.C(n_341),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_SL g416 ( 
.A(n_410),
.B(n_390),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_399),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_412),
.B(n_397),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_416),
.A2(n_410),
.B(n_403),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_398),
.A2(n_381),
.B1(n_379),
.B2(n_392),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_417),
.A2(n_376),
.B1(n_383),
.B2(n_403),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_402),
.A2(n_385),
.B1(n_389),
.B2(n_388),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_419),
.A2(n_420),
.B1(n_12),
.B2(n_11),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_395),
.A2(n_389),
.B1(n_358),
.B2(n_378),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_407),
.B(n_376),
.Y(n_421)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_421),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_425),
.A2(n_434),
.B(n_413),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_426),
.B(n_432),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_427),
.B(n_429),
.Y(n_437)
);

OR2x2_ASAP7_75t_L g428 ( 
.A(n_414),
.B(n_397),
.Y(n_428)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_428),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_419),
.B(n_12),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_431),
.B(n_435),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_418),
.B(n_45),
.Y(n_432)
);

AOI211xp5_ASAP7_75t_L g433 ( 
.A1(n_424),
.A2(n_6),
.B(n_12),
.C(n_2),
.Y(n_433)
);

O2A1O1Ixp33_ASAP7_75t_SL g440 ( 
.A1(n_433),
.A2(n_429),
.B(n_422),
.C(n_411),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_421),
.A2(n_0),
.B(n_1),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_415),
.B(n_1),
.Y(n_435)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_439),
.Y(n_448)
);

NAND3xp33_ASAP7_75t_SL g444 ( 
.A(n_440),
.B(n_414),
.C(n_417),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_430),
.B(n_418),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_441),
.A2(n_442),
.B(n_432),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_428),
.B(n_411),
.Y(n_442)
);

A2O1A1O1Ixp25_ASAP7_75t_L g451 ( 
.A1(n_444),
.A2(n_447),
.B(n_437),
.C(n_3),
.D(n_5),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_445),
.B(n_446),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_436),
.B(n_423),
.C(n_420),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_443),
.A2(n_412),
.B(n_3),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_448),
.B(n_437),
.C(n_438),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_449),
.A2(n_2),
.B(n_3),
.Y(n_453)
);

AOI31xp33_ASAP7_75t_L g452 ( 
.A1(n_451),
.A2(n_5),
.A3(n_2),
.B(n_3),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_452),
.B(n_453),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_454),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_455),
.B(n_450),
.C(n_3),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_456),
.A2(n_5),
.B(n_361),
.Y(n_457)
);


endmodule