module real_aes_6503_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g107 ( .A(n_0), .Y(n_107) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_1), .A2(n_140), .B(n_143), .C(n_218), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_2), .A2(n_168), .B(n_169), .Y(n_167) );
INVx1_ASAP7_75t_L g498 ( .A(n_3), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_4), .B(n_179), .Y(n_178) );
AOI21xp33_ASAP7_75t_L g475 ( .A1(n_5), .A2(n_168), .B(n_476), .Y(n_475) );
AND2x6_ASAP7_75t_L g140 ( .A(n_6), .B(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g243 ( .A(n_7), .Y(n_243) );
INVx1_ASAP7_75t_L g105 ( .A(n_8), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_8), .B(n_40), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_9), .A2(n_267), .B(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_10), .B(n_152), .Y(n_220) );
INVx1_ASAP7_75t_L g480 ( .A(n_11), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_12), .B(n_173), .Y(n_531) );
INVx1_ASAP7_75t_L g132 ( .A(n_13), .Y(n_132) );
INVx1_ASAP7_75t_L g543 ( .A(n_14), .Y(n_543) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_15), .A2(n_187), .B(n_228), .C(n_230), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_16), .B(n_179), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_17), .B(n_469), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_18), .B(n_168), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_19), .B(n_275), .Y(n_274) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_20), .A2(n_173), .B(n_204), .C(n_207), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_21), .B(n_179), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_22), .B(n_152), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_23), .A2(n_206), .B(n_230), .C(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_24), .B(n_152), .Y(n_188) );
CKINVDCx16_ASAP7_75t_R g134 ( .A(n_25), .Y(n_134) );
INVx1_ASAP7_75t_L g185 ( .A(n_26), .Y(n_185) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_27), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_28), .Y(n_216) );
AOI222xp33_ASAP7_75t_L g450 ( .A1(n_29), .A2(n_43), .B1(n_451), .B2(n_739), .C1(n_740), .C2(n_743), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_30), .B(n_152), .Y(n_499) );
INVx1_ASAP7_75t_L g272 ( .A(n_31), .Y(n_272) );
INVx1_ASAP7_75t_L g488 ( .A(n_32), .Y(n_488) );
INVx2_ASAP7_75t_L g138 ( .A(n_33), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_34), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g172 ( .A1(n_35), .A2(n_173), .B(n_174), .C(n_176), .Y(n_172) );
INVxp67_ASAP7_75t_L g273 ( .A(n_36), .Y(n_273) );
CKINVDCx14_ASAP7_75t_R g170 ( .A(n_37), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_L g183 ( .A1(n_38), .A2(n_143), .B(n_184), .C(n_191), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_39), .A2(n_140), .B(n_143), .C(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_40), .B(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g487 ( .A(n_41), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g117 ( .A1(n_42), .A2(n_118), .B1(n_439), .B2(n_440), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_42), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_43), .Y(n_739) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_44), .A2(n_154), .B(n_241), .C(n_242), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_45), .B(n_152), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g193 ( .A(n_46), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_47), .Y(n_269) );
INVx1_ASAP7_75t_L g202 ( .A(n_48), .Y(n_202) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_49), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_50), .B(n_168), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g99 ( .A1(n_51), .A2(n_100), .B1(n_111), .B2(n_747), .Y(n_99) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_52), .A2(n_143), .B1(n_207), .B2(n_486), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_53), .Y(n_514) );
CKINVDCx16_ASAP7_75t_R g495 ( .A(n_54), .Y(n_495) );
CKINVDCx14_ASAP7_75t_R g239 ( .A(n_55), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_56), .A2(n_176), .B(n_241), .C(n_479), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_57), .Y(n_523) );
INVx1_ASAP7_75t_L g477 ( .A(n_58), .Y(n_477) );
INVx1_ASAP7_75t_L g141 ( .A(n_59), .Y(n_141) );
INVx1_ASAP7_75t_L g131 ( .A(n_60), .Y(n_131) );
INVx1_ASAP7_75t_SL g175 ( .A(n_61), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_62), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_63), .B(n_179), .Y(n_209) );
INVx1_ASAP7_75t_L g147 ( .A(n_64), .Y(n_147) );
A2O1A1Ixp33_ASAP7_75t_SL g468 ( .A1(n_65), .A2(n_176), .B(n_469), .C(n_470), .Y(n_468) );
INVxp67_ASAP7_75t_L g471 ( .A(n_66), .Y(n_471) );
INVx1_ASAP7_75t_L g110 ( .A(n_67), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_68), .A2(n_168), .B(n_238), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_69), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_70), .A2(n_168), .B(n_225), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_71), .Y(n_491) );
INVx1_ASAP7_75t_L g517 ( .A(n_72), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_73), .B(n_443), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_74), .A2(n_267), .B(n_268), .Y(n_266) );
CKINVDCx16_ASAP7_75t_R g182 ( .A(n_75), .Y(n_182) );
INVx1_ASAP7_75t_L g226 ( .A(n_76), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_77), .A2(n_140), .B(n_143), .C(n_519), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_78), .A2(n_168), .B(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g229 ( .A(n_79), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_80), .B(n_186), .Y(n_511) );
INVx2_ASAP7_75t_L g129 ( .A(n_81), .Y(n_129) );
INVx1_ASAP7_75t_L g219 ( .A(n_82), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_83), .B(n_469), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_84), .A2(n_140), .B(n_143), .C(n_497), .Y(n_496) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_85), .B(n_107), .C(n_108), .Y(n_106) );
OR2x2_ASAP7_75t_L g444 ( .A(n_85), .B(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g455 ( .A(n_85), .Y(n_455) );
OR2x2_ASAP7_75t_L g738 ( .A(n_85), .B(n_446), .Y(n_738) );
A2O1A1Ixp33_ASAP7_75t_L g142 ( .A1(n_86), .A2(n_143), .B(n_146), .C(n_156), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_87), .B(n_161), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_88), .Y(n_502) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_89), .A2(n_140), .B(n_143), .C(n_529), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_90), .Y(n_535) );
INVx1_ASAP7_75t_L g467 ( .A(n_91), .Y(n_467) );
CKINVDCx16_ASAP7_75t_R g540 ( .A(n_92), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_93), .B(n_186), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_94), .B(n_127), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_95), .B(n_127), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_96), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g205 ( .A(n_97), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_98), .A2(n_168), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx5_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
CKINVDCx9p33_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_103), .Y(n_748) );
OR2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
AND2x2_ASAP7_75t_L g446 ( .A(n_107), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
AO21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_116), .B(n_449), .Y(n_111) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx3_ASAP7_75t_L g746 ( .A(n_113), .Y(n_746) );
INVx2_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OAI21xp5_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_441), .B(n_448), .Y(n_116) );
INVx3_ASAP7_75t_L g440 ( .A(n_118), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_118), .A2(n_453), .B1(n_737), .B2(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_SL g118 ( .A(n_119), .B(n_394), .Y(n_118) );
NOR4xp25_ASAP7_75t_L g119 ( .A(n_120), .B(n_331), .C(n_365), .D(n_381), .Y(n_119) );
NAND4xp25_ASAP7_75t_SL g120 ( .A(n_121), .B(n_257), .C(n_295), .D(n_311), .Y(n_120) );
AOI222xp33_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_194), .B1(n_232), .B2(n_245), .C1(n_250), .C2(n_256), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AOI31xp33_ASAP7_75t_L g427 ( .A1(n_123), .A2(n_428), .A3(n_429), .B(n_431), .Y(n_427) );
OR2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_162), .Y(n_123) );
AND2x2_ASAP7_75t_L g402 ( .A(n_124), .B(n_164), .Y(n_402) );
BUFx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_SL g249 ( .A(n_125), .Y(n_249) );
AND2x2_ASAP7_75t_L g256 ( .A(n_125), .B(n_180), .Y(n_256) );
AND2x2_ASAP7_75t_L g316 ( .A(n_125), .B(n_165), .Y(n_316) );
AO21x2_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_133), .B(n_158), .Y(n_125) );
INVx3_ASAP7_75t_L g179 ( .A(n_126), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_126), .B(n_193), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_126), .B(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_SL g513 ( .A(n_126), .B(n_514), .Y(n_513) );
INVx4_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
HB1xp67_ASAP7_75t_L g166 ( .A(n_127), .Y(n_166) );
OA21x2_ASAP7_75t_L g464 ( .A1(n_127), .A2(n_465), .B(n_472), .Y(n_464) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g265 ( .A(n_128), .Y(n_265) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
AND2x2_ASAP7_75t_SL g161 ( .A(n_129), .B(n_130), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
OAI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_135), .B(n_142), .Y(n_133) );
O2A1O1Ixp33_ASAP7_75t_L g181 ( .A1(n_135), .A2(n_161), .B(n_182), .C(n_183), .Y(n_181) );
OAI21xp5_ASAP7_75t_L g215 ( .A1(n_135), .A2(n_216), .B(n_217), .Y(n_215) );
OAI22xp33_ASAP7_75t_L g484 ( .A1(n_135), .A2(n_157), .B1(n_485), .B2(n_489), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_135), .A2(n_495), .B(n_496), .Y(n_494) );
OAI21xp5_ASAP7_75t_L g516 ( .A1(n_135), .A2(n_517), .B(n_518), .Y(n_516) );
NAND2x1p5_ASAP7_75t_L g135 ( .A(n_136), .B(n_140), .Y(n_135) );
AND2x4_ASAP7_75t_L g168 ( .A(n_136), .B(n_140), .Y(n_168) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
INVx1_ASAP7_75t_L g190 ( .A(n_137), .Y(n_190) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g144 ( .A(n_138), .Y(n_144) );
INVx1_ASAP7_75t_L g208 ( .A(n_138), .Y(n_208) );
INVx1_ASAP7_75t_L g145 ( .A(n_139), .Y(n_145) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_139), .Y(n_150) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_139), .Y(n_152) );
INVx3_ASAP7_75t_L g187 ( .A(n_139), .Y(n_187) );
INVx1_ASAP7_75t_L g469 ( .A(n_139), .Y(n_469) );
INVx4_ASAP7_75t_SL g157 ( .A(n_140), .Y(n_157) );
BUFx3_ASAP7_75t_L g191 ( .A(n_140), .Y(n_191) );
INVx5_ASAP7_75t_L g171 ( .A(n_143), .Y(n_171) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
BUFx3_ASAP7_75t_L g155 ( .A(n_144), .Y(n_155) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_144), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_151), .C(n_153), .Y(n_146) );
O2A1O1Ixp5_ASAP7_75t_L g218 ( .A1(n_148), .A2(n_153), .B(n_219), .C(n_220), .Y(n_218) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
OAI22xp5_ASAP7_75t_SL g486 ( .A1(n_149), .A2(n_150), .B1(n_487), .B2(n_488), .Y(n_486) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx4_ASAP7_75t_L g206 ( .A(n_150), .Y(n_206) );
INVx4_ASAP7_75t_L g173 ( .A(n_152), .Y(n_173) );
INVx2_ASAP7_75t_L g241 ( .A(n_152), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_153), .A2(n_511), .B(n_512), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_153), .A2(n_520), .B(n_521), .Y(n_519) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g230 ( .A(n_155), .Y(n_230) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
O2A1O1Ixp33_ASAP7_75t_L g169 ( .A1(n_157), .A2(n_170), .B(n_171), .C(n_172), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_SL g201 ( .A1(n_157), .A2(n_171), .B(n_202), .C(n_203), .Y(n_201) );
O2A1O1Ixp33_ASAP7_75t_SL g225 ( .A1(n_157), .A2(n_171), .B(n_226), .C(n_227), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_SL g238 ( .A1(n_157), .A2(n_171), .B(n_239), .C(n_240), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_SL g268 ( .A1(n_157), .A2(n_171), .B(n_269), .C(n_270), .Y(n_268) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_157), .A2(n_171), .B(n_467), .C(n_468), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_157), .A2(n_171), .B(n_477), .C(n_478), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g539 ( .A1(n_157), .A2(n_171), .B(n_540), .C(n_541), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
INVx1_ASAP7_75t_L g275 ( .A(n_160), .Y(n_275) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_160), .A2(n_527), .B(n_534), .Y(n_526) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g214 ( .A(n_161), .Y(n_214) );
OA21x2_ASAP7_75t_L g236 ( .A1(n_161), .A2(n_237), .B(n_244), .Y(n_236) );
OA21x2_ASAP7_75t_L g537 ( .A1(n_161), .A2(n_538), .B(n_544), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_162), .B(n_346), .Y(n_345) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_163), .B(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_163), .B(n_260), .Y(n_306) );
AND2x2_ASAP7_75t_L g399 ( .A(n_163), .B(n_339), .Y(n_399) );
OAI321xp33_ASAP7_75t_L g433 ( .A1(n_163), .A2(n_249), .A3(n_406), .B1(n_434), .B2(n_436), .C(n_437), .Y(n_433) );
NAND4xp25_ASAP7_75t_L g437 ( .A(n_163), .B(n_235), .C(n_346), .D(n_438), .Y(n_437) );
AND2x4_ASAP7_75t_L g163 ( .A(n_164), .B(n_180), .Y(n_163) );
AND2x2_ASAP7_75t_L g301 ( .A(n_164), .B(n_247), .Y(n_301) );
AND2x2_ASAP7_75t_L g320 ( .A(n_164), .B(n_249), .Y(n_320) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g248 ( .A(n_165), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g276 ( .A(n_165), .B(n_180), .Y(n_276) );
AND2x2_ASAP7_75t_L g362 ( .A(n_165), .B(n_247), .Y(n_362) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_178), .Y(n_165) );
OA21x2_ASAP7_75t_L g199 ( .A1(n_166), .A2(n_200), .B(n_209), .Y(n_199) );
OA21x2_ASAP7_75t_L g223 ( .A1(n_166), .A2(n_224), .B(n_231), .Y(n_223) );
BUFx2_ASAP7_75t_L g267 ( .A(n_168), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_173), .B(n_175), .Y(n_174) );
INVx3_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_177), .Y(n_532) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_179), .A2(n_475), .B(n_481), .Y(n_474) );
INVx3_ASAP7_75t_SL g247 ( .A(n_180), .Y(n_247) );
AND2x2_ASAP7_75t_L g294 ( .A(n_180), .B(n_281), .Y(n_294) );
OR2x2_ASAP7_75t_L g327 ( .A(n_180), .B(n_249), .Y(n_327) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_180), .Y(n_334) );
AND2x2_ASAP7_75t_L g363 ( .A(n_180), .B(n_248), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_180), .B(n_336), .Y(n_378) );
AND2x2_ASAP7_75t_L g410 ( .A(n_180), .B(n_402), .Y(n_410) );
AND2x2_ASAP7_75t_L g419 ( .A(n_180), .B(n_261), .Y(n_419) );
OR2x6_ASAP7_75t_L g180 ( .A(n_181), .B(n_192), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_188), .C(n_189), .Y(n_184) );
OAI22xp33_ASAP7_75t_L g271 ( .A1(n_186), .A2(n_206), .B1(n_272), .B2(n_273), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_L g497 ( .A1(n_186), .A2(n_498), .B(n_499), .C(n_500), .Y(n_497) );
INVx5_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_187), .B(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_187), .B(n_471), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_187), .B(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_190), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_196), .B(n_210), .Y(n_195) );
INVx1_ASAP7_75t_SL g387 ( .A(n_196), .Y(n_387) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g252 ( .A(n_197), .B(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g234 ( .A(n_198), .B(n_212), .Y(n_234) );
AND2x2_ASAP7_75t_L g323 ( .A(n_198), .B(n_236), .Y(n_323) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g293 ( .A(n_199), .B(n_223), .Y(n_293) );
OR2x2_ASAP7_75t_L g304 ( .A(n_199), .B(n_236), .Y(n_304) );
AND2x2_ASAP7_75t_L g330 ( .A(n_199), .B(n_236), .Y(n_330) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_199), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_206), .B(n_229), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_206), .B(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g500 ( .A(n_207), .Y(n_500) );
INVx3_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_210), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_210), .B(n_387), .Y(n_386) );
INVx2_ASAP7_75t_SL g210 ( .A(n_211), .Y(n_210) );
OR2x2_ASAP7_75t_L g303 ( .A(n_211), .B(n_304), .Y(n_303) );
AOI322xp5_ASAP7_75t_L g389 ( .A1(n_211), .A2(n_293), .A3(n_299), .B1(n_330), .B2(n_380), .C1(n_390), .C2(n_392), .Y(n_389) );
OR2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_223), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_212), .B(n_235), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_212), .B(n_236), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_212), .B(n_253), .Y(n_310) );
AND2x2_ASAP7_75t_L g364 ( .A(n_212), .B(n_330), .Y(n_364) );
INVx1_ASAP7_75t_L g368 ( .A(n_212), .Y(n_368) );
AND2x2_ASAP7_75t_L g380 ( .A(n_212), .B(n_223), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_212), .B(n_252), .Y(n_412) );
INVx4_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g277 ( .A(n_213), .B(n_223), .Y(n_277) );
BUFx3_ASAP7_75t_L g291 ( .A(n_213), .Y(n_291) );
AND3x2_ASAP7_75t_L g373 ( .A(n_213), .B(n_353), .C(n_374), .Y(n_373) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_221), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_214), .B(n_502), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_214), .B(n_523), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_214), .B(n_535), .Y(n_534) );
NAND3xp33_ASAP7_75t_L g233 ( .A(n_223), .B(n_234), .C(n_235), .Y(n_233) );
INVx1_ASAP7_75t_SL g253 ( .A(n_223), .Y(n_253) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_223), .Y(n_358) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g352 ( .A(n_234), .B(n_353), .Y(n_352) );
INVxp67_ASAP7_75t_L g359 ( .A(n_234), .Y(n_359) );
AND2x2_ASAP7_75t_L g397 ( .A(n_235), .B(n_375), .Y(n_397) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
BUFx3_ASAP7_75t_L g278 ( .A(n_236), .Y(n_278) );
AND2x2_ASAP7_75t_L g353 ( .A(n_236), .B(n_253), .Y(n_353) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
OR2x2_ASAP7_75t_L g297 ( .A(n_247), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g416 ( .A(n_247), .B(n_316), .Y(n_416) );
AND2x2_ASAP7_75t_L g430 ( .A(n_247), .B(n_249), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_248), .B(n_261), .Y(n_371) );
AND2x2_ASAP7_75t_L g418 ( .A(n_248), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g281 ( .A(n_249), .B(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g298 ( .A(n_249), .B(n_261), .Y(n_298) );
INVx1_ASAP7_75t_L g308 ( .A(n_249), .Y(n_308) );
AND2x2_ASAP7_75t_L g339 ( .A(n_249), .B(n_261), .Y(n_339) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OAI221xp5_ASAP7_75t_L g381 ( .A1(n_251), .A2(n_382), .B1(n_386), .B2(n_388), .C(n_389), .Y(n_381) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_252), .B(n_254), .Y(n_251) );
AND2x2_ASAP7_75t_L g285 ( .A(n_252), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_255), .B(n_292), .Y(n_435) );
AOI322xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_277), .A3(n_278), .B1(n_279), .B2(n_285), .C1(n_287), .C2(n_294), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_276), .Y(n_259) );
NAND2x1p5_ASAP7_75t_L g315 ( .A(n_260), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_260), .B(n_326), .Y(n_325) );
O2A1O1Ixp33_ASAP7_75t_L g349 ( .A1(n_260), .A2(n_276), .B(n_350), .C(n_351), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_260), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_260), .B(n_320), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_260), .B(n_402), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_260), .B(n_430), .Y(n_429) );
BUFx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_261), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_261), .B(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g391 ( .A(n_261), .B(n_278), .Y(n_391) );
OA21x2_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_266), .B(n_274), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AO21x2_ASAP7_75t_L g282 ( .A1(n_263), .A2(n_283), .B(n_284), .Y(n_282) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_263), .A2(n_516), .B(n_522), .Y(n_515) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AOI21xp5_ASAP7_75t_SL g507 ( .A1(n_264), .A2(n_508), .B(n_509), .Y(n_507) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AO21x2_ASAP7_75t_L g483 ( .A1(n_265), .A2(n_484), .B(n_490), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_265), .B(n_491), .Y(n_490) );
AO21x2_ASAP7_75t_L g493 ( .A1(n_265), .A2(n_494), .B(n_501), .Y(n_493) );
INVx1_ASAP7_75t_L g283 ( .A(n_266), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_274), .Y(n_284) );
INVx1_ASAP7_75t_L g366 ( .A(n_276), .Y(n_366) );
OAI31xp33_ASAP7_75t_L g376 ( .A1(n_276), .A2(n_301), .A3(n_377), .B(n_379), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_276), .B(n_282), .Y(n_428) );
INVx1_ASAP7_75t_SL g289 ( .A(n_277), .Y(n_289) );
AND2x2_ASAP7_75t_L g322 ( .A(n_277), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g403 ( .A(n_277), .B(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g288 ( .A(n_278), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g313 ( .A(n_278), .Y(n_313) );
AND2x2_ASAP7_75t_L g340 ( .A(n_278), .B(n_293), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_278), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g432 ( .A(n_278), .B(n_380), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_280), .B(n_350), .Y(n_423) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g319 ( .A(n_282), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_SL g337 ( .A(n_282), .Y(n_337) );
NAND2xp33_ASAP7_75t_SL g287 ( .A(n_288), .B(n_290), .Y(n_287) );
OAI211xp5_ASAP7_75t_SL g331 ( .A1(n_289), .A2(n_332), .B(n_338), .C(n_354), .Y(n_331) );
OR2x2_ASAP7_75t_L g406 ( .A(n_289), .B(n_387), .Y(n_406) );
OR2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
CKINVDCx16_ASAP7_75t_R g343 ( .A(n_291), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_291), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g312 ( .A(n_293), .B(n_313), .Y(n_312) );
O2A1O1Ixp33_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_299), .B(n_302), .C(n_305), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_SL g346 ( .A(n_298), .Y(n_346) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_301), .B(n_339), .Y(n_344) );
INVx1_ASAP7_75t_L g350 ( .A(n_301), .Y(n_350) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g309 ( .A(n_304), .B(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g342 ( .A(n_304), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g404 ( .A(n_304), .Y(n_404) );
AOI21xp33_ASAP7_75t_SL g305 ( .A1(n_306), .A2(n_307), .B(n_309), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_307), .A2(n_318), .B(n_321), .Y(n_317) );
AOI211xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_314), .B(n_317), .C(n_324), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_312), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_315), .B(n_406), .Y(n_405) );
INVx2_ASAP7_75t_SL g328 ( .A(n_316), .Y(n_328) );
OAI21xp5_ASAP7_75t_L g383 ( .A1(n_318), .A2(n_384), .B(n_385), .Y(n_383) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_323), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g348 ( .A(n_323), .Y(n_348) );
AOI21xp33_ASAP7_75t_SL g324 ( .A1(n_325), .A2(n_328), .B(n_329), .Y(n_324) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g379 ( .A(n_330), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_336), .B(n_362), .Y(n_388) );
AND2x2_ASAP7_75t_L g401 ( .A(n_336), .B(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g415 ( .A(n_336), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g425 ( .A(n_336), .B(n_363), .Y(n_425) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AOI211xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_340), .B(n_341), .C(n_349), .Y(n_338) );
INVx1_ASAP7_75t_L g385 ( .A(n_339), .Y(n_385) );
OAI22xp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_344), .B1(n_345), .B2(n_347), .Y(n_341) );
OR2x2_ASAP7_75t_L g347 ( .A(n_343), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_SL g426 ( .A(n_343), .B(n_404), .Y(n_426) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g420 ( .A(n_353), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_360), .B1(n_363), .B2(n_364), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
INVx1_ASAP7_75t_L g438 ( .A(n_358), .Y(n_438) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g384 ( .A(n_362), .Y(n_384) );
OAI211xp5_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_367), .B(n_369), .C(n_376), .Y(n_365) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
INVx2_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
INVxp67_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVxp67_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_384), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NOR5xp2_ASAP7_75t_L g394 ( .A(n_395), .B(n_413), .C(n_421), .D(n_427), .E(n_433), .Y(n_394) );
OAI211xp5_ASAP7_75t_SL g395 ( .A1(n_396), .A2(n_398), .B(n_400), .C(n_407), .Y(n_395) );
INVxp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_403), .B(n_405), .Y(n_400) );
OAI21xp33_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_410), .B(n_411), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_410), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AOI21xp33_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_417), .B(n_420), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_SL g436 ( .A(n_416), .Y(n_436) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_424), .B(n_426), .Y(n_421) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_440), .A2(n_453), .B1(n_456), .B2(n_737), .Y(n_452) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NOR2x2_ASAP7_75t_L g742 ( .A(n_445), .B(n_455), .Y(n_742) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g454 ( .A(n_446), .B(n_455), .Y(n_454) );
AOI21xp33_ASAP7_75t_L g449 ( .A1(n_448), .A2(n_450), .B(n_746), .Y(n_449) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g745 ( .A(n_456), .Y(n_745) );
INVx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND4x1_ASAP7_75t_L g457 ( .A(n_458), .B(n_655), .C(n_702), .D(n_722), .Y(n_457) );
NOR3xp33_ASAP7_75t_SL g458 ( .A(n_459), .B(n_585), .C(n_610), .Y(n_458) );
OAI211xp5_ASAP7_75t_SL g459 ( .A1(n_460), .A2(n_503), .B(n_545), .C(n_575), .Y(n_459) );
INVxp67_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_462), .B(n_482), .Y(n_461) );
INVx3_ASAP7_75t_SL g627 ( .A(n_462), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_462), .B(n_558), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_462), .B(n_492), .Y(n_708) );
AND2x2_ASAP7_75t_L g731 ( .A(n_462), .B(n_597), .Y(n_731) );
AND2x4_ASAP7_75t_L g462 ( .A(n_463), .B(n_473), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g549 ( .A(n_464), .B(n_474), .Y(n_549) );
INVx3_ASAP7_75t_L g562 ( .A(n_464), .Y(n_562) );
AND2x2_ASAP7_75t_L g567 ( .A(n_464), .B(n_473), .Y(n_567) );
OR2x2_ASAP7_75t_L g618 ( .A(n_464), .B(n_559), .Y(n_618) );
BUFx2_ASAP7_75t_L g638 ( .A(n_464), .Y(n_638) );
AND2x2_ASAP7_75t_L g648 ( .A(n_464), .B(n_559), .Y(n_648) );
AND2x2_ASAP7_75t_L g654 ( .A(n_464), .B(n_483), .Y(n_654) );
INVx1_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_474), .B(n_559), .Y(n_573) );
INVx2_ASAP7_75t_L g583 ( .A(n_474), .Y(n_583) );
AND2x2_ASAP7_75t_L g596 ( .A(n_474), .B(n_562), .Y(n_596) );
OR2x2_ASAP7_75t_L g607 ( .A(n_474), .B(n_559), .Y(n_607) );
AND2x2_ASAP7_75t_SL g653 ( .A(n_474), .B(n_654), .Y(n_653) );
BUFx2_ASAP7_75t_L g665 ( .A(n_474), .Y(n_665) );
AND2x2_ASAP7_75t_L g711 ( .A(n_474), .B(n_483), .Y(n_711) );
INVx3_ASAP7_75t_SL g584 ( .A(n_482), .Y(n_584) );
OR2x2_ASAP7_75t_L g637 ( .A(n_482), .B(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_492), .Y(n_482) );
INVx3_ASAP7_75t_L g559 ( .A(n_483), .Y(n_559) );
AND2x2_ASAP7_75t_L g626 ( .A(n_483), .B(n_493), .Y(n_626) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_483), .Y(n_694) );
AOI33xp33_ASAP7_75t_L g698 ( .A1(n_483), .A2(n_627), .A3(n_634), .B1(n_643), .B2(n_699), .B3(n_700), .Y(n_698) );
INVx1_ASAP7_75t_L g547 ( .A(n_492), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_492), .B(n_562), .Y(n_561) );
NOR3xp33_ASAP7_75t_L g621 ( .A(n_492), .B(n_622), .C(n_624), .Y(n_621) );
AND2x2_ASAP7_75t_L g647 ( .A(n_492), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_492), .B(n_654), .Y(n_657) );
AND2x2_ASAP7_75t_L g710 ( .A(n_492), .B(n_711), .Y(n_710) );
INVx3_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx3_ASAP7_75t_L g566 ( .A(n_493), .Y(n_566) );
OR2x2_ASAP7_75t_L g660 ( .A(n_493), .B(n_559), .Y(n_660) );
OR2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_524), .Y(n_503) );
AOI32xp33_ASAP7_75t_L g611 ( .A1(n_504), .A2(n_612), .A3(n_614), .B1(n_616), .B2(n_619), .Y(n_611) );
NOR2xp67_ASAP7_75t_L g684 ( .A(n_504), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g714 ( .A(n_504), .Y(n_714) );
INVx4_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g646 ( .A(n_505), .B(n_630), .Y(n_646) );
AND2x2_ASAP7_75t_L g666 ( .A(n_505), .B(n_592), .Y(n_666) );
AND2x2_ASAP7_75t_L g734 ( .A(n_505), .B(n_652), .Y(n_734) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_515), .Y(n_505) );
INVx3_ASAP7_75t_L g555 ( .A(n_506), .Y(n_555) );
AND2x2_ASAP7_75t_L g569 ( .A(n_506), .B(n_553), .Y(n_569) );
OR2x2_ASAP7_75t_L g574 ( .A(n_506), .B(n_552), .Y(n_574) );
INVx1_ASAP7_75t_L g581 ( .A(n_506), .Y(n_581) );
AND2x2_ASAP7_75t_L g589 ( .A(n_506), .B(n_563), .Y(n_589) );
AND2x2_ASAP7_75t_L g591 ( .A(n_506), .B(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_506), .B(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g644 ( .A(n_506), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_506), .B(n_729), .Y(n_728) );
OR2x6_ASAP7_75t_L g506 ( .A(n_507), .B(n_513), .Y(n_506) );
INVx2_ASAP7_75t_L g553 ( .A(n_515), .Y(n_553) );
AND2x2_ASAP7_75t_L g599 ( .A(n_515), .B(n_525), .Y(n_599) );
AND2x2_ASAP7_75t_L g609 ( .A(n_515), .B(n_537), .Y(n_609) );
INVx2_ASAP7_75t_L g729 ( .A(n_524), .Y(n_729) );
OR2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_536), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_525), .B(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g570 ( .A(n_525), .Y(n_570) );
AND2x2_ASAP7_75t_L g614 ( .A(n_525), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g630 ( .A(n_525), .B(n_593), .Y(n_630) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g578 ( .A(n_526), .Y(n_578) );
AND2x2_ASAP7_75t_L g592 ( .A(n_526), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g643 ( .A(n_526), .B(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_526), .B(n_553), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_533), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B(n_532), .Y(n_529) );
AND2x2_ASAP7_75t_L g554 ( .A(n_536), .B(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g615 ( .A(n_536), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_536), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g652 ( .A(n_536), .Y(n_652) );
INVx1_ASAP7_75t_L g685 ( .A(n_536), .Y(n_685) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g563 ( .A(n_537), .B(n_553), .Y(n_563) );
INVx1_ASAP7_75t_L g593 ( .A(n_537), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_550), .B1(n_556), .B2(n_563), .C(n_564), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_547), .B(n_567), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_547), .B(n_630), .Y(n_707) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_549), .B(n_597), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_549), .B(n_558), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_549), .B(n_572), .Y(n_701) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_554), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g623 ( .A(n_553), .Y(n_623) );
AND2x2_ASAP7_75t_L g598 ( .A(n_554), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g676 ( .A(n_554), .Y(n_676) );
AND2x2_ASAP7_75t_L g608 ( .A(n_555), .B(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_555), .B(n_578), .Y(n_624) );
AND2x2_ASAP7_75t_L g688 ( .A(n_555), .B(n_614), .Y(n_688) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
BUFx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g597 ( .A(n_559), .B(n_566), .Y(n_597) );
AND2x2_ASAP7_75t_L g693 ( .A(n_560), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_562), .B(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_563), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_563), .B(n_570), .Y(n_658) );
AND2x2_ASAP7_75t_L g678 ( .A(n_563), .B(n_578), .Y(n_678) );
AND2x2_ASAP7_75t_L g699 ( .A(n_563), .B(n_643), .Y(n_699) );
OAI32xp33_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_568), .A3(n_570), .B1(n_571), .B2(n_574), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
INVx1_ASAP7_75t_SL g572 ( .A(n_566), .Y(n_572) );
NAND2x1_ASAP7_75t_L g613 ( .A(n_566), .B(n_596), .Y(n_613) );
OR2x2_ASAP7_75t_L g617 ( .A(n_566), .B(n_618), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_566), .B(n_665), .Y(n_718) );
INVx1_ASAP7_75t_L g586 ( .A(n_567), .Y(n_586) );
OAI221xp5_ASAP7_75t_SL g704 ( .A1(n_568), .A2(n_659), .B1(n_705), .B2(n_708), .C(n_709), .Y(n_704) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g576 ( .A(n_569), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g619 ( .A(n_569), .B(n_592), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_569), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g697 ( .A(n_569), .B(n_630), .Y(n_697) );
INVxp67_ASAP7_75t_L g633 ( .A(n_570), .Y(n_633) );
OR2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
AND2x2_ASAP7_75t_L g703 ( .A(n_572), .B(n_690), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_572), .B(n_653), .Y(n_726) );
INVx1_ASAP7_75t_L g601 ( .A(n_574), .Y(n_601) );
NAND2xp5_ASAP7_75t_SL g682 ( .A(n_574), .B(n_683), .Y(n_682) );
OR2x2_ASAP7_75t_L g719 ( .A(n_574), .B(n_720), .Y(n_719) );
OAI21xp5_ASAP7_75t_SL g575 ( .A1(n_576), .A2(n_579), .B(n_582), .Y(n_575) );
AND2x2_ASAP7_75t_L g588 ( .A(n_577), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g672 ( .A(n_581), .B(n_592), .Y(n_672) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
AND2x2_ASAP7_75t_L g690 ( .A(n_583), .B(n_648), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_583), .B(n_647), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_584), .B(n_596), .Y(n_670) );
OAI211xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B(n_590), .C(n_600), .Y(n_585) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_586), .A2(n_621), .B1(n_625), .B2(n_628), .C(n_631), .Y(n_620) );
AOI31xp33_ASAP7_75t_L g715 ( .A1(n_586), .A2(n_716), .A3(n_717), .B(n_719), .Y(n_715) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_594), .B1(n_596), .B2(n_598), .Y(n_590) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
INVx1_ASAP7_75t_L g716 ( .A(n_596), .Y(n_716) );
INVx1_ASAP7_75t_L g679 ( .A(n_597), .Y(n_679) );
O2A1O1Ixp33_ASAP7_75t_L g722 ( .A1(n_599), .A2(n_723), .B(n_725), .C(n_727), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B1(n_604), .B2(n_608), .Y(n_600) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_605), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OAI221xp5_ASAP7_75t_SL g695 ( .A1(n_607), .A2(n_641), .B1(n_660), .B2(n_696), .C(n_698), .Y(n_695) );
INVx1_ASAP7_75t_L g691 ( .A(n_608), .Y(n_691) );
INVx1_ASAP7_75t_L g645 ( .A(n_609), .Y(n_645) );
NAND3xp33_ASAP7_75t_SL g610 ( .A(n_611), .B(n_620), .C(n_635), .Y(n_610) );
OAI21xp33_ASAP7_75t_L g661 ( .A1(n_612), .A2(n_662), .B(n_666), .Y(n_661) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_614), .B(n_714), .Y(n_713) );
INVxp67_ASAP7_75t_L g721 ( .A(n_615), .Y(n_721) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g659 ( .A(n_622), .B(n_642), .Y(n_659) );
INVx1_ASAP7_75t_L g634 ( .A(n_623), .Y(n_634) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx1_ASAP7_75t_L g632 ( .A(n_626), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_626), .B(n_664), .Y(n_663) );
NOR4xp25_ASAP7_75t_L g631 ( .A(n_627), .B(n_632), .C(n_633), .D(n_634), .Y(n_631) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AOI222xp33_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_640), .B1(n_646), .B2(n_647), .C1(n_649), .C2(n_653), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g636 ( .A(n_637), .B(n_639), .Y(n_636) );
INVx1_ASAP7_75t_L g733 ( .A(n_637), .Y(n_733) );
INVx1_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_645), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_649), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OAI21xp5_ASAP7_75t_SL g709 ( .A1(n_654), .A2(n_710), .B(n_712), .Y(n_709) );
NOR4xp25_ASAP7_75t_L g655 ( .A(n_656), .B(n_667), .C(n_680), .D(n_695), .Y(n_655) );
OAI221xp5_ASAP7_75t_SL g656 ( .A1(n_657), .A2(n_658), .B1(n_659), .B2(n_660), .C(n_661), .Y(n_656) );
INVx1_ASAP7_75t_L g736 ( .A(n_657), .Y(n_736) );
INVx1_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_664), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
OAI222xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_671), .B1(n_673), .B2(n_674), .C1(n_677), .C2(n_679), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AOI211xp5_ASAP7_75t_L g702 ( .A1(n_672), .A2(n_703), .B(n_704), .C(n_715), .Y(n_702) );
OR2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
OAI222xp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_686), .B1(n_687), .B2(n_689), .C1(n_691), .C2(n_692), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVxp67_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_697), .A2(n_700), .B1(n_733), .B2(n_734), .Y(n_732) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OAI211xp5_ASAP7_75t_SL g727 ( .A1(n_728), .A2(n_730), .B(n_732), .C(n_735), .Y(n_727) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
endmodule