module fake_netlist_5_1989_n_1782 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1782);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1782;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_88),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_85),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_103),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_28),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_11),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_63),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_87),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_91),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_3),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_52),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_133),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_112),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_69),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_47),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_129),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_63),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_149),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_107),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_54),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_102),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_144),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_111),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_115),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_116),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_31),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_31),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_28),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_73),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_57),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_11),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_148),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_110),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_130),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_46),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_78),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_57),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_37),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_82),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_44),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_96),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_61),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_139),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_118),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_132),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_58),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_143),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_89),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_101),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_56),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_32),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_70),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_14),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_100),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_84),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_108),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_119),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_68),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_122),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_7),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_127),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_76),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_5),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_4),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_26),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_21),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_90),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_35),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_153),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_1),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_125),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_120),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_86),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_18),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_29),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_151),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_43),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_19),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_13),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_37),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_138),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_5),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_3),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_152),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_46),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_4),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_93),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_56),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_29),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_65),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_52),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_136),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_74),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_137),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_71),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_126),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_123),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_27),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_18),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_49),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_33),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_19),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_62),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_154),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_72),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_62),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_97),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_6),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_42),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_75),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_109),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_105),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_79),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_142),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_39),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_6),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_39),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_135),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_14),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_128),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_54),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_58),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_23),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_134),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_38),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_36),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_22),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_117),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_20),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_64),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_12),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_21),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_16),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_114),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_35),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_16),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_92),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_124),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_44),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_59),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_41),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_20),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_131),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_99),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_113),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_104),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_13),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_50),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_146),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_41),
.Y(n_305)
);

BUFx5_ASAP7_75t_L g306 ( 
.A(n_7),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_27),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_306),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_185),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_268),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_306),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_172),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_190),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_306),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_155),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_198),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_161),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_306),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_165),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_306),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_211),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_306),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_306),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_166),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_0),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_169),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_171),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_212),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_175),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_176),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_259),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_306),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_167),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_255),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_178),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_278),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_179),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_183),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_255),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_186),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_255),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_193),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_197),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_252),
.B(n_226),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_202),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_252),
.B(n_0),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_207),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_255),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_255),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_209),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_214),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_229),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_255),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_217),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_159),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_268),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_222),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_159),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_156),
.B(n_1),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_229),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_224),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_231),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_163),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_236),
.Y(n_364)
);

NOR2xp67_ASAP7_75t_L g365 ( 
.A(n_189),
.B(n_2),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_239),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_242),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_245),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_163),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_170),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_170),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_196),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_249),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_196),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_208),
.Y(n_375)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_226),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_226),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_251),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_260),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_228),
.B(n_2),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_265),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_208),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_L g383 ( 
.A(n_189),
.B(n_8),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_308),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_308),
.B(n_228),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_310),
.B(n_156),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_334),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_311),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_311),
.B(n_157),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_314),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_334),
.Y(n_391)
);

BUFx8_ASAP7_75t_L g392 ( 
.A(n_355),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_314),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_318),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_339),
.Y(n_395)
);

INVx5_ASAP7_75t_L g396 ( 
.A(n_309),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_309),
.B(n_192),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_318),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_320),
.B(n_157),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_339),
.B(n_162),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_320),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_346),
.B(n_344),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_322),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_322),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_323),
.B(n_162),
.Y(n_405)
);

OAI21x1_ASAP7_75t_L g406 ( 
.A1(n_323),
.A2(n_187),
.B(n_177),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_341),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_341),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_348),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_348),
.Y(n_410)
);

OA21x2_ASAP7_75t_L g411 ( 
.A1(n_349),
.A2(n_232),
.B(n_215),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_332),
.Y(n_412)
);

INVx5_ASAP7_75t_L g413 ( 
.A(n_332),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_365),
.B(n_278),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_349),
.Y(n_415)
);

AND2x2_ASAP7_75t_SL g416 ( 
.A(n_325),
.B(n_250),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_353),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_353),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_359),
.B(n_177),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_355),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_352),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_358),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_380),
.B(n_187),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_358),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_363),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_365),
.B(n_247),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_363),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_356),
.B(n_188),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_369),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_369),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g431 ( 
.A(n_370),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_370),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_376),
.B(n_188),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_371),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_371),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_377),
.B(n_195),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_372),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_372),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_374),
.Y(n_439)
);

AND2x6_ASAP7_75t_L g440 ( 
.A(n_374),
.B(n_250),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_375),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_375),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_382),
.B(n_195),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_382),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_352),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_315),
.Y(n_446)
);

AND2x6_ASAP7_75t_L g447 ( 
.A(n_383),
.B(n_250),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_383),
.B(n_199),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_317),
.Y(n_449)
);

CKINVDCx8_ASAP7_75t_R g450 ( 
.A(n_336),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_319),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_360),
.B(n_199),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_390),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_384),
.Y(n_454)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_421),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_390),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_390),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_396),
.B(n_324),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_421),
.Y(n_459)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_413),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_390),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_384),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_396),
.B(n_326),
.Y(n_463)
);

INVx5_ASAP7_75t_L g464 ( 
.A(n_440),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_411),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_386),
.B(n_336),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_384),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_396),
.B(n_327),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_449),
.B(n_329),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_390),
.Y(n_470)
);

OR2x6_ASAP7_75t_L g471 ( 
.A(n_446),
.B(n_201),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_390),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_388),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_388),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_388),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_396),
.B(n_330),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_411),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_388),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_384),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_402),
.B(n_337),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_393),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_384),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_402),
.B(n_338),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_393),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_449),
.B(n_342),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_401),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_450),
.Y(n_487)
);

INVx4_ASAP7_75t_L g488 ( 
.A(n_413),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_449),
.B(n_343),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_393),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_393),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_394),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_394),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_413),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_386),
.B(n_345),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_394),
.Y(n_496)
);

BUFx4f_ASAP7_75t_L g497 ( 
.A(n_411),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_386),
.B(n_350),
.Y(n_498)
);

INVx6_ASAP7_75t_L g499 ( 
.A(n_392),
.Y(n_499)
);

XOR2x2_ASAP7_75t_L g500 ( 
.A(n_445),
.B(n_164),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_411),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_401),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_386),
.B(n_354),
.Y(n_503)
);

INVx6_ASAP7_75t_L g504 ( 
.A(n_392),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_394),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_401),
.Y(n_506)
);

NOR3xp33_ASAP7_75t_L g507 ( 
.A(n_414),
.B(n_256),
.C(n_182),
.Y(n_507)
);

AND2x2_ASAP7_75t_SL g508 ( 
.A(n_416),
.B(n_250),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_398),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_445),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_400),
.B(n_201),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_428),
.B(n_357),
.Y(n_512)
);

OAI22xp33_ASAP7_75t_L g513 ( 
.A1(n_419),
.A2(n_168),
.B1(n_246),
.B2(n_218),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_396),
.B(n_362),
.Y(n_514)
);

OR2x6_ASAP7_75t_L g515 ( 
.A(n_446),
.B(n_204),
.Y(n_515)
);

BUFx10_ASAP7_75t_L g516 ( 
.A(n_451),
.Y(n_516)
);

AND3x1_ASAP7_75t_L g517 ( 
.A(n_419),
.B(n_238),
.C(n_192),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_398),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_401),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_451),
.B(n_364),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_398),
.Y(n_521)
);

INVx4_ASAP7_75t_L g522 ( 
.A(n_413),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_398),
.Y(n_523)
);

OR2x6_ASAP7_75t_L g524 ( 
.A(n_446),
.B(n_204),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_396),
.B(n_366),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_403),
.Y(n_526)
);

BUFx4f_ASAP7_75t_L g527 ( 
.A(n_411),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_401),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_403),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_403),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_428),
.B(n_368),
.Y(n_531)
);

INVx6_ASAP7_75t_L g532 ( 
.A(n_392),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_428),
.B(n_378),
.Y(n_533)
);

INVx1_ASAP7_75t_SL g534 ( 
.A(n_397),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_411),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_403),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_428),
.B(n_381),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_416),
.A2(n_238),
.B1(n_290),
.B2(n_276),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_404),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_404),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_404),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_392),
.B(n_203),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_404),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_412),
.Y(n_544)
);

INVx5_ASAP7_75t_L g545 ( 
.A(n_440),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_412),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_448),
.B(n_276),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_412),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_397),
.B(n_414),
.Y(n_549)
);

BUFx4f_ASAP7_75t_L g550 ( 
.A(n_411),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_400),
.B(n_213),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_412),
.Y(n_552)
);

INVxp33_ASAP7_75t_SL g553 ( 
.A(n_452),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_431),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_431),
.Y(n_555)
);

OR2x6_ASAP7_75t_L g556 ( 
.A(n_446),
.B(n_213),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_416),
.A2(n_290),
.B1(n_233),
.B2(n_232),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_415),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_397),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_416),
.A2(n_281),
.B1(n_233),
.B2(n_280),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_400),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_415),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_415),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_392),
.B(n_210),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_415),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_431),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_417),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_396),
.B(n_333),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_417),
.Y(n_569)
);

BUFx8_ASAP7_75t_SL g570 ( 
.A(n_451),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_448),
.B(n_423),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_431),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_392),
.B(n_248),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_SL g574 ( 
.A1(n_419),
.A2(n_235),
.B1(n_191),
.B2(n_230),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_448),
.B(n_216),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_396),
.B(n_379),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_392),
.B(n_275),
.Y(n_577)
);

BUFx10_ASAP7_75t_L g578 ( 
.A(n_416),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_422),
.Y(n_579)
);

BUFx10_ASAP7_75t_L g580 ( 
.A(n_447),
.Y(n_580)
);

BUFx4f_ASAP7_75t_L g581 ( 
.A(n_447),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_448),
.B(n_216),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_417),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_400),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_396),
.B(n_335),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_396),
.B(n_373),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_397),
.B(n_340),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_424),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_417),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_424),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_424),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_387),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_426),
.B(n_347),
.Y(n_593)
);

INVxp33_ASAP7_75t_L g594 ( 
.A(n_452),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_387),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_387),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_426),
.B(n_351),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_391),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_452),
.A2(n_258),
.B1(n_296),
.B2(n_302),
.Y(n_599)
);

INVx4_ASAP7_75t_L g600 ( 
.A(n_413),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_423),
.A2(n_281),
.B1(n_307),
.B2(n_215),
.Y(n_601)
);

NAND3xp33_ASAP7_75t_SL g602 ( 
.A(n_574),
.B(n_313),
.C(n_312),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_584),
.B(n_452),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_584),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_561),
.Y(n_605)
);

BUFx10_ASAP7_75t_L g606 ( 
.A(n_587),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_510),
.B(n_450),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_561),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_510),
.B(n_450),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_480),
.B(n_361),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_549),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_579),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_561),
.Y(n_613)
);

OAI221xp5_ASAP7_75t_L g614 ( 
.A1(n_601),
.A2(n_423),
.B1(n_436),
.B2(n_433),
.C(n_443),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_571),
.B(n_396),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_571),
.B(n_483),
.Y(n_616)
);

AO221x1_ASAP7_75t_L g617 ( 
.A1(n_513),
.A2(n_174),
.B1(n_250),
.B2(n_263),
.C(n_307),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_560),
.A2(n_447),
.B1(n_400),
.B2(n_436),
.Y(n_618)
);

INVxp33_ASAP7_75t_L g619 ( 
.A(n_500),
.Y(n_619)
);

BUFx8_ASAP7_75t_L g620 ( 
.A(n_466),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_511),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_508),
.B(n_444),
.Y(n_622)
);

NOR2xp67_ASAP7_75t_L g623 ( 
.A(n_593),
.B(n_597),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_579),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_592),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_465),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_455),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_508),
.B(n_444),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_553),
.B(n_367),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_L g630 ( 
.A(n_465),
.B(n_447),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_508),
.B(n_450),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_554),
.B(n_444),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_554),
.B(n_444),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_555),
.B(n_444),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_456),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_555),
.B(n_566),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_469),
.B(n_485),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_489),
.B(n_316),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_511),
.B(n_551),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_566),
.B(n_444),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_592),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_459),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_520),
.B(n_321),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_595),
.Y(n_644)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_459),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_572),
.B(n_433),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_578),
.B(n_433),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_572),
.B(n_436),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_594),
.B(n_328),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_495),
.B(n_331),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_595),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_466),
.B(n_443),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_498),
.B(n_158),
.Y(n_653)
);

INVxp33_ASAP7_75t_SL g654 ( 
.A(n_599),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_549),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_465),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_531),
.B(n_160),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_578),
.B(n_389),
.Y(n_658)
);

BUFx8_ASAP7_75t_L g659 ( 
.A(n_559),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_596),
.Y(n_660)
);

NAND3xp33_ASAP7_75t_L g661 ( 
.A(n_507),
.B(n_399),
.C(n_389),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_503),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_487),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_456),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_503),
.A2(n_447),
.B1(n_400),
.B2(n_289),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_533),
.B(n_400),
.Y(n_666)
);

NAND2xp33_ASAP7_75t_L g667 ( 
.A(n_465),
.B(n_447),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_471),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_578),
.B(n_389),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_599),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_596),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_537),
.B(n_575),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_575),
.B(n_399),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_578),
.B(n_399),
.Y(n_674)
);

O2A1O1Ixp5_ASAP7_75t_L g675 ( 
.A1(n_497),
.A2(n_405),
.B(n_385),
.C(n_443),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_471),
.Y(n_676)
);

INVxp67_ASAP7_75t_L g677 ( 
.A(n_512),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_SL g678 ( 
.A(n_534),
.B(n_247),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_582),
.B(n_405),
.Y(n_679)
);

NAND2xp33_ASAP7_75t_L g680 ( 
.A(n_465),
.B(n_447),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_582),
.B(n_405),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_557),
.B(n_447),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_538),
.A2(n_447),
.B1(n_406),
.B2(n_385),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_570),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_598),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_512),
.B(n_447),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_456),
.B(n_447),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_598),
.Y(n_688)
);

BUFx6f_ASAP7_75t_SL g689 ( 
.A(n_516),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_501),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_581),
.B(n_250),
.Y(n_691)
);

OR2x6_ASAP7_75t_L g692 ( 
.A(n_559),
.B(n_406),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_581),
.B(n_385),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_477),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_SL g695 ( 
.A1(n_500),
.A2(n_271),
.B1(n_241),
.B2(n_240),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_547),
.B(n_447),
.Y(n_696)
);

OAI22xp33_ASAP7_75t_L g697 ( 
.A1(n_471),
.A2(n_267),
.B1(n_300),
.B2(n_262),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_581),
.B(n_497),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_547),
.B(n_422),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_477),
.B(n_447),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_497),
.B(n_406),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_516),
.B(n_173),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_477),
.B(n_413),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_516),
.B(n_422),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_516),
.B(n_180),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_477),
.B(n_413),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_477),
.B(n_413),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_453),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_453),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_471),
.B(n_181),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_457),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_501),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_471),
.B(n_184),
.Y(n_713)
);

NOR2x1p5_ASAP7_75t_L g714 ( 
.A(n_542),
.B(n_194),
.Y(n_714)
);

OAI22xp33_ASAP7_75t_L g715 ( 
.A1(n_515),
.A2(n_227),
.B1(n_262),
.B2(n_267),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_527),
.A2(n_413),
.B(n_406),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_457),
.B(n_413),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_535),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_527),
.B(n_424),
.Y(n_719)
);

NOR2xp67_ASAP7_75t_SL g720 ( 
.A(n_499),
.B(n_227),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_527),
.B(n_550),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_535),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_550),
.B(n_424),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_461),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_461),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_470),
.B(n_413),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_470),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_550),
.B(n_424),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_515),
.B(n_200),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_535),
.A2(n_300),
.B1(n_298),
.B2(n_441),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_517),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_472),
.B(n_424),
.Y(n_732)
);

INVxp67_ASAP7_75t_SL g733 ( 
.A(n_490),
.Y(n_733)
);

O2A1O1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_515),
.A2(n_429),
.B(n_438),
.C(n_435),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_472),
.B(n_424),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_515),
.A2(n_266),
.B1(n_299),
.B2(n_304),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_580),
.B(n_424),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_580),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_511),
.Y(n_739)
);

A2O1A1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_511),
.A2(n_551),
.B(n_244),
.C(n_287),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_517),
.B(n_425),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_551),
.B(n_424),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_551),
.B(n_434),
.Y(n_743)
);

INVxp67_ASAP7_75t_L g744 ( 
.A(n_515),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_458),
.A2(n_442),
.B(n_420),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_473),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_580),
.B(n_434),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_473),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_539),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_524),
.B(n_425),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_580),
.B(n_434),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_524),
.B(n_434),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_524),
.B(n_556),
.Y(n_753)
);

NAND2xp33_ASAP7_75t_L g754 ( 
.A(n_564),
.B(n_298),
.Y(n_754)
);

INVxp67_ASAP7_75t_L g755 ( 
.A(n_524),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_558),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_524),
.B(n_434),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_556),
.B(n_434),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_556),
.B(n_434),
.Y(n_759)
);

O2A1O1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_556),
.A2(n_573),
.B(n_577),
.C(n_568),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_576),
.B(n_585),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_556),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_490),
.B(n_434),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_490),
.B(n_434),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_586),
.B(n_425),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_463),
.B(n_205),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_474),
.A2(n_437),
.B1(n_441),
.B2(n_434),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_468),
.B(n_206),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_530),
.B(n_437),
.Y(n_769)
);

INVxp67_ASAP7_75t_L g770 ( 
.A(n_474),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_530),
.B(n_536),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_476),
.B(n_219),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_475),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_637),
.B(n_530),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_616),
.B(n_672),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_626),
.B(n_588),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_607),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_673),
.B(n_679),
.Y(n_778)
);

AO22x1_ASAP7_75t_L g779 ( 
.A1(n_654),
.A2(n_295),
.B1(n_305),
.B2(n_303),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_612),
.Y(n_780)
);

AOI21x1_ASAP7_75t_L g781 ( 
.A1(n_719),
.A2(n_525),
.B(n_514),
.Y(n_781)
);

INVx11_ASAP7_75t_L g782 ( 
.A(n_620),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_693),
.A2(n_488),
.B(n_460),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_652),
.B(n_427),
.Y(n_784)
);

A2O1A1Ixp33_ASAP7_75t_L g785 ( 
.A1(n_623),
.A2(n_244),
.B(n_254),
.C(n_263),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_612),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_L g787 ( 
.A1(n_675),
.A2(n_478),
.B(n_475),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_681),
.B(n_536),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_662),
.B(n_536),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_626),
.B(n_588),
.Y(n_790)
);

NOR3xp33_ASAP7_75t_L g791 ( 
.A(n_602),
.B(n_429),
.C(n_427),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_611),
.B(n_478),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_693),
.A2(n_488),
.B(n_460),
.Y(n_793)
);

A2O1A1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_614),
.A2(n_287),
.B(n_280),
.C(n_254),
.Y(n_794)
);

NOR4xp25_ASAP7_75t_SL g795 ( 
.A(n_631),
.B(n_294),
.C(n_264),
.D(n_261),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_611),
.B(n_481),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_655),
.B(n_481),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_655),
.B(n_484),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_624),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_626),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_647),
.A2(n_677),
.B1(n_631),
.B2(n_686),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_646),
.B(n_484),
.Y(n_802)
);

NOR2x1p5_ASAP7_75t_L g803 ( 
.A(n_684),
.B(n_220),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_627),
.B(n_427),
.Y(n_804)
);

O2A1O1Ixp5_ASAP7_75t_L g805 ( 
.A1(n_761),
.A2(n_519),
.B(n_462),
.C(n_467),
.Y(n_805)
);

OAI21xp33_ASAP7_75t_SL g806 ( 
.A1(n_658),
.A2(n_492),
.B(n_491),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_648),
.B(n_699),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_L g808 ( 
.A1(n_658),
.A2(n_532),
.B1(n_504),
.B2(n_499),
.Y(n_808)
);

A2O1A1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_653),
.A2(n_429),
.B(n_435),
.C(n_438),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_738),
.A2(n_488),
.B(n_460),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_647),
.A2(n_610),
.B1(n_661),
.B2(n_603),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_738),
.A2(n_488),
.B(n_460),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_738),
.A2(n_522),
.B(n_494),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_704),
.B(n_491),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_669),
.A2(n_532),
.B1(n_504),
.B2(n_499),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_657),
.B(n_492),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_738),
.A2(n_674),
.B(n_669),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_624),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_666),
.B(n_493),
.Y(n_819)
);

AND2x2_ASAP7_75t_SL g820 ( 
.A(n_754),
.B(n_588),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_674),
.A2(n_522),
.B(n_494),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_708),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_639),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_603),
.B(n_493),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_603),
.B(n_496),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_625),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_690),
.B(n_496),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_625),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_709),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_630),
.A2(n_522),
.B(n_494),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_609),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_741),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_626),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_630),
.A2(n_522),
.B(n_494),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_667),
.A2(n_600),
.B(n_509),
.Y(n_835)
);

O2A1O1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_740),
.A2(n_628),
.B(n_622),
.C(n_744),
.Y(n_836)
);

OAI21xp5_ASAP7_75t_L g837 ( 
.A1(n_615),
.A2(n_509),
.B(n_505),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_667),
.A2(n_600),
.B(n_518),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_710),
.A2(n_438),
.B(n_435),
.C(n_505),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_711),
.Y(n_840)
);

O2A1O1Ixp5_ASAP7_75t_SL g841 ( 
.A1(n_761),
.A2(n_552),
.B(n_548),
.C(n_546),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_656),
.B(n_588),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_690),
.A2(n_532),
.B1(n_499),
.B2(n_504),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_641),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_712),
.B(n_518),
.Y(n_845)
);

NOR2xp67_ASAP7_75t_L g846 ( 
.A(n_642),
.B(n_269),
.Y(n_846)
);

BUFx8_ASAP7_75t_L g847 ( 
.A(n_689),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_680),
.A2(n_600),
.B(n_521),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_680),
.A2(n_600),
.B(n_521),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_656),
.B(n_588),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_700),
.A2(n_548),
.B(n_529),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_654),
.A2(n_540),
.B1(n_546),
.B2(n_523),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_639),
.B(n_420),
.Y(n_853)
);

NOR3xp33_ASAP7_75t_L g854 ( 
.A(n_649),
.B(n_284),
.C(n_282),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_656),
.B(n_590),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_656),
.A2(n_552),
.B(n_529),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_694),
.B(n_590),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_650),
.B(n_523),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_712),
.B(n_718),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_694),
.A2(n_526),
.B(n_540),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_638),
.B(n_221),
.Y(n_861)
);

OAI22xp5_ASAP7_75t_L g862 ( 
.A1(n_718),
.A2(n_504),
.B1(n_532),
.B2(n_526),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_714),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_694),
.Y(n_864)
);

O2A1O1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_740),
.A2(n_543),
.B(n_541),
.C(n_544),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_644),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_694),
.B(n_590),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_722),
.B(n_702),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_722),
.B(n_541),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_724),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_668),
.A2(n_676),
.B1(n_762),
.B2(n_755),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_705),
.B(n_543),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_698),
.A2(n_544),
.B(n_545),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_620),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_765),
.B(n_454),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_639),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_698),
.A2(n_545),
.B(n_464),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_737),
.A2(n_545),
.B(n_464),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_SL g879 ( 
.A1(n_643),
.A2(n_247),
.B1(n_301),
.B2(n_286),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_737),
.A2(n_545),
.B(n_464),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_747),
.A2(n_545),
.B(n_464),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_604),
.A2(n_293),
.B1(n_292),
.B2(n_285),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_725),
.Y(n_883)
);

NOR3xp33_ASAP7_75t_L g884 ( 
.A(n_629),
.B(n_234),
.C(n_225),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_750),
.B(n_454),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_747),
.A2(n_464),
.B(n_545),
.Y(n_886)
);

BUFx8_ASAP7_75t_L g887 ( 
.A(n_689),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_696),
.B(n_590),
.Y(n_888)
);

AOI22xp33_ASAP7_75t_L g889 ( 
.A1(n_617),
.A2(n_247),
.B1(n_301),
.B2(n_462),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_644),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_770),
.B(n_467),
.Y(n_891)
);

NOR2x2_ASAP7_75t_L g892 ( 
.A(n_619),
.B(n_301),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_751),
.A2(n_464),
.B(n_479),
.Y(n_893)
);

OAI21xp5_ASAP7_75t_L g894 ( 
.A1(n_701),
.A2(n_479),
.B(n_486),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_751),
.A2(n_482),
.B(n_486),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_721),
.A2(n_502),
.B(n_482),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_721),
.A2(n_506),
.B(n_502),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_730),
.B(n_506),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_636),
.B(n_519),
.Y(n_899)
);

INVxp67_ASAP7_75t_L g900 ( 
.A(n_678),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_618),
.B(n_528),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_605),
.B(n_528),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_727),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_621),
.Y(n_904)
);

OAI22xp5_ASAP7_75t_L g905 ( 
.A1(n_668),
.A2(n_283),
.B1(n_279),
.B2(n_273),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_701),
.A2(n_591),
.B(n_590),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_651),
.Y(n_907)
);

A2O1A1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_713),
.A2(n_729),
.B(n_731),
.C(n_760),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_676),
.B(n_621),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_608),
.B(n_558),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_613),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_620),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_739),
.Y(n_913)
);

BUFx4f_ASAP7_75t_L g914 ( 
.A(n_692),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_635),
.Y(n_915)
);

INVx1_ASAP7_75t_SL g916 ( 
.A(n_663),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_719),
.A2(n_591),
.B(n_589),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_723),
.A2(n_591),
.B(n_589),
.Y(n_918)
);

NOR3xp33_ASAP7_75t_L g919 ( 
.A(n_645),
.B(n_223),
.C(n_237),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_664),
.B(n_562),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_723),
.A2(n_591),
.B(n_583),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_753),
.B(n_420),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_606),
.B(n_243),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_651),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_733),
.B(n_562),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_606),
.B(n_253),
.Y(n_926)
);

O2A1O1Ixp33_ASAP7_75t_SL g927 ( 
.A1(n_697),
.A2(n_583),
.B(n_569),
.C(n_567),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_659),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_660),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_728),
.A2(n_591),
.B(n_569),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_660),
.B(n_671),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_728),
.A2(n_706),
.B(n_707),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_671),
.B(n_685),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_606),
.Y(n_934)
);

O2A1O1Ixp5_ASAP7_75t_L g935 ( 
.A1(n_691),
.A2(n_567),
.B(n_565),
.C(n_563),
.Y(n_935)
);

NOR2xp67_ASAP7_75t_L g936 ( 
.A(n_766),
.B(n_66),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_659),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_685),
.B(n_563),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_703),
.A2(n_565),
.B(n_442),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_762),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_716),
.A2(n_442),
.B(n_420),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_683),
.A2(n_407),
.B(n_391),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_688),
.B(n_437),
.Y(n_943)
);

AOI21xp33_ASAP7_75t_L g944 ( 
.A1(n_768),
.A2(n_270),
.B(n_257),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_746),
.B(n_437),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_689),
.B(n_272),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_695),
.B(n_274),
.Y(n_947)
);

NAND2x1p5_ASAP7_75t_L g948 ( 
.A(n_771),
.B(n_442),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_734),
.A2(n_432),
.B(n_430),
.C(n_291),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_748),
.B(n_441),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_742),
.B(n_430),
.Y(n_951)
);

AOI21x1_ASAP7_75t_L g952 ( 
.A1(n_771),
.A2(n_410),
.B(n_409),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_743),
.A2(n_430),
.B(n_432),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_692),
.A2(n_301),
.B1(n_432),
.B2(n_430),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_773),
.B(n_432),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_772),
.A2(n_410),
.B1(n_395),
.B2(n_407),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_749),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_749),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_756),
.B(n_441),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_756),
.B(n_441),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_754),
.A2(n_418),
.B(n_410),
.C(n_409),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_786),
.Y(n_962)
);

AND3x1_ASAP7_75t_SL g963 ( 
.A(n_803),
.B(n_619),
.C(n_670),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_778),
.B(n_632),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_944),
.A2(n_715),
.B(n_691),
.C(n_634),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_804),
.B(n_670),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_777),
.B(n_659),
.Y(n_967)
);

BUFx4f_ASAP7_75t_L g968 ( 
.A(n_904),
.Y(n_968)
);

AOI22xp33_ASAP7_75t_L g969 ( 
.A1(n_854),
.A2(n_692),
.B1(n_682),
.B2(n_665),
.Y(n_969)
);

NOR2x1_ASAP7_75t_SL g970 ( 
.A(n_800),
.B(n_692),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_831),
.B(n_736),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_775),
.B(n_633),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_861),
.B(n_277),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_823),
.B(n_687),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_908),
.A2(n_640),
.B(n_758),
.C(n_752),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_780),
.Y(n_976)
);

NAND3xp33_ASAP7_75t_L g977 ( 
.A(n_879),
.B(n_288),
.C(n_297),
.Y(n_977)
);

NOR2x1_ASAP7_75t_L g978 ( 
.A(n_807),
.B(n_757),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_799),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_847),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_800),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_819),
.A2(n_745),
.B(n_759),
.Y(n_982)
);

INVx4_ASAP7_75t_L g983 ( 
.A(n_904),
.Y(n_983)
);

NAND2xp33_ASAP7_75t_SL g984 ( 
.A(n_934),
.B(n_720),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_811),
.A2(n_717),
.B1(n_726),
.B2(n_735),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_831),
.B(n_900),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_801),
.A2(n_732),
.B1(n_769),
.B2(n_764),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_908),
.A2(n_763),
.B1(n_767),
.B2(n_441),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_868),
.A2(n_441),
.B1(n_439),
.B2(n_437),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_914),
.A2(n_441),
.B1(n_439),
.B2(n_437),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_900),
.B(n_8),
.Y(n_991)
);

NAND2x1_ASAP7_75t_L g992 ( 
.A(n_800),
.B(n_409),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_914),
.A2(n_441),
.B1(n_439),
.B2(n_437),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_818),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_822),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_859),
.A2(n_441),
.B(n_437),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_904),
.B(n_439),
.Y(n_997)
);

INVx4_ASAP7_75t_L g998 ( 
.A(n_904),
.Y(n_998)
);

AO21x1_ASAP7_75t_L g999 ( 
.A1(n_817),
.A2(n_418),
.B(n_408),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_837),
.A2(n_408),
.B(n_395),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_802),
.A2(n_408),
.B(n_395),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_940),
.Y(n_1002)
);

OA22x2_ASAP7_75t_L g1003 ( 
.A1(n_947),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_1003)
);

NAND3xp33_ASAP7_75t_SL g1004 ( 
.A(n_884),
.B(n_418),
.C(n_407),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_774),
.A2(n_391),
.B(n_439),
.Y(n_1005)
);

OR2x2_ASAP7_75t_L g1006 ( 
.A(n_832),
.B(n_439),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_913),
.B(n_439),
.Y(n_1007)
);

BUFx4f_ASAP7_75t_L g1008 ( 
.A(n_874),
.Y(n_1008)
);

AOI221xp5_ASAP7_75t_L g1009 ( 
.A1(n_794),
.A2(n_439),
.B1(n_437),
.B2(n_15),
.C(n_17),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_923),
.B(n_9),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_829),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_SL g1012 ( 
.A1(n_916),
.A2(n_937),
.B1(n_940),
.B2(n_912),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_923),
.B(n_10),
.Y(n_1013)
);

INVx4_ASAP7_75t_L g1014 ( 
.A(n_800),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_788),
.A2(n_439),
.B(n_437),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_784),
.B(n_439),
.Y(n_1016)
);

CKINVDCx14_ASAP7_75t_R g1017 ( 
.A(n_928),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_853),
.Y(n_1018)
);

AO32x2_ASAP7_75t_L g1019 ( 
.A1(n_871),
.A2(n_15),
.A3(n_17),
.B1(n_22),
.B2(n_23),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_840),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_816),
.A2(n_440),
.B(n_150),
.Y(n_1021)
);

AO21x1_ASAP7_75t_L g1022 ( 
.A1(n_836),
.A2(n_24),
.B(n_25),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_926),
.B(n_24),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_853),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_858),
.A2(n_147),
.B1(n_141),
.B2(n_140),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_858),
.A2(n_25),
.B(n_26),
.C(n_30),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_913),
.B(n_106),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_872),
.A2(n_98),
.B1(n_95),
.B2(n_94),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_870),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_814),
.B(n_440),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_843),
.A2(n_83),
.B(n_81),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_852),
.A2(n_80),
.B1(n_77),
.B2(n_67),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_852),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_875),
.B(n_440),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_833),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_901),
.A2(n_440),
.B(n_36),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_794),
.A2(n_34),
.B(n_38),
.C(n_40),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_926),
.B(n_34),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_946),
.B(n_40),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_936),
.A2(n_42),
.B(n_43),
.C(n_45),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_847),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_946),
.B(n_45),
.Y(n_1042)
);

INVxp67_ASAP7_75t_L g1043 ( 
.A(n_863),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_932),
.A2(n_440),
.B(n_48),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_779),
.B(n_47),
.Y(n_1045)
);

INVx4_ASAP7_75t_L g1046 ( 
.A(n_833),
.Y(n_1046)
);

O2A1O1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_785),
.A2(n_48),
.B(n_49),
.C(n_50),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_913),
.B(n_51),
.Y(n_1048)
);

OR2x2_ASAP7_75t_L g1049 ( 
.A(n_883),
.B(n_51),
.Y(n_1049)
);

INVx4_ASAP7_75t_L g1050 ( 
.A(n_833),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_833),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_789),
.A2(n_53),
.B(n_55),
.C(n_59),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_864),
.A2(n_53),
.B1(n_55),
.B2(n_60),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_864),
.A2(n_60),
.B1(n_61),
.B2(n_440),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_789),
.B(n_440),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_913),
.B(n_440),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_785),
.A2(n_440),
.B(n_884),
.C(n_854),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_942),
.A2(n_440),
.B(n_906),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_903),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_885),
.B(n_440),
.Y(n_1060)
);

AOI221xp5_ASAP7_75t_L g1061 ( 
.A1(n_919),
.A2(n_954),
.B1(n_791),
.B2(n_889),
.C(n_809),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_862),
.A2(n_899),
.B(n_888),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_919),
.B(n_846),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_957),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_823),
.B(n_876),
.Y(n_1065)
);

NAND3xp33_ASAP7_75t_SL g1066 ( 
.A(n_795),
.B(n_791),
.C(n_954),
.Y(n_1066)
);

BUFx12f_ASAP7_75t_L g1067 ( 
.A(n_887),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_824),
.B(n_825),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_776),
.A2(n_850),
.B(n_867),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_876),
.B(n_911),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_826),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_864),
.B(n_882),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_864),
.B(n_911),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_776),
.A2(n_790),
.B(n_850),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_790),
.A2(n_842),
.B(n_867),
.Y(n_1075)
);

BUFx3_ASAP7_75t_L g1076 ( 
.A(n_887),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_922),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_842),
.A2(n_857),
.B(n_855),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_839),
.A2(n_809),
.B(n_949),
.C(n_798),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_SL g1080 ( 
.A(n_782),
.Y(n_1080)
);

AO32x2_ASAP7_75t_L g1081 ( 
.A1(n_841),
.A2(n_808),
.A3(n_815),
.B1(n_905),
.B2(n_839),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_915),
.B(n_792),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_909),
.A2(n_922),
.B1(n_820),
.B2(n_955),
.Y(n_1083)
);

AOI22x1_ASAP7_75t_L g1084 ( 
.A1(n_851),
.A2(n_939),
.B1(n_948),
.B2(n_873),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_924),
.Y(n_1085)
);

O2A1O1Ixp5_ASAP7_75t_L g1086 ( 
.A1(n_781),
.A2(n_949),
.B(n_941),
.C(n_787),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_929),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_909),
.B(n_955),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_828),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_951),
.B(n_796),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_R g1091 ( 
.A(n_952),
.B(n_820),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_958),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_806),
.A2(n_805),
.B(n_888),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_951),
.A2(n_866),
.B1(n_907),
.B2(n_890),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_898),
.A2(n_855),
.B1(n_857),
.B2(n_797),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_844),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_865),
.A2(n_953),
.B(n_897),
.C(n_896),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_948),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_931),
.B(n_933),
.Y(n_1099)
);

OAI22x1_ASAP7_75t_L g1100 ( 
.A1(n_892),
.A2(n_956),
.B1(n_889),
.B2(n_891),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_910),
.B(n_902),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_869),
.A2(n_827),
.B(n_845),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_925),
.B(n_920),
.Y(n_1103)
);

AND2x2_ASAP7_75t_SL g1104 ( 
.A(n_945),
.B(n_950),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_894),
.B(n_938),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_856),
.B(n_860),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_917),
.A2(n_930),
.B1(n_921),
.B2(n_918),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_835),
.A2(n_848),
.B(n_849),
.Y(n_1108)
);

AOI21x1_ASAP7_75t_L g1109 ( 
.A1(n_1000),
.A2(n_943),
.B(n_960),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_964),
.B(n_959),
.Y(n_1110)
);

AO31x2_ASAP7_75t_L g1111 ( 
.A1(n_999),
.A2(n_895),
.A3(n_838),
.B(n_893),
.Y(n_1111)
);

O2A1O1Ixp33_ASAP7_75t_SL g1112 ( 
.A1(n_1040),
.A2(n_961),
.B(n_821),
.C(n_783),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_983),
.Y(n_1113)
);

AO32x2_ASAP7_75t_L g1114 ( 
.A1(n_1033),
.A2(n_927),
.A3(n_935),
.B1(n_793),
.B2(n_877),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_966),
.B(n_986),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_995),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1011),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_SL g1118 ( 
.A1(n_1010),
.A2(n_878),
.B(n_886),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_964),
.B(n_972),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1020),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_1013),
.B(n_881),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1108),
.A2(n_1102),
.B(n_972),
.Y(n_1122)
);

AOI21x1_ASAP7_75t_SL g1123 ( 
.A1(n_1063),
.A2(n_927),
.B(n_880),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_1108),
.A2(n_830),
.B(n_834),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_SL g1125 ( 
.A1(n_1061),
.A2(n_810),
.B(n_812),
.C(n_813),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_1023),
.A2(n_1061),
.B(n_1039),
.C(n_1042),
.Y(n_1126)
);

AO31x2_ASAP7_75t_L g1127 ( 
.A1(n_1022),
.A2(n_1097),
.A3(n_1107),
.B(n_988),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_SL g1128 ( 
.A1(n_1044),
.A2(n_965),
.B(n_970),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_1084),
.A2(n_1015),
.B(n_1069),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_1015),
.A2(n_1074),
.B(n_1075),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1078),
.A2(n_982),
.B(n_1093),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_982),
.A2(n_1058),
.B(n_996),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1058),
.A2(n_1086),
.B(n_1106),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_968),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1102),
.A2(n_1062),
.B(n_1103),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_971),
.A2(n_1057),
.B(n_1038),
.C(n_1066),
.Y(n_1136)
);

AOI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1000),
.A2(n_1062),
.B(n_987),
.Y(n_1137)
);

INVx3_ASAP7_75t_L g1138 ( 
.A(n_983),
.Y(n_1138)
);

AOI221x1_ASAP7_75t_L g1139 ( 
.A1(n_1100),
.A2(n_1026),
.B1(n_1032),
.B2(n_1052),
.C(n_1036),
.Y(n_1139)
);

AO31x2_ASAP7_75t_L g1140 ( 
.A1(n_1095),
.A2(n_985),
.A3(n_1106),
.B(n_989),
.Y(n_1140)
);

NAND3xp33_ASAP7_75t_L g1141 ( 
.A(n_1045),
.B(n_977),
.C(n_991),
.Y(n_1141)
);

NOR2xp67_ASAP7_75t_L g1142 ( 
.A(n_1043),
.B(n_1059),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_998),
.Y(n_1143)
);

INVx1_ASAP7_75t_SL g1144 ( 
.A(n_1049),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1079),
.A2(n_975),
.B(n_1005),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1099),
.A2(n_1068),
.B(n_1016),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1037),
.A2(n_1048),
.B(n_967),
.C(n_1053),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1099),
.A2(n_1068),
.B(n_1016),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1101),
.A2(n_1105),
.B(n_1072),
.Y(n_1149)
);

INVx4_ASAP7_75t_L g1150 ( 
.A(n_968),
.Y(n_1150)
);

O2A1O1Ixp5_ASAP7_75t_L g1151 ( 
.A1(n_1031),
.A2(n_1027),
.B(n_1028),
.C(n_1021),
.Y(n_1151)
);

AO31x2_ASAP7_75t_L g1152 ( 
.A1(n_1005),
.A2(n_1021),
.A3(n_990),
.B(n_993),
.Y(n_1152)
);

AO21x2_ASAP7_75t_L g1153 ( 
.A1(n_1091),
.A2(n_1001),
.B(n_1004),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_969),
.A2(n_978),
.B(n_1030),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_SL g1155 ( 
.A1(n_1009),
.A2(n_1073),
.B(n_1065),
.C(n_1056),
.Y(n_1155)
);

OR2x2_ASAP7_75t_L g1156 ( 
.A(n_973),
.B(n_1029),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_SL g1157 ( 
.A1(n_1047),
.A2(n_1083),
.B(n_1090),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1090),
.B(n_1082),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_1098),
.A2(n_1001),
.B(n_992),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1009),
.A2(n_1003),
.B1(n_962),
.B2(n_1094),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1104),
.A2(n_1070),
.B(n_1030),
.Y(n_1161)
);

CKINVDCx20_ASAP7_75t_R g1162 ( 
.A(n_963),
.Y(n_1162)
);

OA21x2_ASAP7_75t_L g1163 ( 
.A1(n_1055),
.A2(n_1060),
.B(n_1034),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1085),
.Y(n_1164)
);

AOI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1007),
.A2(n_997),
.B(n_1055),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_SL g1166 ( 
.A1(n_1025),
.A2(n_1054),
.B(n_1088),
.Y(n_1166)
);

OAI21xp33_ASAP7_75t_L g1167 ( 
.A1(n_1003),
.A2(n_1018),
.B(n_1024),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1034),
.A2(n_1060),
.B(n_974),
.Y(n_1168)
);

CKINVDCx11_ASAP7_75t_R g1169 ( 
.A(n_1067),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1087),
.A2(n_1092),
.B1(n_1077),
.B2(n_1088),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1077),
.A2(n_994),
.B(n_976),
.C(n_1018),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_1008),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_974),
.B(n_979),
.Y(n_1173)
);

INVx2_ASAP7_75t_SL g1174 ( 
.A(n_1008),
.Y(n_1174)
);

INVx2_ASAP7_75t_SL g1175 ( 
.A(n_980),
.Y(n_1175)
);

A2O1A1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_984),
.A2(n_1024),
.B(n_1096),
.C(n_1064),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1006),
.A2(n_1089),
.B(n_1071),
.Y(n_1177)
);

AND2x6_ASAP7_75t_L g1178 ( 
.A(n_981),
.B(n_1035),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1089),
.Y(n_1179)
);

INVxp67_ASAP7_75t_L g1180 ( 
.A(n_1012),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1089),
.Y(n_1181)
);

INVx4_ASAP7_75t_L g1182 ( 
.A(n_981),
.Y(n_1182)
);

AO31x2_ASAP7_75t_L g1183 ( 
.A1(n_1081),
.A2(n_1050),
.A3(n_1014),
.B(n_1046),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1081),
.A2(n_1051),
.B(n_998),
.Y(n_1184)
);

INVx3_ASAP7_75t_L g1185 ( 
.A(n_1014),
.Y(n_1185)
);

O2A1O1Ixp5_ASAP7_75t_SL g1186 ( 
.A1(n_1051),
.A2(n_1019),
.B(n_981),
.C(n_1035),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1017),
.B(n_1019),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_1035),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1041),
.A2(n_1076),
.B(n_1080),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1080),
.A2(n_637),
.B(n_1108),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1108),
.A2(n_637),
.B(n_775),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1108),
.A2(n_932),
.B(n_1084),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1108),
.A2(n_637),
.B(n_775),
.Y(n_1193)
);

BUFx2_ASAP7_75t_L g1194 ( 
.A(n_1002),
.Y(n_1194)
);

AO31x2_ASAP7_75t_L g1195 ( 
.A1(n_999),
.A2(n_809),
.A3(n_1022),
.B(n_839),
.Y(n_1195)
);

AO31x2_ASAP7_75t_L g1196 ( 
.A1(n_999),
.A2(n_809),
.A3(n_1022),
.B(n_839),
.Y(n_1196)
);

OR2x2_ASAP7_75t_L g1197 ( 
.A(n_966),
.B(n_455),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1062),
.A2(n_637),
.B(n_675),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1010),
.A2(n_637),
.B(n_623),
.C(n_1013),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1010),
.A2(n_637),
.B1(n_643),
.B2(n_638),
.Y(n_1200)
);

INVx3_ASAP7_75t_SL g1201 ( 
.A(n_980),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_964),
.A2(n_637),
.B1(n_778),
.B2(n_508),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1108),
.A2(n_932),
.B(n_1084),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_983),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_966),
.B(n_637),
.Y(n_1205)
);

AO31x2_ASAP7_75t_L g1206 ( 
.A1(n_999),
.A2(n_809),
.A3(n_1022),
.B(n_839),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1108),
.A2(n_932),
.B(n_1084),
.Y(n_1207)
);

OAI22x1_ASAP7_75t_L g1208 ( 
.A1(n_1010),
.A2(n_637),
.B1(n_1023),
.B2(n_1013),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_995),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1108),
.A2(n_637),
.B(n_775),
.Y(n_1210)
);

AO31x2_ASAP7_75t_L g1211 ( 
.A1(n_999),
.A2(n_809),
.A3(n_1022),
.B(n_839),
.Y(n_1211)
);

INVx1_ASAP7_75t_SL g1212 ( 
.A(n_966),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_995),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1062),
.A2(n_637),
.B(n_675),
.Y(n_1214)
);

OR2x6_ASAP7_75t_L g1215 ( 
.A(n_1002),
.B(n_874),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_995),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1108),
.A2(n_637),
.B(n_775),
.Y(n_1217)
);

O2A1O1Ixp33_ASAP7_75t_SL g1218 ( 
.A1(n_1040),
.A2(n_794),
.B(n_908),
.C(n_1061),
.Y(n_1218)
);

BUFx2_ASAP7_75t_R g1219 ( 
.A(n_980),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1010),
.A2(n_637),
.B1(n_654),
.B2(n_1013),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1108),
.A2(n_637),
.B(n_775),
.Y(n_1221)
);

A2O1A1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1010),
.A2(n_637),
.B(n_623),
.C(n_1013),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_995),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_983),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1108),
.A2(n_932),
.B(n_1084),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1108),
.A2(n_932),
.B(n_1084),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_968),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1108),
.A2(n_932),
.B(n_1084),
.Y(n_1228)
);

AO31x2_ASAP7_75t_L g1229 ( 
.A1(n_999),
.A2(n_809),
.A3(n_1022),
.B(n_839),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_966),
.B(n_637),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_966),
.B(n_637),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_966),
.B(n_637),
.Y(n_1232)
);

OR2x6_ASAP7_75t_L g1233 ( 
.A(n_1002),
.B(n_874),
.Y(n_1233)
);

OAI221xp5_ASAP7_75t_L g1234 ( 
.A1(n_1010),
.A2(n_637),
.B1(n_1023),
.B2(n_1013),
.C(n_1039),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_995),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_995),
.Y(n_1236)
);

AO31x2_ASAP7_75t_L g1237 ( 
.A1(n_999),
.A2(n_809),
.A3(n_1022),
.B(n_839),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_968),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_995),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_1067),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_995),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1108),
.A2(n_932),
.B(n_1084),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1108),
.A2(n_738),
.B(n_656),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_966),
.B(n_637),
.Y(n_1244)
);

AOI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1010),
.A2(n_637),
.B1(n_643),
.B2(n_638),
.Y(n_1245)
);

AO22x1_ASAP7_75t_L g1246 ( 
.A1(n_1010),
.A2(n_637),
.B1(n_619),
.B2(n_1013),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_995),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1108),
.A2(n_932),
.B(n_1084),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1108),
.A2(n_932),
.B(n_1084),
.Y(n_1249)
);

AND2x4_ASAP7_75t_L g1250 ( 
.A(n_1018),
.B(n_1024),
.Y(n_1250)
);

O2A1O1Ixp33_ASAP7_75t_SL g1251 ( 
.A1(n_1040),
.A2(n_794),
.B(n_908),
.C(n_1061),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_SL g1252 ( 
.A1(n_1234),
.A2(n_1232),
.B1(n_1230),
.B2(n_1205),
.Y(n_1252)
);

BUFx12f_ASAP7_75t_L g1253 ( 
.A(n_1169),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1234),
.A2(n_1220),
.B1(n_1245),
.B2(n_1200),
.Y(n_1254)
);

INVx6_ASAP7_75t_L g1255 ( 
.A(n_1150),
.Y(n_1255)
);

OAI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1208),
.A2(n_1119),
.B1(n_1158),
.B2(n_1212),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1231),
.B(n_1115),
.Y(n_1257)
);

OAI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1119),
.A2(n_1158),
.B1(n_1212),
.B2(n_1141),
.Y(n_1258)
);

CKINVDCx11_ASAP7_75t_R g1259 ( 
.A(n_1201),
.Y(n_1259)
);

CKINVDCx16_ASAP7_75t_R g1260 ( 
.A(n_1162),
.Y(n_1260)
);

CKINVDCx20_ASAP7_75t_R g1261 ( 
.A(n_1240),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_SL g1262 ( 
.A1(n_1126),
.A2(n_1141),
.B(n_1199),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1134),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1194),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1120),
.Y(n_1265)
);

OAI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1144),
.A2(n_1202),
.B1(n_1197),
.B2(n_1160),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1244),
.A2(n_1157),
.B1(n_1167),
.B2(n_1144),
.Y(n_1267)
);

INVx6_ASAP7_75t_L g1268 ( 
.A(n_1150),
.Y(n_1268)
);

INVx2_ASAP7_75t_SL g1269 ( 
.A(n_1172),
.Y(n_1269)
);

OAI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1202),
.A2(n_1160),
.B1(n_1156),
.B2(n_1139),
.Y(n_1270)
);

INVx5_ASAP7_75t_L g1271 ( 
.A(n_1178),
.Y(n_1271)
);

BUFx12f_ASAP7_75t_L g1272 ( 
.A(n_1175),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_SL g1273 ( 
.A1(n_1187),
.A2(n_1246),
.B1(n_1145),
.B2(n_1180),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1209),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1222),
.A2(n_1136),
.B1(n_1142),
.B2(n_1233),
.Y(n_1275)
);

INVx6_ASAP7_75t_L g1276 ( 
.A(n_1134),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_SL g1277 ( 
.A1(n_1145),
.A2(n_1214),
.B1(n_1198),
.B2(n_1221),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_1174),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1213),
.Y(n_1279)
);

INVx6_ASAP7_75t_L g1280 ( 
.A(n_1134),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1227),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1215),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_SL g1283 ( 
.A1(n_1198),
.A2(n_1214),
.B1(n_1210),
.B2(n_1193),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1215),
.Y(n_1284)
);

BUFx8_ASAP7_75t_L g1285 ( 
.A(n_1227),
.Y(n_1285)
);

INVx4_ASAP7_75t_L g1286 ( 
.A(n_1227),
.Y(n_1286)
);

OAI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1121),
.A2(n_1170),
.B1(n_1149),
.B2(n_1190),
.Y(n_1287)
);

BUFx2_ASAP7_75t_SL g1288 ( 
.A(n_1238),
.Y(n_1288)
);

OAI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1166),
.A2(n_1116),
.B1(n_1235),
.B2(n_1247),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1215),
.A2(n_1233),
.B1(n_1128),
.B2(n_1176),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_SL g1291 ( 
.A(n_1219),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1117),
.Y(n_1292)
);

CKINVDCx6p67_ASAP7_75t_R g1293 ( 
.A(n_1238),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1216),
.Y(n_1294)
);

INVx6_ASAP7_75t_L g1295 ( 
.A(n_1238),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1233),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1190),
.A2(n_1154),
.B1(n_1153),
.B2(n_1168),
.Y(n_1297)
);

CKINVDCx11_ASAP7_75t_R g1298 ( 
.A(n_1219),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1154),
.A2(n_1153),
.B1(n_1168),
.B2(n_1250),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1223),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1173),
.B(n_1146),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1250),
.A2(n_1170),
.B1(n_1173),
.B2(n_1161),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1183),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1236),
.Y(n_1304)
);

CKINVDCx20_ASAP7_75t_R g1305 ( 
.A(n_1189),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_SL g1306 ( 
.A1(n_1191),
.A2(n_1221),
.B1(n_1193),
.B2(n_1210),
.Y(n_1306)
);

CKINVDCx11_ASAP7_75t_R g1307 ( 
.A(n_1188),
.Y(n_1307)
);

CKINVDCx20_ASAP7_75t_R g1308 ( 
.A(n_1189),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1166),
.A2(n_1239),
.B1(n_1241),
.B2(n_1164),
.Y(n_1309)
);

INVx4_ASAP7_75t_SL g1310 ( 
.A(n_1178),
.Y(n_1310)
);

BUFx10_ASAP7_75t_L g1311 ( 
.A(n_1179),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1181),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1191),
.A2(n_1217),
.B1(n_1163),
.B2(n_1135),
.Y(n_1313)
);

CKINVDCx11_ASAP7_75t_R g1314 ( 
.A(n_1188),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_SL g1315 ( 
.A1(n_1217),
.A2(n_1186),
.B1(n_1251),
.B2(n_1218),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_SL g1316 ( 
.A1(n_1131),
.A2(n_1122),
.B1(n_1110),
.B2(n_1148),
.Y(n_1316)
);

INVx4_ASAP7_75t_L g1317 ( 
.A(n_1178),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_SL g1318 ( 
.A1(n_1110),
.A2(n_1184),
.B1(n_1124),
.B2(n_1147),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1171),
.A2(n_1118),
.B1(n_1177),
.B2(n_1243),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1188),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1118),
.A2(n_1155),
.B1(n_1224),
.B2(n_1143),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1163),
.A2(n_1184),
.B1(n_1224),
.B2(n_1204),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1113),
.A2(n_1143),
.B1(n_1204),
.B2(n_1138),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1182),
.Y(n_1324)
);

OAI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1137),
.A2(n_1138),
.B1(n_1185),
.B2(n_1165),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1133),
.A2(n_1185),
.B1(n_1159),
.B2(n_1182),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1132),
.A2(n_1130),
.B1(n_1178),
.B2(n_1249),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1123),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1183),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_1127),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1192),
.A2(n_1248),
.B1(n_1242),
.B2(n_1207),
.Y(n_1331)
);

NAND2x1p5_ASAP7_75t_L g1332 ( 
.A(n_1203),
.B(n_1225),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1226),
.A2(n_1228),
.B1(n_1129),
.B2(n_1151),
.Y(n_1333)
);

OAI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1109),
.A2(n_1127),
.B1(n_1140),
.B2(n_1237),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1127),
.B(n_1140),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1140),
.B(n_1237),
.Y(n_1336)
);

OAI22x1_ASAP7_75t_SL g1337 ( 
.A1(n_1195),
.A2(n_1196),
.B1(n_1229),
.B2(n_1211),
.Y(n_1337)
);

CKINVDCx20_ASAP7_75t_R g1338 ( 
.A(n_1125),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_SL g1339 ( 
.A1(n_1112),
.A2(n_1206),
.B1(n_1229),
.B2(n_1211),
.Y(n_1339)
);

OAI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1196),
.A2(n_1206),
.B1(n_1211),
.B2(n_1229),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1206),
.A2(n_1237),
.B1(n_1114),
.B2(n_1152),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1114),
.A2(n_1234),
.B1(n_1220),
.B2(n_637),
.Y(n_1342)
);

BUFx8_ASAP7_75t_L g1343 ( 
.A(n_1114),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1111),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_1111),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1152),
.A2(n_1234),
.B1(n_637),
.B2(n_1220),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1152),
.A2(n_1234),
.B1(n_1245),
.B2(n_1200),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1111),
.A2(n_1234),
.B1(n_637),
.B2(n_1220),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1234),
.A2(n_637),
.B1(n_1220),
.B2(n_1200),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1234),
.A2(n_637),
.B1(n_1220),
.B2(n_1200),
.Y(n_1350)
);

INVx6_ASAP7_75t_L g1351 ( 
.A(n_1150),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1120),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1234),
.A2(n_637),
.B1(n_1220),
.B2(n_1200),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_SL g1354 ( 
.A1(n_1234),
.A2(n_637),
.B1(n_421),
.B2(n_445),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_SL g1355 ( 
.A1(n_1234),
.A2(n_637),
.B1(n_421),
.B2(n_445),
.Y(n_1355)
);

CKINVDCx20_ASAP7_75t_R g1356 ( 
.A(n_1169),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1234),
.A2(n_637),
.B1(n_421),
.B2(n_445),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1234),
.A2(n_637),
.B1(n_1220),
.B2(n_1200),
.Y(n_1358)
);

CKINVDCx11_ASAP7_75t_R g1359 ( 
.A(n_1169),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1234),
.A2(n_1200),
.B1(n_1245),
.B2(n_637),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1169),
.Y(n_1361)
);

BUFx4f_ASAP7_75t_L g1362 ( 
.A(n_1134),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_1169),
.Y(n_1363)
);

INVx6_ASAP7_75t_L g1364 ( 
.A(n_1150),
.Y(n_1364)
);

INVx6_ASAP7_75t_L g1365 ( 
.A(n_1150),
.Y(n_1365)
);

OAI21xp33_ASAP7_75t_L g1366 ( 
.A1(n_1200),
.A2(n_637),
.B(n_1245),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1234),
.A2(n_1200),
.B1(n_1245),
.B2(n_637),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1120),
.Y(n_1368)
);

OAI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1234),
.A2(n_1245),
.B1(n_1200),
.B2(n_637),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1120),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1120),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1234),
.A2(n_637),
.B1(n_1220),
.B2(n_1200),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1120),
.Y(n_1373)
);

AOI22x1_ASAP7_75t_SL g1374 ( 
.A1(n_1240),
.A2(n_934),
.B1(n_670),
.B2(n_937),
.Y(n_1374)
);

BUFx4f_ASAP7_75t_SL g1375 ( 
.A(n_1172),
.Y(n_1375)
);

BUFx12f_ASAP7_75t_L g1376 ( 
.A(n_1169),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1120),
.Y(n_1377)
);

INVx6_ASAP7_75t_L g1378 ( 
.A(n_1150),
.Y(n_1378)
);

OAI21xp33_ASAP7_75t_L g1379 ( 
.A1(n_1200),
.A2(n_637),
.B(n_1245),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1120),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1339),
.B(n_1273),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1332),
.A2(n_1333),
.B(n_1331),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1257),
.B(n_1252),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1344),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1299),
.B(n_1345),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_1282),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_1359),
.Y(n_1387)
);

AO21x1_ASAP7_75t_L g1388 ( 
.A1(n_1360),
.A2(n_1367),
.B(n_1369),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1339),
.B(n_1273),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1332),
.A2(n_1327),
.B(n_1313),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1329),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1336),
.B(n_1335),
.Y(n_1392)
);

INVx4_ASAP7_75t_L g1393 ( 
.A(n_1271),
.Y(n_1393)
);

OAI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1366),
.A2(n_1379),
.B(n_1369),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1318),
.B(n_1330),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_1284),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1303),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1303),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1343),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1338),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1330),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1301),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1337),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1341),
.B(n_1340),
.Y(n_1404)
);

AO21x2_ASAP7_75t_L g1405 ( 
.A1(n_1325),
.A2(n_1334),
.B(n_1340),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_1328),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1300),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1319),
.A2(n_1326),
.B(n_1297),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_SL g1409 ( 
.A(n_1296),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1304),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1292),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_SL g1412 ( 
.A(n_1252),
.B(n_1349),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1294),
.Y(n_1413)
);

AND2x4_ASAP7_75t_L g1414 ( 
.A(n_1321),
.B(n_1322),
.Y(n_1414)
);

OA21x2_ASAP7_75t_L g1415 ( 
.A1(n_1262),
.A2(n_1342),
.B(n_1348),
.Y(n_1415)
);

OAI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1350),
.A2(n_1358),
.B(n_1353),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1334),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1372),
.A2(n_1354),
.B(n_1355),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1309),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1254),
.A2(n_1354),
.B1(n_1355),
.B2(n_1357),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1312),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1318),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1290),
.A2(n_1302),
.B(n_1275),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1277),
.B(n_1347),
.Y(n_1424)
);

AO21x2_ASAP7_75t_L g1425 ( 
.A1(n_1325),
.A2(n_1289),
.B(n_1270),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1316),
.A2(n_1277),
.B(n_1306),
.Y(n_1426)
);

BUFx8_ASAP7_75t_SL g1427 ( 
.A(n_1253),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1287),
.Y(n_1428)
);

INVx3_ASAP7_75t_L g1429 ( 
.A(n_1271),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1265),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_1259),
.Y(n_1431)
);

INVx3_ASAP7_75t_L g1432 ( 
.A(n_1271),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1274),
.Y(n_1433)
);

NAND2xp33_ASAP7_75t_R g1434 ( 
.A(n_1374),
.B(n_1361),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_1311),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1279),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1352),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1371),
.Y(n_1438)
);

CKINVDCx20_ASAP7_75t_R g1439 ( 
.A(n_1356),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1342),
.B(n_1283),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1377),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1283),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1310),
.B(n_1380),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1306),
.Y(n_1444)
);

BUFx3_ASAP7_75t_L g1445 ( 
.A(n_1255),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1357),
.B(n_1258),
.Y(n_1446)
);

OR2x6_ASAP7_75t_L g1447 ( 
.A(n_1317),
.B(n_1255),
.Y(n_1447)
);

BUFx6f_ASAP7_75t_L g1448 ( 
.A(n_1311),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1258),
.B(n_1256),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1316),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1346),
.A2(n_1266),
.B1(n_1270),
.B2(n_1267),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1368),
.A2(n_1373),
.B(n_1370),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1289),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1315),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1315),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1264),
.B(n_1320),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1324),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1256),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1266),
.B(n_1305),
.Y(n_1459)
);

AND2x4_ASAP7_75t_L g1460 ( 
.A(n_1310),
.B(n_1286),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1263),
.B(n_1281),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1323),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1263),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1260),
.B(n_1269),
.Y(n_1464)
);

NAND2x1p5_ASAP7_75t_L g1465 ( 
.A(n_1286),
.B(n_1281),
.Y(n_1465)
);

OAI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1308),
.A2(n_1362),
.B(n_1278),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1298),
.A2(n_1378),
.B1(n_1351),
.B2(n_1268),
.Y(n_1467)
);

OAI21xp33_ASAP7_75t_SL g1468 ( 
.A1(n_1291),
.A2(n_1362),
.B(n_1288),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1351),
.Y(n_1469)
);

OR2x6_ASAP7_75t_L g1470 ( 
.A(n_1364),
.B(n_1378),
.Y(n_1470)
);

AOI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1420),
.A2(n_1291),
.B1(n_1365),
.B2(n_1378),
.Y(n_1471)
);

AND2x4_ASAP7_75t_L g1472 ( 
.A(n_1386),
.B(n_1261),
.Y(n_1472)
);

A2O1A1Ixp33_ASAP7_75t_L g1473 ( 
.A1(n_1420),
.A2(n_1418),
.B(n_1416),
.C(n_1394),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1427),
.Y(n_1474)
);

OR2x6_ASAP7_75t_L g1475 ( 
.A(n_1423),
.B(n_1365),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1386),
.B(n_1314),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1442),
.B(n_1293),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1396),
.B(n_1307),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1411),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1412),
.A2(n_1363),
.B(n_1375),
.Y(n_1480)
);

O2A1O1Ixp33_ASAP7_75t_SL g1481 ( 
.A1(n_1446),
.A2(n_1285),
.B(n_1376),
.C(n_1375),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1413),
.B(n_1285),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1451),
.A2(n_1276),
.B1(n_1280),
.B2(n_1295),
.Y(n_1483)
);

AO32x2_ASAP7_75t_L g1484 ( 
.A1(n_1435),
.A2(n_1276),
.A3(n_1280),
.B1(n_1295),
.B2(n_1272),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_1439),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1442),
.B(n_1276),
.Y(n_1486)
);

AOI211xp5_ASAP7_75t_L g1487 ( 
.A1(n_1388),
.A2(n_1280),
.B(n_1295),
.C(n_1383),
.Y(n_1487)
);

O2A1O1Ixp33_ASAP7_75t_SL g1488 ( 
.A1(n_1459),
.A2(n_1466),
.B(n_1435),
.C(n_1403),
.Y(n_1488)
);

AO32x2_ASAP7_75t_L g1489 ( 
.A1(n_1393),
.A2(n_1404),
.A3(n_1392),
.B1(n_1403),
.B2(n_1458),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1444),
.B(n_1402),
.Y(n_1490)
);

INVx5_ASAP7_75t_L g1491 ( 
.A(n_1447),
.Y(n_1491)
);

O2A1O1Ixp33_ASAP7_75t_L g1492 ( 
.A1(n_1388),
.A2(n_1426),
.B(n_1428),
.C(n_1449),
.Y(n_1492)
);

AOI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1415),
.A2(n_1424),
.B1(n_1440),
.B2(n_1381),
.Y(n_1493)
);

OAI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1423),
.A2(n_1424),
.B(n_1428),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1400),
.A2(n_1406),
.B1(n_1449),
.B2(n_1467),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1387),
.Y(n_1496)
);

O2A1O1Ixp33_ASAP7_75t_L g1497 ( 
.A1(n_1453),
.A2(n_1422),
.B(n_1444),
.C(n_1458),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1421),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1456),
.B(n_1399),
.Y(n_1499)
);

A2O1A1Ixp33_ASAP7_75t_L g1500 ( 
.A1(n_1440),
.A2(n_1453),
.B(n_1414),
.C(n_1389),
.Y(n_1500)
);

A2O1A1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1414),
.A2(n_1381),
.B(n_1389),
.C(n_1408),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1400),
.A2(n_1406),
.B1(n_1415),
.B2(n_1422),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1402),
.B(n_1437),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1457),
.Y(n_1504)
);

OA21x2_ASAP7_75t_L g1505 ( 
.A1(n_1408),
.A2(n_1382),
.B(n_1390),
.Y(n_1505)
);

INVx1_ASAP7_75t_SL g1506 ( 
.A(n_1463),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1407),
.Y(n_1507)
);

BUFx3_ASAP7_75t_L g1508 ( 
.A(n_1464),
.Y(n_1508)
);

AOI221xp5_ASAP7_75t_L g1509 ( 
.A1(n_1419),
.A2(n_1450),
.B1(n_1454),
.B2(n_1455),
.C(n_1462),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1441),
.B(n_1461),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1464),
.B(n_1431),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1410),
.B(n_1450),
.Y(n_1512)
);

NOR4xp25_ASAP7_75t_SL g1513 ( 
.A(n_1434),
.B(n_1455),
.C(n_1454),
.D(n_1419),
.Y(n_1513)
);

A2O1A1Ixp33_ASAP7_75t_L g1514 ( 
.A1(n_1414),
.A2(n_1468),
.B(n_1395),
.C(n_1385),
.Y(n_1514)
);

OAI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1415),
.A2(n_1390),
.B(n_1468),
.Y(n_1515)
);

OAI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1452),
.A2(n_1382),
.B(n_1395),
.Y(n_1516)
);

OR2x6_ASAP7_75t_L g1517 ( 
.A(n_1447),
.B(n_1470),
.Y(n_1517)
);

AO32x2_ASAP7_75t_L g1518 ( 
.A1(n_1393),
.A2(n_1425),
.A3(n_1397),
.B1(n_1398),
.B2(n_1405),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_SL g1519 ( 
.A1(n_1470),
.A2(n_1447),
.B1(n_1443),
.B2(n_1469),
.Y(n_1519)
);

AOI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1425),
.A2(n_1409),
.B1(n_1443),
.B2(n_1447),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1489),
.Y(n_1521)
);

CKINVDCx20_ASAP7_75t_R g1522 ( 
.A(n_1474),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1507),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1516),
.B(n_1505),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_1473),
.B(n_1448),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1498),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1516),
.B(n_1505),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1471),
.A2(n_1405),
.B1(n_1417),
.B2(n_1409),
.Y(n_1528)
);

NOR2x1_ASAP7_75t_R g1529 ( 
.A(n_1496),
.B(n_1460),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_1485),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1518),
.B(n_1405),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1479),
.Y(n_1532)
);

BUFx6f_ASAP7_75t_L g1533 ( 
.A(n_1518),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1493),
.B(n_1417),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1518),
.B(n_1405),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_SL g1536 ( 
.A1(n_1502),
.A2(n_1409),
.B1(n_1432),
.B2(n_1429),
.Y(n_1536)
);

NAND3xp33_ASAP7_75t_L g1537 ( 
.A(n_1487),
.B(n_1430),
.C(n_1433),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_1484),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1512),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1471),
.A2(n_1409),
.B1(n_1430),
.B2(n_1433),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1490),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1489),
.B(n_1384),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1480),
.A2(n_1493),
.B1(n_1494),
.B2(n_1509),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1487),
.A2(n_1470),
.B1(n_1438),
.B2(n_1436),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1503),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1506),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1510),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1515),
.B(n_1384),
.Y(n_1548)
);

OAI221xp5_ASAP7_75t_L g1549 ( 
.A1(n_1543),
.A2(n_1480),
.B1(n_1492),
.B2(n_1501),
.C(n_1500),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1548),
.B(n_1491),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_SL g1551 ( 
.A1(n_1537),
.A2(n_1495),
.B1(n_1515),
.B2(n_1508),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1545),
.B(n_1504),
.Y(n_1552)
);

BUFx2_ASAP7_75t_L g1553 ( 
.A(n_1538),
.Y(n_1553)
);

OAI221xp5_ASAP7_75t_L g1554 ( 
.A1(n_1543),
.A2(n_1514),
.B1(n_1488),
.B2(n_1520),
.C(n_1497),
.Y(n_1554)
);

OAI221xp5_ASAP7_75t_L g1555 ( 
.A1(n_1525),
.A2(n_1520),
.B1(n_1477),
.B2(n_1481),
.C(n_1482),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1546),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1525),
.A2(n_1472),
.B1(n_1475),
.B2(n_1486),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1523),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1521),
.B(n_1401),
.Y(n_1559)
);

INVx4_ASAP7_75t_L g1560 ( 
.A(n_1538),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1523),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1542),
.Y(n_1562)
);

AND2x4_ASAP7_75t_SL g1563 ( 
.A(n_1538),
.B(n_1517),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1523),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1521),
.B(n_1391),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1532),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1546),
.Y(n_1567)
);

NOR2xp67_ASAP7_75t_SL g1568 ( 
.A(n_1537),
.B(n_1432),
.Y(n_1568)
);

BUFx2_ASAP7_75t_L g1569 ( 
.A(n_1538),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1533),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_SL g1571 ( 
.A(n_1529),
.B(n_1519),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1547),
.B(n_1499),
.Y(n_1572)
);

NOR3xp33_ASAP7_75t_SL g1573 ( 
.A(n_1549),
.B(n_1530),
.C(n_1511),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_R g1574 ( 
.A(n_1571),
.B(n_1522),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1556),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1558),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1558),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1561),
.Y(n_1578)
);

INVx4_ASAP7_75t_L g1579 ( 
.A(n_1560),
.Y(n_1579)
);

AND2x2_ASAP7_75t_SL g1580 ( 
.A(n_1571),
.B(n_1538),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1556),
.B(n_1539),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1561),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1566),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1564),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1562),
.B(n_1538),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1564),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1567),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1550),
.B(n_1524),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1562),
.B(n_1538),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1567),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1570),
.B(n_1533),
.Y(n_1591)
);

OAI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1551),
.A2(n_1528),
.B1(n_1536),
.B2(n_1540),
.C(n_1544),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1562),
.B(n_1538),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1570),
.B(n_1533),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1565),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1555),
.B(n_1549),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1562),
.B(n_1538),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1550),
.B(n_1524),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1552),
.B(n_1539),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1551),
.B(n_1544),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1552),
.B(n_1539),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1553),
.B(n_1524),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1553),
.B(n_1527),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1553),
.B(n_1569),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1566),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1570),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1569),
.B(n_1527),
.Y(n_1607)
);

INVx2_ASAP7_75t_SL g1608 ( 
.A(n_1579),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1580),
.B(n_1588),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1576),
.Y(n_1610)
);

INVxp67_ASAP7_75t_SL g1611 ( 
.A(n_1575),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1576),
.Y(n_1612)
);

NOR2x1_ASAP7_75t_L g1613 ( 
.A(n_1579),
.B(n_1522),
.Y(n_1613)
);

OAI21xp33_ASAP7_75t_L g1614 ( 
.A1(n_1596),
.A2(n_1554),
.B(n_1531),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1596),
.A2(n_1554),
.B1(n_1555),
.B2(n_1568),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1599),
.B(n_1570),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1591),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1591),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1577),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1577),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1600),
.B(n_1526),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1599),
.B(n_1559),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1578),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_SL g1624 ( 
.A(n_1580),
.B(n_1529),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1591),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1580),
.B(n_1569),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1588),
.B(n_1560),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1578),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1582),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1594),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1582),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1584),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1584),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1586),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1586),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1601),
.B(n_1526),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1601),
.B(n_1541),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1575),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1573),
.B(n_1541),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1573),
.B(n_1541),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1587),
.Y(n_1641)
);

OAI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1592),
.A2(n_1568),
.B(n_1557),
.Y(n_1642)
);

OAI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1592),
.A2(n_1568),
.B(n_1557),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1581),
.B(n_1559),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1587),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1581),
.B(n_1572),
.Y(n_1646)
);

INVx2_ASAP7_75t_SL g1647 ( 
.A(n_1579),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1590),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1590),
.B(n_1572),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1611),
.B(n_1594),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1610),
.Y(n_1651)
);

NAND3xp33_ASAP7_75t_L g1652 ( 
.A(n_1615),
.B(n_1533),
.C(n_1560),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1610),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1609),
.B(n_1604),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1638),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1609),
.B(n_1604),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1626),
.B(n_1604),
.Y(n_1657)
);

AOI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1614),
.A2(n_1534),
.B(n_1530),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1621),
.B(n_1574),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1626),
.B(n_1579),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1642),
.B(n_1560),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1645),
.B(n_1594),
.Y(n_1662)
);

OAI21xp33_ASAP7_75t_L g1663 ( 
.A1(n_1643),
.A2(n_1624),
.B(n_1639),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1619),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1613),
.B(n_1579),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1619),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1627),
.B(n_1588),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1640),
.B(n_1472),
.Y(n_1668)
);

NAND3xp33_ASAP7_75t_L g1669 ( 
.A(n_1648),
.B(n_1533),
.C(n_1560),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1627),
.B(n_1588),
.Y(n_1670)
);

CKINVDCx16_ASAP7_75t_R g1671 ( 
.A(n_1608),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1638),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1636),
.B(n_1602),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1620),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1649),
.B(n_1646),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1641),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1620),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1648),
.B(n_1602),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1617),
.B(n_1595),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1608),
.B(n_1588),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1617),
.B(n_1595),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1647),
.B(n_1598),
.Y(n_1682)
);

INVx3_ASAP7_75t_SL g1683 ( 
.A(n_1647),
.Y(n_1683)
);

AND2x4_ASAP7_75t_SL g1684 ( 
.A(n_1641),
.B(n_1476),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1655),
.Y(n_1685)
);

OAI21xp33_ASAP7_75t_L g1686 ( 
.A1(n_1663),
.A2(n_1534),
.B(n_1531),
.Y(n_1686)
);

NOR4xp25_ASAP7_75t_L g1687 ( 
.A(n_1663),
.B(n_1618),
.C(n_1625),
.D(n_1630),
.Y(n_1687)
);

AOI32xp33_ASAP7_75t_L g1688 ( 
.A1(n_1661),
.A2(n_1602),
.A3(n_1603),
.B1(n_1607),
.B2(n_1598),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1658),
.B(n_1618),
.Y(n_1689)
);

OAI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1652),
.A2(n_1665),
.B(n_1659),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1668),
.B(n_1625),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1665),
.B(n_1671),
.Y(n_1692)
);

AOI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1652),
.A2(n_1563),
.B1(n_1535),
.B2(n_1598),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1672),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1676),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1650),
.Y(n_1696)
);

AOI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1669),
.A2(n_1533),
.B1(n_1630),
.B2(n_1607),
.C(n_1603),
.Y(n_1697)
);

AOI21xp33_ASAP7_75t_L g1698 ( 
.A1(n_1650),
.A2(n_1616),
.B(n_1623),
.Y(n_1698)
);

OAI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1660),
.A2(n_1628),
.B(n_1612),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1651),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1651),
.Y(n_1701)
);

INVxp67_ASAP7_75t_L g1702 ( 
.A(n_1653),
.Y(n_1702)
);

NOR2x1_ASAP7_75t_L g1703 ( 
.A(n_1653),
.B(n_1623),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1684),
.B(n_1637),
.Y(n_1704)
);

AOI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1660),
.A2(n_1563),
.B1(n_1535),
.B2(n_1598),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1684),
.B(n_1616),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1664),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1657),
.B(n_1598),
.Y(n_1708)
);

OAI21xp33_ASAP7_75t_L g1709 ( 
.A1(n_1657),
.A2(n_1535),
.B(n_1603),
.Y(n_1709)
);

O2A1O1Ixp5_ASAP7_75t_SL g1710 ( 
.A1(n_1702),
.A2(n_1677),
.B(n_1674),
.C(n_1666),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1696),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1696),
.Y(n_1712)
);

OAI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1687),
.A2(n_1662),
.B(n_1678),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1708),
.B(n_1671),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1703),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1700),
.Y(n_1716)
);

OAI31xp33_ASAP7_75t_L g1717 ( 
.A1(n_1686),
.A2(n_1682),
.A3(n_1680),
.B(n_1656),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1685),
.B(n_1654),
.Y(n_1718)
);

OAI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1693),
.A2(n_1683),
.B1(n_1654),
.B2(n_1656),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1701),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1694),
.Y(n_1721)
);

NOR3xp33_ASAP7_75t_SL g1722 ( 
.A(n_1692),
.B(n_1673),
.C(n_1666),
.Y(n_1722)
);

AOI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1706),
.A2(n_1682),
.B1(n_1680),
.B2(n_1670),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1690),
.B(n_1689),
.Y(n_1724)
);

NAND4xp25_ASAP7_75t_SL g1725 ( 
.A(n_1688),
.B(n_1667),
.C(n_1670),
.D(n_1675),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1695),
.B(n_1667),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1707),
.Y(n_1727)
);

OAI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1699),
.A2(n_1662),
.B(n_1681),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1711),
.Y(n_1729)
);

XOR2xp5_ASAP7_75t_L g1730 ( 
.A(n_1719),
.B(n_1691),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1726),
.B(n_1706),
.Y(n_1731)
);

INVxp67_ASAP7_75t_SL g1732 ( 
.A(n_1712),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1714),
.B(n_1704),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1718),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1721),
.B(n_1702),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1721),
.Y(n_1736)
);

XNOR2x1_ASAP7_75t_L g1737 ( 
.A(n_1726),
.B(n_1478),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1728),
.B(n_1675),
.Y(n_1738)
);

AOI211xp5_ASAP7_75t_SL g1739 ( 
.A1(n_1715),
.A2(n_1698),
.B(n_1697),
.C(n_1709),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1724),
.B(n_1683),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_SL g1741 ( 
.A(n_1740),
.B(n_1714),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1732),
.Y(n_1742)
);

AOI21xp33_ASAP7_75t_SL g1743 ( 
.A1(n_1731),
.A2(n_1724),
.B(n_1683),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1737),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1738),
.B(n_1713),
.Y(n_1745)
);

NAND4xp25_ASAP7_75t_L g1746 ( 
.A(n_1733),
.B(n_1723),
.C(n_1726),
.D(n_1717),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1734),
.B(n_1722),
.Y(n_1747)
);

AO21x1_ASAP7_75t_L g1748 ( 
.A1(n_1735),
.A2(n_1710),
.B(n_1716),
.Y(n_1748)
);

AOI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1735),
.A2(n_1727),
.B(n_1720),
.Y(n_1749)
);

HB1xp67_ASAP7_75t_L g1750 ( 
.A(n_1736),
.Y(n_1750)
);

NOR4xp25_ASAP7_75t_L g1751 ( 
.A(n_1745),
.B(n_1729),
.C(n_1725),
.D(n_1710),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1744),
.B(n_1730),
.Y(n_1752)
);

AOI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1746),
.A2(n_1741),
.B1(n_1747),
.B2(n_1748),
.Y(n_1753)
);

AOI221xp5_ASAP7_75t_L g1754 ( 
.A1(n_1743),
.A2(n_1742),
.B1(n_1749),
.B2(n_1750),
.C(n_1739),
.Y(n_1754)
);

AOI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1749),
.A2(n_1739),
.B(n_1677),
.Y(n_1755)
);

O2A1O1Ixp33_ASAP7_75t_L g1756 ( 
.A1(n_1755),
.A2(n_1674),
.B(n_1664),
.C(n_1679),
.Y(n_1756)
);

XNOR2xp5_ASAP7_75t_L g1757 ( 
.A(n_1753),
.B(n_1705),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1752),
.Y(n_1758)
);

AOI32xp33_ASAP7_75t_L g1759 ( 
.A1(n_1754),
.A2(n_1751),
.A3(n_1607),
.B1(n_1597),
.B2(n_1593),
.Y(n_1759)
);

OAI211xp5_ASAP7_75t_L g1760 ( 
.A1(n_1751),
.A2(n_1681),
.B(n_1679),
.C(n_1513),
.Y(n_1760)
);

OAI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1753),
.A2(n_1644),
.B1(n_1635),
.B2(n_1634),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1756),
.Y(n_1762)
);

NOR2xp67_ASAP7_75t_L g1763 ( 
.A(n_1758),
.B(n_1761),
.Y(n_1763)
);

NAND2x1p5_ASAP7_75t_L g1764 ( 
.A(n_1759),
.B(n_1445),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1757),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1760),
.Y(n_1766)
);

AND4x1_ASAP7_75t_L g1767 ( 
.A(n_1765),
.B(n_1540),
.C(n_1528),
.D(n_1633),
.Y(n_1767)
);

NAND3xp33_ASAP7_75t_SL g1768 ( 
.A(n_1762),
.B(n_1513),
.C(n_1536),
.Y(n_1768)
);

INVx1_ASAP7_75t_SL g1769 ( 
.A(n_1764),
.Y(n_1769)
);

XNOR2x1_ASAP7_75t_L g1770 ( 
.A(n_1769),
.B(n_1763),
.Y(n_1770)
);

AOI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1770),
.A2(n_1766),
.B1(n_1763),
.B2(n_1768),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1771),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1771),
.A2(n_1767),
.B1(n_1629),
.B2(n_1633),
.Y(n_1773)
);

NOR3x1_ASAP7_75t_L g1774 ( 
.A(n_1772),
.B(n_1629),
.C(n_1644),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1773),
.B(n_1606),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1775),
.A2(n_1606),
.B1(n_1632),
.B2(n_1631),
.Y(n_1776)
);

XNOR2xp5_ASAP7_75t_L g1777 ( 
.A(n_1774),
.B(n_1460),
.Y(n_1777)
);

AOI221x1_ASAP7_75t_L g1778 ( 
.A1(n_1777),
.A2(n_1776),
.B1(n_1583),
.B2(n_1605),
.C(n_1597),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1778),
.B(n_1622),
.Y(n_1779)
);

AOI22x1_ASAP7_75t_L g1780 ( 
.A1(n_1779),
.A2(n_1465),
.B1(n_1460),
.B2(n_1622),
.Y(n_1780)
);

OAI221xp5_ASAP7_75t_R g1781 ( 
.A1(n_1780),
.A2(n_1589),
.B1(n_1597),
.B2(n_1593),
.C(n_1585),
.Y(n_1781)
);

AOI211xp5_ASAP7_75t_L g1782 ( 
.A1(n_1781),
.A2(n_1483),
.B(n_1460),
.C(n_1445),
.Y(n_1782)
);


endmodule