module fake_jpeg_11408_n_476 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_476);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_476;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_9),
.B(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_SL g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_1),
.B(n_6),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_7),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_55),
.B(n_103),
.Y(n_130)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_56),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_57),
.Y(n_132)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_24),
.B(n_6),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_59),
.B(n_89),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_60),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_61),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_62),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_63),
.Y(n_172)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_65),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_66),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_68),
.B(n_82),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_69),
.Y(n_173)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_71),
.Y(n_144)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_73),
.Y(n_174)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_74),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_75),
.Y(n_161)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_76),
.Y(n_163)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_50),
.Y(n_77)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_78),
.Y(n_183)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_79),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_80),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_81),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_27),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g166 ( 
.A(n_83),
.Y(n_166)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_84),
.Y(n_194)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

BUFx10_ASAP7_75t_L g168 ( 
.A(n_86),
.Y(n_168)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_88),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_18),
.B(n_9),
.Y(n_89)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_91),
.Y(n_157)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_92),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g191 ( 
.A(n_93),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_94),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_19),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_95),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_48),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_102),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_97),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_98),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_41),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_46),
.B1(n_28),
.B2(n_25),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_31),
.B(n_16),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_37),
.B(n_36),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_115),
.Y(n_137)
);

BUFx16f_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_110),
.Y(n_134)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_106),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_21),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_1),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_29),
.B(n_36),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_108),
.B(n_13),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_30),
.Y(n_109)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_109),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_43),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_30),
.Y(n_111)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_111),
.Y(n_188)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_19),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_114),
.Y(n_135)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_32),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_113),
.A2(n_67),
.B1(n_90),
.B2(n_95),
.Y(n_120)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_43),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_39),
.Y(n_115)
);

INVx6_ASAP7_75t_SL g116 ( 
.A(n_32),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_9),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_39),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_3),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_115),
.A2(n_53),
.B1(n_34),
.B2(n_46),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_119),
.A2(n_192),
.B1(n_171),
.B2(n_167),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_120),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_121),
.A2(n_141),
.B1(n_158),
.B2(n_184),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_53),
.C(n_34),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_136),
.B(n_143),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_138),
.B(n_151),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_59),
.A2(n_28),
.B1(n_25),
.B2(n_21),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_142),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_89),
.B(n_10),
.C(n_14),
.Y(n_143)
);

OR2x4_ASAP7_75t_SL g147 ( 
.A(n_101),
.B(n_1),
.Y(n_147)
);

AO22x1_ASAP7_75t_L g240 ( 
.A1(n_147),
.A2(n_185),
.B1(n_165),
.B2(n_175),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_150),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_16),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_137),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_88),
.B(n_14),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_154),
.B(n_155),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_93),
.B(n_10),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_57),
.A2(n_13),
.B1(n_4),
.B2(n_5),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_94),
.B(n_5),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_159),
.B(n_160),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_98),
.B(n_99),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_113),
.A2(n_111),
.B1(n_109),
.B2(n_62),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_167),
.A2(n_171),
.B1(n_187),
.B2(n_189),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_65),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_73),
.B(n_75),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_179),
.B(n_191),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_66),
.A2(n_69),
.B1(n_117),
.B2(n_81),
.Y(n_184)
);

OA22x2_ASAP7_75t_L g185 ( 
.A1(n_77),
.A2(n_68),
.B1(n_91),
.B2(n_58),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_102),
.A2(n_35),
.B1(n_116),
.B2(n_41),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_116),
.A2(n_35),
.B1(n_41),
.B2(n_80),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_59),
.B(n_55),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_193),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_59),
.A2(n_55),
.B1(n_103),
.B2(n_68),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_59),
.B(n_55),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_187),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_195),
.B(n_200),
.Y(n_268)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_132),
.Y(n_197)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_197),
.Y(n_270)
);

BUFx12_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_198),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_147),
.A2(n_169),
.B1(n_126),
.B2(n_189),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_SL g275 ( 
.A1(n_202),
.A2(n_240),
.B(n_252),
.C(n_172),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_130),
.B(n_127),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_203),
.B(n_208),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_163),
.Y(n_204)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_204),
.Y(n_266)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_125),
.Y(n_205)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_205),
.Y(n_267)
);

NAND3xp33_ASAP7_75t_L g206 ( 
.A(n_134),
.B(n_122),
.C(n_135),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_206),
.B(n_210),
.Y(n_264)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_207),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_168),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_144),
.Y(n_209)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_209),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_168),
.Y(n_210)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_161),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_212),
.Y(n_284)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_149),
.Y(n_213)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_213),
.Y(n_289)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_178),
.Y(n_215)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_215),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_132),
.Y(n_216)
);

INVx8_ASAP7_75t_L g262 ( 
.A(n_216),
.Y(n_262)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_217),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_128),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_218),
.B(n_220),
.Y(n_271)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_152),
.Y(n_219)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_219),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_156),
.B(n_118),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_221),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_150),
.B(n_157),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_223),
.B(n_227),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_140),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_224),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_225),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_131),
.Y(n_226)
);

NAND2xp33_ASAP7_75t_SL g303 ( 
.A(n_226),
.B(n_230),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_185),
.B(n_123),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_184),
.A2(n_173),
.B1(n_186),
.B2(n_148),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_228),
.A2(n_254),
.B1(n_258),
.B2(n_252),
.Y(n_278)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_177),
.Y(n_231)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_231),
.Y(n_291)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_164),
.Y(n_232)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_232),
.Y(n_269)
);

A2O1A1Ixp33_ASAP7_75t_L g233 ( 
.A1(n_147),
.A2(n_188),
.B(n_120),
.C(n_139),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_256),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_183),
.Y(n_234)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_234),
.Y(n_279)
);

BUFx12f_ASAP7_75t_L g235 ( 
.A(n_129),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_235),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_145),
.B(n_165),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_236),
.Y(n_286)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_133),
.Y(n_237)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_237),
.Y(n_294)
);

INVx11_ASAP7_75t_L g238 ( 
.A(n_139),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_238),
.Y(n_293)
);

INVx3_ASAP7_75t_SL g239 ( 
.A(n_174),
.Y(n_239)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_239),
.Y(n_295)
);

OR2x2_ASAP7_75t_SL g241 ( 
.A(n_124),
.B(n_162),
.Y(n_241)
);

AND2x2_ASAP7_75t_SL g263 ( 
.A(n_241),
.B(n_257),
.Y(n_263)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_145),
.Y(n_243)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_243),
.Y(n_297)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_176),
.Y(n_244)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_244),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_140),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_245),
.B(n_247),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_174),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_246),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_146),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_148),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_248),
.B(n_253),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_169),
.B(n_129),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_249),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_182),
.A2(n_173),
.B1(n_170),
.B2(n_172),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_186),
.B(n_182),
.Y(n_253)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_191),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_255),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_191),
.Y(n_256)
);

BUFx12f_ASAP7_75t_L g257 ( 
.A(n_166),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_180),
.B(n_170),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_242),
.A2(n_196),
.B1(n_228),
.B2(n_202),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_260),
.A2(n_277),
.B1(n_278),
.B2(n_285),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_226),
.A2(n_211),
.B1(n_240),
.B2(n_200),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_273),
.A2(n_288),
.B1(n_296),
.B2(n_293),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_275),
.A2(n_198),
.B1(n_235),
.B2(n_277),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_196),
.A2(n_180),
.B1(n_211),
.B2(n_214),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_214),
.A2(n_251),
.B(n_206),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_281),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_222),
.A2(n_199),
.B1(n_250),
.B2(n_233),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_229),
.A2(n_241),
.B1(n_239),
.B2(n_237),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_201),
.A2(n_197),
.B1(n_248),
.B2(n_245),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_292),
.A2(n_263),
.B1(n_295),
.B2(n_279),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_204),
.A2(n_234),
.B1(n_224),
.B2(n_216),
.Y(n_296)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_297),
.Y(n_308)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_308),
.Y(n_350)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_294),
.Y(n_309)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_309),
.Y(n_344)
);

O2A1O1Ixp33_ASAP7_75t_L g310 ( 
.A1(n_259),
.A2(n_238),
.B(n_257),
.C(n_256),
.Y(n_310)
);

OA22x2_ASAP7_75t_L g355 ( 
.A1(n_310),
.A2(n_318),
.B1(n_333),
.B2(n_291),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_271),
.B(n_235),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_311),
.Y(n_345)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_297),
.Y(n_312)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_312),
.Y(n_362)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_280),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_301),
.Y(n_315)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_315),
.Y(n_366)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_301),
.Y(n_316)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_316),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_263),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_317),
.A2(n_320),
.B(n_293),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_260),
.A2(n_231),
.B1(n_207),
.B2(n_212),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_R g319 ( 
.A1(n_282),
.A2(n_257),
.B(n_217),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_319),
.B(n_276),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_273),
.B(n_255),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_284),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_321),
.B(n_324),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_322),
.A2(n_326),
.B(n_276),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_281),
.B(n_198),
.Y(n_323)
);

BUFx24_ASAP7_75t_SL g363 ( 
.A(n_323),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_259),
.B(n_286),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_303),
.A2(n_268),
.B1(n_288),
.B2(n_275),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_325),
.A2(n_334),
.B1(n_343),
.B2(n_317),
.Y(n_359)
);

AOI32xp33_ASAP7_75t_L g326 ( 
.A1(n_286),
.A2(n_304),
.A3(n_275),
.B1(n_263),
.B2(n_305),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_261),
.B(n_289),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_327),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_290),
.B(n_264),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_328),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_299),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_329),
.B(n_332),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_300),
.B(n_306),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_330),
.Y(n_371)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_295),
.Y(n_331)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_331),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_298),
.B(n_279),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_275),
.A2(n_296),
.B1(n_266),
.B2(n_302),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_266),
.Y(n_335)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_335),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_275),
.B(n_269),
.C(n_294),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_336),
.B(n_325),
.C(n_343),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_269),
.Y(n_337)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_337),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_274),
.B(n_287),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_338),
.B(n_340),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_287),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_339),
.B(n_272),
.Y(n_370)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_283),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_283),
.B(n_267),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_341),
.B(n_342),
.Y(n_367)
);

NOR2x1p5_ASAP7_75t_L g342 ( 
.A(n_302),
.B(n_280),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_347),
.B(n_348),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_313),
.A2(n_270),
.B1(n_262),
.B2(n_291),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_351),
.A2(n_356),
.B1(n_368),
.B2(n_334),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_321),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_354),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_355),
.B(n_310),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_313),
.A2(n_270),
.B1(n_262),
.B2(n_265),
.Y(n_356)
);

OAI22x1_ASAP7_75t_L g391 ( 
.A1(n_359),
.A2(n_319),
.B1(n_333),
.B2(n_342),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_364),
.A2(n_323),
.B(n_320),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_365),
.A2(n_307),
.B(n_320),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_324),
.A2(n_265),
.B1(n_272),
.B2(n_267),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_370),
.B(n_337),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_371),
.B(n_329),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_372),
.B(n_373),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_361),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_349),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_375),
.Y(n_396)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_349),
.Y(n_376)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_376),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_365),
.A2(n_336),
.B(n_322),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_377),
.B(n_378),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_359),
.A2(n_307),
.B(n_326),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_361),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_379),
.Y(n_401)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_352),
.Y(n_380)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_380),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_381),
.A2(n_382),
.B1(n_385),
.B2(n_387),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_345),
.B(n_314),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_383),
.Y(n_408)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_352),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_386),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_353),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_350),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_362),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_389),
.B(n_393),
.Y(n_411)
);

OA21x2_ASAP7_75t_L g403 ( 
.A1(n_390),
.A2(n_391),
.B(n_367),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_364),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_392),
.A2(n_395),
.B1(n_368),
.B2(n_347),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_353),
.A2(n_308),
.B(n_312),
.Y(n_393)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_366),
.Y(n_395)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_397),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_394),
.B(n_348),
.C(n_357),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_400),
.C(n_402),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_394),
.B(n_357),
.C(n_363),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_378),
.B(n_358),
.C(n_360),
.Y(n_402)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_403),
.Y(n_421)
);

OA22x2_ASAP7_75t_L g404 ( 
.A1(n_381),
.A2(n_355),
.B1(n_367),
.B2(n_354),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_404),
.B(n_342),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_390),
.A2(n_356),
.B1(n_351),
.B2(n_355),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_406),
.A2(n_412),
.B1(n_413),
.B2(n_382),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_390),
.A2(n_355),
.B1(n_360),
.B2(n_358),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_392),
.A2(n_393),
.B1(n_391),
.B2(n_389),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_398),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_416),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_417),
.B(n_427),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_399),
.B(n_377),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_419),
.B(n_422),
.C(n_423),
.Y(n_434)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_398),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_420),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_402),
.B(n_400),
.C(n_405),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_405),
.B(n_375),
.C(n_344),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_397),
.B(n_411),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_424),
.B(n_426),
.C(n_415),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_396),
.A2(n_388),
.B(n_374),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_425),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_411),
.B(n_370),
.Y(n_426)
);

CKINVDCx14_ASAP7_75t_R g427 ( 
.A(n_414),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_428),
.A2(n_412),
.B1(n_413),
.B2(n_406),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_401),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_429),
.B(n_395),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_426),
.B(n_410),
.Y(n_431)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_431),
.Y(n_451)
);

CKINVDCx14_ASAP7_75t_R g432 ( 
.A(n_428),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_432),
.B(n_439),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_418),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_437),
.A2(n_441),
.B1(n_417),
.B2(n_421),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_425),
.B(n_408),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_440),
.B(n_424),
.Y(n_442)
);

INVx13_ASAP7_75t_L g441 ( 
.A(n_421),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_442),
.B(n_449),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_443),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_435),
.B(n_415),
.C(n_419),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_444),
.B(n_445),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_434),
.B(n_435),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_437),
.A2(n_433),
.B1(n_430),
.B2(n_418),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_447),
.A2(n_436),
.B1(n_440),
.B2(n_430),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_434),
.B(n_422),
.C(n_423),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_448),
.B(n_450),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_434),
.B(n_403),
.C(n_404),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_449),
.B(n_433),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_452),
.B(n_457),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_448),
.A2(n_431),
.B(n_439),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_458),
.B(n_459),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_450),
.A2(n_438),
.B(n_388),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_453),
.B(n_451),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_460),
.B(n_463),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_454),
.B(n_444),
.Y(n_461)
);

AOI21x1_ASAP7_75t_L g469 ( 
.A1(n_461),
.A2(n_456),
.B(n_369),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_455),
.B(n_346),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_456),
.B(n_446),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_464),
.B(n_462),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_467),
.B(n_468),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_462),
.B(n_438),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_469),
.B(n_465),
.C(n_403),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_470),
.B(n_404),
.C(n_438),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_472),
.A2(n_471),
.B1(n_438),
.B2(n_466),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_473),
.A2(n_432),
.B(n_441),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_474),
.A2(n_409),
.B(n_407),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_475),
.B(n_346),
.Y(n_476)
);


endmodule