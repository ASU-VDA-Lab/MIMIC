module fake_jpeg_7746_n_179 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_6),
.B(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx2_ASAP7_75t_SL g31 ( 
.A(n_29),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_0),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_33),
.A2(n_17),
.B1(n_20),
.B2(n_23),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_41),
.A2(n_27),
.B1(n_26),
.B2(n_25),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_16),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_42),
.B(n_14),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_21),
.C(n_15),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_18),
.C(n_3),
.Y(n_75)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_20),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_15),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_24),
.Y(n_68)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_63),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_19),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_57),
.B(n_68),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_19),
.B1(n_16),
.B2(n_28),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_47),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_70),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_20),
.B1(n_23),
.B2(n_19),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_60),
.A2(n_62),
.B1(n_65),
.B2(n_69),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_49),
.A2(n_35),
.B1(n_30),
.B2(n_23),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_61),
.A2(n_64),
.B1(n_44),
.B2(n_40),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_16),
.B1(n_25),
.B2(n_28),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_53),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_35),
.B1(n_30),
.B2(n_46),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_14),
.B1(n_27),
.B2(n_26),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_75),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_67),
.A2(n_48),
.B1(n_4),
.B2(n_5),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_50),
.A2(n_24),
.B1(n_18),
.B2(n_22),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_22),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_72),
.Y(n_93)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_80),
.Y(n_98)
);

AND2x6_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_0),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_SL g87 ( 
.A(n_74),
.B(n_76),
.C(n_57),
.Y(n_87)
);

NOR2x1_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_39),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_39),
.C(n_38),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_51),
.C(n_52),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_38),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_52),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_53),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_32),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_2),
.Y(n_82)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_87),
.B(n_94),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_77),
.C(n_100),
.Y(n_114)
);

OAI22x1_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_105),
.B1(n_96),
.B2(n_85),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_92),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_99),
.B(n_80),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_40),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_102),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_101),
.A2(n_73),
.B1(n_63),
.B2(n_72),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_44),
.Y(n_102)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_58),
.B(n_3),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_65),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_84),
.B(n_68),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_110),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_84),
.B(n_66),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_85),
.A2(n_76),
.B1(n_55),
.B2(n_61),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_119),
.B1(n_122),
.B2(n_90),
.Y(n_137)
);

OAI32xp33_ASAP7_75t_L g113 ( 
.A1(n_102),
.A2(n_74),
.A3(n_62),
.B1(n_70),
.B2(n_79),
.Y(n_113)
);

A2O1A1O1Ixp25_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_91),
.B(n_93),
.C(n_98),
.D(n_99),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_115),
.C(n_123),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_75),
.C(n_81),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_86),
.B(n_97),
.Y(n_116)
);

BUFx24_ASAP7_75t_SL g133 ( 
.A(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_97),
.B(n_89),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_83),
.B(n_82),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_101),
.B(n_5),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_88),
.Y(n_129)
);

NOR3xp33_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_96),
.C(n_91),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_127),
.Y(n_148)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

AO221x1_ASAP7_75t_L g140 ( 
.A1(n_128),
.A2(n_130),
.B1(n_135),
.B2(n_139),
.C(n_123),
.Y(n_140)
);

XOR2x1_ASAP7_75t_SL g142 ( 
.A(n_129),
.B(n_131),
.Y(n_142)
);

INVxp33_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

NAND3xp33_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_91),
.C(n_104),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_132),
.A2(n_134),
.B(n_90),
.Y(n_146)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_137),
.A2(n_109),
.B1(n_115),
.B2(n_94),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_143),
.B1(n_144),
.B2(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_139),
.A2(n_124),
.B1(n_109),
.B2(n_111),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_136),
.A2(n_106),
.B(n_114),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_145),
.A2(n_149),
.B(n_133),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_129),
.C(n_136),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_147),
.Y(n_155)
);

XOR2x2_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_121),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_126),
.A2(n_108),
.B1(n_120),
.B2(n_72),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_153),
.C(n_154),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_95),
.C(n_92),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_95),
.B(n_92),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_158),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_32),
.C(n_7),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_144),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_159),
.B(n_7),
.Y(n_165)
);

AOI31xp67_ASAP7_75t_L g160 ( 
.A1(n_157),
.A2(n_149),
.A3(n_142),
.B(n_146),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_160),
.B(n_164),
.Y(n_169)
);

AO21x1_ASAP7_75t_L g162 ( 
.A1(n_151),
.A2(n_148),
.B(n_143),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_163),
.Y(n_170)
);

BUFx4f_ASAP7_75t_SL g163 ( 
.A(n_156),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_150),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_165),
.B(n_8),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_161),
.B(n_153),
.Y(n_167)
);

AOI322xp5_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_168),
.A3(n_166),
.B1(n_154),
.B2(n_11),
.C1(n_12),
.C2(n_10),
.Y(n_174)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_152),
.B(n_158),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_165),
.Y(n_172)
);

AO21x1_ASAP7_75t_L g176 ( 
.A1(n_172),
.A2(n_173),
.B(n_174),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_169),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_SL g175 ( 
.A1(n_174),
.A2(n_168),
.B(n_10),
.C(n_11),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_12),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_8),
.C(n_12),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_178),
.Y(n_179)
);


endmodule