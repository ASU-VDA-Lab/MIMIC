module fake_jpeg_17874_n_59 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_8),
.Y(n_9)
);

BUFx12_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_3),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_16),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_21)
);

NOR3xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_25),
.C(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_23),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_16),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_5),
.B1(n_12),
.B2(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NAND3xp33_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_10),
.C(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_31),
.A2(n_10),
.B1(n_17),
.B2(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_11),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_17),
.Y(n_40)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_37),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_41),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_32),
.B1(n_36),
.B2(n_28),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_29),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_47),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_48),
.B(n_39),
.Y(n_52)
);

INVxp33_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_50),
.A2(n_48),
.B(n_38),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_28),
.B(n_27),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_40),
.B1(n_45),
.B2(n_41),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_56),
.C(n_27),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_57),
.A2(n_44),
.B1(n_34),
.B2(n_51),
.Y(n_58)
);

AOI31xp33_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_42),
.A3(n_44),
.B(n_10),
.Y(n_59)
);


endmodule