module fake_jpeg_30512_n_247 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_247);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_3),
.B(n_17),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_23),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_56),
.Y(n_73)
);

CKINVDCx9p33_ASAP7_75t_R g52 ( 
.A(n_23),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_53),
.Y(n_72)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_61),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_23),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_8),
.Y(n_59)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_65),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_28),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_26),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_36),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_52),
.A2(n_37),
.B1(n_26),
.B2(n_40),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_67),
.A2(n_87),
.B1(n_88),
.B2(n_66),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_44),
.A2(n_29),
.B1(n_43),
.B2(n_35),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_21),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_34),
.B1(n_41),
.B2(n_40),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_71),
.A2(n_77),
.B1(n_48),
.B2(n_47),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_46),
.A2(n_32),
.B1(n_41),
.B2(n_30),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_43),
.C(n_35),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_83),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_57),
.B(n_30),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_79),
.B(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_61),
.B(n_25),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_34),
.B1(n_32),
.B2(n_31),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_60),
.A2(n_31),
.B1(n_25),
.B2(n_38),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_95),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_68),
.A2(n_60),
.B(n_50),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_76),
.C(n_90),
.Y(n_124)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

AO22x1_ASAP7_75t_L g98 ( 
.A1(n_68),
.A2(n_53),
.B1(n_56),
.B2(n_49),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_112),
.B1(n_114),
.B2(n_116),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_89),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_99),
.B(n_106),
.Y(n_123)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

NOR2xp67_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_38),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_103),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_42),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_42),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_108),
.Y(n_133)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_83),
.A2(n_53),
.B(n_49),
.C(n_55),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_21),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_68),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_119),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_72),
.B(n_15),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_110),
.B(n_122),
.Y(n_128)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_53),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_118),
.Y(n_140)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_81),
.A2(n_63),
.B1(n_56),
.B2(n_42),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_117),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_66),
.A2(n_21),
.B(n_42),
.C(n_2),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_21),
.Y(n_119)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_120),
.Y(n_135)
);

CKINVDCx6p67_ASAP7_75t_R g121 ( 
.A(n_69),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_121),
.Y(n_143)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_107),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_94),
.B(n_92),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_142),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_94),
.B(n_76),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_101),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_144),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_114),
.B1(n_94),
.B2(n_98),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_145),
.A2(n_154),
.B1(n_135),
.B2(n_137),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_96),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_147),
.C(n_141),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_126),
.A2(n_106),
.B1(n_113),
.B2(n_95),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_127),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_122),
.B1(n_75),
.B2(n_82),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_140),
.A2(n_75),
.B1(n_82),
.B2(n_90),
.Y(n_150)
);

AOI21xp33_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_121),
.B(n_118),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_155),
.Y(n_162)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_136),
.Y(n_153)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_116),
.B1(n_115),
.B2(n_120),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_133),
.B(n_13),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_159),
.Y(n_160)
);

NAND2x1p5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_121),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_157),
.A2(n_124),
.B(n_138),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_130),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_158),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_129),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_161),
.B(n_166),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_137),
.C(n_139),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_168),
.A2(n_150),
.B1(n_157),
.B2(n_156),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_128),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_170),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_139),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_135),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_172),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_143),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_143),
.Y(n_173)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_173),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_174),
.A2(n_145),
.B1(n_154),
.B2(n_157),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_129),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_175),
.B(n_131),
.Y(n_181)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_167),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_177),
.A2(n_168),
.B1(n_174),
.B2(n_165),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_166),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_131),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_179),
.B(n_183),
.Y(n_193)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_181),
.Y(n_198)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_159),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_127),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_186),
.B(n_188),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_160),
.Y(n_188)
);

AOI21x1_ASAP7_75t_SL g190 ( 
.A1(n_179),
.A2(n_164),
.B(n_171),
.Y(n_190)
);

INVx13_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

FAx1_ASAP7_75t_SL g191 ( 
.A(n_185),
.B(n_161),
.CI(n_170),
.CON(n_191),
.SN(n_191)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_7),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_192),
.A2(n_189),
.B1(n_132),
.B2(n_117),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_187),
.B(n_162),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_196),
.B(n_189),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_197),
.A2(n_100),
.B1(n_93),
.B2(n_2),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_185),
.B(n_160),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_202),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_165),
.C(n_132),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_180),
.C(n_178),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_121),
.Y(n_202)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_203),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_198),
.B(n_184),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_212),
.Y(n_217)
);

AO221x1_ASAP7_75t_L g205 ( 
.A1(n_200),
.A2(n_187),
.B1(n_176),
.B2(n_188),
.C(n_130),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_211),
.Y(n_215)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_199),
.C(n_201),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_210),
.A2(n_197),
.B1(n_194),
.B2(n_191),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_190),
.A2(n_66),
.B(n_1),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_195),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_213),
.B(n_195),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_9),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_212),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_208),
.C(n_211),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_207),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_221),
.B(n_220),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_6),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_223),
.B(n_224),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_209),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_225),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_227),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_228),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_222),
.A2(n_208),
.B1(n_11),
.B2(n_4),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_230),
.B(n_231),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_5),
.C(n_16),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_229),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_229),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_237),
.A2(n_239),
.B(n_240),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_219),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_238),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_232),
.A2(n_215),
.B1(n_228),
.B2(n_217),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_233),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_242),
.A2(n_236),
.B1(n_238),
.B2(n_18),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_243),
.A2(n_244),
.B(n_0),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_19),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_245),
.B(n_0),
.C(n_1),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_1),
.Y(n_247)
);


endmodule