module fake_ariane_2986_n_121 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_17, n_4, n_2, n_18, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_121);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_121;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_119;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_120;
wire n_106;
wire n_53;
wire n_111;
wire n_115;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_49;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_107;
wire n_72;
wire n_105;
wire n_44;
wire n_30;
wire n_82;
wire n_42;
wire n_31;
wire n_57;
wire n_70;
wire n_117;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_112;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_118;
wire n_93;
wire n_61;
wire n_108;
wire n_102;
wire n_43;
wire n_87;
wire n_81;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_116;
wire n_104;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_35;
wire n_54;

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVxp67_ASAP7_75t_SL g31 ( 
.A(n_4),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_24),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVxp33_ASAP7_75t_SL g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_28),
.B(n_0),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVxp33_ASAP7_75t_SL g57 ( 
.A(n_27),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_35),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NAND2x1p5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_39),
.Y(n_64)
);

NAND2x1p5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_42),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_60),
.A2(n_41),
.B1(n_33),
.B2(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

AO22x2_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_44),
.B1(n_43),
.B2(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

AO22x2_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_34),
.B1(n_38),
.B2(n_36),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_57),
.B(n_59),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_64),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_59),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_66),
.A2(n_57),
.B1(n_58),
.B2(n_35),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_52),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_49),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_49),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_63),
.B(n_62),
.C(n_69),
.Y(n_83)
);

CKINVDCx5p33_ASAP7_75t_R g84 ( 
.A(n_79),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_72),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_68),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

AND2x4_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_74),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_81),
.B1(n_82),
.B2(n_80),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

AOI221x1_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_85),
.B1(n_68),
.B2(n_72),
.C(n_86),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_89),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_84),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_93),
.A2(n_91),
.B(n_88),
.Y(n_97)
);

OA21x2_ASAP7_75t_L g98 ( 
.A1(n_93),
.A2(n_91),
.B(n_92),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

BUFx4f_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_50),
.Y(n_103)
);

OR2x6_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_72),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

AND2x4_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_99),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_4),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_104),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_103),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_106),
.B(n_100),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);

CKINVDCx5p33_ASAP7_75t_R g112 ( 
.A(n_110),
.Y(n_112)
);

NOR2x1p5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_108),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_SL g114 ( 
.A1(n_111),
.A2(n_7),
.B(n_8),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_9),
.Y(n_115)
);

AOI21xp33_ASAP7_75t_L g116 ( 
.A1(n_114),
.A2(n_54),
.B(n_53),
.Y(n_116)
);

NAND4xp25_ASAP7_75t_SL g117 ( 
.A(n_115),
.B(n_14),
.C(n_16),
.D(n_20),
.Y(n_117)
);

NAND4xp25_ASAP7_75t_SL g118 ( 
.A(n_116),
.B(n_21),
.C(n_23),
.D(n_25),
.Y(n_118)
);

NOR3xp33_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_75),
.C(n_78),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_118),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_120),
.Y(n_121)
);


endmodule