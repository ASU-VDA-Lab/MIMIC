module fake_netlist_1_2317_n_693 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_693);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_693;
wire n_117;
wire n_663;
wire n_513;
wire n_361;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_462;
wire n_232;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_529;
wire n_455;
wire n_312;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_466;
wire n_302;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_581;
wire n_458;
wire n_504;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_7), .Y(n_78) );
HB1xp67_ASAP7_75t_L g79 ( .A(n_67), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_22), .Y(n_80) );
INVxp67_ASAP7_75t_L g81 ( .A(n_54), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_27), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_3), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_63), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_40), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_30), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_9), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_11), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_59), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_56), .Y(n_90) );
XNOR2xp5_ASAP7_75t_L g91 ( .A(n_14), .B(n_0), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_1), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_39), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_1), .Y(n_94) );
INVxp67_ASAP7_75t_L g95 ( .A(n_55), .Y(n_95) );
NOR2xp67_ASAP7_75t_L g96 ( .A(n_37), .B(n_4), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_23), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_77), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_32), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_64), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_44), .Y(n_101) );
INVx1_ASAP7_75t_SL g102 ( .A(n_25), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_36), .Y(n_103) );
CKINVDCx16_ASAP7_75t_R g104 ( .A(n_66), .Y(n_104) );
INVxp67_ASAP7_75t_SL g105 ( .A(n_68), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_15), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_18), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_28), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_35), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_52), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_10), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_49), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_4), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_12), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_16), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_71), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_17), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_7), .Y(n_118) );
INVxp33_ASAP7_75t_SL g119 ( .A(n_24), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_29), .Y(n_120) );
INVx1_ASAP7_75t_SL g121 ( .A(n_9), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_10), .Y(n_122) );
NOR2xp67_ASAP7_75t_L g123 ( .A(n_8), .B(n_43), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_75), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_60), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_118), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_104), .Y(n_127) );
AND2x4_ASAP7_75t_L g128 ( .A(n_88), .B(n_0), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_79), .B(n_2), .Y(n_129) );
NOR2xp33_ASAP7_75t_SL g130 ( .A(n_90), .B(n_45), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_85), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_118), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_110), .B(n_2), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_87), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_85), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_80), .B(n_3), .Y(n_136) );
BUFx3_ASAP7_75t_L g137 ( .A(n_86), .Y(n_137) );
HB1xp67_ASAP7_75t_L g138 ( .A(n_87), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_88), .B(n_5), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_116), .Y(n_140) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_92), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_86), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_89), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_89), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_82), .Y(n_145) );
AOI22xp5_ASAP7_75t_L g146 ( .A1(n_119), .A2(n_5), .B1(n_6), .B2(n_8), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_116), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_120), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_84), .B(n_6), .Y(n_149) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_92), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_98), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_94), .B(n_11), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_100), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_120), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_103), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_106), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_125), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_107), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_94), .B(n_12), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_108), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_109), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_78), .B(n_13), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_122), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_112), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_83), .B(n_13), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_122), .Y(n_166) );
OAI22xp5_ASAP7_75t_L g167 ( .A1(n_111), .A2(n_19), .B1(n_20), .B2(n_21), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_115), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_128), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_157), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_128), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_128), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_157), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_138), .B(n_101), .Y(n_174) );
BUFx2_ASAP7_75t_L g175 ( .A(n_134), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_157), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_163), .Y(n_177) );
AND2x2_ASAP7_75t_L g178 ( .A(n_141), .B(n_101), .Y(n_178) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_157), .Y(n_179) );
AND2x6_ASAP7_75t_L g180 ( .A(n_162), .B(n_124), .Y(n_180) );
BUFx10_ASAP7_75t_L g181 ( .A(n_127), .Y(n_181) );
OR2x2_ASAP7_75t_L g182 ( .A(n_150), .B(n_121), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_157), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_134), .A2(n_119), .B1(n_113), .B2(n_114), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_162), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_140), .Y(n_186) );
NAND2x1p5_ASAP7_75t_L g187 ( .A(n_162), .B(n_117), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_165), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_165), .Y(n_189) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_166), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_140), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_165), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_139), .Y(n_193) );
INVx4_ASAP7_75t_L g194 ( .A(n_137), .Y(n_194) );
INVx3_ASAP7_75t_L g195 ( .A(n_147), .Y(n_195) );
BUFx3_ASAP7_75t_L g196 ( .A(n_147), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_145), .B(n_97), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_148), .Y(n_198) );
INVx2_ASAP7_75t_SL g199 ( .A(n_137), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_148), .Y(n_200) );
BUFx2_ASAP7_75t_L g201 ( .A(n_166), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_145), .B(n_97), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_154), .Y(n_203) );
BUFx8_ASAP7_75t_SL g204 ( .A(n_127), .Y(n_204) );
AO22x2_ASAP7_75t_L g205 ( .A1(n_167), .A2(n_105), .B1(n_102), .B2(n_95), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_154), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_151), .B(n_81), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_126), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_151), .B(n_99), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_126), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_126), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_131), .B(n_99), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_131), .B(n_93), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_139), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_132), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_132), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_135), .B(n_96), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_132), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_135), .Y(n_219) );
CKINVDCx5p33_ASAP7_75t_R g220 ( .A(n_152), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_142), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_142), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_143), .Y(n_223) );
CKINVDCx11_ASAP7_75t_R g224 ( .A(n_158), .Y(n_224) );
BUFx3_ASAP7_75t_L g225 ( .A(n_158), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_129), .A2(n_93), .B1(n_90), .B2(n_91), .Y(n_226) );
NAND2x1p5_ASAP7_75t_L g227 ( .A(n_143), .B(n_123), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_212), .B(n_144), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_220), .A2(n_159), .B1(n_133), .B2(n_146), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_213), .B(n_168), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_225), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_176), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_212), .B(n_168), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_225), .Y(n_234) );
OAI22xp5_ASAP7_75t_SL g235 ( .A1(n_177), .A2(n_91), .B1(n_136), .B2(n_149), .Y(n_235) );
BUFx3_ASAP7_75t_L g236 ( .A(n_180), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_171), .A2(n_144), .B(n_155), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_197), .B(n_164), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_202), .B(n_164), .Y(n_239) );
INVx2_ASAP7_75t_SL g240 ( .A(n_174), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_193), .B(n_156), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_216), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_216), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_209), .B(n_156), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_194), .B(n_155), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_176), .Y(n_246) );
INVx3_ASAP7_75t_L g247 ( .A(n_196), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_169), .B(n_153), .Y(n_248) );
NOR3xp33_ASAP7_75t_L g249 ( .A(n_224), .B(n_153), .C(n_160), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_194), .B(n_161), .Y(n_250) );
NOR2x1_ASAP7_75t_L g251 ( .A(n_182), .B(n_161), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_214), .B(n_160), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_180), .A2(n_130), .B1(n_31), .B2(n_33), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_176), .Y(n_254) );
INVx3_ASAP7_75t_L g255 ( .A(n_196), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_194), .B(n_26), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_199), .B(n_34), .Y(n_257) );
NOR2xp33_ASAP7_75t_SL g258 ( .A(n_175), .B(n_38), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_220), .A2(n_184), .B1(n_180), .B2(n_178), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_176), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_216), .Y(n_261) );
BUFx12f_ASAP7_75t_L g262 ( .A(n_224), .Y(n_262) );
OAI22xp5_ASAP7_75t_L g263 ( .A1(n_187), .A2(n_41), .B1(n_42), .B2(n_46), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_216), .Y(n_264) );
BUFx3_ASAP7_75t_L g265 ( .A(n_180), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_180), .A2(n_47), .B1(n_48), .B2(n_50), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_199), .B(n_207), .Y(n_267) );
AND2x4_ASAP7_75t_L g268 ( .A(n_174), .B(n_51), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_216), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_176), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_219), .B(n_53), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_208), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_185), .B(n_57), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_179), .Y(n_274) );
AO21x1_ASAP7_75t_L g275 ( .A1(n_187), .A2(n_58), .B(n_61), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_221), .B(n_62), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_208), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_222), .B(n_65), .Y(n_278) );
BUFx3_ASAP7_75t_L g279 ( .A(n_180), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_188), .B(n_69), .Y(n_280) );
NAND2xp33_ASAP7_75t_L g281 ( .A(n_187), .B(n_70), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_169), .B(n_72), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_210), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_175), .B(n_73), .Y(n_284) );
BUFx2_ASAP7_75t_L g285 ( .A(n_201), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_191), .Y(n_286) );
BUFx3_ASAP7_75t_L g287 ( .A(n_169), .Y(n_287) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_191), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_179), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_223), .B(n_74), .Y(n_290) );
INVxp67_ASAP7_75t_SL g291 ( .A(n_182), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_286), .Y(n_292) );
INVx3_ASAP7_75t_L g293 ( .A(n_287), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_259), .B(n_178), .Y(n_294) );
INVx1_ASAP7_75t_SL g295 ( .A(n_285), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_245), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_248), .Y(n_297) );
INVx4_ASAP7_75t_L g298 ( .A(n_236), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_248), .Y(n_299) );
INVx3_ASAP7_75t_L g300 ( .A(n_287), .Y(n_300) );
BUFx4f_ASAP7_75t_L g301 ( .A(n_262), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_286), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_291), .Y(n_303) );
BUFx3_ASAP7_75t_L g304 ( .A(n_236), .Y(n_304) );
OA22x2_ASAP7_75t_L g305 ( .A1(n_235), .A2(n_226), .B1(n_201), .B2(n_190), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g306 ( .A1(n_240), .A2(n_205), .B1(n_192), .B2(n_189), .Y(n_306) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_265), .Y(n_307) );
BUFx2_ASAP7_75t_L g308 ( .A(n_268), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_250), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_286), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_286), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_288), .Y(n_312) );
NOR2xp33_ASAP7_75t_SL g313 ( .A(n_265), .B(n_204), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_233), .B(n_172), .Y(n_314) );
INVx3_ASAP7_75t_SL g315 ( .A(n_268), .Y(n_315) );
OAI22xp5_ASAP7_75t_L g316 ( .A1(n_279), .A2(n_205), .B1(n_227), .B2(n_217), .Y(n_316) );
OR2x6_ASAP7_75t_L g317 ( .A(n_279), .B(n_205), .Y(n_317) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_288), .Y(n_318) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_247), .Y(n_319) );
INVx2_ASAP7_75t_SL g320 ( .A(n_251), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g321 ( .A1(n_229), .A2(n_205), .B1(n_181), .B2(n_217), .Y(n_321) );
INVx3_ASAP7_75t_L g322 ( .A(n_247), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_288), .Y(n_323) );
NAND2x2_ASAP7_75t_L g324 ( .A(n_228), .B(n_204), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_249), .B(n_217), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_252), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_288), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_272), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_277), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_233), .A2(n_227), .B1(n_206), .B2(n_203), .Y(n_330) );
INVx2_ASAP7_75t_SL g331 ( .A(n_284), .Y(n_331) );
O2A1O1Ixp33_ASAP7_75t_L g332 ( .A1(n_238), .A2(n_227), .B(n_186), .C(n_206), .Y(n_332) );
BUFx8_ASAP7_75t_SL g333 ( .A(n_239), .Y(n_333) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_255), .Y(n_334) );
OR2x6_ASAP7_75t_L g335 ( .A(n_237), .B(n_181), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_241), .B(n_181), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_244), .A2(n_170), .B(n_183), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_241), .B(n_195), .Y(n_338) );
NAND2xp5_ASAP7_75t_SL g339 ( .A(n_275), .B(n_200), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_230), .B(n_195), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_252), .A2(n_195), .B1(n_198), .B2(n_218), .Y(n_341) );
INVx2_ASAP7_75t_SL g342 ( .A(n_255), .Y(n_342) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_295), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_333), .Y(n_344) );
OAI21x1_ASAP7_75t_L g345 ( .A1(n_339), .A2(n_282), .B(n_256), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_328), .Y(n_346) );
AO31x2_ASAP7_75t_L g347 ( .A1(n_316), .A2(n_280), .A3(n_273), .B(n_263), .Y(n_347) );
OAI21x1_ASAP7_75t_L g348 ( .A1(n_339), .A2(n_282), .B(n_257), .Y(n_348) );
INVx8_ASAP7_75t_L g349 ( .A(n_317), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_305), .A2(n_230), .B1(n_177), .B2(n_234), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_303), .B(n_267), .Y(n_351) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_303), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_328), .Y(n_353) );
AOI21xp33_ASAP7_75t_L g354 ( .A1(n_332), .A2(n_273), .B(n_280), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_315), .B(n_231), .Y(n_355) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_333), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_317), .Y(n_357) );
OAI21x1_ASAP7_75t_L g358 ( .A1(n_292), .A2(n_310), .B(n_323), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_326), .B(n_283), .Y(n_359) );
OA21x2_ASAP7_75t_L g360 ( .A1(n_306), .A2(n_290), .B(n_271), .Y(n_360) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_337), .A2(n_276), .B(n_278), .Y(n_361) );
INVx3_ASAP7_75t_L g362 ( .A(n_307), .Y(n_362) );
O2A1O1Ixp33_ASAP7_75t_L g363 ( .A1(n_336), .A2(n_198), .B(n_281), .C(n_210), .Y(n_363) );
INVx3_ASAP7_75t_L g364 ( .A(n_307), .Y(n_364) );
INVx3_ASAP7_75t_L g365 ( .A(n_307), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_296), .B(n_198), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_294), .B(n_218), .Y(n_367) );
INVx4_ASAP7_75t_L g368 ( .A(n_307), .Y(n_368) );
NAND2x1p5_ASAP7_75t_L g369 ( .A(n_304), .B(n_243), .Y(n_369) );
INVx6_ASAP7_75t_L g370 ( .A(n_298), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_317), .Y(n_371) );
INVx4_ASAP7_75t_L g372 ( .A(n_304), .Y(n_372) );
OAI22xp33_ASAP7_75t_L g373 ( .A1(n_315), .A2(n_258), .B1(n_215), .B2(n_211), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_309), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_346), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_346), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_374), .B(n_294), .Y(n_377) );
AO21x2_ASAP7_75t_L g378 ( .A1(n_354), .A2(n_321), .B(n_330), .Y(n_378) );
A2O1A1Ixp33_ASAP7_75t_L g379 ( .A1(n_374), .A2(n_308), .B(n_314), .C(n_331), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_351), .B(n_325), .Y(n_380) );
AOI22xp33_ASAP7_75t_SL g381 ( .A1(n_349), .A2(n_305), .B1(n_313), .B2(n_325), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_353), .Y(n_382) );
AOI222xp33_ASAP7_75t_L g383 ( .A1(n_350), .A2(n_325), .B1(n_301), .B2(n_320), .C1(n_338), .C2(n_340), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_353), .Y(n_384) );
AOI22xp33_ASAP7_75t_SL g385 ( .A1(n_349), .A2(n_324), .B1(n_301), .B2(n_335), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_349), .A2(n_335), .B1(n_319), .B2(n_322), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_352), .B(n_329), .Y(n_387) );
OAI221xp5_ASAP7_75t_L g388 ( .A1(n_343), .A2(n_324), .B1(n_341), .B2(n_335), .C(n_253), .Y(n_388) );
OAI22xp33_ASAP7_75t_L g389 ( .A1(n_349), .A2(n_329), .B1(n_319), .B2(n_342), .Y(n_389) );
AND2x6_ASAP7_75t_SL g390 ( .A(n_344), .B(n_297), .Y(n_390) );
AO21x2_ASAP7_75t_L g391 ( .A1(n_354), .A2(n_292), .B(n_311), .Y(n_391) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_367), .A2(n_341), .B1(n_211), .B2(n_215), .C(n_299), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_358), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_349), .A2(n_371), .B1(n_357), .B2(n_366), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_366), .B(n_203), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_359), .Y(n_396) );
BUFx12f_ASAP7_75t_L g397 ( .A(n_344), .Y(n_397) );
A2O1A1Ixp33_ASAP7_75t_L g398 ( .A1(n_363), .A2(n_322), .B(n_253), .C(n_300), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_359), .B(n_300), .Y(n_399) );
INVx1_ASAP7_75t_SL g400 ( .A(n_355), .Y(n_400) );
INVxp67_ASAP7_75t_L g401 ( .A(n_356), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_355), .A2(n_293), .B1(n_334), .B2(n_298), .Y(n_402) );
INVxp67_ASAP7_75t_L g403 ( .A(n_396), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_375), .Y(n_404) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_396), .B(n_373), .Y(n_405) );
INVx2_ASAP7_75t_SL g406 ( .A(n_375), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_377), .B(n_347), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_387), .B(n_368), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_387), .B(n_368), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_375), .B(n_368), .Y(n_410) );
BUFx2_ASAP7_75t_L g411 ( .A(n_376), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_393), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_376), .B(n_368), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_393), .Y(n_414) );
AOI221xp5_ASAP7_75t_L g415 ( .A1(n_377), .A2(n_186), .B1(n_266), .B2(n_200), .C(n_191), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_376), .B(n_347), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_382), .B(n_362), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_393), .Y(n_418) );
BUFx3_ASAP7_75t_L g419 ( .A(n_382), .Y(n_419) );
INVx1_ASAP7_75t_SL g420 ( .A(n_400), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_382), .Y(n_421) );
OAI33xp33_ASAP7_75t_L g422 ( .A1(n_389), .A2(n_183), .A3(n_170), .B1(n_264), .B2(n_261), .B3(n_269), .Y(n_422) );
INVx2_ASAP7_75t_SL g423 ( .A(n_384), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_400), .B(n_360), .Y(n_424) );
BUFx3_ASAP7_75t_L g425 ( .A(n_384), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_384), .B(n_362), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_395), .B(n_362), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_395), .B(n_364), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_401), .B(n_372), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_399), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_391), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_380), .B(n_364), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_391), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_383), .B(n_364), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_391), .Y(n_435) );
BUFx4f_ASAP7_75t_SL g436 ( .A(n_397), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_412), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_412), .Y(n_438) );
INVx2_ASAP7_75t_SL g439 ( .A(n_410), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_436), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_430), .B(n_383), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_412), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_430), .B(n_381), .Y(n_443) );
BUFx2_ASAP7_75t_L g444 ( .A(n_411), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_414), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_411), .B(n_378), .Y(n_446) );
AND2x4_ASAP7_75t_L g447 ( .A(n_419), .B(n_378), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_403), .B(n_394), .Y(n_448) );
OAI221xp5_ASAP7_75t_L g449 ( .A1(n_429), .A2(n_385), .B1(n_388), .B2(n_379), .C(n_386), .Y(n_449) );
INVx2_ASAP7_75t_SL g450 ( .A(n_410), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_406), .B(n_378), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_406), .B(n_360), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_414), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_403), .B(n_390), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_414), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_420), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_418), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_406), .B(n_360), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_423), .B(n_360), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_420), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_408), .B(n_390), .Y(n_461) );
INVx3_ASAP7_75t_L g462 ( .A(n_419), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_407), .B(n_347), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_408), .B(n_409), .Y(n_464) );
CKINVDCx5p33_ASAP7_75t_R g465 ( .A(n_409), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_418), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_423), .B(n_347), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_423), .B(n_347), .Y(n_468) );
INVx1_ASAP7_75t_SL g469 ( .A(n_413), .Y(n_469) );
INVx1_ASAP7_75t_SL g470 ( .A(n_419), .Y(n_470) );
AND2x4_ASAP7_75t_L g471 ( .A(n_425), .B(n_365), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_434), .A2(n_370), .B1(n_397), .B2(n_402), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_418), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_404), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_434), .A2(n_392), .B1(n_397), .B2(n_370), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_413), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_404), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_421), .Y(n_478) );
AO21x2_ASAP7_75t_L g479 ( .A1(n_431), .A2(n_345), .B(n_398), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_407), .B(n_365), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_424), .B(n_200), .Y(n_481) );
INVx3_ASAP7_75t_L g482 ( .A(n_425), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_421), .Y(n_483) );
BUFx2_ASAP7_75t_L g484 ( .A(n_425), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_417), .B(n_365), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_467), .B(n_416), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_467), .B(n_416), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_468), .B(n_424), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_456), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_460), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_468), .B(n_435), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_465), .B(n_432), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_452), .B(n_435), .Y(n_493) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_476), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_474), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_452), .B(n_431), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_458), .B(n_433), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_441), .A2(n_432), .B1(n_428), .B2(n_427), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_438), .Y(n_499) );
INVx3_ASAP7_75t_L g500 ( .A(n_462), .Y(n_500) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_444), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_458), .B(n_433), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_464), .B(n_427), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_459), .B(n_433), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_474), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_469), .B(n_405), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_474), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_477), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_477), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_477), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_478), .Y(n_511) );
INVx3_ASAP7_75t_L g512 ( .A(n_462), .Y(n_512) );
INVxp67_ASAP7_75t_L g513 ( .A(n_454), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_478), .Y(n_514) );
INVx1_ASAP7_75t_SL g515 ( .A(n_440), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_478), .Y(n_516) );
NAND2x1p5_ASAP7_75t_L g517 ( .A(n_484), .B(n_426), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_484), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_438), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_463), .B(n_444), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_483), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_483), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_483), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_480), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_461), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_437), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_459), .B(n_417), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_437), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_439), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_439), .B(n_428), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_463), .B(n_426), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_449), .A2(n_422), .B1(n_415), .B2(n_370), .Y(n_532) );
INVxp67_ASAP7_75t_SL g533 ( .A(n_462), .Y(n_533) );
INVxp67_ASAP7_75t_SL g534 ( .A(n_462), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_443), .B(n_372), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_442), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_450), .B(n_415), .Y(n_537) );
OR2x4_ASAP7_75t_L g538 ( .A(n_448), .B(n_422), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_451), .B(n_345), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_451), .B(n_348), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_446), .B(n_450), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_470), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_438), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_494), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_524), .B(n_446), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_489), .Y(n_546) );
INVx2_ASAP7_75t_SL g547 ( .A(n_529), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_525), .B(n_475), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_490), .Y(n_549) );
NOR3xp33_ASAP7_75t_L g550 ( .A(n_513), .B(n_475), .C(n_481), .Y(n_550) );
INVx1_ASAP7_75t_SL g551 ( .A(n_529), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_541), .B(n_470), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_520), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_535), .A2(n_472), .B1(n_485), .B2(n_447), .Y(n_554) );
INVx1_ASAP7_75t_SL g555 ( .A(n_515), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_520), .Y(n_556) );
OAI21xp5_ASAP7_75t_L g557 ( .A1(n_532), .A2(n_481), .B(n_485), .Y(n_557) );
INVx2_ASAP7_75t_SL g558 ( .A(n_542), .Y(n_558) );
INVx4_ASAP7_75t_L g559 ( .A(n_517), .Y(n_559) );
INVxp33_ASAP7_75t_L g560 ( .A(n_517), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_503), .B(n_455), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_541), .B(n_482), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_491), .B(n_455), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_526), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_499), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_491), .B(n_466), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_527), .B(n_482), .Y(n_567) );
INVxp67_ASAP7_75t_L g568 ( .A(n_501), .Y(n_568) );
AND2x4_ASAP7_75t_L g569 ( .A(n_500), .B(n_447), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_499), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_500), .B(n_447), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_527), .B(n_482), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_486), .B(n_487), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_486), .B(n_466), .Y(n_574) );
NAND2x1_ASAP7_75t_SL g575 ( .A(n_500), .B(n_482), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_487), .B(n_471), .Y(n_576) );
INVx1_ASAP7_75t_SL g577 ( .A(n_518), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_493), .B(n_442), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_528), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_493), .B(n_445), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_498), .A2(n_447), .B1(n_471), .B2(n_479), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_496), .B(n_453), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_496), .B(n_453), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_531), .B(n_457), .Y(n_584) );
INVx2_ASAP7_75t_SL g585 ( .A(n_517), .Y(n_585) );
AOI322xp5_ASAP7_75t_L g586 ( .A1(n_492), .A2(n_473), .A3(n_457), .B1(n_445), .B2(n_471), .C1(n_266), .C2(n_200), .Y(n_586) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_533), .A2(n_473), .B(n_471), .Y(n_587) );
OAI21x1_ASAP7_75t_L g588 ( .A1(n_512), .A2(n_537), .B(n_534), .Y(n_588) );
NOR2x1_ASAP7_75t_L g589 ( .A(n_512), .B(n_479), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_536), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_531), .B(n_479), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_488), .B(n_191), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_488), .B(n_76), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_530), .B(n_348), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_497), .B(n_191), .Y(n_595) );
NOR2x2_ASAP7_75t_L g596 ( .A(n_519), .B(n_302), .Y(n_596) );
O2A1O1Ixp33_ASAP7_75t_L g597 ( .A1(n_544), .A2(n_506), .B(n_512), .C(n_508), .Y(n_597) );
OAI21xp33_ASAP7_75t_L g598 ( .A1(n_581), .A2(n_506), .B(n_539), .Y(n_598) );
OAI21xp5_ASAP7_75t_L g599 ( .A1(n_587), .A2(n_507), .B(n_508), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_573), .B(n_497), .Y(n_600) );
A2O1A1Ixp33_ASAP7_75t_L g601 ( .A1(n_560), .A2(n_507), .B(n_509), .C(n_510), .Y(n_601) );
INVx2_ASAP7_75t_SL g602 ( .A(n_547), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_544), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_550), .A2(n_539), .B1(n_540), .B2(n_502), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_551), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_553), .B(n_556), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_587), .A2(n_538), .B(n_510), .Y(n_607) );
OAI211xp5_ASAP7_75t_L g608 ( .A1(n_581), .A2(n_540), .B(n_509), .C(n_504), .Y(n_608) );
INVx2_ASAP7_75t_SL g609 ( .A(n_555), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_545), .B(n_538), .Y(n_610) );
INVxp67_ASAP7_75t_L g611 ( .A(n_558), .Y(n_611) );
OAI21xp5_ASAP7_75t_L g612 ( .A1(n_586), .A2(n_505), .B(n_495), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_546), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_549), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_550), .A2(n_538), .B1(n_502), .B2(n_504), .Y(n_615) );
OAI22xp33_ASAP7_75t_L g616 ( .A1(n_559), .A2(n_511), .B1(n_523), .B2(n_514), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_559), .B(n_585), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_561), .B(n_574), .Y(n_618) );
INVx1_ASAP7_75t_SL g619 ( .A(n_596), .Y(n_619) );
AOI31xp33_ASAP7_75t_L g620 ( .A1(n_560), .A2(n_516), .A3(n_522), .B(n_521), .Y(n_620) );
NAND4xp25_ASAP7_75t_SL g621 ( .A(n_554), .B(n_543), .C(n_519), .D(n_361), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_548), .A2(n_543), .B1(n_370), .B2(n_372), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_577), .B(n_372), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_557), .A2(n_593), .B1(n_568), .B2(n_594), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_568), .B(n_200), .Y(n_625) );
AO22x1_ASAP7_75t_L g626 ( .A1(n_596), .A2(n_334), .B1(n_298), .B2(n_293), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_576), .B(n_584), .Y(n_627) );
OAI22xp33_ASAP7_75t_SL g628 ( .A1(n_563), .A2(n_369), .B1(n_173), .B2(n_310), .Y(n_628) );
OAI21xp5_ASAP7_75t_SL g629 ( .A1(n_569), .A2(n_369), .B(n_334), .Y(n_629) );
OAI32xp33_ASAP7_75t_L g630 ( .A1(n_566), .A2(n_369), .A3(n_173), .B1(n_302), .B2(n_327), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_578), .A2(n_334), .B1(n_318), .B2(n_179), .Y(n_631) );
INVx4_ASAP7_75t_L g632 ( .A(n_569), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_565), .Y(n_633) );
NAND4xp25_ASAP7_75t_L g634 ( .A(n_592), .B(n_173), .C(n_242), .D(n_232), .Y(n_634) );
NOR3xp33_ASAP7_75t_L g635 ( .A(n_621), .B(n_595), .C(n_588), .Y(n_635) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_603), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_613), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_633), .Y(n_638) );
XNOR2xp5_ASAP7_75t_L g639 ( .A(n_605), .B(n_602), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_615), .B(n_580), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_614), .Y(n_641) );
NAND3xp33_ASAP7_75t_L g642 ( .A(n_607), .B(n_589), .C(n_591), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_606), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_598), .A2(n_571), .B1(n_569), .B2(n_562), .Y(n_644) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_609), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_600), .Y(n_646) );
AOI211xp5_ASAP7_75t_L g647 ( .A1(n_619), .A2(n_571), .B(n_567), .C(n_572), .Y(n_647) );
NOR4xp25_ASAP7_75t_L g648 ( .A(n_611), .B(n_590), .C(n_579), .D(n_564), .Y(n_648) );
INVxp67_ASAP7_75t_SL g649 ( .A(n_597), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_610), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_618), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_604), .B(n_583), .Y(n_652) );
A2O1A1Ixp33_ASAP7_75t_L g653 ( .A1(n_620), .A2(n_575), .B(n_552), .C(n_571), .Y(n_653) );
AO22x2_ASAP7_75t_L g654 ( .A1(n_608), .A2(n_570), .B1(n_565), .B2(n_582), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_625), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_624), .B(n_570), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_612), .B(n_179), .Y(n_657) );
O2A1O1Ixp5_ASAP7_75t_L g658 ( .A1(n_649), .A2(n_626), .B(n_617), .C(n_632), .Y(n_658) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_649), .A2(n_627), .B1(n_599), .B2(n_616), .C(n_632), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_650), .A2(n_623), .B1(n_634), .B2(n_628), .Y(n_660) );
AOI32xp33_ASAP7_75t_L g661 ( .A1(n_654), .A2(n_631), .A3(n_601), .B1(n_629), .B2(n_634), .Y(n_661) );
NAND5xp2_ASAP7_75t_L g662 ( .A(n_635), .B(n_622), .C(n_630), .D(n_179), .E(n_358), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_636), .Y(n_663) );
AOI211xp5_ASAP7_75t_L g664 ( .A1(n_648), .A2(n_327), .B(n_323), .C(n_312), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_637), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_652), .A2(n_312), .B1(n_311), .B2(n_318), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_640), .A2(n_318), .B1(n_246), .B2(n_254), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_641), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_653), .A2(n_318), .B(n_246), .Y(n_669) );
OAI22xp33_ASAP7_75t_L g670 ( .A1(n_645), .A2(n_232), .B1(n_254), .B2(n_260), .Y(n_670) );
XOR2x2_ASAP7_75t_L g671 ( .A(n_639), .B(n_260), .Y(n_671) );
AOI211xp5_ASAP7_75t_L g672 ( .A1(n_659), .A2(n_635), .B(n_642), .C(n_655), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_665), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_663), .B(n_651), .Y(n_674) );
AOI211xp5_ASAP7_75t_L g675 ( .A1(n_662), .A2(n_647), .B(n_656), .C(n_657), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_660), .A2(n_644), .B1(n_654), .B2(n_643), .Y(n_676) );
OAI311xp33_ASAP7_75t_L g677 ( .A1(n_661), .A2(n_654), .A3(n_646), .B1(n_638), .C1(n_289), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_668), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_671), .A2(n_270), .B1(n_274), .B2(n_289), .Y(n_679) );
INVx1_ASAP7_75t_SL g680 ( .A(n_674), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_678), .Y(n_681) );
NOR3xp33_ASAP7_75t_L g682 ( .A(n_672), .B(n_658), .C(n_670), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_673), .Y(n_683) );
NAND3xp33_ASAP7_75t_SL g684 ( .A(n_682), .B(n_676), .C(n_675), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_681), .Y(n_685) );
XNOR2xp5_ASAP7_75t_L g686 ( .A(n_680), .B(n_679), .Y(n_686) );
NOR3xp33_ASAP7_75t_L g687 ( .A(n_684), .B(n_683), .C(n_677), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_685), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_687), .A2(n_686), .B1(n_664), .B2(n_666), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_689), .A2(n_688), .B1(n_667), .B2(n_669), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_690), .Y(n_691) );
BUFx3_ASAP7_75t_L g692 ( .A(n_691), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_692), .A2(n_270), .B1(n_274), .B2(n_684), .Y(n_693) );
endmodule