module fake_ariane_151_n_748 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_748);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_748;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_677;
wire n_614;
wire n_604;
wire n_222;
wire n_478;
wire n_703;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_655;
wire n_544;
wire n_216;
wire n_692;
wire n_540;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_289;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

INVxp33_ASAP7_75t_L g155 ( 
.A(n_34),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_24),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_19),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_123),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_111),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_113),
.B(n_31),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_97),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_35),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_6),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_103),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_19),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_83),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_44),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_0),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_68),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_7),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_153),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_2),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_14),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_67),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_96),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_110),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_147),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_48),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_40),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_134),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_36),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_93),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_124),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_127),
.B(n_2),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_52),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_14),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_5),
.B(n_74),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_69),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_38),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_128),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_104),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_114),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_26),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_94),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_54),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_118),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_32),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_79),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_84),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_106),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_109),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_16),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_28),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_107),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_177),
.Y(n_211)
);

AND2x4_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_0),
.Y(n_212)
);

OA21x2_ASAP7_75t_L g213 ( 
.A1(n_159),
.A2(n_1),
.B(n_3),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_183),
.B(n_1),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_183),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_157),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_170),
.Y(n_218)
);

AND2x6_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_20),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_168),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_170),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_172),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_170),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_175),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_160),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_156),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g229 ( 
.A(n_208),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_178),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_192),
.Y(n_231)
);

AND2x4_ASAP7_75t_L g232 ( 
.A(n_161),
.B(n_162),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_188),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_173),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_176),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_180),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_170),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_187),
.Y(n_238)
);

OA21x2_ASAP7_75t_L g239 ( 
.A1(n_181),
.A2(n_8),
.B(n_9),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_185),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_206),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_194),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_155),
.B(n_8),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_195),
.B(n_9),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_188),
.Y(n_245)
);

AND2x4_ASAP7_75t_L g246 ( 
.A(n_197),
.B(n_10),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_201),
.B(n_10),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_207),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

AND2x4_ASAP7_75t_L g250 ( 
.A(n_202),
.B(n_11),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_204),
.Y(n_251)
);

OAI21x1_ASAP7_75t_L g252 ( 
.A1(n_209),
.A2(n_80),
.B(n_151),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_170),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_215),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_211),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_L g256 ( 
.A1(n_216),
.A2(n_235),
.B1(n_214),
.B2(n_241),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_211),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_215),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_217),
.Y(n_259)
);

AOI21x1_ASAP7_75t_L g260 ( 
.A1(n_218),
.A2(n_163),
.B(n_171),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_216),
.A2(n_189),
.B1(n_205),
.B2(n_193),
.Y(n_261)
);

NAND2xp33_ASAP7_75t_L g262 ( 
.A(n_219),
.B(n_170),
.Y(n_262)
);

NOR2x1p5_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_158),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_250),
.A2(n_193),
.B1(n_169),
.B2(n_203),
.Y(n_264)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_217),
.Y(n_265)
);

NAND2xp33_ASAP7_75t_L g266 ( 
.A(n_219),
.B(n_199),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_230),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_223),
.Y(n_268)
);

NAND2xp33_ASAP7_75t_L g269 ( 
.A(n_219),
.B(n_199),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_223),
.Y(n_270)
);

NOR2x1p5_ASAP7_75t_L g271 ( 
.A(n_229),
.B(n_164),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_226),
.Y(n_272)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_219),
.Y(n_273)
);

NAND3xp33_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_169),
.C(n_203),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_241),
.B(n_165),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_226),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_215),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_215),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_236),
.B(n_240),
.Y(n_279)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_219),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_238),
.Y(n_281)
);

AND2x6_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_199),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_222),
.B(n_11),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_231),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_231),
.Y(n_285)
);

NAND2xp33_ASAP7_75t_L g286 ( 
.A(n_219),
.B(n_203),
.Y(n_286)
);

INVx2_ASAP7_75t_SL g287 ( 
.A(n_222),
.Y(n_287)
);

INVx2_ASAP7_75t_SL g288 ( 
.A(n_246),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_250),
.B(n_167),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_215),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_225),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_212),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_220),
.Y(n_293)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_219),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_232),
.B(n_174),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_246),
.B(n_179),
.Y(n_296)
);

INVxp33_ASAP7_75t_L g297 ( 
.A(n_238),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_246),
.B(n_182),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_225),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_232),
.B(n_184),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_227),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_232),
.B(n_186),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_268),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_256),
.A2(n_228),
.B1(n_212),
.B2(n_244),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_212),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_281),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_270),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_301),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_227),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_264),
.A2(n_234),
.B1(n_248),
.B2(n_247),
.Y(n_310)
);

A2O1A1Ixp33_ASAP7_75t_L g311 ( 
.A1(n_292),
.A2(n_240),
.B(n_236),
.C(n_242),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_254),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_255),
.Y(n_313)
);

AND2x4_ASAP7_75t_L g314 ( 
.A(n_279),
.B(n_234),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_301),
.B(n_242),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_259),
.B(n_191),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_272),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_257),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_251),
.Y(n_319)
);

NAND3xp33_ASAP7_75t_L g320 ( 
.A(n_261),
.B(n_213),
.C(n_239),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_276),
.Y(n_321)
);

O2A1O1Ixp5_ASAP7_75t_L g322 ( 
.A1(n_292),
.A2(n_220),
.B(n_224),
.C(n_221),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_282),
.B(n_251),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_279),
.Y(n_324)
);

BUFx8_ASAP7_75t_L g325 ( 
.A(n_259),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_254),
.Y(n_326)
);

INVx8_ASAP7_75t_L g327 ( 
.A(n_282),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_258),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_258),
.Y(n_329)
);

NOR2xp67_ASAP7_75t_L g330 ( 
.A(n_287),
.B(n_251),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_284),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_287),
.B(n_196),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_281),
.A2(n_239),
.B1(n_213),
.B2(n_220),
.Y(n_333)
);

NOR3x1_ASAP7_75t_L g334 ( 
.A(n_283),
.B(n_12),
.C(n_13),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_265),
.B(n_198),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_275),
.B(n_218),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_262),
.A2(n_213),
.B1(n_239),
.B2(n_200),
.Y(n_337)
);

AND3x1_ASAP7_75t_L g338 ( 
.A(n_300),
.B(n_253),
.C(n_237),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_295),
.B(n_221),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_302),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_262),
.A2(n_213),
.B1(n_239),
.B2(n_224),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g342 ( 
.A1(n_282),
.A2(n_237),
.B1(n_253),
.B2(n_203),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_265),
.B(n_210),
.Y(n_343)
);

OAI22xp33_ASAP7_75t_L g344 ( 
.A1(n_296),
.A2(n_225),
.B1(n_233),
.B2(n_245),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_282),
.B(n_225),
.Y(n_345)
);

OR2x6_ASAP7_75t_L g346 ( 
.A(n_263),
.B(n_252),
.Y(n_346)
);

NAND3xp33_ASAP7_75t_L g347 ( 
.A(n_266),
.B(n_249),
.C(n_245),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_285),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_298),
.B(n_225),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_297),
.B(n_252),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_277),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_277),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_278),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_282),
.B(n_233),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_282),
.A2(n_245),
.B1(n_233),
.B2(n_249),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_278),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_267),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_293),
.B(n_289),
.Y(n_358)
);

NAND2x1p5_ASAP7_75t_L g359 ( 
.A(n_271),
.B(n_233),
.Y(n_359)
);

OAI22x1_ASAP7_75t_L g360 ( 
.A1(n_297),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_360)
);

NOR3xp33_ASAP7_75t_L g361 ( 
.A(n_274),
.B(n_15),
.C(n_16),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_266),
.B(n_233),
.Y(n_362)
);

A2O1A1Ixp33_ASAP7_75t_L g363 ( 
.A1(n_269),
.A2(n_249),
.B(n_245),
.C(n_17),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_273),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_273),
.B(n_245),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_260),
.B(n_249),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_269),
.A2(n_249),
.B1(n_18),
.B2(n_17),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_305),
.B(n_286),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_339),
.A2(n_286),
.B(n_294),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_325),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_306),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_340),
.B(n_273),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_365),
.A2(n_294),
.B(n_280),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_364),
.A2(n_294),
.B(n_280),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_314),
.B(n_280),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_303),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_307),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_338),
.A2(n_299),
.B1(n_291),
.B2(n_290),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_327),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_317),
.Y(n_380)
);

INVx4_ASAP7_75t_L g381 ( 
.A(n_327),
.Y(n_381)
);

INVxp33_ASAP7_75t_L g382 ( 
.A(n_330),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_314),
.B(n_290),
.Y(n_383)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_324),
.B(n_18),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_308),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_322),
.A2(n_299),
.B(n_291),
.Y(n_386)
);

OAI321xp33_ASAP7_75t_L g387 ( 
.A1(n_304),
.A2(n_21),
.A3(n_22),
.B1(n_23),
.B2(n_25),
.C(n_27),
.Y(n_387)
);

NOR2x1_ASAP7_75t_R g388 ( 
.A(n_316),
.B(n_29),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_304),
.B(n_30),
.Y(n_389)
);

OAI21x1_ASAP7_75t_L g390 ( 
.A1(n_341),
.A2(n_33),
.B(n_37),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_309),
.B(n_338),
.Y(n_391)
);

A2O1A1Ixp33_ASAP7_75t_L g392 ( 
.A1(n_336),
.A2(n_39),
.B(n_41),
.C(n_42),
.Y(n_392)
);

AO21x2_ASAP7_75t_L g393 ( 
.A1(n_337),
.A2(n_43),
.B(n_45),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_325),
.Y(n_394)
);

NAND2xp33_ASAP7_75t_L g395 ( 
.A(n_327),
.B(n_46),
.Y(n_395)
);

NAND2x1p5_ASAP7_75t_L g396 ( 
.A(n_348),
.B(n_47),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_364),
.A2(n_319),
.B(n_358),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_315),
.B(n_49),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_366),
.A2(n_331),
.B(n_321),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_310),
.B(n_50),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_350),
.Y(n_401)
);

A2O1A1Ixp33_ASAP7_75t_L g402 ( 
.A1(n_333),
.A2(n_51),
.B(n_53),
.C(n_55),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_346),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_357),
.B(n_154),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_349),
.A2(n_56),
.B(n_57),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_335),
.B(n_58),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_332),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_359),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_362),
.A2(n_62),
.B(n_63),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_343),
.B(n_64),
.Y(n_410)
);

NOR3xp33_ASAP7_75t_L g411 ( 
.A(n_361),
.B(n_65),
.C(n_66),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_313),
.B(n_149),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_311),
.A2(n_70),
.B(n_71),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_318),
.B(n_72),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_345),
.A2(n_73),
.B(n_75),
.Y(n_415)
);

AO32x2_ASAP7_75t_L g416 ( 
.A1(n_333),
.A2(n_76),
.A3(n_77),
.B1(n_78),
.B2(n_81),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_354),
.A2(n_82),
.B(n_85),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_346),
.A2(n_86),
.B(n_87),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_323),
.B(n_148),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_320),
.B(n_88),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_334),
.B(n_89),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_337),
.B(n_90),
.Y(n_422)
);

AO22x1_ASAP7_75t_L g423 ( 
.A1(n_360),
.A2(n_145),
.B1(n_92),
.B2(n_95),
.Y(n_423)
);

A2O1A1Ixp33_ASAP7_75t_L g424 ( 
.A1(n_367),
.A2(n_91),
.B(n_98),
.C(n_99),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_346),
.A2(n_101),
.B(n_102),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_342),
.A2(n_105),
.B1(n_108),
.B2(n_112),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_312),
.B(n_115),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_312),
.B(n_143),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_326),
.A2(n_328),
.B(n_329),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_347),
.B(n_116),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_352),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_353),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_312),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_351),
.B(n_142),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_351),
.B(n_117),
.Y(n_435)
);

A2O1A1Ixp33_ASAP7_75t_L g436 ( 
.A1(n_363),
.A2(n_119),
.B(n_120),
.C(n_121),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_351),
.A2(n_122),
.B(n_125),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_371),
.Y(n_438)
);

AO22x2_ASAP7_75t_L g439 ( 
.A1(n_389),
.A2(n_344),
.B1(n_355),
.B2(n_356),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_399),
.A2(n_355),
.B(n_356),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_401),
.B(n_356),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_376),
.B(n_126),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_377),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_380),
.B(n_129),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_400),
.B(n_130),
.Y(n_445)
);

AOI21x1_ASAP7_75t_L g446 ( 
.A1(n_422),
.A2(n_131),
.B(n_132),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_379),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_370),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_374),
.A2(n_133),
.B(n_135),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_385),
.Y(n_450)
);

OAI21x1_ASAP7_75t_L g451 ( 
.A1(n_390),
.A2(n_136),
.B(n_137),
.Y(n_451)
);

BUFx4_ASAP7_75t_SL g452 ( 
.A(n_403),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_384),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_432),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_398),
.A2(n_140),
.B1(n_141),
.B2(n_375),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_372),
.B(n_368),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_397),
.A2(n_369),
.B(n_373),
.Y(n_457)
);

OR2x2_ASAP7_75t_L g458 ( 
.A(n_394),
.B(n_408),
.Y(n_458)
);

NAND2x1_ASAP7_75t_L g459 ( 
.A(n_381),
.B(n_379),
.Y(n_459)
);

A2O1A1Ixp33_ASAP7_75t_L g460 ( 
.A1(n_420),
.A2(n_391),
.B(n_406),
.C(n_424),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_381),
.A2(n_402),
.B(n_434),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_382),
.B(n_421),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_404),
.A2(n_386),
.B(n_395),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_431),
.B(n_383),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_433),
.B(n_379),
.Y(n_465)
);

AO22x2_ASAP7_75t_L g466 ( 
.A1(n_416),
.A2(n_393),
.B1(n_423),
.B2(n_387),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_396),
.A2(n_410),
.B1(n_425),
.B2(n_418),
.Y(n_467)
);

NOR2xp67_ASAP7_75t_L g468 ( 
.A(n_378),
.B(n_412),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_413),
.A2(n_436),
.B(n_411),
.Y(n_469)
);

OAI21x1_ASAP7_75t_L g470 ( 
.A1(n_419),
.A2(n_429),
.B(n_435),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_433),
.B(n_388),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_416),
.Y(n_472)
);

OAI21x1_ASAP7_75t_L g473 ( 
.A1(n_427),
.A2(n_428),
.B(n_414),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_392),
.A2(n_405),
.B(n_409),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_415),
.A2(n_417),
.B(n_407),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_416),
.B(n_396),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_433),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_393),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_430),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_426),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_437),
.A2(n_322),
.B(n_399),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_376),
.Y(n_482)
);

OAI21x1_ASAP7_75t_L g483 ( 
.A1(n_390),
.A2(n_386),
.B(n_419),
.Y(n_483)
);

OAI21x1_ASAP7_75t_L g484 ( 
.A1(n_390),
.A2(n_386),
.B(n_419),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_401),
.B(n_308),
.Y(n_485)
);

NAND3xp33_ASAP7_75t_SL g486 ( 
.A(n_370),
.B(n_304),
.C(n_281),
.Y(n_486)
);

BUFx4f_ASAP7_75t_L g487 ( 
.A(n_396),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_374),
.A2(n_364),
.B(n_397),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_374),
.A2(n_364),
.B(n_397),
.Y(n_489)
);

OAI21x1_ASAP7_75t_L g490 ( 
.A1(n_390),
.A2(n_386),
.B(n_419),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_401),
.B(n_308),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_389),
.A2(n_304),
.B1(n_288),
.B2(n_422),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_472),
.B(n_482),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_438),
.Y(n_494)
);

AO31x2_ASAP7_75t_L g495 ( 
.A1(n_478),
.A2(n_460),
.A3(n_492),
.B(n_467),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_447),
.Y(n_496)
);

AOI21x1_ASAP7_75t_L g497 ( 
.A1(n_463),
.A2(n_457),
.B(n_490),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_443),
.Y(n_498)
);

OA21x2_ASAP7_75t_L g499 ( 
.A1(n_470),
.A2(n_474),
.B(n_473),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_454),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_446),
.Y(n_501)
);

OAI21x1_ASAP7_75t_L g502 ( 
.A1(n_451),
.A2(n_474),
.B(n_475),
.Y(n_502)
);

AO21x2_ASAP7_75t_L g503 ( 
.A1(n_476),
.A2(n_481),
.B(n_475),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_442),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_444),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_456),
.A2(n_488),
.B(n_489),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_480),
.A2(n_481),
.B(n_468),
.Y(n_507)
);

OA21x2_ASAP7_75t_L g508 ( 
.A1(n_469),
.A2(n_440),
.B(n_445),
.Y(n_508)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_492),
.B(n_453),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_469),
.A2(n_467),
.B(n_440),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_466),
.Y(n_511)
);

BUFx2_ASAP7_75t_SL g512 ( 
.A(n_479),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_477),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_449),
.A2(n_461),
.B(n_479),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_441),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_447),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_464),
.B(n_462),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_450),
.Y(n_518)
);

NOR2xp67_ASAP7_75t_L g519 ( 
.A(n_465),
.B(n_447),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_485),
.A2(n_491),
.B(n_455),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_487),
.A2(n_466),
.B(n_459),
.Y(n_521)
);

OAI21x1_ASAP7_75t_L g522 ( 
.A1(n_471),
.A2(n_486),
.B(n_439),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_439),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g524 ( 
.A1(n_487),
.A2(n_458),
.B(n_452),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_448),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_485),
.B(n_308),
.Y(n_526)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_483),
.A2(n_490),
.B(n_484),
.Y(n_527)
);

OAI21x1_ASAP7_75t_SL g528 ( 
.A1(n_469),
.A2(n_467),
.B(n_474),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_466),
.A2(n_261),
.B1(n_492),
.B2(n_400),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_454),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_443),
.Y(n_531)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_438),
.B(n_443),
.Y(n_532)
);

AOI21xp33_ASAP7_75t_SL g533 ( 
.A1(n_450),
.A2(n_306),
.B(n_228),
.Y(n_533)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_438),
.B(n_443),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_493),
.B(n_517),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_516),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_493),
.B(n_509),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_503),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_498),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_516),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_517),
.B(n_509),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_498),
.Y(n_542)
);

AO21x2_ASAP7_75t_L g543 ( 
.A1(n_501),
.A2(n_528),
.B(n_510),
.Y(n_543)
);

OR2x6_ASAP7_75t_L g544 ( 
.A(n_521),
.B(n_512),
.Y(n_544)
);

OAI21x1_ASAP7_75t_L g545 ( 
.A1(n_527),
.A2(n_497),
.B(n_502),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_531),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_531),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_523),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_503),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_523),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_495),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_495),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_500),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_529),
.B(n_515),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_500),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_530),
.Y(n_556)
);

OAI21x1_ASAP7_75t_SL g557 ( 
.A1(n_507),
.A2(n_506),
.B(n_504),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_494),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_494),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_515),
.B(n_512),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_516),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_495),
.Y(n_562)
);

AO31x2_ASAP7_75t_L g563 ( 
.A1(n_511),
.A2(n_505),
.A3(n_504),
.B(n_495),
.Y(n_563)
);

OR2x2_ASAP7_75t_L g564 ( 
.A(n_532),
.B(n_534),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_524),
.Y(n_565)
);

INVx1_ASAP7_75t_SL g566 ( 
.A(n_564),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_564),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_539),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_539),
.Y(n_569)
);

AO21x2_ASAP7_75t_L g570 ( 
.A1(n_557),
.A2(n_522),
.B(n_511),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_541),
.B(n_522),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_535),
.B(n_534),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_535),
.B(n_508),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_542),
.Y(n_574)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_537),
.B(n_532),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_559),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_537),
.B(n_508),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_565),
.B(n_496),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_559),
.B(n_518),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_548),
.B(n_508),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_558),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_546),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_543),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_547),
.B(n_554),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_556),
.Y(n_585)
);

OR2x2_ASAP7_75t_SL g586 ( 
.A(n_547),
.B(n_525),
.Y(n_586)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_536),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_554),
.A2(n_505),
.B1(n_520),
.B2(n_525),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_560),
.B(n_553),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_563),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_536),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_536),
.Y(n_592)
);

NAND2x1p5_ASAP7_75t_L g593 ( 
.A(n_565),
.B(n_514),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_565),
.A2(n_533),
.B1(n_526),
.B2(n_496),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_543),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_548),
.B(n_524),
.Y(n_596)
);

INVx2_ASAP7_75t_SL g597 ( 
.A(n_536),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_553),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_543),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_536),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_550),
.B(n_499),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_555),
.B(n_513),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_550),
.B(n_499),
.Y(n_603)
);

AOI221xp5_ASAP7_75t_L g604 ( 
.A1(n_551),
.A2(n_533),
.B1(n_513),
.B2(n_496),
.C(n_519),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_566),
.B(n_555),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_567),
.B(n_563),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_578),
.Y(n_607)
);

INVxp33_ASAP7_75t_L g608 ( 
.A(n_572),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_580),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_573),
.B(n_562),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_573),
.B(n_552),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_568),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_577),
.B(n_552),
.Y(n_613)
);

NAND2x1_ASAP7_75t_L g614 ( 
.A(n_592),
.B(n_557),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_585),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_580),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_569),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_577),
.B(n_552),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_571),
.B(n_551),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g620 ( 
.A(n_575),
.B(n_551),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_576),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_571),
.B(n_584),
.Y(n_622)
);

NAND2xp67_ASAP7_75t_L g623 ( 
.A(n_584),
.B(n_538),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_596),
.Y(n_624)
);

INVxp67_ASAP7_75t_SL g625 ( 
.A(n_581),
.Y(n_625)
);

NOR2xp67_ASAP7_75t_L g626 ( 
.A(n_592),
.B(n_549),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_574),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_582),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_598),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_589),
.B(n_549),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_575),
.B(n_563),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_601),
.B(n_603),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_579),
.B(n_602),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_601),
.B(n_538),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_588),
.B(n_563),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_603),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_621),
.B(n_594),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_617),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_633),
.B(n_596),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_617),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_607),
.B(n_578),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_628),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_628),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_625),
.B(n_597),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_622),
.B(n_597),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_615),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_607),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_612),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_627),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_632),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_624),
.B(n_578),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_629),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_622),
.B(n_600),
.Y(n_653)
);

AOI21xp33_ASAP7_75t_L g654 ( 
.A1(n_635),
.A2(n_570),
.B(n_590),
.Y(n_654)
);

HB1xp67_ASAP7_75t_SL g655 ( 
.A(n_620),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_610),
.B(n_600),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_605),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_620),
.Y(n_658)
);

OR2x2_ASAP7_75t_L g659 ( 
.A(n_619),
.B(n_586),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_609),
.Y(n_660)
);

OR2x2_ASAP7_75t_L g661 ( 
.A(n_619),
.B(n_586),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_631),
.B(n_599),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_624),
.B(n_544),
.Y(n_663)
);

OAI31xp33_ASAP7_75t_L g664 ( 
.A1(n_608),
.A2(n_583),
.A3(n_599),
.B(n_595),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_609),
.Y(n_665)
);

NAND2xp33_ASAP7_75t_L g666 ( 
.A(n_616),
.B(n_536),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_638),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_647),
.B(n_632),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_650),
.B(n_616),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_662),
.B(n_636),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_653),
.B(n_610),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_644),
.B(n_592),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_656),
.B(n_611),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_640),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_651),
.B(n_636),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_642),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_651),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_651),
.B(n_611),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_645),
.B(n_618),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_660),
.B(n_665),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_643),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_648),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_637),
.B(n_630),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_639),
.B(n_613),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_646),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_676),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_682),
.B(n_637),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_682),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_668),
.Y(n_689)
);

AOI21xp33_ASAP7_75t_L g690 ( 
.A1(n_683),
.A2(n_664),
.B(n_657),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_676),
.Y(n_691)
);

NOR4xp25_ASAP7_75t_L g692 ( 
.A(n_669),
.B(n_649),
.C(n_652),
.D(n_654),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_672),
.A2(n_666),
.B(n_641),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_679),
.B(n_658),
.Y(n_694)
);

NOR2x1_ASAP7_75t_L g695 ( 
.A(n_677),
.B(n_681),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_681),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_689),
.B(n_668),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_695),
.Y(n_698)
);

AOI221xp5_ASAP7_75t_L g699 ( 
.A1(n_692),
.A2(n_667),
.B1(n_674),
.B2(n_680),
.C(n_684),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_693),
.A2(n_641),
.B(n_666),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_686),
.Y(n_701)
);

INVxp67_ASAP7_75t_L g702 ( 
.A(n_687),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_688),
.Y(n_703)
);

NAND3xp33_ASAP7_75t_L g704 ( 
.A(n_699),
.B(n_690),
.C(n_691),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_699),
.A2(n_690),
.B(n_696),
.Y(n_705)
);

OAI21xp33_ASAP7_75t_L g706 ( 
.A1(n_702),
.A2(n_694),
.B(n_680),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_700),
.A2(n_659),
.B1(n_661),
.B2(n_655),
.Y(n_707)
);

OAI21xp33_ASAP7_75t_L g708 ( 
.A1(n_698),
.A2(n_668),
.B(n_670),
.Y(n_708)
);

NOR4xp25_ASAP7_75t_L g709 ( 
.A(n_704),
.B(n_701),
.C(n_697),
.D(n_670),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_706),
.B(n_703),
.Y(n_710)
);

NOR3x1_ASAP7_75t_L g711 ( 
.A(n_705),
.B(n_677),
.C(n_614),
.Y(n_711)
);

NAND3xp33_ASAP7_75t_SL g712 ( 
.A(n_707),
.B(n_614),
.C(n_678),
.Y(n_712)
);

OAI21xp33_ASAP7_75t_L g713 ( 
.A1(n_708),
.A2(n_675),
.B(n_679),
.Y(n_713)
);

NOR3xp33_ASAP7_75t_L g714 ( 
.A(n_712),
.B(n_604),
.C(n_496),
.Y(n_714)
);

NOR2x1_ASAP7_75t_L g715 ( 
.A(n_710),
.B(n_671),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_711),
.B(n_671),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_715),
.B(n_709),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_714),
.Y(n_718)
);

NOR2x1_ASAP7_75t_L g719 ( 
.A(n_716),
.B(n_713),
.Y(n_719)
);

NAND2x1_ASAP7_75t_L g720 ( 
.A(n_716),
.B(n_675),
.Y(n_720)
);

AND2x2_ASAP7_75t_SL g721 ( 
.A(n_717),
.B(n_675),
.Y(n_721)
);

AND3x4_ASAP7_75t_L g722 ( 
.A(n_719),
.B(n_663),
.C(n_655),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_720),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_718),
.Y(n_724)
);

OAI21xp5_ASAP7_75t_L g725 ( 
.A1(n_717),
.A2(n_678),
.B(n_673),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_717),
.A2(n_544),
.B1(n_663),
.B2(n_606),
.Y(n_726)
);

OA22x2_ASAP7_75t_L g727 ( 
.A1(n_722),
.A2(n_673),
.B1(n_663),
.B2(n_544),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_SL g728 ( 
.A1(n_724),
.A2(n_544),
.B1(n_540),
.B2(n_561),
.Y(n_728)
);

NAND4xp25_ASAP7_75t_L g729 ( 
.A(n_725),
.B(n_519),
.C(n_591),
.D(n_587),
.Y(n_729)
);

XOR2xp5_ASAP7_75t_L g730 ( 
.A(n_721),
.B(n_561),
.Y(n_730)
);

OR2x6_ASAP7_75t_L g731 ( 
.A(n_723),
.B(n_540),
.Y(n_731)
);

BUFx12f_ASAP7_75t_L g732 ( 
.A(n_726),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_724),
.Y(n_733)
);

OAI21x1_ASAP7_75t_L g734 ( 
.A1(n_733),
.A2(n_685),
.B(n_591),
.Y(n_734)
);

AOI21xp33_ASAP7_75t_L g735 ( 
.A1(n_730),
.A2(n_561),
.B(n_570),
.Y(n_735)
);

OAI21x1_ASAP7_75t_L g736 ( 
.A1(n_727),
.A2(n_685),
.B(n_591),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_729),
.B(n_731),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_732),
.Y(n_738)
);

OAI21xp5_ASAP7_75t_SL g739 ( 
.A1(n_738),
.A2(n_728),
.B(n_561),
.Y(n_739)
);

OAI21xp5_ASAP7_75t_L g740 ( 
.A1(n_737),
.A2(n_544),
.B(n_626),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_735),
.A2(n_570),
.B1(n_583),
.B2(n_595),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_734),
.B(n_623),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_739),
.A2(n_736),
.B1(n_593),
.B2(n_561),
.Y(n_743)
);

OAI22xp33_ASAP7_75t_L g744 ( 
.A1(n_742),
.A2(n_561),
.B1(n_593),
.B2(n_634),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_744),
.B(n_743),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_743),
.B(n_740),
.Y(n_746)
);

AO21x2_ASAP7_75t_L g747 ( 
.A1(n_745),
.A2(n_741),
.B(n_545),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_747),
.A2(n_746),
.B1(n_593),
.B2(n_634),
.Y(n_748)
);


endmodule