module fake_netlist_6_3867_n_1846 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1846);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1846;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1832;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_93),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_163),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_100),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_54),
.Y(n_169)
);

BUFx10_ASAP7_75t_L g170 ( 
.A(n_117),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_83),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_54),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_39),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_146),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_142),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_154),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_127),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_33),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_35),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_24),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_123),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_133),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_121),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_33),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_62),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_92),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_69),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_126),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_106),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_143),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_118),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_101),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_109),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_76),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_72),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_113),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_61),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_2),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_152),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_42),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_51),
.Y(n_201)
);

BUFx10_ASAP7_75t_L g202 ( 
.A(n_124),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_162),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_79),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_148),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_27),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_20),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_2),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_112),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_84),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_14),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_132),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_125),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_32),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_14),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_20),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_16),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_56),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_150),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_139),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_122),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_80),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_59),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_63),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_48),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_49),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_5),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_19),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_145),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_85),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_21),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_8),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_120),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_107),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_28),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_65),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_11),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_114),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_157),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_24),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_4),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_13),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_45),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_141),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_40),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_45),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_158),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_67),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_55),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g250 ( 
.A(n_86),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_95),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_131),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_156),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_165),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_47),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_74),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_30),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_129),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_19),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_151),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_149),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_135),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_81),
.Y(n_263)
);

BUFx2_ASAP7_75t_SL g264 ( 
.A(n_1),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_17),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_42),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_164),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_153),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_137),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_90),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_6),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_71),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_136),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_160),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_111),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_25),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_105),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_4),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_48),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_35),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_9),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_13),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_22),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_88),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_68),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_60),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_36),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_51),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_9),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_31),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_108),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_116),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_66),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_94),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_17),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_30),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_144),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_89),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_70),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_78),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_26),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_52),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_140),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_31),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_82),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_87),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_29),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_38),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_34),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_91),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_15),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_57),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_32),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_138),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_53),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_15),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_41),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_115),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_10),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_6),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_37),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_102),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_16),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_50),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_56),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_130),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_43),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_77),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_147),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_104),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_40),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_27),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_245),
.B(n_256),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_198),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_271),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_271),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_271),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_271),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_271),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_282),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_282),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_203),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_206),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_207),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_282),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_282),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_267),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_282),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_184),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_184),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_217),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_217),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_225),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_205),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_318),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_225),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_243),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_240),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_277),
.B(n_0),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_208),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_310),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_243),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_194),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_250),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_240),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_200),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_201),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_226),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_250),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_211),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_214),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_256),
.B(n_0),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_235),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_215),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_195),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_237),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_216),
.Y(n_377)
);

CKINVDCx14_ASAP7_75t_R g378 ( 
.A(n_240),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_218),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_227),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_228),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_231),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_196),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_232),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_266),
.B(n_1),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_264),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_241),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_246),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_255),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_265),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_279),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_244),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_209),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_210),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_257),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_242),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_220),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_280),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_221),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_283),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_287),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_304),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_319),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_250),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_320),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_223),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_249),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_257),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_169),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_308),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_308),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_229),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_170),
.Y(n_413)
);

INVxp33_ASAP7_75t_SL g414 ( 
.A(n_169),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_346),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_348),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_364),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_335),
.B(n_336),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_346),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_348),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_333),
.B(n_204),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_364),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_337),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_338),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_339),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_334),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_409),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_340),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_392),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_369),
.Y(n_430)
);

AND3x2_ASAP7_75t_L g431 ( 
.A(n_372),
.B(n_229),
.C(n_189),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_369),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_341),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_404),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_404),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_345),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_412),
.B(n_166),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_412),
.B(n_166),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_359),
.B(n_204),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_349),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_349),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_350),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_350),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_392),
.B(n_167),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_351),
.B(n_204),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_366),
.B(n_167),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_413),
.B(n_172),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_351),
.Y(n_448)
);

INVx6_ASAP7_75t_L g449 ( 
.A(n_354),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_352),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_352),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_353),
.B(n_244),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_353),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_356),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_356),
.Y(n_455)
);

NOR2x1_ASAP7_75t_L g456 ( 
.A(n_363),
.B(n_258),
.Y(n_456)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_334),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_357),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_357),
.Y(n_459)
);

BUFx8_ASAP7_75t_L g460 ( 
.A(n_367),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_362),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_343),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_362),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_395),
.B(n_258),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_395),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_343),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_408),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_408),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_410),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_410),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_411),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_411),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_344),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_368),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_373),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_376),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_387),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_388),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_389),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_390),
.B(n_322),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_344),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_391),
.B(n_168),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_398),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_400),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_401),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_402),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_403),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_405),
.B(n_322),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_422),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_417),
.Y(n_490)
);

BUFx8_ASAP7_75t_SL g491 ( 
.A(n_426),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_479),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_421),
.B(n_360),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_422),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_479),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_417),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_429),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_479),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_422),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_456),
.B(n_360),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_422),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_430),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_421),
.B(n_370),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_445),
.B(n_386),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_429),
.Y(n_505)
);

NAND2x1p5_ASAP7_75t_L g506 ( 
.A(n_479),
.B(n_181),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_444),
.Y(n_507)
);

BUFx4f_ASAP7_75t_L g508 ( 
.A(n_475),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_479),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_423),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_430),
.Y(n_511)
);

NAND3xp33_ASAP7_75t_L g512 ( 
.A(n_439),
.B(n_213),
.C(n_193),
.Y(n_512)
);

INVx5_ASAP7_75t_L g513 ( 
.A(n_417),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_452),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_452),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_439),
.B(n_370),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_423),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_425),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_445),
.B(n_378),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_456),
.B(n_371),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_444),
.B(n_371),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_425),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_428),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_447),
.B(n_374),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_466),
.A2(n_383),
.B1(n_375),
.B2(n_406),
.Y(n_525)
);

BUFx4f_ASAP7_75t_L g526 ( 
.A(n_475),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_452),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_445),
.B(n_480),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_430),
.Y(n_529)
);

AND3x1_ASAP7_75t_L g530 ( 
.A(n_447),
.B(n_385),
.C(n_222),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_417),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_417),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_480),
.B(n_374),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_466),
.B(n_377),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_473),
.B(n_377),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_431),
.B(n_379),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_430),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_473),
.A2(n_295),
.B1(n_311),
.B2(n_332),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_480),
.B(n_379),
.Y(n_539)
);

INVx6_ASAP7_75t_L g540 ( 
.A(n_460),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_431),
.Y(n_541)
);

INVx5_ASAP7_75t_L g542 ( 
.A(n_417),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_432),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_428),
.Y(n_544)
);

BUFx10_ASAP7_75t_L g545 ( 
.A(n_449),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_452),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_427),
.Y(n_547)
);

INVx5_ASAP7_75t_L g548 ( 
.A(n_417),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_417),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_432),
.Y(n_550)
);

INVxp67_ASAP7_75t_SL g551 ( 
.A(n_417),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_432),
.Y(n_552)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_427),
.Y(n_553)
);

BUFx6f_ASAP7_75t_SL g554 ( 
.A(n_480),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_434),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_426),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_432),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_436),
.Y(n_558)
);

INVxp67_ASAP7_75t_SL g559 ( 
.A(n_434),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_480),
.B(n_488),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_446),
.B(n_414),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_418),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_418),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_416),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_452),
.B(n_380),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_452),
.B(n_380),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_464),
.B(n_381),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_436),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_480),
.A2(n_185),
.B1(n_199),
.B2(n_212),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_416),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_416),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_420),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_420),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_464),
.B(n_381),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_426),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_464),
.B(n_460),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_420),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_488),
.A2(n_185),
.B1(n_199),
.B2(n_212),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_488),
.A2(n_185),
.B1(n_199),
.B2(n_212),
.Y(n_579)
);

AND2x6_ASAP7_75t_L g580 ( 
.A(n_434),
.B(n_185),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_457),
.B(n_382),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_457),
.B(n_382),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_449),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_424),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_434),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_424),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_436),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_457),
.B(n_384),
.Y(n_588)
);

BUFx6f_ASAP7_75t_SL g589 ( 
.A(n_488),
.Y(n_589)
);

AND3x2_ASAP7_75t_L g590 ( 
.A(n_462),
.B(n_365),
.C(n_358),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_464),
.B(n_460),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_462),
.B(n_384),
.Y(n_592)
);

CKINVDCx11_ASAP7_75t_R g593 ( 
.A(n_462),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_449),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_481),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_446),
.B(n_393),
.Y(n_596)
);

BUFx8_ASAP7_75t_SL g597 ( 
.A(n_481),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_481),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_482),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_460),
.B(n_396),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_424),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_449),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_434),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_L g604 ( 
.A(n_482),
.B(n_407),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_433),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_460),
.B(n_396),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_434),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_433),
.Y(n_608)
);

BUFx10_ASAP7_75t_L g609 ( 
.A(n_449),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_460),
.B(n_407),
.Y(n_610)
);

INVx5_ASAP7_75t_L g611 ( 
.A(n_434),
.Y(n_611)
);

OR2x2_ASAP7_75t_L g612 ( 
.A(n_437),
.B(n_259),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_433),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_436),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_434),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_474),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_415),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_464),
.B(n_197),
.Y(n_618)
);

CKINVDCx6p67_ASAP7_75t_R g619 ( 
.A(n_437),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_415),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_438),
.B(n_394),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_434),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_SL g623 ( 
.A(n_449),
.B(n_361),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_415),
.Y(n_624)
);

INVx5_ASAP7_75t_L g625 ( 
.A(n_435),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_474),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_474),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_415),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_488),
.B(n_397),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_419),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_419),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_419),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_464),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_474),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_435),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_438),
.B(n_276),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_419),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_435),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_512),
.A2(n_185),
.B1(n_298),
.B2(n_254),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_L g640 ( 
.A1(n_507),
.A2(n_399),
.B1(n_449),
.B2(n_355),
.Y(n_640)
);

NOR2x2_ASAP7_75t_L g641 ( 
.A(n_530),
.B(n_385),
.Y(n_641)
);

OR2x6_ASAP7_75t_L g642 ( 
.A(n_547),
.B(n_483),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_599),
.B(n_168),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_507),
.B(n_299),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_528),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_491),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_528),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_514),
.Y(n_648)
);

OR2x2_ASAP7_75t_L g649 ( 
.A(n_547),
.B(n_483),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_584),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_514),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_514),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_515),
.Y(n_653)
);

INVxp33_ASAP7_75t_L g654 ( 
.A(n_597),
.Y(n_654)
);

NAND2x1p5_ASAP7_75t_L g655 ( 
.A(n_583),
.B(n_594),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_515),
.B(n_199),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_556),
.Y(n_657)
);

OAI22xp33_ASAP7_75t_L g658 ( 
.A1(n_516),
.A2(n_342),
.B1(n_347),
.B2(n_300),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_515),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_497),
.B(n_484),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_562),
.B(n_435),
.Y(n_661)
);

NOR3xp33_ASAP7_75t_L g662 ( 
.A(n_525),
.B(n_484),
.C(n_477),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_561),
.B(n_171),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_562),
.B(n_435),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_563),
.B(n_493),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_527),
.B(n_199),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_503),
.B(n_171),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_527),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_497),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_584),
.Y(n_670)
);

NAND2xp33_ASAP7_75t_R g671 ( 
.A(n_595),
.B(n_172),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_563),
.B(n_435),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_551),
.A2(n_230),
.B(n_219),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_521),
.B(n_435),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_586),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_618),
.B(n_435),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_560),
.B(n_435),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_527),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_546),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_560),
.B(n_475),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_546),
.B(n_212),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_504),
.B(n_475),
.Y(n_682)
);

NOR2xp67_ASAP7_75t_L g683 ( 
.A(n_553),
.B(n_477),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_559),
.B(n_475),
.Y(n_684)
);

OR2x2_ASAP7_75t_L g685 ( 
.A(n_505),
.B(n_477),
.Y(n_685)
);

NOR2xp67_ASAP7_75t_L g686 ( 
.A(n_596),
.B(n_476),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_586),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_505),
.B(n_472),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_546),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_633),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_L g691 ( 
.A1(n_619),
.A2(n_247),
.B1(n_261),
.B2(n_238),
.Y(n_691)
);

BUFx5_ASAP7_75t_L g692 ( 
.A(n_580),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_633),
.Y(n_693)
);

NOR2xp67_ASAP7_75t_SL g694 ( 
.A(n_540),
.B(n_512),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_633),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_SL g696 ( 
.A(n_623),
.B(n_595),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_621),
.B(n_174),
.Y(n_697)
);

OAI22xp5_ASAP7_75t_L g698 ( 
.A1(n_619),
.A2(n_236),
.B1(n_234),
.B2(n_233),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_510),
.B(n_475),
.Y(n_699)
);

AO22x2_ASAP7_75t_L g700 ( 
.A1(n_541),
.A2(n_270),
.B1(n_286),
.B2(n_285),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_510),
.B(n_517),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_519),
.B(n_612),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_517),
.B(n_475),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_519),
.B(n_174),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_518),
.B(n_475),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_601),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_612),
.B(n_175),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_518),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_522),
.B(n_475),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_565),
.B(n_212),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_566),
.B(n_254),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_522),
.Y(n_712)
);

NAND2x1p5_ASAP7_75t_L g713 ( 
.A(n_583),
.B(n_272),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_636),
.B(n_175),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_636),
.B(n_176),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_533),
.B(n_176),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_523),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_567),
.B(n_177),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_533),
.B(n_177),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_539),
.B(n_574),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_500),
.B(n_182),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_523),
.B(n_544),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_601),
.Y(n_723)
);

INVx8_ASAP7_75t_L g724 ( 
.A(n_554),
.Y(n_724)
);

NAND3xp33_ASAP7_75t_L g725 ( 
.A(n_604),
.B(n_281),
.C(n_278),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_569),
.A2(n_254),
.B1(n_298),
.B2(n_250),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_605),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_544),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_564),
.B(n_487),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_539),
.B(n_182),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_605),
.Y(n_731)
);

NAND2xp33_ASAP7_75t_L g732 ( 
.A(n_576),
.B(n_591),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_608),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_564),
.B(n_487),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_608),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_629),
.B(n_183),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_629),
.A2(n_291),
.B1(n_224),
.B2(n_239),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_541),
.B(n_183),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_613),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_600),
.B(n_186),
.Y(n_740)
);

NOR2x1p5_ASAP7_75t_L g741 ( 
.A(n_536),
.B(n_173),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_490),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_545),
.B(n_254),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_520),
.B(n_186),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_570),
.B(n_487),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_613),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_575),
.B(n_472),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_578),
.A2(n_254),
.B1(n_298),
.B2(n_250),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_570),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_571),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_571),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_524),
.A2(n_602),
.B1(n_594),
.B2(n_534),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_535),
.B(n_187),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_572),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_572),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_573),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_602),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_573),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_606),
.B(n_187),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_577),
.B(n_487),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_577),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_593),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_598),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_492),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_492),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_610),
.B(n_188),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_495),
.B(n_487),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_489),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_495),
.B(n_487),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_545),
.B(n_188),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_581),
.B(n_190),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_489),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_554),
.A2(n_262),
.B1(n_248),
.B2(n_251),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_582),
.B(n_190),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_498),
.B(n_487),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_545),
.B(n_191),
.Y(n_776)
);

OAI221xp5_ASAP7_75t_L g777 ( 
.A1(n_538),
.A2(n_476),
.B1(n_486),
.B2(n_485),
.C(n_478),
.Y(n_777)
);

OAI22xp33_ASAP7_75t_L g778 ( 
.A1(n_538),
.A2(n_575),
.B1(n_540),
.B2(n_598),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_498),
.B(n_487),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_494),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_509),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_509),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_490),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_494),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_588),
.B(n_476),
.Y(n_785)
);

OAI22xp5_ASAP7_75t_L g786 ( 
.A1(n_540),
.A2(n_326),
.B1(n_305),
.B2(n_273),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_496),
.B(n_487),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_554),
.A2(n_260),
.B1(n_252),
.B2(n_253),
.Y(n_788)
);

A2O1A1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_616),
.A2(n_297),
.B(n_328),
.C(n_455),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_592),
.B(n_191),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_530),
.B(n_486),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_545),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_496),
.B(n_549),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_616),
.Y(n_794)
);

OAI22xp33_ASAP7_75t_L g795 ( 
.A1(n_540),
.A2(n_506),
.B1(n_180),
.B2(n_179),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_496),
.B(n_549),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_626),
.Y(n_797)
);

NOR3xp33_ASAP7_75t_L g798 ( 
.A(n_626),
.B(n_289),
.C(n_288),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_627),
.Y(n_799)
);

BUFx2_ASAP7_75t_L g800 ( 
.A(n_590),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_627),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_609),
.B(n_506),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_634),
.B(n_192),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_634),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_496),
.B(n_455),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_499),
.Y(n_806)
);

BUFx5_ASAP7_75t_L g807 ( 
.A(n_580),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_549),
.B(n_455),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_609),
.B(n_298),
.Y(n_809)
);

NAND2xp33_ASAP7_75t_L g810 ( 
.A(n_792),
.B(n_506),
.Y(n_810)
);

NOR3xp33_ASAP7_75t_L g811 ( 
.A(n_640),
.B(n_329),
.C(n_192),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_802),
.A2(n_526),
.B(n_508),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_802),
.A2(n_526),
.B(n_508),
.Y(n_813)
);

O2A1O1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_665),
.A2(n_557),
.B(n_550),
.C(n_478),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_686),
.B(n_609),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_644),
.B(n_549),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_644),
.B(n_585),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_677),
.A2(n_526),
.B(n_508),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_682),
.A2(n_555),
.B(n_531),
.Y(n_819)
);

NOR2x1p5_ASAP7_75t_L g820 ( 
.A(n_762),
.B(n_173),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_752),
.A2(n_579),
.B1(n_589),
.B2(n_622),
.Y(n_821)
);

AND2x2_ASAP7_75t_SL g822 ( 
.A(n_696),
.B(n_298),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_642),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_650),
.Y(n_824)
);

OAI21xp5_ASAP7_75t_L g825 ( 
.A1(n_661),
.A2(n_622),
.B(n_532),
.Y(n_825)
);

AOI33xp33_ASAP7_75t_L g826 ( 
.A1(n_657),
.A2(n_451),
.A3(n_461),
.B1(n_459),
.B2(n_454),
.B3(n_440),
.Y(n_826)
);

BUFx8_ASAP7_75t_SL g827 ( 
.A(n_646),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_697),
.B(n_585),
.Y(n_828)
);

INVx4_ASAP7_75t_L g829 ( 
.A(n_724),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_669),
.B(n_609),
.Y(n_830)
);

INVx4_ASAP7_75t_L g831 ( 
.A(n_724),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_676),
.A2(n_555),
.B(n_531),
.Y(n_832)
);

AOI21x1_ASAP7_75t_L g833 ( 
.A1(n_743),
.A2(n_557),
.B(n_550),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_663),
.B(n_531),
.Y(n_834)
);

AO21x1_ASAP7_75t_L g835 ( 
.A1(n_673),
.A2(n_555),
.B(n_531),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_708),
.B(n_607),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_712),
.B(n_607),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_717),
.B(n_728),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_664),
.A2(n_622),
.B(n_532),
.Y(n_839)
);

NOR2x1_ASAP7_75t_L g840 ( 
.A(n_651),
.B(n_555),
.Y(n_840)
);

NAND2xp33_ASAP7_75t_SL g841 ( 
.A(n_741),
.B(n_589),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_674),
.A2(n_532),
.B(n_607),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_680),
.A2(n_635),
.B(n_607),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_718),
.B(n_635),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_645),
.B(n_476),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_647),
.A2(n_589),
.B1(n_635),
.B2(n_638),
.Y(n_846)
);

AND2x6_ASAP7_75t_L g847 ( 
.A(n_791),
.B(n_635),
.Y(n_847)
);

NOR2xp67_ASAP7_75t_L g848 ( 
.A(n_725),
.B(n_478),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_R g849 ( 
.A(n_763),
.B(n_329),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_672),
.A2(n_638),
.B(n_501),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_724),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_718),
.B(n_638),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_754),
.Y(n_853)
);

OAI321xp33_ASAP7_75t_L g854 ( 
.A1(n_715),
.A2(n_461),
.A3(n_459),
.B1(n_440),
.B2(n_451),
.C(n_454),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_778),
.B(n_330),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_702),
.B(n_715),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_688),
.B(n_638),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_684),
.A2(n_501),
.B(n_499),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_651),
.A2(n_615),
.B1(n_490),
.B2(n_603),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_720),
.A2(n_511),
.B(n_502),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_642),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_747),
.B(n_660),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_771),
.A2(n_529),
.B(n_502),
.C(n_537),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_701),
.B(n_490),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_722),
.B(n_490),
.Y(n_865)
);

AOI21x1_ASAP7_75t_L g866 ( 
.A1(n_743),
.A2(n_809),
.B(n_711),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_735),
.B(n_603),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_732),
.A2(n_529),
.B(n_511),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_746),
.B(n_603),
.Y(n_869)
);

NOR3xp33_ASAP7_75t_L g870 ( 
.A(n_658),
.B(n_330),
.C(n_478),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_749),
.B(n_603),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_652),
.A2(n_603),
.B1(n_615),
.B2(n_263),
.Y(n_872)
);

AOI21x1_ASAP7_75t_L g873 ( 
.A1(n_809),
.A2(n_537),
.B(n_543),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_649),
.B(n_485),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_642),
.Y(n_875)
);

O2A1O1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_777),
.A2(n_486),
.B(n_485),
.C(n_552),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_750),
.B(n_615),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_710),
.A2(n_543),
.B(n_552),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_751),
.B(n_615),
.Y(n_879)
);

O2A1O1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_667),
.A2(n_485),
.B(n_486),
.C(n_568),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_755),
.B(n_615),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_643),
.B(n_290),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_710),
.A2(n_587),
.B(n_568),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_711),
.A2(n_558),
.B(n_614),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_754),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_785),
.A2(n_284),
.B1(n_268),
.B2(n_269),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_756),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_683),
.B(n_753),
.Y(n_888)
);

INVx4_ASAP7_75t_L g889 ( 
.A(n_652),
.Y(n_889)
);

A2O1A1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_771),
.A2(n_455),
.B(n_458),
.C(n_470),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_761),
.B(n_558),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_648),
.A2(n_292),
.B1(n_274),
.B2(n_275),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_804),
.B(n_587),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_793),
.A2(n_614),
.B(n_632),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_753),
.B(n_293),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_685),
.B(n_178),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_670),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_670),
.Y(n_898)
);

NAND3xp33_ASAP7_75t_L g899 ( 
.A(n_774),
.B(n_301),
.C(n_296),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_796),
.A2(n_624),
.B(n_632),
.Y(n_900)
);

OAI21xp5_ASAP7_75t_L g901 ( 
.A1(n_794),
.A2(n_637),
.B(n_631),
.Y(n_901)
);

O2A1O1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_707),
.A2(n_459),
.B(n_440),
.C(n_451),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_675),
.B(n_617),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_805),
.A2(n_631),
.B(n_630),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_653),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_808),
.A2(n_637),
.B(n_630),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_756),
.Y(n_907)
);

OAI22xp5_ASAP7_75t_L g908 ( 
.A1(n_653),
.A2(n_294),
.B1(n_303),
.B2(n_306),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_675),
.B(n_617),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_687),
.B(n_620),
.Y(n_910)
);

BUFx8_ASAP7_75t_L g911 ( 
.A(n_800),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_774),
.B(n_302),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_L g913 ( 
.A1(n_764),
.A2(n_628),
.B(n_624),
.Y(n_913)
);

AOI21xp33_ASAP7_75t_L g914 ( 
.A1(n_790),
.A2(n_321),
.B(n_317),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_790),
.B(n_714),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_706),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_659),
.A2(n_314),
.B1(n_455),
.B2(n_458),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_668),
.A2(n_580),
.B1(n_470),
.B2(n_458),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_783),
.A2(n_625),
.B(n_611),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_758),
.Y(n_920)
);

O2A1O1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_740),
.A2(n_454),
.B(n_461),
.C(n_628),
.Y(n_921)
);

NAND2x1p5_ASAP7_75t_L g922 ( 
.A(n_757),
.B(n_513),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_783),
.A2(n_625),
.B(n_513),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_721),
.Y(n_924)
);

O2A1O1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_759),
.A2(n_620),
.B(n_458),
.C(n_470),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_699),
.A2(n_625),
.B(n_611),
.Y(n_926)
);

A2O1A1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_721),
.A2(n_458),
.B(n_470),
.C(n_453),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_706),
.B(n_470),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_678),
.A2(n_313),
.B1(n_312),
.B2(n_323),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_723),
.B(n_441),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_744),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_679),
.B(n_441),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_689),
.B(n_441),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_703),
.A2(n_625),
.B(n_611),
.Y(n_934)
);

AO21x1_ASAP7_75t_L g935 ( 
.A1(n_656),
.A2(n_453),
.B(n_471),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_723),
.B(n_727),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_727),
.Y(n_937)
);

OAI21x1_ASAP7_75t_L g938 ( 
.A1(n_787),
.A2(n_467),
.B(n_441),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_705),
.A2(n_625),
.B(n_611),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_709),
.A2(n_625),
.B(n_611),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_744),
.B(n_170),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_731),
.B(n_442),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_795),
.B(n_737),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_704),
.B(n_178),
.Y(n_944)
);

AOI22xp33_ASAP7_75t_L g945 ( 
.A1(n_690),
.A2(n_250),
.B1(n_580),
.B2(n_443),
.Y(n_945)
);

INVxp67_ASAP7_75t_L g946 ( 
.A(n_671),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_731),
.B(n_442),
.Y(n_947)
);

BUFx4f_ASAP7_75t_L g948 ( 
.A(n_713),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_738),
.B(n_307),
.Y(n_949)
);

NOR3xp33_ASAP7_75t_L g950 ( 
.A(n_736),
.B(n_309),
.C(n_316),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_733),
.B(n_442),
.Y(n_951)
);

AOI22xp33_ASAP7_75t_L g952 ( 
.A1(n_693),
.A2(n_250),
.B1(n_580),
.B2(n_443),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_729),
.A2(n_611),
.B(n_513),
.Y(n_953)
);

AND2x2_ASAP7_75t_SL g954 ( 
.A(n_726),
.B(n_170),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_716),
.B(n_179),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_758),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_719),
.B(n_315),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_730),
.B(n_766),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_695),
.B(n_442),
.Y(n_959)
);

NAND2xp33_ASAP7_75t_L g960 ( 
.A(n_692),
.B(n_250),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_733),
.B(n_448),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_757),
.A2(n_180),
.B1(n_324),
.B2(n_325),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_783),
.Y(n_963)
);

INVx1_ASAP7_75t_SL g964 ( 
.A(n_641),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_734),
.A2(n_513),
.B(n_548),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_662),
.B(n_202),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_739),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_739),
.B(n_448),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_768),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_765),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_655),
.A2(n_325),
.B1(n_327),
.B2(n_331),
.Y(n_971)
);

A2O1A1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_803),
.A2(n_782),
.B(n_781),
.C(n_801),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_L g973 ( 
.A1(n_745),
.A2(n_580),
.B(n_548),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_797),
.B(n_799),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_768),
.B(n_772),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_691),
.B(n_698),
.Y(n_976)
);

INVx4_ASAP7_75t_L g977 ( 
.A(n_783),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_772),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_780),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_784),
.B(n_450),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_784),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_773),
.B(n_324),
.Y(n_982)
);

INVxp67_ASAP7_75t_L g983 ( 
.A(n_671),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_806),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_798),
.B(n_202),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_760),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_655),
.B(n_742),
.Y(n_987)
);

OR2x2_ASAP7_75t_L g988 ( 
.A(n_654),
.B(n_327),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_742),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_R g990 ( 
.A(n_767),
.B(n_331),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_769),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_656),
.A2(n_513),
.B(n_548),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_666),
.A2(n_513),
.B(n_548),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_713),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_666),
.A2(n_681),
.B1(n_694),
.B2(n_788),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_815),
.A2(n_770),
.B(n_776),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_827),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_912),
.B(n_946),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_824),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_864),
.A2(n_681),
.B(n_786),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_851),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_856),
.B(n_700),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_897),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_963),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_823),
.Y(n_1005)
);

BUFx2_ASAP7_75t_L g1006 ( 
.A(n_861),
.Y(n_1006)
);

INVxp67_ASAP7_75t_L g1007 ( 
.A(n_875),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_983),
.B(n_924),
.Y(n_1008)
);

OR2x2_ASAP7_75t_L g1009 ( 
.A(n_862),
.B(n_775),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_931),
.B(n_692),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_898),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_896),
.B(n_700),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_865),
.A2(n_748),
.B(n_726),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_812),
.A2(n_748),
.B(n_779),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_976),
.A2(n_639),
.B(n_789),
.C(n_453),
.Y(n_1015)
);

NAND2xp33_ASAP7_75t_SL g1016 ( 
.A(n_851),
.B(n_639),
.Y(n_1016)
);

A2O1A1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_958),
.A2(n_467),
.B(n_465),
.C(n_450),
.Y(n_1017)
);

CKINVDCx11_ASAP7_75t_R g1018 ( 
.A(n_964),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_914),
.B(n_202),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_853),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_R g1021 ( 
.A(n_841),
.B(n_807),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_982),
.B(n_807),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_882),
.A2(n_468),
.B(n_450),
.C(n_453),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_916),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_874),
.B(n_955),
.Y(n_1025)
);

O2A1O1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_943),
.A2(n_471),
.B(n_469),
.C(n_468),
.Y(n_1026)
);

NOR2x1_ASAP7_75t_R g1027 ( 
.A(n_851),
.B(n_807),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_885),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_944),
.B(n_988),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_954),
.A2(n_469),
.B1(n_463),
.B2(n_465),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_937),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_888),
.B(n_807),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_812),
.A2(n_542),
.B(n_548),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_957),
.B(n_807),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_963),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_838),
.B(n_807),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_949),
.A2(n_468),
.B(n_463),
.C(n_465),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_991),
.B(n_692),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_822),
.B(n_692),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_887),
.Y(n_1040)
);

NOR3xp33_ASAP7_75t_SL g1041 ( 
.A(n_971),
.B(n_3),
.C(n_5),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_813),
.A2(n_542),
.B(n_548),
.Y(n_1042)
);

O2A1O1Ixp5_ASAP7_75t_SL g1043 ( 
.A1(n_941),
.A2(n_580),
.B(n_7),
.C(n_8),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_907),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_899),
.B(n_692),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_813),
.A2(n_542),
.B(n_692),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_920),
.Y(n_1047)
);

O2A1O1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_855),
.A2(n_471),
.B(n_469),
.C(n_468),
.Y(n_1048)
);

NAND2xp33_ASAP7_75t_L g1049 ( 
.A(n_994),
.B(n_443),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_895),
.B(n_962),
.Y(n_1050)
);

NAND3xp33_ASAP7_75t_SL g1051 ( 
.A(n_811),
.B(n_471),
.C(n_469),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_870),
.A2(n_467),
.B(n_465),
.C(n_463),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_948),
.B(n_467),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_995),
.A2(n_463),
.B(n_443),
.C(n_542),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_970),
.B(n_443),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_844),
.A2(n_542),
.B(n_443),
.Y(n_1056)
);

OR2x4_ASAP7_75t_L g1057 ( 
.A(n_994),
.B(n_443),
.Y(n_1057)
);

AO21x1_ASAP7_75t_L g1058 ( 
.A1(n_828),
.A2(n_3),
.B(n_7),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_956),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_852),
.A2(n_542),
.B(n_443),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_963),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_843),
.A2(n_443),
.B(n_161),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_966),
.B(n_10),
.Y(n_1063)
);

NAND2x1p5_ASAP7_75t_L g1064 ( 
.A(n_905),
.B(n_159),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_911),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_986),
.B(n_11),
.Y(n_1066)
);

OAI22x1_ASAP7_75t_L g1067 ( 
.A1(n_985),
.A2(n_12),
.B1(n_18),
.B2(n_21),
.Y(n_1067)
);

INVx1_ASAP7_75t_SL g1068 ( 
.A(n_990),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_845),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_889),
.B(n_12),
.Y(n_1070)
);

INVx4_ASAP7_75t_L g1071 ( 
.A(n_829),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_829),
.B(n_155),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_905),
.A2(n_134),
.B1(n_128),
.B2(n_119),
.Y(n_1073)
);

INVx2_ASAP7_75t_SL g1074 ( 
.A(n_849),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_967),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_948),
.B(n_110),
.Y(n_1076)
);

NAND2x1p5_ASAP7_75t_L g1077 ( 
.A(n_831),
.B(n_103),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_845),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_857),
.B(n_893),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_972),
.A2(n_889),
.B1(n_817),
.B2(n_816),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_832),
.A2(n_99),
.B(n_98),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_974),
.B(n_22),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_826),
.B(n_23),
.Y(n_1083)
);

O2A1O1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_950),
.A2(n_23),
.B(n_25),
.C(n_26),
.Y(n_1084)
);

NAND3xp33_ASAP7_75t_SL g1085 ( 
.A(n_886),
.B(n_28),
.C(n_29),
.Y(n_1085)
);

O2A1O1Ixp5_ASAP7_75t_L g1086 ( 
.A1(n_835),
.A2(n_97),
.B(n_96),
.C(n_75),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_936),
.B(n_34),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_978),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_977),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_994),
.B(n_73),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_892),
.B(n_64),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_819),
.A2(n_58),
.B(n_38),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_834),
.B(n_37),
.Y(n_1093)
);

INVx6_ASAP7_75t_L g1094 ( 
.A(n_911),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_854),
.B(n_39),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_977),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_821),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_831),
.B(n_44),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_819),
.A2(n_818),
.B(n_839),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_932),
.B(n_46),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_SL g1101 ( 
.A(n_847),
.Y(n_1101)
);

OR2x6_ASAP7_75t_L g1102 ( 
.A(n_820),
.B(n_46),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_932),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_933),
.B(n_47),
.Y(n_1104)
);

NOR3xp33_ASAP7_75t_L g1105 ( 
.A(n_929),
.B(n_49),
.C(n_50),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_933),
.B(n_52),
.Y(n_1106)
);

O2A1O1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_902),
.A2(n_890),
.B(n_810),
.C(n_927),
.Y(n_1107)
);

CKINVDCx8_ASAP7_75t_R g1108 ( 
.A(n_847),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_969),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_908),
.B(n_53),
.Y(n_1110)
);

OR2x6_ASAP7_75t_L g1111 ( 
.A(n_922),
.B(n_55),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_818),
.A2(n_57),
.B(n_825),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_959),
.B(n_848),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_959),
.B(n_989),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_867),
.A2(n_869),
.B1(n_877),
.B2(n_879),
.Y(n_1115)
);

AOI21xp33_ASAP7_75t_L g1116 ( 
.A1(n_836),
.A2(n_837),
.B(n_891),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_880),
.A2(n_925),
.B(n_921),
.C(n_860),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_979),
.B(n_981),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_987),
.A2(n_859),
.B(n_842),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_984),
.B(n_847),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_863),
.A2(n_917),
.B(n_846),
.C(n_814),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_847),
.B(n_975),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_871),
.B(n_881),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_847),
.B(n_910),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_840),
.A2(n_922),
.B1(n_909),
.B2(n_903),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_843),
.B(n_942),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_842),
.A2(n_960),
.B(n_830),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_860),
.A2(n_876),
.B(n_884),
.C(n_883),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_SL g1129 ( 
.A1(n_918),
.A2(n_952),
.B1(n_945),
.B2(n_928),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_SL g1130 ( 
.A1(n_973),
.A2(n_913),
.B(n_901),
.C(n_868),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_872),
.A2(n_930),
.B(n_968),
.C(n_951),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_947),
.Y(n_1132)
);

INVx1_ASAP7_75t_SL g1133 ( 
.A(n_961),
.Y(n_1133)
);

OR2x6_ASAP7_75t_L g1134 ( 
.A(n_992),
.B(n_993),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_980),
.Y(n_1135)
);

INVx5_ASAP7_75t_L g1136 ( 
.A(n_935),
.Y(n_1136)
);

NOR2xp67_ASAP7_75t_SL g1137 ( 
.A(n_992),
.B(n_993),
.Y(n_1137)
);

AOI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_883),
.A2(n_884),
.B1(n_850),
.B2(n_894),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_850),
.B(n_858),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_894),
.A2(n_900),
.B(n_904),
.C(n_878),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_858),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_904),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_866),
.A2(n_868),
.B1(n_833),
.B2(n_900),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_906),
.B(n_965),
.Y(n_1144)
);

NOR3xp33_ASAP7_75t_SL g1145 ( 
.A(n_878),
.B(n_965),
.C(n_953),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_953),
.B(n_934),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_938),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_998),
.B(n_926),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1025),
.B(n_926),
.Y(n_1149)
);

AOI21x1_ASAP7_75t_L g1150 ( 
.A1(n_1137),
.A2(n_1144),
.B(n_1146),
.Y(n_1150)
);

HB1xp67_ASAP7_75t_L g1151 ( 
.A(n_1006),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_1005),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1112),
.A2(n_934),
.B(n_939),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1088),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1046),
.A2(n_873),
.B(n_939),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1033),
.A2(n_940),
.B(n_919),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_1001),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_1050),
.A2(n_923),
.B(n_940),
.C(n_1019),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1034),
.A2(n_1099),
.B(n_1130),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_1068),
.B(n_1029),
.Y(n_1160)
);

AO31x2_ASAP7_75t_L g1161 ( 
.A1(n_1143),
.A2(n_1054),
.A3(n_1140),
.B(n_1147),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1022),
.A2(n_1127),
.B(n_1139),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1126),
.A2(n_1000),
.B(n_1080),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_1008),
.B(n_1068),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1119),
.A2(n_1013),
.B(n_1123),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1014),
.A2(n_1131),
.B(n_1116),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1062),
.A2(n_1079),
.B(n_996),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1042),
.A2(n_1056),
.B(n_1060),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1009),
.B(n_1133),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_SL g1170 ( 
.A1(n_1095),
.A2(n_1091),
.B(n_1076),
.C(n_1093),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1133),
.B(n_1012),
.Y(n_1171)
);

INVx5_ASAP7_75t_L g1172 ( 
.A(n_1001),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1138),
.A2(n_1141),
.B(n_1142),
.Y(n_1173)
);

AO32x2_ASAP7_75t_L g1174 ( 
.A1(n_1097),
.A2(n_1030),
.A3(n_1115),
.B1(n_1125),
.B2(n_1129),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1062),
.A2(n_1128),
.B(n_1117),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1036),
.A2(n_1107),
.B(n_1039),
.Y(n_1176)
);

BUFx3_ASAP7_75t_L g1177 ( 
.A(n_1001),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_1074),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1015),
.A2(n_1121),
.B(n_1052),
.Y(n_1179)
);

AO31x2_ASAP7_75t_L g1180 ( 
.A1(n_1030),
.A2(n_1058),
.A3(n_1017),
.B(n_1037),
.Y(n_1180)
);

INVx3_ASAP7_75t_L g1181 ( 
.A(n_1108),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1049),
.A2(n_1038),
.B(n_1122),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_1069),
.B(n_1078),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_999),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1124),
.A2(n_1045),
.B(n_1032),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1134),
.A2(n_1016),
.B(n_1027),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1101),
.A2(n_1057),
.B1(n_1110),
.B2(n_1083),
.Y(n_1187)
);

NAND2x1p5_ASAP7_75t_L g1188 ( 
.A(n_1071),
.B(n_1089),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1134),
.A2(n_1113),
.B(n_1081),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1135),
.B(n_1132),
.Y(n_1190)
);

AOI221xp5_ASAP7_75t_L g1191 ( 
.A1(n_1063),
.A2(n_1085),
.B1(n_1105),
.B2(n_1084),
.C(n_1067),
.Y(n_1191)
);

AOI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1134),
.A2(n_1087),
.B(n_1053),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_997),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1026),
.A2(n_1055),
.B(n_1120),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_1101),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1007),
.B(n_1041),
.Y(n_1196)
);

AO31x2_ASAP7_75t_L g1197 ( 
.A1(n_1023),
.A2(n_1092),
.A3(n_1118),
.B(n_1066),
.Y(n_1197)
);

NAND2xp33_ASAP7_75t_R g1198 ( 
.A(n_1021),
.B(n_1145),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1103),
.B(n_1104),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1103),
.A2(n_1135),
.B1(n_1003),
.B2(n_1011),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1082),
.B(n_1100),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1109),
.Y(n_1202)
);

INVx3_ASAP7_75t_SL g1203 ( 
.A(n_1094),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1024),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_SL g1205 ( 
.A1(n_1090),
.A2(n_1010),
.B(n_1098),
.C(n_1106),
.Y(n_1205)
);

NOR4xp25_ASAP7_75t_L g1206 ( 
.A(n_1051),
.B(n_1070),
.C(n_1031),
.D(n_1048),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1102),
.B(n_1020),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1114),
.A2(n_1136),
.B(n_1096),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1040),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1044),
.B(n_1075),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1086),
.A2(n_1064),
.B(n_1047),
.Y(n_1211)
);

OA21x2_ASAP7_75t_L g1212 ( 
.A1(n_1059),
.A2(n_1028),
.B(n_1136),
.Y(n_1212)
);

AOI221x1_ASAP7_75t_L g1213 ( 
.A1(n_1073),
.A2(n_1043),
.B1(n_1072),
.B2(n_1004),
.C(n_1089),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_1018),
.Y(n_1214)
);

CKINVDCx8_ASAP7_75t_R g1215 ( 
.A(n_1035),
.Y(n_1215)
);

INVx1_ASAP7_75t_SL g1216 ( 
.A(n_1035),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1072),
.B(n_1004),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1057),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1136),
.A2(n_1111),
.B(n_1077),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1035),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1102),
.B(n_1111),
.Y(n_1221)
);

AOI21xp33_ASAP7_75t_L g1222 ( 
.A1(n_1111),
.A2(n_1102),
.B(n_1061),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1061),
.A2(n_1094),
.B(n_1065),
.Y(n_1223)
);

AOI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1061),
.A2(n_915),
.B1(n_1019),
.B2(n_912),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1046),
.A2(n_938),
.B(n_1033),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1022),
.A2(n_954),
.B1(n_822),
.B2(n_665),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1034),
.A2(n_802),
.B(n_732),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1034),
.A2(n_802),
.B(n_732),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_1069),
.B(n_829),
.Y(n_1229)
);

O2A1O1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1019),
.A2(n_912),
.B(n_915),
.C(n_697),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1034),
.A2(n_802),
.B(n_732),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1046),
.A2(n_938),
.B(n_1033),
.Y(n_1232)
);

A2O1A1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1050),
.A2(n_915),
.B(n_856),
.C(n_912),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1019),
.A2(n_915),
.B1(n_912),
.B2(n_976),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_998),
.B(n_862),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1034),
.A2(n_802),
.B(n_732),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1108),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1088),
.Y(n_1238)
);

NAND3x1_ASAP7_75t_L g1239 ( 
.A(n_1019),
.B(n_538),
.C(n_912),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1088),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1143),
.A2(n_1054),
.A3(n_835),
.B(n_1099),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1046),
.A2(n_938),
.B(n_1033),
.Y(n_1242)
);

O2A1O1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1019),
.A2(n_912),
.B(n_915),
.C(n_697),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_998),
.B(n_342),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1022),
.A2(n_915),
.B1(n_856),
.B2(n_912),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1034),
.A2(n_802),
.B(n_732),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_998),
.B(n_862),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_998),
.B(n_862),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1019),
.A2(n_915),
.B1(n_912),
.B2(n_976),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_998),
.B(n_342),
.Y(n_1250)
);

AO31x2_ASAP7_75t_L g1251 ( 
.A1(n_1143),
.A2(n_1054),
.A3(n_835),
.B(n_1099),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1088),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_998),
.B(n_862),
.Y(n_1253)
);

AO31x2_ASAP7_75t_L g1254 ( 
.A1(n_1143),
.A2(n_1054),
.A3(n_835),
.B(n_1099),
.Y(n_1254)
);

AOI221xp5_ASAP7_75t_L g1255 ( 
.A1(n_1019),
.A2(n_658),
.B1(n_914),
.B2(n_530),
.C(n_915),
.Y(n_1255)
);

A2O1A1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1050),
.A2(n_915),
.B(n_856),
.C(n_912),
.Y(n_1256)
);

NOR2xp67_ASAP7_75t_L g1257 ( 
.A(n_996),
.B(n_507),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1034),
.A2(n_802),
.B(n_732),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1046),
.A2(n_938),
.B(n_1033),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_997),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1034),
.A2(n_802),
.B(n_732),
.Y(n_1261)
);

BUFx12f_ASAP7_75t_L g1262 ( 
.A(n_1018),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1005),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1046),
.A2(n_938),
.B(n_1033),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1050),
.A2(n_915),
.B(n_856),
.C(n_912),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1046),
.A2(n_938),
.B(n_1033),
.Y(n_1266)
);

AO31x2_ASAP7_75t_L g1267 ( 
.A1(n_1143),
.A2(n_1054),
.A3(n_835),
.B(n_1099),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1034),
.A2(n_802),
.B(n_732),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1034),
.A2(n_802),
.B(n_732),
.Y(n_1269)
);

AOI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1019),
.A2(n_915),
.B1(n_912),
.B2(n_976),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1088),
.Y(n_1271)
);

NOR4xp25_ASAP7_75t_L g1272 ( 
.A(n_1084),
.B(n_1085),
.C(n_1097),
.D(n_1019),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1034),
.A2(n_802),
.B(n_732),
.Y(n_1273)
);

O2A1O1Ixp33_ASAP7_75t_SL g1274 ( 
.A1(n_1095),
.A2(n_943),
.B(n_1091),
.C(n_1076),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1034),
.A2(n_802),
.B(n_732),
.Y(n_1275)
);

O2A1O1Ixp33_ASAP7_75t_SL g1276 ( 
.A1(n_1095),
.A2(n_943),
.B(n_1091),
.C(n_1076),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1088),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_997),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_998),
.B(n_696),
.Y(n_1279)
);

NAND3xp33_ASAP7_75t_L g1280 ( 
.A(n_1019),
.B(n_912),
.C(n_697),
.Y(n_1280)
);

AOI221xp5_ASAP7_75t_SL g1281 ( 
.A1(n_1097),
.A2(n_1083),
.B1(n_1110),
.B2(n_1095),
.C(n_1002),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1034),
.A2(n_802),
.B(n_732),
.Y(n_1282)
);

A2O1A1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1050),
.A2(n_915),
.B(n_856),
.C(n_912),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_1108),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1034),
.A2(n_802),
.B(n_732),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1005),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1046),
.A2(n_938),
.B(n_1033),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1046),
.A2(n_938),
.B(n_1033),
.Y(n_1288)
);

AOI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1137),
.A2(n_1144),
.B(n_1146),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1112),
.A2(n_1014),
.B(n_1062),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1109),
.Y(n_1291)
);

INVx5_ASAP7_75t_L g1292 ( 
.A(n_1001),
.Y(n_1292)
);

AOI221x1_ASAP7_75t_L g1293 ( 
.A1(n_1019),
.A2(n_1112),
.B1(n_912),
.B2(n_1105),
.C(n_1099),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_1069),
.B(n_829),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1034),
.A2(n_802),
.B(n_732),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1034),
.A2(n_802),
.B(n_732),
.Y(n_1296)
);

O2A1O1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1019),
.A2(n_912),
.B(n_915),
.C(n_697),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1088),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1034),
.A2(n_802),
.B(n_732),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_SL g1300 ( 
.A1(n_1107),
.A2(n_1083),
.B(n_1058),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1034),
.A2(n_802),
.B(n_732),
.Y(n_1301)
);

O2A1O1Ixp5_ASAP7_75t_SL g1302 ( 
.A1(n_1146),
.A2(n_941),
.B(n_1144),
.C(n_966),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_1172),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1260),
.Y(n_1304)
);

OAI22xp33_ASAP7_75t_SL g1305 ( 
.A1(n_1234),
.A2(n_1249),
.B1(n_1270),
.B2(n_1245),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1234),
.A2(n_1249),
.B1(n_1270),
.B2(n_1255),
.Y(n_1306)
);

AOI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1239),
.A2(n_1280),
.B1(n_1250),
.B2(n_1244),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1280),
.A2(n_1191),
.B1(n_1226),
.B2(n_1201),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1184),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1226),
.A2(n_1175),
.B1(n_1224),
.B2(n_1279),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_1193),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1278),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_1262),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1175),
.A2(n_1224),
.B1(n_1300),
.B2(n_1253),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1152),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1204),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1235),
.B(n_1247),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1248),
.A2(n_1290),
.B1(n_1179),
.B2(n_1196),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_SL g1319 ( 
.A1(n_1230),
.A2(n_1297),
.B(n_1243),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1151),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1202),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1290),
.A2(n_1179),
.B1(n_1187),
.B2(n_1169),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1291),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1238),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1240),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_SL g1326 ( 
.A1(n_1221),
.A2(n_1233),
.B1(n_1265),
.B2(n_1256),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1286),
.Y(n_1327)
);

INVx1_ASAP7_75t_SL g1328 ( 
.A(n_1160),
.Y(n_1328)
);

OAI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1171),
.A2(n_1293),
.B1(n_1190),
.B2(n_1298),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1252),
.Y(n_1330)
);

OAI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1271),
.A2(n_1277),
.B1(n_1187),
.B2(n_1209),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1210),
.Y(n_1332)
);

BUFx2_ASAP7_75t_SL g1333 ( 
.A(n_1292),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1283),
.B(n_1164),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1167),
.A2(n_1149),
.B1(n_1199),
.B2(n_1207),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1218),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1181),
.A2(n_1284),
.B1(n_1237),
.B2(n_1217),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_1215),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1183),
.B(n_1272),
.Y(n_1339)
);

INVx4_ASAP7_75t_L g1340 ( 
.A(n_1203),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1148),
.A2(n_1163),
.B1(n_1176),
.B2(n_1166),
.Y(n_1341)
);

BUFx8_ASAP7_75t_L g1342 ( 
.A(n_1178),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1200),
.A2(n_1165),
.B1(n_1222),
.B2(n_1272),
.Y(n_1343)
);

CKINVDCx11_ASAP7_75t_R g1344 ( 
.A(n_1157),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_SL g1345 ( 
.A1(n_1219),
.A2(n_1186),
.B1(n_1195),
.B2(n_1237),
.Y(n_1345)
);

BUFx3_ASAP7_75t_L g1346 ( 
.A(n_1263),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_SL g1347 ( 
.A1(n_1195),
.A2(n_1284),
.B1(n_1181),
.B2(n_1162),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1212),
.Y(n_1348)
);

CKINVDCx6p67_ASAP7_75t_R g1349 ( 
.A(n_1177),
.Y(n_1349)
);

BUFx8_ASAP7_75t_SL g1350 ( 
.A(n_1214),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1183),
.A2(n_1158),
.B1(n_1229),
.B2(n_1294),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1159),
.A2(n_1185),
.B1(n_1257),
.B2(n_1173),
.Y(n_1352)
);

INVx1_ASAP7_75t_SL g1353 ( 
.A(n_1216),
.Y(n_1353)
);

BUFx12f_ASAP7_75t_L g1354 ( 
.A(n_1229),
.Y(n_1354)
);

BUFx12f_ASAP7_75t_L g1355 ( 
.A(n_1294),
.Y(n_1355)
);

CKINVDCx11_ASAP7_75t_R g1356 ( 
.A(n_1216),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1220),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1257),
.A2(n_1189),
.B1(n_1281),
.B2(n_1273),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_1208),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1281),
.A2(n_1269),
.B1(n_1282),
.B2(n_1236),
.Y(n_1360)
);

BUFx6f_ASAP7_75t_L g1361 ( 
.A(n_1223),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_SL g1362 ( 
.A1(n_1227),
.A2(n_1246),
.B(n_1275),
.Y(n_1362)
);

INVx1_ASAP7_75t_SL g1363 ( 
.A(n_1188),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1228),
.A2(n_1285),
.B1(n_1261),
.B2(n_1301),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1205),
.B(n_1274),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1276),
.B(n_1170),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1231),
.A2(n_1268),
.B1(n_1258),
.B2(n_1299),
.Y(n_1367)
);

OAI21xp33_ASAP7_75t_L g1368 ( 
.A1(n_1206),
.A2(n_1302),
.B(n_1192),
.Y(n_1368)
);

INVx3_ASAP7_75t_L g1369 ( 
.A(n_1150),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_1182),
.Y(n_1370)
);

OAI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1198),
.A2(n_1213),
.B1(n_1295),
.B2(n_1296),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1289),
.Y(n_1372)
);

AOI21xp33_ASAP7_75t_L g1373 ( 
.A1(n_1153),
.A2(n_1194),
.B(n_1211),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_SL g1374 ( 
.A1(n_1206),
.A2(n_1153),
.B1(n_1174),
.B2(n_1197),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1161),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1168),
.A2(n_1156),
.B1(n_1155),
.B2(n_1287),
.Y(n_1376)
);

BUFx8_ASAP7_75t_L g1377 ( 
.A(n_1174),
.Y(n_1377)
);

BUFx12f_ASAP7_75t_L g1378 ( 
.A(n_1197),
.Y(n_1378)
);

BUFx12f_ASAP7_75t_L g1379 ( 
.A(n_1197),
.Y(n_1379)
);

INVx5_ASAP7_75t_L g1380 ( 
.A(n_1241),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1174),
.A2(n_1288),
.B1(n_1225),
.B2(n_1232),
.Y(n_1381)
);

CKINVDCx20_ASAP7_75t_R g1382 ( 
.A(n_1241),
.Y(n_1382)
);

CKINVDCx11_ASAP7_75t_R g1383 ( 
.A(n_1180),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1180),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1242),
.A2(n_1259),
.B1(n_1264),
.B2(n_1266),
.Y(n_1385)
);

AOI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1180),
.A2(n_1251),
.B1(n_1254),
.B2(n_1267),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1251),
.B(n_1254),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1254),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_SL g1389 ( 
.A1(n_1267),
.A2(n_1245),
.B1(n_696),
.B2(n_1280),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1154),
.Y(n_1390)
);

OAI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1234),
.A2(n_1249),
.B1(n_1270),
.B2(n_1245),
.Y(n_1391)
);

INVx2_ASAP7_75t_SL g1392 ( 
.A(n_1152),
.Y(n_1392)
);

BUFx10_ASAP7_75t_L g1393 ( 
.A(n_1214),
.Y(n_1393)
);

CKINVDCx11_ASAP7_75t_R g1394 ( 
.A(n_1262),
.Y(n_1394)
);

BUFx8_ASAP7_75t_L g1395 ( 
.A(n_1262),
.Y(n_1395)
);

BUFx10_ASAP7_75t_L g1396 ( 
.A(n_1214),
.Y(n_1396)
);

INVx1_ASAP7_75t_SL g1397 ( 
.A(n_1151),
.Y(n_1397)
);

OAI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1234),
.A2(n_1249),
.B1(n_1270),
.B2(n_1245),
.Y(n_1398)
);

OAI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1234),
.A2(n_1249),
.B1(n_1270),
.B2(n_1245),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1154),
.Y(n_1400)
);

BUFx8_ASAP7_75t_L g1401 ( 
.A(n_1262),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1154),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1234),
.A2(n_1270),
.B1(n_1249),
.B2(n_1255),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1234),
.A2(n_1249),
.B1(n_1270),
.B2(n_1256),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1260),
.Y(n_1405)
);

BUFx10_ASAP7_75t_L g1406 ( 
.A(n_1214),
.Y(n_1406)
);

INVx2_ASAP7_75t_SL g1407 ( 
.A(n_1152),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_1260),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1154),
.Y(n_1409)
);

INVx1_ASAP7_75t_SL g1410 ( 
.A(n_1151),
.Y(n_1410)
);

INVx6_ASAP7_75t_L g1411 ( 
.A(n_1172),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1202),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1154),
.Y(n_1413)
);

CKINVDCx8_ASAP7_75t_R g1414 ( 
.A(n_1214),
.Y(n_1414)
);

CKINVDCx6p67_ASAP7_75t_R g1415 ( 
.A(n_1262),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1154),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_1260),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1154),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1234),
.A2(n_1270),
.B1(n_1249),
.B2(n_1255),
.Y(n_1419)
);

CKINVDCx11_ASAP7_75t_R g1420 ( 
.A(n_1262),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1234),
.A2(n_1270),
.B1(n_1249),
.B2(n_1255),
.Y(n_1421)
);

BUFx8_ASAP7_75t_L g1422 ( 
.A(n_1262),
.Y(n_1422)
);

BUFx2_ASAP7_75t_SL g1423 ( 
.A(n_1172),
.Y(n_1423)
);

BUFx10_ASAP7_75t_L g1424 ( 
.A(n_1214),
.Y(n_1424)
);

INVx5_ASAP7_75t_L g1425 ( 
.A(n_1172),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1234),
.B(n_1249),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1154),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1234),
.A2(n_1270),
.B1(n_1249),
.B2(n_1255),
.Y(n_1428)
);

BUFx3_ASAP7_75t_L g1429 ( 
.A(n_1152),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_SL g1430 ( 
.A1(n_1245),
.A2(n_696),
.B1(n_1280),
.B2(n_954),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1385),
.A2(n_1376),
.B(n_1367),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1320),
.Y(n_1432)
);

INVx3_ASAP7_75t_L g1433 ( 
.A(n_1378),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1397),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_1361),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1348),
.Y(n_1436)
);

OR2x6_ASAP7_75t_L g1437 ( 
.A(n_1379),
.B(n_1362),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1306),
.A2(n_1403),
.B1(n_1428),
.B2(n_1419),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1388),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1382),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1385),
.A2(n_1364),
.B(n_1381),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1339),
.B(n_1426),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1381),
.A2(n_1352),
.B(n_1358),
.Y(n_1443)
);

BUFx3_ASAP7_75t_L g1444 ( 
.A(n_1359),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1384),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1352),
.A2(n_1358),
.B(n_1360),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1317),
.B(n_1334),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1375),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1372),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1410),
.Y(n_1450)
);

AO21x2_ASAP7_75t_L g1451 ( 
.A1(n_1371),
.A2(n_1373),
.B(n_1391),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1387),
.Y(n_1452)
);

INVx4_ASAP7_75t_L g1453 ( 
.A(n_1425),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1318),
.B(n_1332),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1374),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1360),
.A2(n_1341),
.B(n_1369),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1341),
.A2(n_1366),
.B(n_1365),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1386),
.A2(n_1343),
.B(n_1322),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1328),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1318),
.B(n_1322),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1389),
.B(n_1310),
.Y(n_1461)
);

INVxp67_ASAP7_75t_L g1462 ( 
.A(n_1346),
.Y(n_1462)
);

AO31x2_ASAP7_75t_L g1463 ( 
.A1(n_1404),
.A2(n_1371),
.A3(n_1368),
.B(n_1351),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1380),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1380),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1380),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1335),
.B(n_1324),
.Y(n_1467)
);

OA21x2_ASAP7_75t_L g1468 ( 
.A1(n_1319),
.A2(n_1343),
.B(n_1310),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1335),
.A2(n_1314),
.B(n_1409),
.Y(n_1469)
);

AOI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1391),
.A2(n_1398),
.B(n_1399),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1306),
.A2(n_1403),
.B1(n_1428),
.B2(n_1419),
.Y(n_1471)
);

INVx1_ASAP7_75t_SL g1472 ( 
.A(n_1356),
.Y(n_1472)
);

AOI221xp5_ASAP7_75t_L g1473 ( 
.A1(n_1398),
.A2(n_1399),
.B1(n_1305),
.B2(n_1308),
.C(n_1421),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1421),
.A2(n_1430),
.B1(n_1308),
.B2(n_1307),
.Y(n_1474)
);

NAND2x1p5_ASAP7_75t_L g1475 ( 
.A(n_1370),
.B(n_1425),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1309),
.Y(n_1476)
);

CKINVDCx11_ASAP7_75t_R g1477 ( 
.A(n_1414),
.Y(n_1477)
);

OA21x2_ASAP7_75t_L g1478 ( 
.A1(n_1314),
.A2(n_1416),
.B(n_1390),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1389),
.B(n_1326),
.Y(n_1479)
);

OAI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1430),
.A2(n_1326),
.B1(n_1347),
.B2(n_1345),
.Y(n_1480)
);

OR2x6_ASAP7_75t_L g1481 ( 
.A(n_1333),
.B(n_1423),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1383),
.B(n_1325),
.Y(n_1482)
);

OA21x2_ASAP7_75t_L g1483 ( 
.A1(n_1316),
.A2(n_1400),
.B(n_1418),
.Y(n_1483)
);

INVx3_ASAP7_75t_L g1484 ( 
.A(n_1377),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1329),
.B(n_1412),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1329),
.B(n_1321),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1425),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1330),
.B(n_1402),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1413),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_1377),
.Y(n_1490)
);

INVx2_ASAP7_75t_SL g1491 ( 
.A(n_1411),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1427),
.A2(n_1337),
.B(n_1336),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1323),
.Y(n_1493)
);

INVxp67_ASAP7_75t_SL g1494 ( 
.A(n_1357),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1331),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1353),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_1354),
.Y(n_1497)
);

OA21x2_ASAP7_75t_L g1498 ( 
.A1(n_1331),
.A2(n_1347),
.B(n_1345),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1355),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1411),
.Y(n_1500)
);

BUFx6f_ASAP7_75t_L g1501 ( 
.A(n_1303),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_1350),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1363),
.B(n_1340),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1349),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1392),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1407),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_SL g1507 ( 
.A1(n_1340),
.A2(n_1342),
.B(n_1344),
.Y(n_1507)
);

INVx3_ASAP7_75t_L g1508 ( 
.A(n_1338),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1338),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1315),
.A2(n_1429),
.B1(n_1327),
.B2(n_1415),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1338),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1342),
.Y(n_1512)
);

BUFx2_ASAP7_75t_L g1513 ( 
.A(n_1311),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1393),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1304),
.B(n_1312),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1393),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1433),
.B(n_1417),
.Y(n_1517)
);

OAI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1471),
.A2(n_1405),
.B1(n_1408),
.B2(n_1313),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1440),
.B(n_1406),
.Y(n_1519)
);

INVx1_ASAP7_75t_SL g1520 ( 
.A(n_1513),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1474),
.A2(n_1406),
.B1(n_1424),
.B2(n_1396),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1483),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1431),
.A2(n_1395),
.B(n_1401),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1440),
.B(n_1396),
.Y(n_1524)
);

OAI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1470),
.A2(n_1424),
.B(n_1395),
.Y(n_1525)
);

O2A1O1Ixp33_ASAP7_75t_L g1526 ( 
.A1(n_1438),
.A2(n_1401),
.B(n_1422),
.C(n_1420),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1476),
.B(n_1394),
.Y(n_1527)
);

AND2x4_ASAP7_75t_L g1528 ( 
.A(n_1433),
.B(n_1422),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1482),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1483),
.Y(n_1530)
);

NAND4xp25_ASAP7_75t_L g1531 ( 
.A(n_1473),
.B(n_1447),
.C(n_1442),
.D(n_1454),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1442),
.B(n_1480),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_R g1533 ( 
.A(n_1477),
.B(n_1502),
.Y(n_1533)
);

BUFx12f_ASAP7_75t_L g1534 ( 
.A(n_1513),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1432),
.B(n_1434),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1483),
.Y(n_1536)
);

AOI221xp5_ASAP7_75t_L g1537 ( 
.A1(n_1479),
.A2(n_1460),
.B1(n_1455),
.B2(n_1461),
.C(n_1495),
.Y(n_1537)
);

INVxp67_ASAP7_75t_L g1538 ( 
.A(n_1496),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1492),
.Y(n_1539)
);

OAI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_1458),
.A2(n_1460),
.B(n_1468),
.Y(n_1540)
);

NOR2x1_ASAP7_75t_SL g1541 ( 
.A(n_1437),
.B(n_1481),
.Y(n_1541)
);

A2O1A1Ixp33_ASAP7_75t_L g1542 ( 
.A1(n_1479),
.A2(n_1458),
.B(n_1461),
.C(n_1446),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1489),
.B(n_1449),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1450),
.B(n_1459),
.Y(n_1544)
);

AO21x2_ASAP7_75t_L g1545 ( 
.A1(n_1464),
.A2(n_1466),
.B(n_1465),
.Y(n_1545)
);

OAI22x1_ASAP7_75t_SL g1546 ( 
.A1(n_1472),
.A2(n_1516),
.B1(n_1514),
.B2(n_1512),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1488),
.B(n_1494),
.Y(n_1547)
);

OR2x6_ASAP7_75t_L g1548 ( 
.A(n_1437),
.B(n_1446),
.Y(n_1548)
);

OR2x6_ASAP7_75t_L g1549 ( 
.A(n_1437),
.B(n_1475),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1503),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1482),
.Y(n_1551)
);

AOI221xp5_ASAP7_75t_L g1552 ( 
.A1(n_1495),
.A2(n_1485),
.B1(n_1486),
.B2(n_1467),
.C(n_1451),
.Y(n_1552)
);

AOI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1475),
.A2(n_1468),
.B(n_1498),
.Y(n_1553)
);

AOI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1468),
.A2(n_1444),
.B1(n_1437),
.B2(n_1498),
.Y(n_1554)
);

AOI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1468),
.A2(n_1444),
.B1(n_1498),
.B2(n_1516),
.Y(n_1555)
);

OAI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1457),
.A2(n_1469),
.B(n_1492),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1478),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1451),
.B(n_1452),
.Y(n_1558)
);

A2O1A1Ixp33_ASAP7_75t_L g1559 ( 
.A1(n_1469),
.A2(n_1444),
.B(n_1443),
.C(n_1484),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1467),
.B(n_1493),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1451),
.B(n_1452),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1451),
.B(n_1452),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1467),
.B(n_1436),
.Y(n_1563)
);

NAND2xp33_ASAP7_75t_L g1564 ( 
.A(n_1475),
.B(n_1487),
.Y(n_1564)
);

AO32x2_ASAP7_75t_L g1565 ( 
.A1(n_1435),
.A2(n_1491),
.A3(n_1500),
.B1(n_1453),
.B2(n_1478),
.Y(n_1565)
);

AO21x2_ASAP7_75t_L g1566 ( 
.A1(n_1464),
.A2(n_1465),
.B(n_1466),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1498),
.A2(n_1457),
.B(n_1456),
.Y(n_1567)
);

OAI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1456),
.A2(n_1443),
.B(n_1431),
.Y(n_1568)
);

NOR2x1_ASAP7_75t_L g1569 ( 
.A(n_1514),
.B(n_1481),
.Y(n_1569)
);

OR2x2_ASAP7_75t_SL g1570 ( 
.A(n_1557),
.B(n_1478),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1565),
.B(n_1441),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1522),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1530),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_1533),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1558),
.B(n_1561),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_SL g1576 ( 
.A1(n_1532),
.A2(n_1490),
.B1(n_1484),
.B2(n_1507),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1536),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1561),
.B(n_1463),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1565),
.B(n_1441),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1565),
.B(n_1448),
.Y(n_1580)
);

NOR2xp33_ASAP7_75t_L g1581 ( 
.A(n_1531),
.B(n_1511),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1543),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1562),
.B(n_1439),
.Y(n_1583)
);

INVxp67_ASAP7_75t_L g1584 ( 
.A(n_1545),
.Y(n_1584)
);

INVx2_ASAP7_75t_SL g1585 ( 
.A(n_1545),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1562),
.B(n_1439),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1568),
.B(n_1445),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1566),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1552),
.B(n_1463),
.Y(n_1589)
);

BUFx6f_ASAP7_75t_L g1590 ( 
.A(n_1523),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1548),
.B(n_1541),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1540),
.B(n_1445),
.Y(n_1592)
);

INVxp67_ASAP7_75t_SL g1593 ( 
.A(n_1539),
.Y(n_1593)
);

INVx4_ASAP7_75t_L g1594 ( 
.A(n_1549),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1532),
.B(n_1509),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1575),
.B(n_1563),
.Y(n_1596)
);

AOI33xp33_ASAP7_75t_L g1597 ( 
.A1(n_1576),
.A2(n_1537),
.A3(n_1520),
.B1(n_1555),
.B2(n_1505),
.B3(n_1554),
.Y(n_1597)
);

AOI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1581),
.A2(n_1521),
.B1(n_1589),
.B2(n_1595),
.Y(n_1598)
);

AND2x2_ASAP7_75t_SL g1599 ( 
.A(n_1589),
.B(n_1564),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1583),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_SL g1601 ( 
.A(n_1576),
.B(n_1517),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1573),
.Y(n_1602)
);

BUFx2_ASAP7_75t_L g1603 ( 
.A(n_1591),
.Y(n_1603)
);

INVxp67_ASAP7_75t_L g1604 ( 
.A(n_1581),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1583),
.Y(n_1605)
);

OAI21xp33_ASAP7_75t_SL g1606 ( 
.A1(n_1589),
.A2(n_1569),
.B(n_1549),
.Y(n_1606)
);

INVx1_ASAP7_75t_SL g1607 ( 
.A(n_1583),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1572),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1572),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_SL g1610 ( 
.A(n_1574),
.B(n_1517),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1572),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1592),
.B(n_1538),
.Y(n_1612)
);

AO21x2_ASAP7_75t_L g1613 ( 
.A1(n_1584),
.A2(n_1556),
.B(n_1567),
.Y(n_1613)
);

INVx1_ASAP7_75t_SL g1614 ( 
.A(n_1583),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1595),
.A2(n_1527),
.B1(n_1534),
.B2(n_1524),
.Y(n_1615)
);

NAND3xp33_ASAP7_75t_L g1616 ( 
.A(n_1588),
.B(n_1542),
.C(n_1553),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1594),
.A2(n_1527),
.B1(n_1534),
.B2(n_1524),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1577),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1582),
.B(n_1529),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1577),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1575),
.B(n_1560),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1592),
.B(n_1547),
.Y(n_1622)
);

BUFx6f_ASAP7_75t_L g1623 ( 
.A(n_1590),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1594),
.A2(n_1519),
.B1(n_1551),
.B2(n_1549),
.Y(n_1624)
);

AOI221xp5_ASAP7_75t_L g1625 ( 
.A1(n_1578),
.A2(n_1542),
.B1(n_1559),
.B2(n_1546),
.C(n_1544),
.Y(n_1625)
);

NAND4xp25_ASAP7_75t_SL g1626 ( 
.A(n_1578),
.B(n_1526),
.C(n_1525),
.D(n_1559),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1582),
.B(n_1566),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1594),
.A2(n_1519),
.B1(n_1549),
.B2(n_1550),
.Y(n_1628)
);

OAI221xp5_ASAP7_75t_L g1629 ( 
.A1(n_1578),
.A2(n_1510),
.B1(n_1518),
.B2(n_1535),
.C(n_1564),
.Y(n_1629)
);

INVxp67_ASAP7_75t_SL g1630 ( 
.A(n_1588),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1602),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1603),
.B(n_1571),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1608),
.Y(n_1633)
);

NAND2x1p5_ASAP7_75t_L g1634 ( 
.A(n_1599),
.B(n_1594),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1608),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1603),
.B(n_1571),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1600),
.B(n_1571),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1609),
.Y(n_1638)
);

NAND2xp33_ASAP7_75t_R g1639 ( 
.A(n_1612),
.B(n_1533),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1600),
.B(n_1571),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1610),
.B(n_1574),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1598),
.B(n_1586),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1607),
.B(n_1579),
.Y(n_1643)
);

INVx4_ASAP7_75t_L g1644 ( 
.A(n_1623),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1609),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1598),
.B(n_1586),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1623),
.B(n_1591),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1622),
.B(n_1586),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1604),
.B(n_1575),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1607),
.B(n_1614),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1611),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1614),
.B(n_1579),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1621),
.B(n_1592),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1629),
.B(n_1528),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1602),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1605),
.B(n_1579),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1611),
.Y(n_1657)
);

INVx2_ASAP7_75t_SL g1658 ( 
.A(n_1623),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1627),
.B(n_1580),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1627),
.B(n_1580),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1621),
.B(n_1592),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1626),
.A2(n_1490),
.B1(n_1484),
.B2(n_1528),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1599),
.B(n_1580),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1618),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1620),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1620),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1633),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1649),
.B(n_1625),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1633),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1649),
.B(n_1597),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1663),
.B(n_1599),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1653),
.B(n_1661),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1642),
.B(n_1619),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1631),
.Y(n_1674)
);

INVxp67_ASAP7_75t_L g1675 ( 
.A(n_1639),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1638),
.Y(n_1676)
);

INVxp67_ASAP7_75t_L g1677 ( 
.A(n_1654),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1642),
.B(n_1619),
.Y(n_1678)
);

OAI21xp5_ASAP7_75t_SL g1679 ( 
.A1(n_1662),
.A2(n_1601),
.B(n_1616),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1653),
.B(n_1616),
.Y(n_1680)
);

INVx1_ASAP7_75t_SL g1681 ( 
.A(n_1641),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1638),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1663),
.B(n_1591),
.Y(n_1683)
);

AND2x4_ASAP7_75t_L g1684 ( 
.A(n_1647),
.B(n_1591),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1663),
.B(n_1591),
.Y(n_1685)
);

AOI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1662),
.A2(n_1606),
.B1(n_1528),
.B2(n_1484),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1651),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1651),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1631),
.Y(n_1689)
);

INVxp67_ASAP7_75t_SL g1690 ( 
.A(n_1634),
.Y(n_1690)
);

NAND2x1_ASAP7_75t_L g1691 ( 
.A(n_1644),
.B(n_1647),
.Y(n_1691)
);

NOR2x1_ASAP7_75t_L g1692 ( 
.A(n_1644),
.B(n_1517),
.Y(n_1692)
);

NOR3x1_ASAP7_75t_L g1693 ( 
.A(n_1646),
.B(n_1504),
.C(n_1515),
.Y(n_1693)
);

OR2x6_ASAP7_75t_L g1694 ( 
.A(n_1634),
.B(n_1623),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1634),
.B(n_1591),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1646),
.B(n_1587),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1634),
.B(n_1647),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1647),
.B(n_1591),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1631),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1665),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1665),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1661),
.B(n_1587),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_SL g1703 ( 
.A(n_1647),
.B(n_1606),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1655),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1655),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1632),
.B(n_1623),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1648),
.B(n_1587),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1655),
.Y(n_1708)
);

AOI32xp33_ASAP7_75t_SL g1709 ( 
.A1(n_1635),
.A2(n_1630),
.A3(n_1505),
.B1(n_1593),
.B2(n_1504),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1700),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1667),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1680),
.B(n_1648),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_SL g1713 ( 
.A(n_1675),
.B(n_1594),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1670),
.B(n_1615),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1667),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1668),
.B(n_1587),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1699),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1669),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1692),
.B(n_1644),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1671),
.B(n_1632),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1669),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1671),
.B(n_1632),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1692),
.B(n_1636),
.Y(n_1723)
);

OR2x6_ASAP7_75t_L g1724 ( 
.A(n_1691),
.B(n_1507),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1680),
.B(n_1673),
.Y(n_1725)
);

NAND2x1p5_ASAP7_75t_L g1726 ( 
.A(n_1691),
.B(n_1644),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1697),
.B(n_1636),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1697),
.B(n_1636),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1677),
.B(n_1596),
.Y(n_1729)
);

INVxp67_ASAP7_75t_SL g1730 ( 
.A(n_1693),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1676),
.Y(n_1731)
);

INVxp67_ASAP7_75t_L g1732 ( 
.A(n_1681),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1699),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1679),
.B(n_1515),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1676),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1682),
.Y(n_1736)
);

OAI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1679),
.A2(n_1617),
.B(n_1624),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1682),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1687),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1693),
.B(n_1596),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_SL g1741 ( 
.A(n_1690),
.B(n_1594),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1683),
.B(n_1656),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1678),
.B(n_1637),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1672),
.B(n_1650),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1696),
.B(n_1637),
.Y(n_1745)
);

AOI221xp5_ASAP7_75t_SL g1746 ( 
.A1(n_1737),
.A2(n_1703),
.B1(n_1706),
.B2(n_1683),
.C(n_1685),
.Y(n_1746)
);

OAI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1730),
.A2(n_1686),
.B1(n_1694),
.B2(n_1709),
.Y(n_1747)
);

OAI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1714),
.A2(n_1686),
.B1(n_1694),
.B2(n_1709),
.Y(n_1748)
);

AOI21xp33_ASAP7_75t_L g1749 ( 
.A1(n_1732),
.A2(n_1694),
.B(n_1688),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1734),
.B(n_1685),
.Y(n_1750)
);

OAI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1716),
.A2(n_1694),
.B1(n_1628),
.B2(n_1570),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1726),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1711),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1725),
.B(n_1672),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1720),
.B(n_1695),
.Y(n_1755)
);

AND2x4_ASAP7_75t_SL g1756 ( 
.A(n_1724),
.B(n_1694),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1711),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1724),
.A2(n_1570),
.B1(n_1684),
.B2(n_1695),
.Y(n_1758)
);

NOR2x1_ASAP7_75t_L g1759 ( 
.A(n_1724),
.B(n_1687),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1725),
.B(n_1512),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1720),
.B(n_1698),
.Y(n_1761)
);

OAI21xp33_ASAP7_75t_L g1762 ( 
.A1(n_1713),
.A2(n_1706),
.B(n_1702),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1726),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1710),
.B(n_1512),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1718),
.Y(n_1765)
);

OAI21xp5_ASAP7_75t_SL g1766 ( 
.A1(n_1740),
.A2(n_1684),
.B(n_1698),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_SL g1767 ( 
.A(n_1719),
.B(n_1623),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1729),
.B(n_1707),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1722),
.B(n_1684),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1718),
.Y(n_1770)
);

OAI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1719),
.A2(n_1701),
.B(n_1688),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1753),
.Y(n_1772)
);

OAI322xp33_ASAP7_75t_L g1773 ( 
.A1(n_1747),
.A2(n_1710),
.A3(n_1715),
.B1(n_1731),
.B2(n_1736),
.C1(n_1735),
.C2(n_1739),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1757),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1764),
.B(n_1722),
.Y(n_1775)
);

HB1xp67_ASAP7_75t_L g1776 ( 
.A(n_1765),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1769),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1770),
.Y(n_1778)
);

O2A1O1Ixp33_ASAP7_75t_L g1779 ( 
.A1(n_1747),
.A2(n_1738),
.B(n_1721),
.C(n_1724),
.Y(n_1779)
);

AOI222xp33_ASAP7_75t_L g1780 ( 
.A1(n_1748),
.A2(n_1723),
.B1(n_1721),
.B2(n_1743),
.C1(n_1741),
.C2(n_1745),
.Y(n_1780)
);

OAI211xp5_ASAP7_75t_L g1781 ( 
.A1(n_1749),
.A2(n_1723),
.B(n_1712),
.C(n_1744),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1750),
.B(n_1712),
.Y(n_1782)
);

INVxp67_ASAP7_75t_L g1783 ( 
.A(n_1764),
.Y(n_1783)
);

AOI21xp33_ASAP7_75t_L g1784 ( 
.A1(n_1748),
.A2(n_1719),
.B(n_1744),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1754),
.Y(n_1785)
);

OAI32xp33_ASAP7_75t_L g1786 ( 
.A1(n_1771),
.A2(n_1726),
.A3(n_1701),
.B1(n_1728),
.B2(n_1727),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1768),
.B(n_1717),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1755),
.B(n_1761),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1759),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1760),
.B(n_1727),
.Y(n_1790)
);

AOI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1746),
.A2(n_1728),
.B1(n_1684),
.B2(n_1613),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1780),
.A2(n_1760),
.B1(n_1754),
.B2(n_1762),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1776),
.Y(n_1793)
);

INVx1_ASAP7_75t_SL g1794 ( 
.A(n_1787),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1789),
.Y(n_1795)
);

AOI31xp33_ASAP7_75t_L g1796 ( 
.A1(n_1785),
.A2(n_1752),
.A3(n_1763),
.B(n_1751),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1776),
.Y(n_1797)
);

OAI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1779),
.A2(n_1766),
.B1(n_1756),
.B2(n_1758),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1787),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1777),
.B(n_1742),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1788),
.B(n_1777),
.Y(n_1801)
);

XNOR2x1_ASAP7_75t_L g1802 ( 
.A(n_1789),
.B(n_1497),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1772),
.Y(n_1803)
);

NAND4xp25_ASAP7_75t_L g1804 ( 
.A(n_1792),
.B(n_1801),
.C(n_1798),
.D(n_1794),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1801),
.B(n_1788),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1793),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1799),
.B(n_1783),
.Y(n_1807)
);

NAND3xp33_ASAP7_75t_L g1808 ( 
.A(n_1802),
.B(n_1784),
.C(n_1781),
.Y(n_1808)
);

AOI221xp5_ASAP7_75t_L g1809 ( 
.A1(n_1796),
.A2(n_1773),
.B1(n_1786),
.B2(n_1774),
.C(n_1778),
.Y(n_1809)
);

NAND3xp33_ASAP7_75t_L g1810 ( 
.A(n_1802),
.B(n_1791),
.C(n_1775),
.Y(n_1810)
);

NAND4xp25_ASAP7_75t_L g1811 ( 
.A(n_1800),
.B(n_1782),
.C(n_1790),
.D(n_1767),
.Y(n_1811)
);

AOI211xp5_ASAP7_75t_L g1812 ( 
.A1(n_1797),
.A2(n_1767),
.B(n_1717),
.C(n_1733),
.Y(n_1812)
);

NAND3xp33_ASAP7_75t_L g1813 ( 
.A(n_1795),
.B(n_1733),
.C(n_1644),
.Y(n_1813)
);

NOR3xp33_ASAP7_75t_L g1814 ( 
.A(n_1803),
.B(n_1499),
.C(n_1497),
.Y(n_1814)
);

AND4x1_ASAP7_75t_L g1815 ( 
.A(n_1808),
.B(n_1795),
.C(n_1511),
.D(n_1509),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1805),
.B(n_1742),
.Y(n_1816)
);

AOI322xp5_ASAP7_75t_L g1817 ( 
.A1(n_1809),
.A2(n_1660),
.A3(n_1659),
.B1(n_1652),
.B2(n_1643),
.C1(n_1640),
.C2(n_1637),
.Y(n_1817)
);

NAND4xp25_ASAP7_75t_L g1818 ( 
.A(n_1804),
.B(n_1497),
.C(n_1499),
.D(n_1503),
.Y(n_1818)
);

AOI221xp5_ASAP7_75t_L g1819 ( 
.A1(n_1810),
.A2(n_1756),
.B1(n_1658),
.B2(n_1704),
.C(n_1699),
.Y(n_1819)
);

NAND3x1_ASAP7_75t_SL g1820 ( 
.A(n_1819),
.B(n_1814),
.C(n_1807),
.Y(n_1820)
);

AND4x1_ASAP7_75t_L g1821 ( 
.A(n_1816),
.B(n_1806),
.C(n_1813),
.D(n_1812),
.Y(n_1821)
);

OAI31xp33_ASAP7_75t_L g1822 ( 
.A1(n_1818),
.A2(n_1811),
.A3(n_1658),
.B(n_1503),
.Y(n_1822)
);

AND2x4_ASAP7_75t_L g1823 ( 
.A(n_1815),
.B(n_1462),
.Y(n_1823)
);

NOR2x1_ASAP7_75t_L g1824 ( 
.A(n_1817),
.B(n_1499),
.Y(n_1824)
);

AOI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1818),
.A2(n_1658),
.B(n_1704),
.Y(n_1825)
);

INVx2_ASAP7_75t_SL g1826 ( 
.A(n_1823),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1821),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1820),
.Y(n_1828)
);

XOR2x1_ASAP7_75t_L g1829 ( 
.A(n_1824),
.B(n_1506),
.Y(n_1829)
);

NAND4xp75_ASAP7_75t_L g1830 ( 
.A(n_1822),
.B(n_1704),
.C(n_1705),
.D(n_1708),
.Y(n_1830)
);

NOR3xp33_ASAP7_75t_L g1831 ( 
.A(n_1827),
.B(n_1825),
.C(n_1508),
.Y(n_1831)
);

AOI221xp5_ASAP7_75t_L g1832 ( 
.A1(n_1828),
.A2(n_1708),
.B1(n_1705),
.B2(n_1689),
.C(n_1674),
.Y(n_1832)
);

AOI222xp33_ASAP7_75t_L g1833 ( 
.A1(n_1826),
.A2(n_1674),
.B1(n_1689),
.B2(n_1584),
.C1(n_1585),
.C2(n_1660),
.Y(n_1833)
);

HB1xp67_ASAP7_75t_L g1834 ( 
.A(n_1831),
.Y(n_1834)
);

AOI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1834),
.A2(n_1830),
.B1(n_1832),
.B2(n_1833),
.Y(n_1835)
);

XNOR2xp5_ASAP7_75t_L g1836 ( 
.A(n_1835),
.B(n_1829),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1835),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1836),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1837),
.Y(n_1839)
);

AO21x2_ASAP7_75t_L g1840 ( 
.A1(n_1839),
.A2(n_1659),
.B(n_1660),
.Y(n_1840)
);

OAI21x1_ASAP7_75t_L g1841 ( 
.A1(n_1838),
.A2(n_1508),
.B(n_1659),
.Y(n_1841)
);

XNOR2xp5_ASAP7_75t_L g1842 ( 
.A(n_1841),
.B(n_1508),
.Y(n_1842)
);

OAI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1842),
.A2(n_1840),
.B1(n_1650),
.B2(n_1508),
.Y(n_1843)
);

OAI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1843),
.A2(n_1840),
.B1(n_1650),
.B2(n_1481),
.Y(n_1844)
);

AOI221xp5_ASAP7_75t_L g1845 ( 
.A1(n_1844),
.A2(n_1666),
.B1(n_1664),
.B2(n_1645),
.C(n_1657),
.Y(n_1845)
);

AOI211xp5_ASAP7_75t_L g1846 ( 
.A1(n_1845),
.A2(n_1501),
.B(n_1500),
.C(n_1491),
.Y(n_1846)
);


endmodule