module fake_ariane_2766_n_1934 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_172, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1934);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1934;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_177;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_110),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_145),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_28),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_14),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_63),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_18),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_109),
.Y(n_181)
);

BUFx10_ASAP7_75t_L g182 ( 
.A(n_124),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_115),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_5),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_130),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_31),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_83),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_139),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_0),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_19),
.Y(n_191)
);

INVxp67_ASAP7_75t_SL g192 ( 
.A(n_50),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_67),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_8),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_102),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_69),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_74),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_78),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_132),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_25),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g201 ( 
.A(n_65),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_63),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_168),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_55),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_25),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_113),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_73),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_103),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_93),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_31),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_125),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_37),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_87),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_112),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_39),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_33),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_97),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_164),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_69),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_35),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_94),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_171),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_151),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_100),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_162),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_67),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_138),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_126),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_15),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_8),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_54),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_150),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_59),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_172),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_118),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_146),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_56),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_36),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_33),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_143),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_17),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_64),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_159),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_3),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_77),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_128),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_5),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_44),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_58),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_104),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_14),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_80),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_88),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_99),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_27),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_59),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_161),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_117),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_55),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_147),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_89),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_70),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_6),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_34),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_81),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_141),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_20),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_51),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_92),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_58),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_131),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_2),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_160),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_107),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_170),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_163),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_167),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_10),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_0),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_12),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_111),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_37),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_28),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_96),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_101),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_56),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_54),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_62),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_35),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_136),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_165),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_27),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_119),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_7),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_60),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_15),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_127),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_66),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_72),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_48),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_142),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_106),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_135),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_157),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_51),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_66),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_2),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_46),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_90),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_4),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_53),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_3),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_169),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_133),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_79),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_45),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_155),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_72),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_57),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_6),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_60),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_137),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_86),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_84),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_120),
.Y(n_325)
);

BUFx10_ASAP7_75t_L g326 ( 
.A(n_30),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_16),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_166),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_34),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_18),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_68),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_17),
.Y(n_332)
);

BUFx10_ASAP7_75t_L g333 ( 
.A(n_50),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_19),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_1),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_11),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_121),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_62),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_71),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_11),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_22),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_41),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_148),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_95),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_181),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_175),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_280),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_201),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_201),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_201),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_195),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_201),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_198),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_245),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_258),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_201),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_314),
.B(n_1),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_175),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_201),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_201),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_271),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_303),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_280),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_180),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_179),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_205),
.Y(n_366)
);

INVxp33_ASAP7_75t_SL g367 ( 
.A(n_184),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_190),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_R g369 ( 
.A(n_173),
.B(n_158),
.Y(n_369)
);

INVxp33_ASAP7_75t_SL g370 ( 
.A(n_191),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_200),
.Y(n_371)
);

NOR2xp67_ASAP7_75t_L g372 ( 
.A(n_212),
.B(n_4),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_201),
.Y(n_373)
);

NOR2xp67_ASAP7_75t_L g374 ( 
.A(n_212),
.B(n_7),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_202),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_201),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_204),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_176),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_207),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_216),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_242),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_176),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_219),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_213),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_220),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_213),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_177),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_299),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_308),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_214),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_214),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_312),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_233),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_221),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_221),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_240),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_177),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_240),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_237),
.Y(n_399)
);

OR2x2_ASAP7_75t_L g400 ( 
.A(n_248),
.B(n_9),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_241),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_318),
.Y(n_402)
);

NOR2xp67_ASAP7_75t_L g403 ( 
.A(n_248),
.B(n_9),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_244),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_314),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_257),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_186),
.B(n_10),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_186),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_187),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_187),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_247),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_257),
.B(n_12),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_260),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_260),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_186),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_187),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_251),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_255),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_276),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_276),
.Y(n_420)
);

NOR2xp67_ASAP7_75t_L g421 ( 
.A(n_248),
.B(n_283),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_277),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_256),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_259),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_262),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_264),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_277),
.B(n_13),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_302),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_188),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_302),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_365),
.B(n_218),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_348),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_348),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_351),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_378),
.B(n_223),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_349),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_407),
.B(n_378),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_354),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_349),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_350),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_371),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_350),
.Y(n_442)
);

OR2x6_ASAP7_75t_L g443 ( 
.A(n_400),
.B(n_283),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_382),
.B(n_297),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_352),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_357),
.B(n_300),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_352),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_366),
.Y(n_448)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_407),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_356),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_356),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_355),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_359),
.Y(n_453)
);

BUFx8_ASAP7_75t_L g454 ( 
.A(n_400),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_359),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_360),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_360),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_373),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_373),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_376),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_409),
.B(n_182),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_408),
.B(n_309),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_376),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_382),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_362),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_345),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_384),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_384),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_381),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_386),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_386),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_390),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_353),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_390),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_388),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_389),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_391),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_347),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_391),
.B(n_304),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_394),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_394),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_361),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_395),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_364),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_395),
.B(n_226),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_396),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_368),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_396),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_375),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_377),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_398),
.B(n_226),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_398),
.B(n_304),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_406),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_379),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_406),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_413),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_380),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_404),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_383),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_413),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_414),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_414),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_385),
.B(n_182),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_419),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_419),
.B(n_226),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_393),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_399),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_464),
.Y(n_508)
);

NAND3xp33_ASAP7_75t_L g509 ( 
.A(n_462),
.B(n_357),
.C(n_401),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_432),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_464),
.Y(n_511)
);

NAND3xp33_ASAP7_75t_L g512 ( 
.A(n_462),
.B(n_417),
.C(n_411),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_449),
.B(n_415),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_449),
.B(n_420),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_449),
.B(n_437),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_445),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_441),
.B(n_347),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_468),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_468),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_432),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_477),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_449),
.B(n_420),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_437),
.B(n_422),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_437),
.B(n_422),
.Y(n_524)
);

AND2x6_ASAP7_75t_L g525 ( 
.A(n_437),
.B(n_252),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_441),
.B(n_363),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_445),
.Y(n_527)
);

AND2x6_ASAP7_75t_L g528 ( 
.A(n_437),
.B(n_252),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_486),
.B(n_428),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_477),
.Y(n_530)
);

OAI22xp33_ASAP7_75t_L g531 ( 
.A1(n_443),
.A2(n_374),
.B1(n_372),
.B2(n_405),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_467),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_481),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_481),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_445),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_467),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_448),
.Y(n_537)
);

NAND2x1p5_ASAP7_75t_L g538 ( 
.A(n_503),
.B(n_372),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_443),
.B(n_374),
.Y(n_539)
);

AND2x6_ASAP7_75t_L g540 ( 
.A(n_491),
.B(n_252),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_478),
.Y(n_541)
);

NAND2x1p5_ASAP7_75t_L g542 ( 
.A(n_491),
.B(n_428),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_436),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_486),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_447),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_443),
.B(n_346),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_436),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_443),
.B(n_358),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_439),
.Y(n_549)
);

INVx1_ASAP7_75t_SL g550 ( 
.A(n_469),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_434),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_439),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_486),
.B(n_367),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_498),
.B(n_478),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_438),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_443),
.A2(n_430),
.B1(n_412),
.B2(n_427),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_498),
.B(n_418),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_486),
.B(n_370),
.Y(n_558)
);

NAND2x1_ASAP7_75t_L g559 ( 
.A(n_443),
.B(n_430),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_452),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_484),
.Y(n_561)
);

AND2x6_ASAP7_75t_L g562 ( 
.A(n_491),
.B(n_253),
.Y(n_562)
);

BUFx4f_ASAP7_75t_L g563 ( 
.A(n_467),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_467),
.B(n_423),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_483),
.Y(n_565)
);

OAI221xp5_ASAP7_75t_L g566 ( 
.A1(n_435),
.A2(n_387),
.B1(n_397),
.B2(n_403),
.C(n_230),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_454),
.A2(n_424),
.B1(n_426),
.B2(n_425),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_465),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_467),
.B(n_470),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_483),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_466),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_467),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_467),
.B(n_470),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_491),
.B(n_421),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_502),
.B(n_429),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_487),
.B(n_410),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_491),
.B(n_421),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_447),
.Y(n_578)
);

OAI22xp33_ASAP7_75t_L g579 ( 
.A1(n_461),
.A2(n_249),
.B1(n_267),
.B2(n_286),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_489),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_502),
.B(n_416),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_447),
.Y(n_582)
);

NAND2x1p5_ASAP7_75t_L g583 ( 
.A(n_505),
.B(n_403),
.Y(n_583)
);

INVx6_ASAP7_75t_L g584 ( 
.A(n_505),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_454),
.A2(n_319),
.B1(n_334),
.B2(n_283),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_488),
.Y(n_586)
);

INVx5_ASAP7_75t_L g587 ( 
.A(n_470),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_488),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_470),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_502),
.B(n_317),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_501),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_490),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_501),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_470),
.B(n_502),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_494),
.B(n_326),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_505),
.B(n_193),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_504),
.B(n_183),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_473),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_L g599 ( 
.A1(n_454),
.A2(n_319),
.B1(n_334),
.B2(n_194),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_450),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_505),
.B(n_193),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_504),
.B(n_317),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_470),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_497),
.Y(n_604)
);

AND2x6_ASAP7_75t_L g605 ( 
.A(n_505),
.B(n_253),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_471),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_454),
.B(n_328),
.Y(n_607)
);

AND2x6_ASAP7_75t_L g608 ( 
.A(n_485),
.B(n_253),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_454),
.B(n_440),
.Y(n_609)
);

OR2x2_ASAP7_75t_L g610 ( 
.A(n_499),
.B(n_194),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_440),
.B(n_451),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_506),
.Y(n_612)
);

INVx6_ASAP7_75t_L g613 ( 
.A(n_470),
.Y(n_613)
);

INVxp67_ASAP7_75t_SL g614 ( 
.A(n_433),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_433),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_451),
.B(n_453),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_471),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_471),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_453),
.B(n_328),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_450),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_472),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_507),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_435),
.A2(n_192),
.B1(n_272),
.B2(n_270),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_SL g624 ( 
.A(n_461),
.B(n_182),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_450),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_472),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_458),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_456),
.B(n_273),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_472),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_474),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_485),
.B(n_196),
.Y(n_631)
);

NOR2x1p5_ASAP7_75t_L g632 ( 
.A(n_444),
.B(n_196),
.Y(n_632)
);

BUFx10_ASAP7_75t_L g633 ( 
.A(n_482),
.Y(n_633)
);

INVxp33_ASAP7_75t_SL g634 ( 
.A(n_431),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_485),
.B(n_210),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_444),
.B(n_210),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_458),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_475),
.Y(n_638)
);

CKINVDCx16_ASAP7_75t_R g639 ( 
.A(n_476),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_458),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_459),
.B(n_273),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_474),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_456),
.B(n_211),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_433),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_474),
.Y(n_645)
);

NOR2x1p5_ASAP7_75t_L g646 ( 
.A(n_479),
.B(n_215),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_480),
.Y(n_647)
);

OR2x6_ASAP7_75t_L g648 ( 
.A(n_479),
.B(n_319),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_480),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_492),
.B(n_215),
.Y(n_650)
);

INVx4_ASAP7_75t_L g651 ( 
.A(n_433),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_480),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_431),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_459),
.B(n_300),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_446),
.A2(n_268),
.B1(n_278),
.B2(n_279),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_433),
.Y(n_656)
);

BUFx10_ASAP7_75t_L g657 ( 
.A(n_460),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_493),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_460),
.B(n_188),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_493),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_575),
.B(n_581),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_546),
.A2(n_446),
.B1(n_496),
.B2(n_495),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_510),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_553),
.B(n_493),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_553),
.B(n_558),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_541),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_546),
.A2(n_500),
.B1(n_496),
.B2(n_495),
.Y(n_667)
);

AND2x2_ASAP7_75t_SL g668 ( 
.A(n_624),
.B(n_492),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_585),
.A2(n_463),
.B1(n_459),
.B2(n_495),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_510),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_558),
.B(n_496),
.Y(n_671)
);

O2A1O1Ixp5_ASAP7_75t_L g672 ( 
.A1(n_594),
.A2(n_463),
.B(n_500),
.C(n_334),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_513),
.B(n_500),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_650),
.B(n_463),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_650),
.B(n_433),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_650),
.B(n_433),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_657),
.B(n_442),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_516),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_514),
.B(n_442),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_509),
.B(n_442),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_657),
.Y(n_681)
);

NAND2x1_ASAP7_75t_L g682 ( 
.A(n_525),
.B(n_442),
.Y(n_682)
);

OAI22xp33_ASAP7_75t_L g683 ( 
.A1(n_567),
.A2(n_231),
.B1(n_229),
.B2(n_230),
.Y(n_683)
);

A2O1A1Ixp33_ASAP7_75t_L g684 ( 
.A1(n_590),
.A2(n_231),
.B(n_229),
.C(n_238),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_546),
.B(n_548),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_522),
.B(n_442),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_554),
.B(n_392),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_515),
.B(n_442),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_520),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_643),
.B(n_556),
.Y(n_690)
);

A2O1A1Ixp33_ASAP7_75t_L g691 ( 
.A1(n_590),
.A2(n_310),
.B(n_238),
.C(n_239),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_520),
.Y(n_692)
);

NAND2xp33_ASAP7_75t_L g693 ( 
.A(n_525),
.B(n_457),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_643),
.B(n_442),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_556),
.B(n_455),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_SL g696 ( 
.A1(n_548),
.A2(n_402),
.B1(n_326),
.B2(n_333),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_548),
.B(n_455),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_597),
.B(n_455),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_523),
.B(n_455),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_557),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_524),
.B(n_455),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_526),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_516),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_543),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_574),
.B(n_577),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_525),
.A2(n_227),
.B1(n_203),
.B2(n_344),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_543),
.Y(n_707)
);

NOR2x1p5_ASAP7_75t_L g708 ( 
.A(n_551),
.B(n_282),
.Y(n_708)
);

AO22x1_ASAP7_75t_L g709 ( 
.A1(n_517),
.A2(n_306),
.B1(n_307),
.B2(n_342),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_574),
.B(n_455),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_527),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_585),
.A2(n_243),
.B1(n_182),
.B2(n_333),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_657),
.B(n_457),
.Y(n_713)
);

A2O1A1Ixp33_ASAP7_75t_SL g714 ( 
.A1(n_616),
.A2(n_311),
.B(n_263),
.C(n_340),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_527),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_547),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_576),
.Y(n_717)
);

O2A1O1Ixp5_ASAP7_75t_L g718 ( 
.A1(n_594),
.A2(n_239),
.B(n_327),
.C(n_263),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_574),
.B(n_455),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_535),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_577),
.B(n_457),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_577),
.B(n_457),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_539),
.B(n_288),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_648),
.B(n_457),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_584),
.B(n_457),
.Y(n_725)
);

AO22x1_ASAP7_75t_L g726 ( 
.A1(n_551),
.A2(n_329),
.B1(n_316),
.B2(n_341),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_584),
.B(n_457),
.Y(n_727)
);

OAI22x1_ASAP7_75t_L g728 ( 
.A1(n_571),
.A2(n_287),
.B1(n_298),
.B2(n_320),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_648),
.B(n_288),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_525),
.A2(n_206),
.B1(n_343),
.B2(n_224),
.Y(n_730)
);

OR2x6_ASAP7_75t_L g731 ( 
.A(n_559),
.B(n_294),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_544),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_547),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_584),
.B(n_289),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_549),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_648),
.B(n_294),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_539),
.B(n_296),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_531),
.B(n_292),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_512),
.B(n_544),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_610),
.Y(n_740)
);

NOR2x1p5_ASAP7_75t_L g741 ( 
.A(n_555),
.B(n_295),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_544),
.B(n_178),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_599),
.A2(n_243),
.B1(n_326),
.B2(n_333),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_539),
.B(n_178),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_561),
.B(n_580),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_538),
.B(n_542),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_525),
.A2(n_189),
.B1(n_208),
.B2(n_209),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_535),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_508),
.B(n_296),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_511),
.B(n_305),
.Y(n_750)
);

NOR2xp67_ASAP7_75t_L g751 ( 
.A(n_604),
.B(n_174),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_550),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_518),
.B(n_305),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_519),
.B(n_310),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_528),
.A2(n_290),
.B1(n_199),
.B2(n_217),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_521),
.B(n_530),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_549),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_552),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_609),
.B(n_178),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_638),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_538),
.B(n_321),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_533),
.B(n_311),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_592),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_545),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_528),
.A2(n_608),
.B1(n_562),
.B2(n_605),
.Y(n_765)
);

OR2x2_ASAP7_75t_SL g766 ( 
.A(n_639),
.B(n_327),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_552),
.B(n_178),
.Y(n_767)
);

BUFx8_ASAP7_75t_L g768 ( 
.A(n_612),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_555),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_534),
.B(n_331),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_565),
.B(n_331),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_570),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_586),
.B(n_332),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_588),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_542),
.B(n_330),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_528),
.A2(n_281),
.B1(n_232),
.B2(n_234),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_595),
.B(n_326),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_591),
.B(n_332),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_593),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_630),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_528),
.B(n_339),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_528),
.B(n_339),
.Y(n_782)
);

INVxp67_ASAP7_75t_L g783 ( 
.A(n_622),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_596),
.B(n_340),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_658),
.B(n_336),
.Y(n_785)
);

NOR2x1p5_ASAP7_75t_L g786 ( 
.A(n_560),
.B(n_338),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_616),
.B(n_185),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_608),
.B(n_222),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_608),
.B(n_225),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_545),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_SL g791 ( 
.A(n_560),
.B(n_243),
.Y(n_791)
);

BUFx3_ASAP7_75t_L g792 ( 
.A(n_568),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_608),
.A2(n_275),
.B1(n_337),
.B2(n_235),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_578),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_578),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_608),
.B(n_228),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_614),
.A2(n_284),
.B(n_236),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_630),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_568),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_529),
.B(n_246),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_582),
.Y(n_801)
);

NAND2xp33_ASAP7_75t_L g802 ( 
.A(n_540),
.B(n_300),
.Y(n_802)
);

BUFx5_ASAP7_75t_L g803 ( 
.A(n_540),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_599),
.A2(n_243),
.B1(n_333),
.B2(n_335),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_540),
.A2(n_291),
.B1(n_250),
.B2(n_325),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_582),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_633),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_656),
.Y(n_808)
);

OAI22xp33_ASAP7_75t_L g809 ( 
.A1(n_636),
.A2(n_335),
.B1(n_300),
.B2(n_285),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_540),
.A2(n_254),
.B1(n_261),
.B2(n_324),
.Y(n_810)
);

INVx8_ASAP7_75t_L g811 ( 
.A(n_540),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_656),
.B(n_178),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_646),
.A2(n_335),
.B1(n_300),
.B2(n_188),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_606),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_607),
.B(n_265),
.Y(n_815)
);

NOR2xp67_ASAP7_75t_L g816 ( 
.A(n_571),
.B(n_266),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_596),
.B(n_269),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_596),
.B(n_274),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_562),
.A2(n_335),
.B1(n_300),
.B2(n_285),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_601),
.B(n_315),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_601),
.B(n_313),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_601),
.B(n_323),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_611),
.A2(n_293),
.B(n_301),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_600),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_562),
.A2(n_335),
.B1(n_285),
.B2(n_369),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_600),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_620),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_583),
.B(n_631),
.Y(n_828)
);

AND2x6_ASAP7_75t_SL g829 ( 
.A(n_598),
.B(n_13),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_631),
.B(n_16),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_620),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_656),
.B(n_197),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_763),
.Y(n_833)
);

NAND2x1p5_ASAP7_75t_L g834 ( 
.A(n_685),
.B(n_587),
.Y(n_834)
);

AO22x1_ASAP7_75t_L g835 ( 
.A1(n_768),
.A2(n_598),
.B1(n_634),
.B2(n_769),
.Y(n_835)
);

INVx1_ASAP7_75t_SL g836 ( 
.A(n_752),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_685),
.A2(n_605),
.B1(n_562),
.B2(n_579),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_763),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_772),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_665),
.B(n_583),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_705),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_811),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_774),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_690),
.A2(n_668),
.B1(n_738),
.B2(n_661),
.Y(n_844)
);

AND2x4_ASAP7_75t_SL g845 ( 
.A(n_830),
.B(n_633),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_811),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_661),
.B(n_632),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_678),
.Y(n_848)
);

NOR3xp33_ASAP7_75t_SL g849 ( 
.A(n_683),
.B(n_623),
.C(n_653),
.Y(n_849)
);

BUFx3_ASAP7_75t_L g850 ( 
.A(n_769),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_678),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_779),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_807),
.B(n_631),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_756),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_702),
.B(n_564),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_830),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_703),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_681),
.B(n_635),
.Y(n_858)
);

BUFx12f_ASAP7_75t_SL g859 ( 
.A(n_745),
.Y(n_859)
);

CKINVDCx20_ASAP7_75t_R g860 ( 
.A(n_768),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_814),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_681),
.B(n_635),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_792),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_668),
.A2(n_605),
.B1(n_562),
.B2(n_564),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_811),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_811),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_738),
.A2(n_605),
.B1(n_635),
.B2(n_566),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_703),
.Y(n_868)
);

BUFx4f_ASAP7_75t_L g869 ( 
.A(n_666),
.Y(n_869)
);

OAI21xp33_ASAP7_75t_L g870 ( 
.A1(n_791),
.A2(n_655),
.B(n_602),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_664),
.B(n_605),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_803),
.B(n_656),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_792),
.Y(n_873)
);

INVx5_ASAP7_75t_L g874 ( 
.A(n_808),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_780),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_830),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_807),
.B(n_537),
.Y(n_877)
);

OR2x6_ASAP7_75t_L g878 ( 
.A(n_799),
.B(n_633),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_687),
.B(n_653),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_711),
.Y(n_880)
);

NAND2xp33_ASAP7_75t_SL g881 ( 
.A(n_732),
.B(n_619),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_803),
.B(n_532),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_711),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_671),
.B(n_659),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_787),
.B(n_659),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_715),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_715),
.Y(n_887)
);

OR2x6_ASAP7_75t_L g888 ( 
.A(n_799),
.B(n_537),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_723),
.B(n_617),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_803),
.B(n_532),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_723),
.B(n_737),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_720),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_723),
.B(n_618),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_768),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_760),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_828),
.Y(n_896)
);

INVx1_ASAP7_75t_SL g897 ( 
.A(n_700),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_697),
.Y(n_898)
);

NOR3xp33_ASAP7_75t_SL g899 ( 
.A(n_684),
.B(n_641),
.C(n_322),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_808),
.Y(n_900)
);

NAND3xp33_ASAP7_75t_SL g901 ( 
.A(n_783),
.B(n_628),
.C(n_621),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_798),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_737),
.B(n_626),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_740),
.Y(n_904)
);

INVx1_ASAP7_75t_SL g905 ( 
.A(n_766),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_675),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_717),
.Y(n_907)
);

NOR2xp67_ASAP7_75t_L g908 ( 
.A(n_816),
.B(n_641),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_737),
.B(n_629),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_720),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_676),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_748),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_784),
.B(n_642),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_674),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_777),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_803),
.B(n_532),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_748),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_804),
.A2(n_743),
.B1(n_712),
.B2(n_784),
.Y(n_918)
);

CKINVDCx16_ASAP7_75t_R g919 ( 
.A(n_784),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_746),
.A2(n_613),
.B1(n_569),
.B2(n_573),
.Y(n_920)
);

OR2x6_ASAP7_75t_L g921 ( 
.A(n_708),
.B(n_569),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_663),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_710),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_670),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_764),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_731),
.B(n_645),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_726),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_775),
.B(n_647),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_746),
.A2(n_613),
.B1(n_573),
.B2(n_651),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_689),
.Y(n_930)
);

BUFx4f_ASAP7_75t_L g931 ( 
.A(n_731),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_764),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_731),
.B(n_649),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_775),
.B(n_652),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_790),
.Y(n_935)
);

AND3x1_ASAP7_75t_SL g936 ( 
.A(n_741),
.B(n_634),
.C(n_21),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_786),
.Y(n_937)
);

AOI22xp5_ASAP7_75t_L g938 ( 
.A1(n_739),
.A2(n_613),
.B1(n_651),
.B2(n_644),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_729),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_731),
.B(n_660),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_790),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_808),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_734),
.B(n_625),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_692),
.Y(n_944)
);

INVx3_ASAP7_75t_SL g945 ( 
.A(n_803),
.Y(n_945)
);

OR2x2_ASAP7_75t_L g946 ( 
.A(n_736),
.B(n_625),
.Y(n_946)
);

AOI22xp33_ASAP7_75t_L g947 ( 
.A1(n_744),
.A2(n_637),
.B1(n_627),
.B2(n_640),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_803),
.B(n_532),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_704),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_707),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_716),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_719),
.Y(n_952)
);

NAND2xp33_ASAP7_75t_L g953 ( 
.A(n_803),
.B(n_732),
.Y(n_953)
);

OR2x6_ASAP7_75t_L g954 ( 
.A(n_682),
.B(n_627),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_733),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_734),
.B(n_637),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_808),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_794),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_765),
.B(n_640),
.Y(n_959)
);

INVx5_ASAP7_75t_L g960 ( 
.A(n_732),
.Y(n_960)
);

OR2x6_ASAP7_75t_L g961 ( 
.A(n_709),
.B(n_744),
.Y(n_961)
);

AOI22x1_ASAP7_75t_L g962 ( 
.A1(n_823),
.A2(n_572),
.B1(n_651),
.B2(n_644),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_735),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_794),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_739),
.B(n_644),
.Y(n_965)
);

NAND3xp33_ASAP7_75t_L g966 ( 
.A(n_761),
.B(n_615),
.C(n_603),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_R g967 ( 
.A(n_802),
.B(n_572),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_757),
.Y(n_968)
);

BUFx2_ASAP7_75t_L g969 ( 
.A(n_781),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_758),
.B(n_615),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_SL g971 ( 
.A1(n_761),
.A2(n_335),
.B1(n_197),
.B2(n_178),
.Y(n_971)
);

NOR3xp33_ASAP7_75t_SL g972 ( 
.A(n_684),
.B(n_654),
.C(n_21),
.Y(n_972)
);

OAI22xp33_ASAP7_75t_L g973 ( 
.A1(n_667),
.A2(n_572),
.B1(n_615),
.B2(n_603),
.Y(n_973)
);

OR2x2_ASAP7_75t_L g974 ( 
.A(n_749),
.B(n_654),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_795),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_R g976 ( 
.A(n_802),
.B(n_603),
.Y(n_976)
);

NAND2xp33_ASAP7_75t_SL g977 ( 
.A(n_677),
.B(n_713),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_795),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_R g979 ( 
.A(n_693),
.B(n_603),
.Y(n_979)
);

INVxp67_ASAP7_75t_L g980 ( 
.A(n_785),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_801),
.Y(n_981)
);

OR2x6_ASAP7_75t_L g982 ( 
.A(n_751),
.B(n_782),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_721),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_801),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_722),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_679),
.A2(n_563),
.B(n_589),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_806),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_677),
.B(n_589),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_728),
.Y(n_989)
);

AND2x2_ASAP7_75t_SL g990 ( 
.A(n_693),
.B(n_563),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_817),
.B(n_589),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_818),
.B(n_589),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_673),
.B(n_536),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_694),
.B(n_536),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_829),
.Y(n_995)
);

OR2x6_ASAP7_75t_L g996 ( 
.A(n_724),
.B(n_536),
.Y(n_996)
);

BUFx12f_ASAP7_75t_L g997 ( 
.A(n_696),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_806),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_L g999 ( 
.A1(n_695),
.A2(n_536),
.B1(n_587),
.B2(n_197),
.Y(n_999)
);

NOR3xp33_ASAP7_75t_SL g1000 ( 
.A(n_691),
.B(n_20),
.C(n_22),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_824),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_824),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_750),
.B(n_587),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_826),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_753),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_826),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_754),
.B(n_587),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_827),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_713),
.B(n_23),
.Y(n_1009)
);

AND3x1_ASAP7_75t_SL g1010 ( 
.A(n_714),
.B(n_23),
.C(n_24),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_827),
.Y(n_1011)
);

BUFx12f_ASAP7_75t_L g1012 ( 
.A(n_714),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_831),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_831),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_762),
.Y(n_1015)
);

NOR2x1p5_ASAP7_75t_L g1016 ( 
.A(n_820),
.B(n_821),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_770),
.B(n_24),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_771),
.B(n_26),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_725),
.Y(n_1019)
);

NAND3xp33_ASAP7_75t_L g1020 ( 
.A(n_815),
.B(n_197),
.C(n_29),
.Y(n_1020)
);

NOR3xp33_ASAP7_75t_SL g1021 ( 
.A(n_691),
.B(n_26),
.C(n_29),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_725),
.A2(n_197),
.B1(n_32),
.B2(n_36),
.Y(n_1022)
);

INVx2_ASAP7_75t_SL g1023 ( 
.A(n_773),
.Y(n_1023)
);

BUFx2_ASAP7_75t_L g1024 ( 
.A(n_822),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_778),
.Y(n_1025)
);

OA22x2_ASAP7_75t_L g1026 ( 
.A1(n_844),
.A2(n_891),
.B1(n_989),
.B2(n_905),
.Y(n_1026)
);

A2O1A1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_840),
.A2(n_680),
.B(n_662),
.C(n_727),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_L g1028 ( 
.A1(n_986),
.A2(n_759),
.B(n_672),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_846),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_953),
.A2(n_686),
.B(n_688),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_962),
.A2(n_759),
.B(n_832),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_L g1032 ( 
.A1(n_872),
.A2(n_832),
.B(n_812),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_840),
.A2(n_800),
.B1(n_706),
.B2(n_730),
.Y(n_1033)
);

BUFx8_ASAP7_75t_L g1034 ( 
.A(n_877),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_856),
.A2(n_776),
.B1(n_747),
.B2(n_755),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_SL g1036 ( 
.A1(n_928),
.A2(n_699),
.B(n_701),
.Y(n_1036)
);

AOI21xp33_ASAP7_75t_L g1037 ( 
.A1(n_870),
.A2(n_680),
.B(n_793),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_872),
.A2(n_812),
.B(n_698),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_882),
.A2(n_916),
.B(n_890),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_847),
.A2(n_742),
.B(n_727),
.C(n_718),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_960),
.B(n_805),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_854),
.B(n_813),
.Y(n_1042)
);

INVx6_ASAP7_75t_L g1043 ( 
.A(n_838),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_888),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_839),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1005),
.B(n_669),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_843),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_884),
.A2(n_742),
.B(n_796),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_882),
.A2(n_767),
.B(n_819),
.Y(n_1049)
);

OA22x2_ASAP7_75t_L g1050 ( 
.A1(n_891),
.A2(n_867),
.B1(n_888),
.B2(n_879),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_852),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_846),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_L g1053 ( 
.A1(n_890),
.A2(n_767),
.B(n_789),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1015),
.B(n_825),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_885),
.A2(n_810),
.B(n_788),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_916),
.A2(n_797),
.B(n_809),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_1025),
.B(n_30),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_L g1058 ( 
.A1(n_948),
.A2(n_197),
.B(n_156),
.Y(n_1058)
);

O2A1O1Ixp5_ASAP7_75t_L g1059 ( 
.A1(n_977),
.A2(n_32),
.B(n_38),
.C(n_39),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_856),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_919),
.B(n_40),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_876),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_965),
.A2(n_75),
.B(n_152),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_881),
.A2(n_153),
.B(n_149),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_948),
.A2(n_140),
.B(n_134),
.Y(n_1065)
);

NAND2x1p5_ASAP7_75t_L g1066 ( 
.A(n_931),
.B(n_846),
.Y(n_1066)
);

AO31x2_ASAP7_75t_L g1067 ( 
.A1(n_943),
.A2(n_42),
.A3(n_43),
.B(n_45),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_873),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_861),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_860),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_841),
.B(n_46),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_876),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_1072)
);

OR2x2_ASAP7_75t_L g1073 ( 
.A(n_836),
.B(n_47),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_848),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_848),
.Y(n_1075)
);

AOI21x1_ASAP7_75t_L g1076 ( 
.A1(n_988),
.A2(n_76),
.B(n_123),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_841),
.B(n_49),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_1000),
.A2(n_52),
.B(n_53),
.C(n_57),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_858),
.A2(n_52),
.B(n_61),
.C(n_64),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_994),
.A2(n_988),
.B(n_993),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1023),
.B(n_61),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_939),
.B(n_65),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_881),
.A2(n_91),
.B(n_122),
.Y(n_1083)
);

NOR2xp67_ASAP7_75t_L g1084 ( 
.A(n_833),
.B(n_85),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_915),
.B(n_68),
.Y(n_1085)
);

AO31x2_ASAP7_75t_L g1086 ( 
.A1(n_956),
.A2(n_70),
.A3(n_71),
.B(n_73),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_999),
.A2(n_82),
.B(n_98),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_896),
.B(n_105),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_999),
.A2(n_108),
.B(n_116),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_960),
.B(n_129),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_918),
.A2(n_837),
.B1(n_862),
.B2(n_934),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_896),
.B(n_914),
.Y(n_1092)
);

NOR2x1_ASAP7_75t_L g1093 ( 
.A(n_888),
.B(n_894),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_871),
.A2(n_938),
.B(n_991),
.Y(n_1094)
);

INVx1_ASAP7_75t_SL g1095 ( 
.A(n_897),
.Y(n_1095)
);

AOI21xp33_ASAP7_75t_L g1096 ( 
.A1(n_855),
.A2(n_961),
.B(n_893),
.Y(n_1096)
);

AOI211x1_ASAP7_75t_L g1097 ( 
.A1(n_875),
.A2(n_902),
.B(n_901),
.C(n_1018),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_991),
.A2(n_992),
.B(n_929),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_977),
.A2(n_990),
.B(n_1007),
.Y(n_1099)
);

AOI21xp33_ASAP7_75t_L g1100 ( 
.A1(n_855),
.A2(n_961),
.B(n_889),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_891),
.B(n_913),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_918),
.A2(n_1019),
.B1(n_864),
.B2(n_931),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_838),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_913),
.B(n_1024),
.Y(n_1104)
);

AO31x2_ASAP7_75t_L g1105 ( 
.A1(n_992),
.A2(n_910),
.A3(n_958),
.B(n_912),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_859),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_1003),
.A2(n_932),
.B(n_935),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_SL g1108 ( 
.A1(n_1022),
.A2(n_1017),
.B(n_970),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_851),
.A2(n_932),
.B(n_964),
.Y(n_1109)
);

CKINVDCx11_ASAP7_75t_R g1110 ( 
.A(n_878),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_851),
.A2(n_964),
.B(n_886),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_990),
.A2(n_973),
.B(n_960),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_973),
.A2(n_960),
.B(n_1019),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_853),
.B(n_898),
.Y(n_1114)
);

AOI21x1_ASAP7_75t_L g1115 ( 
.A1(n_966),
.A2(n_954),
.B(n_978),
.Y(n_1115)
);

O2A1O1Ixp5_ASAP7_75t_L g1116 ( 
.A1(n_1020),
.A2(n_942),
.B(n_957),
.C(n_1009),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_980),
.A2(n_959),
.B(n_954),
.Y(n_1117)
);

AOI21x1_ASAP7_75t_L g1118 ( 
.A1(n_954),
.A2(n_998),
.B(n_1006),
.Y(n_1118)
);

BUFx8_ASAP7_75t_L g1119 ( 
.A(n_877),
.Y(n_1119)
);

AOI21xp33_ASAP7_75t_L g1120 ( 
.A1(n_961),
.A2(n_903),
.B(n_909),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_922),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_857),
.A2(n_917),
.B(n_958),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_850),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_924),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_853),
.B(n_898),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_857),
.A2(n_917),
.B(n_910),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_868),
.A2(n_912),
.B(n_892),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_907),
.B(n_845),
.Y(n_1128)
);

AO32x2_ASAP7_75t_L g1129 ( 
.A1(n_1012),
.A2(n_1010),
.A3(n_899),
.B1(n_972),
.B2(n_1021),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_868),
.A2(n_975),
.B(n_892),
.Y(n_1130)
);

NOR4xp25_ASAP7_75t_L g1131 ( 
.A(n_930),
.B(n_944),
.C(n_963),
.D(n_951),
.Y(n_1131)
);

OAI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_920),
.A2(n_911),
.B(n_906),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_853),
.B(n_923),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_880),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_949),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_923),
.B(n_952),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_880),
.A2(n_925),
.B(n_935),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_845),
.B(n_849),
.Y(n_1138)
);

INVxp67_ASAP7_75t_L g1139 ( 
.A(n_904),
.Y(n_1139)
);

NAND3xp33_ASAP7_75t_L g1140 ( 
.A(n_927),
.B(n_971),
.C(n_835),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_952),
.B(n_969),
.Y(n_1141)
);

A2O1A1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_1009),
.A2(n_959),
.B(n_974),
.C(n_1016),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_877),
.B(n_863),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_959),
.A2(n_926),
.B(n_957),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_883),
.A2(n_941),
.B(n_1011),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_883),
.A2(n_941),
.B(n_1011),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_926),
.A2(n_942),
.B(n_940),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_886),
.A2(n_925),
.B(n_887),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_850),
.B(n_863),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_887),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_975),
.Y(n_1151)
);

INVx4_ASAP7_75t_L g1152 ( 
.A(n_874),
.Y(n_1152)
);

AOI21xp33_ASAP7_75t_L g1153 ( 
.A1(n_946),
.A2(n_985),
.B(n_968),
.Y(n_1153)
);

INVx6_ASAP7_75t_L g1154 ( 
.A(n_878),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_SL g1155 ( 
.A1(n_950),
.A2(n_955),
.B(n_1001),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1001),
.A2(n_947),
.B(n_1013),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_947),
.A2(n_1014),
.B(n_1008),
.Y(n_1157)
);

NOR3xp33_ASAP7_75t_L g1158 ( 
.A(n_937),
.B(n_908),
.C(n_895),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_985),
.Y(n_1159)
);

HB1xp67_ASAP7_75t_L g1160 ( 
.A(n_983),
.Y(n_1160)
);

OR2x2_ASAP7_75t_L g1161 ( 
.A(n_878),
.B(n_921),
.Y(n_1161)
);

NOR4xp25_ASAP7_75t_L g1162 ( 
.A(n_1010),
.B(n_936),
.C(n_984),
.D(n_981),
.Y(n_1162)
);

AOI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_933),
.A2(n_940),
.B1(n_997),
.B2(n_926),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_983),
.B(n_933),
.Y(n_1164)
);

AOI221x1_ASAP7_75t_L g1165 ( 
.A1(n_1009),
.A2(n_983),
.B1(n_1002),
.B2(n_1004),
.C(n_900),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_983),
.B(n_987),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_846),
.B(n_866),
.Y(n_1167)
);

INVx4_ASAP7_75t_L g1168 ( 
.A(n_874),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_987),
.B(n_921),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_834),
.A2(n_842),
.B(n_865),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_894),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_869),
.A2(n_866),
.B(n_874),
.C(n_900),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_834),
.A2(n_945),
.B(n_1012),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_945),
.A2(n_976),
.B(n_979),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_921),
.B(n_869),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_979),
.A2(n_874),
.B(n_967),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_967),
.A2(n_900),
.B(n_976),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_900),
.A2(n_982),
.B(n_996),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_982),
.A2(n_996),
.B(n_866),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_996),
.A2(n_982),
.B(n_866),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_995),
.B(n_936),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_997),
.B(n_919),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_953),
.A2(n_884),
.B(n_840),
.Y(n_1183)
);

NAND2x1p5_ASAP7_75t_L g1184 ( 
.A(n_931),
.B(n_846),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_840),
.A2(n_665),
.B(n_885),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_840),
.B(n_844),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_854),
.B(n_665),
.Y(n_1187)
);

AOI221xp5_ASAP7_75t_L g1188 ( 
.A1(n_1091),
.A2(n_1085),
.B1(n_1186),
.B2(n_1187),
.C(n_1162),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1026),
.A2(n_1050),
.B1(n_1046),
.B2(n_1186),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1068),
.B(n_1139),
.Y(n_1190)
);

NAND3xp33_ASAP7_75t_L g1191 ( 
.A(n_1078),
.B(n_1097),
.C(n_1185),
.Y(n_1191)
);

AO21x2_ASAP7_75t_L g1192 ( 
.A1(n_1036),
.A2(n_1037),
.B(n_1094),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1031),
.A2(n_1028),
.B(n_1107),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1142),
.A2(n_1085),
.B1(n_1078),
.B2(n_1102),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1045),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1123),
.B(n_1149),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1026),
.A2(n_1050),
.B1(n_1120),
.B2(n_1140),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1074),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1031),
.A2(n_1028),
.B(n_1107),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1092),
.B(n_1136),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1074),
.Y(n_1201)
);

BUFx2_ASAP7_75t_L g1202 ( 
.A(n_1160),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1096),
.A2(n_1100),
.B1(n_1182),
.B2(n_1153),
.Y(n_1203)
);

AOI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1099),
.A2(n_1115),
.B(n_1112),
.Y(n_1204)
);

NOR2xp67_ASAP7_75t_SL g1205 ( 
.A(n_1183),
.B(n_1064),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1047),
.Y(n_1206)
);

BUFx2_ASAP7_75t_L g1207 ( 
.A(n_1160),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_1174),
.Y(n_1208)
);

INVxp67_ASAP7_75t_L g1209 ( 
.A(n_1095),
.Y(n_1209)
);

AOI21xp33_ASAP7_75t_SL g1210 ( 
.A1(n_1068),
.A2(n_1070),
.B(n_1175),
.Y(n_1210)
);

OR2x6_ASAP7_75t_L g1211 ( 
.A(n_1174),
.B(n_1176),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1109),
.Y(n_1212)
);

INVx4_ASAP7_75t_L g1213 ( 
.A(n_1152),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1038),
.A2(n_1039),
.B(n_1032),
.Y(n_1214)
);

OA21x2_ASAP7_75t_L g1215 ( 
.A1(n_1080),
.A2(n_1038),
.B(n_1098),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_1043),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_1043),
.Y(n_1217)
);

AO21x2_ASAP7_75t_L g1218 ( 
.A1(n_1108),
.A2(n_1048),
.B(n_1118),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_1104),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1032),
.A2(n_1053),
.B(n_1058),
.Y(n_1220)
);

OR2x2_ASAP7_75t_L g1221 ( 
.A(n_1114),
.B(n_1125),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1055),
.A2(n_1027),
.B(n_1113),
.Y(n_1222)
);

AOI221xp5_ASAP7_75t_L g1223 ( 
.A1(n_1131),
.A2(n_1079),
.B1(n_1033),
.B2(n_1035),
.C(n_1060),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_1152),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_SL g1225 ( 
.A1(n_1155),
.A2(n_1144),
.B(n_1132),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1142),
.A2(n_1116),
.B(n_1117),
.C(n_1027),
.Y(n_1226)
);

AO21x2_ASAP7_75t_L g1227 ( 
.A1(n_1156),
.A2(n_1157),
.B(n_1030),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1133),
.A2(n_1077),
.B1(n_1071),
.B2(n_1057),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_1123),
.B(n_1103),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1101),
.B(n_1051),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1141),
.B(n_1128),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1053),
.A2(n_1058),
.B(n_1156),
.Y(n_1232)
);

BUFx12f_ASAP7_75t_L g1233 ( 
.A(n_1110),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1069),
.B(n_1129),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1157),
.A2(n_1065),
.B(n_1087),
.Y(n_1235)
);

AO21x2_ASAP7_75t_L g1236 ( 
.A1(n_1109),
.A2(n_1146),
.B(n_1122),
.Y(n_1236)
);

OAI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1040),
.A2(n_1081),
.B(n_1082),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1075),
.Y(n_1238)
);

AND3x2_ASAP7_75t_L g1239 ( 
.A(n_1138),
.B(n_1106),
.C(n_1158),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_1070),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1075),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1134),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1111),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1159),
.Y(n_1244)
);

AO21x2_ASAP7_75t_L g1245 ( 
.A1(n_1111),
.A2(n_1126),
.B(n_1130),
.Y(n_1245)
);

AO31x2_ASAP7_75t_L g1246 ( 
.A1(n_1165),
.A2(n_1134),
.A3(n_1151),
.B(n_1150),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1083),
.A2(n_1041),
.B(n_1063),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1147),
.A2(n_1163),
.B1(n_1154),
.B2(n_1044),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1122),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1129),
.B(n_1143),
.Y(n_1250)
);

CKINVDCx6p67_ASAP7_75t_R g1251 ( 
.A(n_1110),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1150),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1151),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1159),
.B(n_1164),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1166),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1126),
.Y(n_1256)
);

CKINVDCx20_ASAP7_75t_R g1257 ( 
.A(n_1034),
.Y(n_1257)
);

INVx1_ASAP7_75t_SL g1258 ( 
.A(n_1043),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1168),
.Y(n_1259)
);

INVx4_ASAP7_75t_L g1260 ( 
.A(n_1168),
.Y(n_1260)
);

AO21x2_ASAP7_75t_L g1261 ( 
.A1(n_1127),
.A2(n_1145),
.B(n_1148),
.Y(n_1261)
);

OR2x6_ASAP7_75t_L g1262 ( 
.A(n_1177),
.B(n_1178),
.Y(n_1262)
);

O2A1O1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1062),
.A2(n_1072),
.B(n_1059),
.C(n_1073),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1034),
.A2(n_1119),
.B1(n_1042),
.B2(n_1054),
.Y(n_1264)
);

CKINVDCx6p67_ASAP7_75t_R g1265 ( 
.A(n_1103),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1041),
.A2(n_1173),
.B(n_1056),
.Y(n_1266)
);

OAI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1173),
.A2(n_1056),
.B(n_1088),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1121),
.Y(n_1268)
);

INVx8_ASAP7_75t_L g1269 ( 
.A(n_1167),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1154),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1089),
.A2(n_1130),
.B(n_1137),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1154),
.A2(n_1161),
.B1(n_1169),
.B2(n_1172),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_1171),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_SL g1274 ( 
.A(n_1034),
.B(n_1119),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1172),
.A2(n_1124),
.B1(n_1135),
.B2(n_1093),
.Y(n_1275)
);

INVx4_ASAP7_75t_L g1276 ( 
.A(n_1167),
.Y(n_1276)
);

AO21x2_ASAP7_75t_L g1277 ( 
.A1(n_1127),
.A2(n_1137),
.B(n_1148),
.Y(n_1277)
);

OAI222xp33_ASAP7_75t_L g1278 ( 
.A1(n_1061),
.A2(n_1181),
.B1(n_1184),
.B2(n_1066),
.C1(n_1090),
.C2(n_1179),
.Y(n_1278)
);

AO31x2_ASAP7_75t_L g1279 ( 
.A1(n_1105),
.A2(n_1086),
.A3(n_1067),
.B(n_1145),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1146),
.A2(n_1076),
.B(n_1170),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1129),
.B(n_1184),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1067),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1066),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1170),
.A2(n_1049),
.B(n_1180),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1067),
.Y(n_1285)
);

OA21x2_ASAP7_75t_L g1286 ( 
.A1(n_1049),
.A2(n_1090),
.B(n_1180),
.Y(n_1286)
);

INVx4_ASAP7_75t_L g1287 ( 
.A(n_1167),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1029),
.B(n_1052),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1067),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1181),
.A2(n_1029),
.B1(n_1052),
.B2(n_1084),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1129),
.B(n_1181),
.Y(n_1291)
);

A2O1A1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1052),
.A2(n_1086),
.B(n_1119),
.C(n_1105),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1105),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_1105),
.B(n_1086),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1086),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1187),
.B(n_1005),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1074),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_1110),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1109),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1095),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1031),
.A2(n_1028),
.B(n_1107),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1068),
.B(n_551),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1109),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1183),
.A2(n_953),
.B(n_1185),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1074),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_SL g1306 ( 
.A1(n_1099),
.A2(n_1036),
.B(n_1183),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1031),
.A2(n_1028),
.B(n_1107),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_1123),
.B(n_1149),
.Y(n_1308)
);

OAI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1050),
.A2(n_791),
.B1(n_624),
.B2(n_844),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1074),
.Y(n_1310)
);

INVx4_ASAP7_75t_L g1311 ( 
.A(n_1152),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1185),
.B(n_844),
.Y(n_1312)
);

INVx1_ASAP7_75t_SL g1313 ( 
.A(n_1095),
.Y(n_1313)
);

AND2x4_ASAP7_75t_SL g1314 ( 
.A(n_1128),
.B(n_878),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1074),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1183),
.A2(n_953),
.B(n_1185),
.Y(n_1316)
);

INVx4_ASAP7_75t_L g1317 ( 
.A(n_1152),
.Y(n_1317)
);

INVxp67_ASAP7_75t_SL g1318 ( 
.A(n_1174),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_R g1319 ( 
.A1(n_1060),
.A2(n_1072),
.B(n_1062),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1045),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1123),
.B(n_1149),
.Y(n_1321)
);

AO21x2_ASAP7_75t_L g1322 ( 
.A1(n_1036),
.A2(n_1037),
.B(n_1094),
.Y(n_1322)
);

INVx1_ASAP7_75t_SL g1323 ( 
.A(n_1095),
.Y(n_1323)
);

AOI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1099),
.A2(n_1115),
.B(n_1186),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1109),
.Y(n_1325)
);

INVx3_ASAP7_75t_L g1326 ( 
.A(n_1152),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1045),
.Y(n_1327)
);

CKINVDCx20_ASAP7_75t_R g1328 ( 
.A(n_1110),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1045),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1026),
.A2(n_461),
.B1(n_624),
.B2(n_345),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1185),
.B(n_844),
.Y(n_1331)
);

INVx1_ASAP7_75t_SL g1332 ( 
.A(n_1095),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1160),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1123),
.B(n_1149),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1031),
.A2(n_1028),
.B(n_1107),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_1068),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1026),
.A2(n_461),
.B1(n_579),
.B2(n_624),
.Y(n_1337)
);

NOR2xp67_ASAP7_75t_L g1338 ( 
.A(n_1139),
.B(n_561),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1185),
.A2(n_665),
.B(n_840),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1160),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1031),
.A2(n_1028),
.B(n_1107),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_1068),
.Y(n_1342)
);

AO21x2_ASAP7_75t_L g1343 ( 
.A1(n_1036),
.A2(n_1037),
.B(n_1094),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1031),
.A2(n_1028),
.B(n_1107),
.Y(n_1344)
);

OR2x6_ASAP7_75t_L g1345 ( 
.A(n_1174),
.B(n_1176),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1045),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1187),
.B(n_1005),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1031),
.A2(n_1028),
.B(n_1107),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1031),
.A2(n_1028),
.B(n_1107),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1043),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1109),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1045),
.Y(n_1352)
);

OAI21xp33_ASAP7_75t_SL g1353 ( 
.A1(n_1185),
.A2(n_844),
.B(n_690),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1312),
.B(n_1331),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1254),
.B(n_1244),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1195),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1276),
.B(n_1287),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1200),
.B(n_1296),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1206),
.Y(n_1359)
);

CKINVDCx12_ASAP7_75t_R g1360 ( 
.A(n_1221),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1336),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1312),
.B(n_1331),
.Y(n_1362)
);

NOR3xp33_ASAP7_75t_SL g1363 ( 
.A(n_1240),
.B(n_1342),
.C(n_1336),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1246),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1319),
.A2(n_1188),
.B1(n_1194),
.B2(n_1337),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1234),
.B(n_1250),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1268),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1193),
.A2(n_1301),
.B(n_1199),
.Y(n_1368)
);

NAND2x1_ASAP7_75t_L g1369 ( 
.A(n_1225),
.B(n_1306),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1191),
.A2(n_1223),
.B1(n_1347),
.B2(n_1339),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1330),
.A2(n_1309),
.B1(n_1189),
.B2(n_1197),
.Y(n_1371)
);

BUFx12f_ASAP7_75t_L g1372 ( 
.A(n_1240),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1203),
.A2(n_1228),
.B1(n_1264),
.B2(n_1291),
.Y(n_1373)
);

BUFx10_ASAP7_75t_L g1374 ( 
.A(n_1302),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1246),
.Y(n_1375)
);

INVxp33_ASAP7_75t_SL g1376 ( 
.A(n_1342),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1246),
.Y(n_1377)
);

INVx4_ASAP7_75t_R g1378 ( 
.A(n_1216),
.Y(n_1378)
);

AND2x6_ASAP7_75t_L g1379 ( 
.A(n_1281),
.B(n_1208),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_SL g1380 ( 
.A1(n_1237),
.A2(n_1290),
.B(n_1263),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_1229),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1291),
.A2(n_1226),
.B1(n_1222),
.B2(n_1273),
.Y(n_1382)
);

CKINVDCx20_ASAP7_75t_R g1383 ( 
.A(n_1298),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1234),
.B(n_1250),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1246),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1353),
.A2(n_1248),
.B1(n_1281),
.B2(n_1300),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1230),
.B(n_1221),
.Y(n_1387)
);

INVx2_ASAP7_75t_SL g1388 ( 
.A(n_1196),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1273),
.A2(n_1251),
.B1(n_1298),
.B2(n_1328),
.Y(n_1389)
);

OAI221xp5_ASAP7_75t_L g1390 ( 
.A1(n_1338),
.A2(n_1247),
.B1(n_1231),
.B2(n_1274),
.C(n_1267),
.Y(n_1390)
);

INVx1_ASAP7_75t_SL g1391 ( 
.A(n_1313),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_SL g1392 ( 
.A1(n_1275),
.A2(n_1272),
.B1(n_1257),
.B2(n_1233),
.Y(n_1392)
);

INVx3_ASAP7_75t_L g1393 ( 
.A(n_1208),
.Y(n_1393)
);

OAI221xp5_ASAP7_75t_L g1394 ( 
.A1(n_1209),
.A2(n_1190),
.B1(n_1332),
.B2(n_1323),
.C(n_1352),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1230),
.A2(n_1255),
.B1(n_1294),
.B2(n_1219),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1233),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1320),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1202),
.B(n_1207),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1327),
.Y(n_1399)
);

INVx4_ASAP7_75t_L g1400 ( 
.A(n_1265),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1329),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1246),
.Y(n_1402)
);

AOI221xp5_ASAP7_75t_L g1403 ( 
.A1(n_1346),
.A2(n_1295),
.B1(n_1282),
.B2(n_1285),
.C(n_1289),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1328),
.A2(n_1316),
.B1(n_1304),
.B2(n_1257),
.Y(n_1404)
);

CKINVDCx11_ASAP7_75t_R g1405 ( 
.A(n_1265),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1198),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_1269),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1255),
.A2(n_1294),
.B1(n_1293),
.B2(n_1196),
.Y(n_1408)
);

O2A1O1Ixp5_ASAP7_75t_L g1409 ( 
.A1(n_1205),
.A2(n_1324),
.B(n_1266),
.C(n_1318),
.Y(n_1409)
);

NAND2xp33_ASAP7_75t_SL g1410 ( 
.A(n_1205),
.B(n_1213),
.Y(n_1410)
);

NAND2xp33_ASAP7_75t_R g1411 ( 
.A(n_1239),
.B(n_1229),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1201),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1308),
.B(n_1321),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1293),
.A2(n_1321),
.B1(n_1308),
.B2(n_1334),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1201),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1334),
.A2(n_1305),
.B1(n_1253),
.B2(n_1252),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_1269),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1269),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1216),
.B(n_1350),
.Y(n_1419)
);

AOI221xp5_ASAP7_75t_L g1420 ( 
.A1(n_1210),
.A2(n_1278),
.B1(n_1292),
.B2(n_1343),
.C(n_1192),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1238),
.Y(n_1421)
);

OR2x6_ASAP7_75t_L g1422 ( 
.A(n_1262),
.B(n_1211),
.Y(n_1422)
);

BUFx12f_ASAP7_75t_L g1423 ( 
.A(n_1217),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1241),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1350),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1258),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1241),
.Y(n_1427)
);

NAND3xp33_ASAP7_75t_SL g1428 ( 
.A(n_1202),
.B(n_1340),
.C(n_1333),
.Y(n_1428)
);

INVx3_ASAP7_75t_L g1429 ( 
.A(n_1208),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1314),
.A2(n_1217),
.B1(n_1276),
.B2(n_1287),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1242),
.Y(n_1431)
);

AOI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1314),
.A2(n_1270),
.B1(n_1287),
.B2(n_1276),
.Y(n_1432)
);

INVx3_ASAP7_75t_L g1433 ( 
.A(n_1208),
.Y(n_1433)
);

BUFx6f_ASAP7_75t_L g1434 ( 
.A(n_1269),
.Y(n_1434)
);

INVx4_ASAP7_75t_L g1435 ( 
.A(n_1288),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1288),
.B(n_1270),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1242),
.Y(n_1437)
);

AOI221xp5_ASAP7_75t_L g1438 ( 
.A1(n_1192),
.A2(n_1343),
.B1(n_1322),
.B2(n_1225),
.C(n_1340),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1252),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1253),
.A2(n_1310),
.B1(n_1297),
.B2(n_1305),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1297),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1310),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1315),
.A2(n_1192),
.B1(n_1343),
.B2(n_1322),
.Y(n_1443)
);

NAND2xp33_ASAP7_75t_R g1444 ( 
.A(n_1288),
.B(n_1286),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1279),
.B(n_1322),
.Y(n_1445)
);

CKINVDCx20_ASAP7_75t_R g1446 ( 
.A(n_1283),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1315),
.A2(n_1283),
.B1(n_1262),
.B2(n_1286),
.Y(n_1447)
);

NOR2xp67_ASAP7_75t_SL g1448 ( 
.A(n_1213),
.B(n_1311),
.Y(n_1448)
);

CKINVDCx11_ASAP7_75t_R g1449 ( 
.A(n_1208),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_1262),
.Y(n_1450)
);

AO31x2_ASAP7_75t_L g1451 ( 
.A1(n_1212),
.A2(n_1351),
.A3(n_1325),
.B(n_1243),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_SL g1452 ( 
.A(n_1224),
.B(n_1259),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1236),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_SL g1454 ( 
.A1(n_1213),
.A2(n_1311),
.B1(n_1260),
.B2(n_1317),
.Y(n_1454)
);

AOI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1218),
.A2(n_1262),
.B1(n_1286),
.B2(n_1211),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_1260),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1279),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1224),
.A2(n_1326),
.B1(n_1259),
.B2(n_1260),
.Y(n_1458)
);

INVx3_ASAP7_75t_L g1459 ( 
.A(n_1311),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1218),
.A2(n_1211),
.B1(n_1345),
.B2(n_1325),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1236),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1193),
.A2(n_1199),
.B(n_1301),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1236),
.Y(n_1463)
);

NOR2xp67_ASAP7_75t_L g1464 ( 
.A(n_1317),
.B(n_1326),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1279),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1279),
.B(n_1215),
.Y(n_1466)
);

A2O1A1Ixp33_ASAP7_75t_SL g1467 ( 
.A1(n_1256),
.A2(n_1351),
.B(n_1303),
.C(n_1212),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1279),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1211),
.A2(n_1345),
.B1(n_1303),
.B2(n_1299),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1243),
.Y(n_1470)
);

INVxp67_ASAP7_75t_SL g1471 ( 
.A(n_1215),
.Y(n_1471)
);

OAI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1214),
.A2(n_1349),
.B(n_1348),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1204),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1345),
.B(n_1317),
.Y(n_1474)
);

CKINVDCx6p67_ASAP7_75t_R g1475 ( 
.A(n_1204),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1249),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1284),
.B(n_1299),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1284),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_SL g1479 ( 
.A1(n_1235),
.A2(n_1227),
.B1(n_1232),
.B2(n_1220),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1227),
.A2(n_1277),
.B1(n_1261),
.B2(n_1245),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1245),
.A2(n_1261),
.B1(n_1277),
.B2(n_1271),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1245),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1261),
.Y(n_1483)
);

BUFx8_ASAP7_75t_L g1484 ( 
.A(n_1280),
.Y(n_1484)
);

INVx4_ASAP7_75t_L g1485 ( 
.A(n_1277),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1271),
.A2(n_1232),
.B1(n_1280),
.B2(n_1307),
.Y(n_1486)
);

INVx3_ASAP7_75t_L g1487 ( 
.A(n_1335),
.Y(n_1487)
);

AO221x2_ASAP7_75t_L g1488 ( 
.A1(n_1341),
.A2(n_1194),
.B1(n_1191),
.B2(n_1309),
.C(n_1353),
.Y(n_1488)
);

INVx4_ASAP7_75t_L g1489 ( 
.A(n_1344),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1195),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1195),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1246),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1312),
.B(n_1331),
.Y(n_1493)
);

INVx4_ASAP7_75t_L g1494 ( 
.A(n_1265),
.Y(n_1494)
);

AND2x2_ASAP7_75t_SL g1495 ( 
.A(n_1337),
.B(n_931),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1246),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1244),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1246),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1410),
.A2(n_1380),
.B(n_1365),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1354),
.B(n_1362),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1356),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1371),
.A2(n_1370),
.B1(n_1488),
.B2(n_1495),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1400),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1359),
.Y(n_1504)
);

NAND3xp33_ASAP7_75t_L g1505 ( 
.A(n_1438),
.B(n_1420),
.C(n_1373),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1392),
.A2(n_1404),
.B1(n_1382),
.B2(n_1386),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1367),
.Y(n_1507)
);

AOI222xp33_ASAP7_75t_L g1508 ( 
.A1(n_1495),
.A2(n_1358),
.B1(n_1493),
.B2(n_1354),
.C1(n_1362),
.C2(n_1394),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1397),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1493),
.B(n_1387),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1426),
.A2(n_1425),
.B1(n_1400),
.B2(n_1494),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1366),
.B(n_1384),
.Y(n_1512)
);

INVx8_ASAP7_75t_L g1513 ( 
.A(n_1423),
.Y(n_1513)
);

OAI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1355),
.A2(n_1413),
.B1(n_1411),
.B2(n_1383),
.Y(n_1514)
);

BUFx3_ASAP7_75t_L g1515 ( 
.A(n_1423),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1366),
.B(n_1384),
.Y(n_1516)
);

OA21x2_ASAP7_75t_L g1517 ( 
.A1(n_1472),
.A2(n_1462),
.B(n_1368),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1398),
.B(n_1381),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1497),
.B(n_1398),
.Y(n_1519)
);

AOI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1488),
.A2(n_1369),
.B(n_1409),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1399),
.A2(n_1401),
.B1(n_1491),
.B2(n_1490),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1390),
.B(n_1400),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1391),
.A2(n_1445),
.B1(n_1395),
.B2(n_1446),
.Y(n_1523)
);

OAI221xp5_ASAP7_75t_L g1524 ( 
.A1(n_1443),
.A2(n_1480),
.B1(n_1460),
.B2(n_1419),
.C(n_1426),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1445),
.A2(n_1446),
.B1(n_1405),
.B2(n_1383),
.Y(n_1525)
);

AOI222xp33_ASAP7_75t_L g1526 ( 
.A1(n_1406),
.A2(n_1412),
.B1(n_1427),
.B2(n_1441),
.C1(n_1415),
.C2(n_1442),
.Y(n_1526)
);

AOI221xp5_ASAP7_75t_L g1527 ( 
.A1(n_1466),
.A2(n_1403),
.B1(n_1457),
.B2(n_1468),
.C(n_1465),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1363),
.Y(n_1528)
);

OA21x2_ASAP7_75t_L g1529 ( 
.A1(n_1481),
.A2(n_1486),
.B(n_1471),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1405),
.A2(n_1374),
.B1(n_1416),
.B2(n_1372),
.Y(n_1530)
);

OAI221xp5_ASAP7_75t_L g1531 ( 
.A1(n_1389),
.A2(n_1432),
.B1(n_1455),
.B2(n_1469),
.C(n_1494),
.Y(n_1531)
);

OAI22xp33_ASAP7_75t_SL g1532 ( 
.A1(n_1450),
.A2(n_1494),
.B1(n_1388),
.B2(n_1422),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_SL g1533 ( 
.A1(n_1379),
.A2(n_1484),
.B1(n_1466),
.B2(n_1430),
.Y(n_1533)
);

OAI221xp5_ASAP7_75t_L g1534 ( 
.A1(n_1414),
.A2(n_1479),
.B1(n_1447),
.B2(n_1396),
.C(n_1418),
.Y(n_1534)
);

AOI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1360),
.A2(n_1436),
.B1(n_1418),
.B2(n_1425),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1436),
.B(n_1435),
.Y(n_1536)
);

OAI221xp5_ASAP7_75t_L g1537 ( 
.A1(n_1396),
.A2(n_1485),
.B1(n_1473),
.B2(n_1408),
.C(n_1463),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1436),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_SL g1539 ( 
.A1(n_1376),
.A2(n_1372),
.B1(n_1361),
.B2(n_1360),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1376),
.A2(n_1361),
.B1(n_1357),
.B2(n_1464),
.Y(n_1540)
);

AOI221xp5_ASAP7_75t_L g1541 ( 
.A1(n_1428),
.A2(n_1461),
.B1(n_1483),
.B2(n_1453),
.C(n_1482),
.Y(n_1541)
);

AOI221xp5_ASAP7_75t_L g1542 ( 
.A1(n_1482),
.A2(n_1476),
.B1(n_1470),
.B2(n_1440),
.C(n_1485),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1357),
.A2(n_1454),
.B1(n_1459),
.B2(n_1452),
.Y(n_1543)
);

OR2x6_ASAP7_75t_L g1544 ( 
.A(n_1422),
.B(n_1474),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1459),
.A2(n_1456),
.B1(n_1458),
.B2(n_1417),
.Y(n_1545)
);

AOI221xp5_ASAP7_75t_L g1546 ( 
.A1(n_1364),
.A2(n_1498),
.B1(n_1375),
.B2(n_1377),
.C(n_1496),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1374),
.A2(n_1437),
.B1(n_1439),
.B2(n_1421),
.Y(n_1547)
);

OAI332xp33_ASAP7_75t_L g1548 ( 
.A1(n_1374),
.A2(n_1478),
.A3(n_1477),
.B1(n_1437),
.B2(n_1431),
.B3(n_1424),
.C1(n_1385),
.C2(n_1498),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1456),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1424),
.A2(n_1431),
.B1(n_1434),
.B2(n_1417),
.Y(n_1550)
);

AOI221xp5_ASAP7_75t_L g1551 ( 
.A1(n_1364),
.A2(n_1375),
.B1(n_1377),
.B2(n_1492),
.C(n_1496),
.Y(n_1551)
);

INVx2_ASAP7_75t_SL g1552 ( 
.A(n_1378),
.Y(n_1552)
);

OAI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1407),
.A2(n_1417),
.B1(n_1434),
.B2(n_1456),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1407),
.A2(n_1434),
.B1(n_1417),
.B2(n_1379),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1379),
.A2(n_1385),
.B1(n_1492),
.B2(n_1402),
.Y(n_1555)
);

OAI211xp5_ASAP7_75t_L g1556 ( 
.A1(n_1449),
.A2(n_1489),
.B(n_1487),
.C(n_1459),
.Y(n_1556)
);

AOI221xp5_ASAP7_75t_L g1557 ( 
.A1(n_1402),
.A2(n_1467),
.B1(n_1429),
.B2(n_1433),
.C(n_1393),
.Y(n_1557)
);

AOI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1444),
.A2(n_1449),
.B1(n_1448),
.B2(n_1475),
.Y(n_1558)
);

OAI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1475),
.A2(n_1393),
.B1(n_1429),
.B2(n_1433),
.Y(n_1559)
);

OAI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1393),
.A2(n_1429),
.B1(n_1433),
.B2(n_1489),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1484),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1451),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1451),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1451),
.B(n_1487),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1354),
.B(n_1362),
.Y(n_1565)
);

INVx3_ASAP7_75t_L g1566 ( 
.A(n_1435),
.Y(n_1566)
);

A2O1A1Ixp33_ASAP7_75t_L g1567 ( 
.A1(n_1365),
.A2(n_844),
.B(n_1194),
.C(n_1188),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1365),
.A2(n_1330),
.B1(n_1194),
.B2(n_1050),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1365),
.A2(n_1330),
.B1(n_1194),
.B2(n_1050),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1365),
.A2(n_1330),
.B1(n_1194),
.B2(n_1050),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1354),
.B(n_1362),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1355),
.B(n_1366),
.Y(n_1572)
);

AOI221xp5_ASAP7_75t_L g1573 ( 
.A1(n_1365),
.A2(n_579),
.B1(n_1370),
.B2(n_683),
.C(n_738),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1365),
.A2(n_1330),
.B1(n_1194),
.B2(n_1050),
.Y(n_1574)
);

BUFx6f_ASAP7_75t_L g1575 ( 
.A(n_1407),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1358),
.B(n_1354),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1355),
.B(n_1366),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1365),
.A2(n_1330),
.B1(n_1194),
.B2(n_1050),
.Y(n_1578)
);

OAI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1365),
.A2(n_1319),
.B1(n_1194),
.B2(n_844),
.Y(n_1579)
);

NAND3xp33_ASAP7_75t_L g1580 ( 
.A(n_1370),
.B(n_1365),
.C(n_1188),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1358),
.B(n_1354),
.Y(n_1581)
);

OAI221xp5_ASAP7_75t_L g1582 ( 
.A1(n_1365),
.A2(n_791),
.B1(n_624),
.B2(n_849),
.C(n_461),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1365),
.A2(n_1330),
.B1(n_1194),
.B2(n_1050),
.Y(n_1583)
);

AOI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1410),
.A2(n_1247),
.B(n_1304),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1354),
.B(n_1362),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1354),
.B(n_1362),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1354),
.B(n_1362),
.Y(n_1587)
);

AOI321xp33_ASAP7_75t_L g1588 ( 
.A1(n_1365),
.A2(n_1194),
.A3(n_1370),
.B1(n_1188),
.B2(n_1337),
.C(n_1371),
.Y(n_1588)
);

AOI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1365),
.A2(n_624),
.B1(n_1194),
.B2(n_791),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_SL g1590 ( 
.A1(n_1365),
.A2(n_1194),
.B1(n_1026),
.B2(n_1050),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1365),
.A2(n_1330),
.B1(n_1194),
.B2(n_1050),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1497),
.Y(n_1592)
);

OAI211xp5_ASAP7_75t_SL g1593 ( 
.A1(n_1363),
.A2(n_783),
.B(n_717),
.C(n_1370),
.Y(n_1593)
);

OAI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1365),
.A2(n_1194),
.B1(n_844),
.B2(n_1370),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1365),
.A2(n_1319),
.B1(n_1194),
.B2(n_844),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1356),
.Y(n_1596)
);

BUFx6f_ASAP7_75t_L g1597 ( 
.A(n_1407),
.Y(n_1597)
);

INVx3_ASAP7_75t_L g1598 ( 
.A(n_1435),
.Y(n_1598)
);

NAND3xp33_ASAP7_75t_L g1599 ( 
.A(n_1370),
.B(n_1365),
.C(n_1188),
.Y(n_1599)
);

OAI221xp5_ASAP7_75t_L g1600 ( 
.A1(n_1573),
.A2(n_1588),
.B1(n_1580),
.B2(n_1599),
.C(n_1589),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1512),
.B(n_1516),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1500),
.B(n_1565),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1564),
.B(n_1571),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1585),
.B(n_1586),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1563),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1592),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1587),
.B(n_1548),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1517),
.Y(n_1608)
);

BUFx2_ASAP7_75t_L g1609 ( 
.A(n_1517),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1576),
.B(n_1581),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1572),
.B(n_1577),
.Y(n_1611)
);

OAI33xp33_ASAP7_75t_L g1612 ( 
.A1(n_1594),
.A2(n_1595),
.A3(n_1579),
.B1(n_1506),
.B2(n_1505),
.B3(n_1519),
.Y(n_1612)
);

BUFx3_ASAP7_75t_L g1613 ( 
.A(n_1561),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1562),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1529),
.B(n_1517),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1529),
.B(n_1518),
.Y(n_1616)
);

INVx3_ASAP7_75t_L g1617 ( 
.A(n_1529),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1510),
.B(n_1521),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1521),
.B(n_1526),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1544),
.B(n_1554),
.Y(n_1620)
);

NAND2x1_ASAP7_75t_L g1621 ( 
.A(n_1558),
.B(n_1520),
.Y(n_1621)
);

BUFx3_ASAP7_75t_L g1622 ( 
.A(n_1538),
.Y(n_1622)
);

INVx4_ASAP7_75t_R g1623 ( 
.A(n_1552),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1501),
.B(n_1504),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1507),
.B(n_1509),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1596),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1555),
.B(n_1557),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_SL g1628 ( 
.A(n_1499),
.B(n_1594),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1555),
.B(n_1533),
.Y(n_1629)
);

AOI221xp5_ASAP7_75t_L g1630 ( 
.A1(n_1567),
.A2(n_1502),
.B1(n_1582),
.B2(n_1568),
.C(n_1570),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_SL g1631 ( 
.A(n_1567),
.B(n_1522),
.Y(n_1631)
);

BUFx2_ASAP7_75t_L g1632 ( 
.A(n_1560),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1537),
.B(n_1524),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1546),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1527),
.B(n_1584),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_L g1636 ( 
.A(n_1522),
.B(n_1593),
.Y(n_1636)
);

AO21x2_ASAP7_75t_L g1637 ( 
.A1(n_1559),
.A2(n_1534),
.B(n_1514),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1531),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1614),
.Y(n_1639)
);

INVx5_ASAP7_75t_L g1640 ( 
.A(n_1617),
.Y(n_1640)
);

OAI322xp33_ASAP7_75t_L g1641 ( 
.A1(n_1631),
.A2(n_1514),
.A3(n_1511),
.B1(n_1535),
.B2(n_1502),
.C1(n_1540),
.C2(n_1543),
.Y(n_1641)
);

OA21x2_ASAP7_75t_L g1642 ( 
.A1(n_1608),
.A2(n_1541),
.B(n_1542),
.Y(n_1642)
);

NAND3xp33_ASAP7_75t_L g1643 ( 
.A(n_1631),
.B(n_1570),
.C(n_1591),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1611),
.B(n_1606),
.Y(n_1644)
);

CKINVDCx16_ASAP7_75t_R g1645 ( 
.A(n_1622),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1605),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1605),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1606),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1608),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1630),
.A2(n_1590),
.B1(n_1569),
.B2(n_1578),
.Y(n_1650)
);

INVx1_ASAP7_75t_SL g1651 ( 
.A(n_1613),
.Y(n_1651)
);

AOI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1630),
.A2(n_1578),
.B1(n_1583),
.B2(n_1569),
.Y(n_1652)
);

OAI21x1_ASAP7_75t_SL g1653 ( 
.A1(n_1607),
.A2(n_1525),
.B(n_1530),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1628),
.A2(n_1591),
.B1(n_1583),
.B2(n_1574),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1608),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_R g1656 ( 
.A(n_1636),
.B(n_1528),
.Y(n_1656)
);

AOI321xp33_ASAP7_75t_L g1657 ( 
.A1(n_1600),
.A2(n_1568),
.A3(n_1574),
.B1(n_1523),
.B2(n_1525),
.C(n_1530),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1603),
.B(n_1547),
.Y(n_1658)
);

OAI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1600),
.A2(n_1508),
.B1(n_1523),
.B2(n_1547),
.C(n_1550),
.Y(n_1659)
);

OAI31xp33_ASAP7_75t_L g1660 ( 
.A1(n_1628),
.A2(n_1532),
.A3(n_1553),
.B(n_1556),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1635),
.B(n_1559),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1633),
.A2(n_1550),
.B1(n_1551),
.B2(n_1515),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1626),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1626),
.Y(n_1664)
);

NAND4xp25_ASAP7_75t_L g1665 ( 
.A(n_1636),
.B(n_1635),
.C(n_1607),
.D(n_1638),
.Y(n_1665)
);

NAND3xp33_ASAP7_75t_L g1666 ( 
.A(n_1638),
.B(n_1528),
.C(n_1503),
.Y(n_1666)
);

BUFx2_ASAP7_75t_L g1667 ( 
.A(n_1632),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1609),
.Y(n_1668)
);

OR2x6_ASAP7_75t_L g1669 ( 
.A(n_1620),
.B(n_1513),
.Y(n_1669)
);

OAI221xp5_ASAP7_75t_L g1670 ( 
.A1(n_1633),
.A2(n_1515),
.B1(n_1539),
.B2(n_1545),
.C(n_1536),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1609),
.Y(n_1671)
);

INVxp67_ASAP7_75t_SL g1672 ( 
.A(n_1609),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1603),
.B(n_1566),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1603),
.B(n_1598),
.Y(n_1674)
);

OAI33xp33_ASAP7_75t_L g1675 ( 
.A1(n_1619),
.A2(n_1618),
.A3(n_1634),
.B1(n_1625),
.B2(n_1610),
.B3(n_1626),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_R g1676 ( 
.A(n_1613),
.B(n_1513),
.Y(n_1676)
);

AOI221xp5_ASAP7_75t_L g1677 ( 
.A1(n_1612),
.A2(n_1553),
.B1(n_1513),
.B2(n_1575),
.C(n_1597),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1611),
.B(n_1549),
.Y(n_1678)
);

BUFx3_ASAP7_75t_L g1679 ( 
.A(n_1613),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1667),
.B(n_1632),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1667),
.B(n_1615),
.Y(n_1681)
);

INVxp67_ASAP7_75t_L g1682 ( 
.A(n_1648),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1646),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1646),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1640),
.B(n_1615),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1640),
.B(n_1615),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1647),
.Y(n_1687)
);

INVx1_ASAP7_75t_SL g1688 ( 
.A(n_1640),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1640),
.B(n_1616),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1640),
.B(n_1616),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1640),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1644),
.B(n_1616),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1640),
.B(n_1601),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1665),
.B(n_1612),
.Y(n_1694)
);

BUFx3_ASAP7_75t_L g1695 ( 
.A(n_1669),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1672),
.B(n_1635),
.Y(n_1696)
);

INVx1_ASAP7_75t_SL g1697 ( 
.A(n_1649),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1658),
.B(n_1673),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1658),
.B(n_1673),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1658),
.B(n_1601),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1639),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1639),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1674),
.B(n_1601),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1663),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1644),
.B(n_1611),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1663),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1672),
.B(n_1604),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1661),
.B(n_1618),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1649),
.B(n_1617),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1655),
.B(n_1617),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1661),
.B(n_1617),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1655),
.B(n_1617),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1664),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1668),
.B(n_1604),
.Y(n_1714)
);

INVx1_ASAP7_75t_SL g1715 ( 
.A(n_1708),
.Y(n_1715)
);

INVxp67_ASAP7_75t_SL g1716 ( 
.A(n_1696),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1695),
.B(n_1669),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1705),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1696),
.B(n_1648),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1683),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1683),
.Y(n_1721)
);

NOR3x1_ASAP7_75t_L g1722 ( 
.A(n_1696),
.B(n_1665),
.C(n_1670),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1683),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1695),
.B(n_1669),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1680),
.B(n_1668),
.Y(n_1725)
);

AND2x2_ASAP7_75t_SL g1726 ( 
.A(n_1680),
.B(n_1642),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1700),
.B(n_1645),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1684),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1708),
.B(n_1705),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1700),
.B(n_1645),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1701),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1701),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1705),
.Y(n_1733)
);

INVxp67_ASAP7_75t_L g1734 ( 
.A(n_1694),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1708),
.B(n_1678),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1684),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1684),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1680),
.B(n_1671),
.Y(n_1738)
);

AND2x4_ASAP7_75t_L g1739 ( 
.A(n_1695),
.B(n_1669),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1708),
.B(n_1678),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1680),
.B(n_1671),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1700),
.B(n_1698),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1694),
.A2(n_1643),
.B1(n_1675),
.B2(n_1654),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1705),
.B(n_1602),
.Y(n_1744)
);

INVx1_ASAP7_75t_SL g1745 ( 
.A(n_1711),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1700),
.B(n_1624),
.Y(n_1746)
);

AOI322xp5_ASAP7_75t_L g1747 ( 
.A1(n_1681),
.A2(n_1652),
.A3(n_1650),
.B1(n_1619),
.B2(n_1629),
.C1(n_1677),
.C2(n_1675),
.Y(n_1747)
);

AOI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1711),
.A2(n_1660),
.B(n_1654),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1687),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1711),
.B(n_1624),
.Y(n_1750)
);

INVx2_ASAP7_75t_SL g1751 ( 
.A(n_1693),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1698),
.B(n_1679),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1687),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1715),
.B(n_1711),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1729),
.B(n_1735),
.Y(n_1755)
);

NAND2x1p5_ASAP7_75t_L g1756 ( 
.A(n_1726),
.B(n_1695),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_L g1757 ( 
.A(n_1734),
.B(n_1670),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1742),
.B(n_1698),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1726),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1748),
.B(n_1698),
.Y(n_1760)
);

NAND4xp25_ASAP7_75t_L g1761 ( 
.A(n_1722),
.B(n_1657),
.C(n_1643),
.D(n_1652),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1720),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1729),
.B(n_1692),
.Y(n_1763)
);

AND4x1_ASAP7_75t_L g1764 ( 
.A(n_1743),
.B(n_1660),
.C(n_1677),
.D(n_1666),
.Y(n_1764)
);

INVx1_ASAP7_75t_SL g1765 ( 
.A(n_1735),
.Y(n_1765)
);

INVxp67_ASAP7_75t_SL g1766 ( 
.A(n_1725),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1740),
.B(n_1692),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1731),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1744),
.B(n_1602),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1744),
.B(n_1703),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1731),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1740),
.B(n_1692),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1747),
.B(n_1699),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1742),
.B(n_1699),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1727),
.B(n_1699),
.Y(n_1775)
);

INVx1_ASAP7_75t_SL g1776 ( 
.A(n_1727),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1745),
.B(n_1746),
.Y(n_1777)
);

CKINVDCx20_ASAP7_75t_R g1778 ( 
.A(n_1730),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1732),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1720),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1716),
.B(n_1699),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1730),
.B(n_1681),
.Y(n_1782)
);

AOI221x1_ASAP7_75t_L g1783 ( 
.A1(n_1717),
.A2(n_1653),
.B1(n_1666),
.B2(n_1634),
.C(n_1704),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1752),
.B(n_1681),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1719),
.B(n_1692),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1752),
.B(n_1681),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1717),
.B(n_1695),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1718),
.B(n_1693),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1733),
.B(n_1682),
.Y(n_1789)
);

OAI31xp33_ASAP7_75t_L g1790 ( 
.A1(n_1719),
.A2(n_1659),
.A3(n_1627),
.B(n_1629),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1750),
.B(n_1707),
.Y(n_1791)
);

INVxp33_ASAP7_75t_SL g1792 ( 
.A(n_1738),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1721),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1751),
.B(n_1693),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1721),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1723),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1757),
.B(n_1717),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1755),
.Y(n_1798)
);

INVxp67_ASAP7_75t_SL g1799 ( 
.A(n_1756),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1760),
.B(n_1714),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1775),
.B(n_1693),
.Y(n_1801)
);

INVx2_ASAP7_75t_SL g1802 ( 
.A(n_1756),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1762),
.Y(n_1803)
);

NAND3x2_ASAP7_75t_L g1804 ( 
.A(n_1755),
.B(n_1686),
.C(n_1685),
.Y(n_1804)
);

INVx1_ASAP7_75t_SL g1805 ( 
.A(n_1778),
.Y(n_1805)
);

AOI21xp33_ASAP7_75t_SL g1806 ( 
.A1(n_1756),
.A2(n_1751),
.B(n_1741),
.Y(n_1806)
);

NOR4xp25_ASAP7_75t_L g1807 ( 
.A(n_1761),
.B(n_1697),
.C(n_1641),
.D(n_1682),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1762),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1780),
.Y(n_1809)
);

OAI221xp5_ASAP7_75t_L g1810 ( 
.A1(n_1764),
.A2(n_1657),
.B1(n_1659),
.B2(n_1642),
.C(n_1662),
.Y(n_1810)
);

OAI21xp33_ASAP7_75t_L g1811 ( 
.A1(n_1773),
.A2(n_1709),
.B(n_1710),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1768),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1780),
.Y(n_1813)
);

INVxp67_ASAP7_75t_SL g1814 ( 
.A(n_1764),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1793),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1775),
.B(n_1703),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1793),
.Y(n_1817)
);

INVx1_ASAP7_75t_SL g1818 ( 
.A(n_1776),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1795),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1795),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1796),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1790),
.B(n_1714),
.Y(n_1822)
);

AOI31xp33_ASAP7_75t_L g1823 ( 
.A1(n_1776),
.A2(n_1688),
.A3(n_1689),
.B(n_1690),
.Y(n_1823)
);

AOI211xp5_ASAP7_75t_L g1824 ( 
.A1(n_1759),
.A2(n_1641),
.B(n_1656),
.C(n_1688),
.Y(n_1824)
);

A2O1A1Ixp33_ASAP7_75t_L g1825 ( 
.A1(n_1790),
.A2(n_1689),
.B(n_1690),
.C(n_1686),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1768),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1765),
.B(n_1769),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1765),
.B(n_1714),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1796),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1766),
.B(n_1792),
.Y(n_1830)
);

OAI21xp33_ASAP7_75t_L g1831 ( 
.A1(n_1759),
.A2(n_1754),
.B(n_1761),
.Y(n_1831)
);

OAI21xp33_ASAP7_75t_L g1832 ( 
.A1(n_1759),
.A2(n_1709),
.B(n_1710),
.Y(n_1832)
);

OAI32xp33_ASAP7_75t_L g1833 ( 
.A1(n_1822),
.A2(n_1754),
.A3(n_1783),
.B1(n_1785),
.B2(n_1781),
.Y(n_1833)
);

AOI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1814),
.A2(n_1810),
.B1(n_1807),
.B2(n_1831),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1805),
.B(n_1783),
.Y(n_1835)
);

OAI21xp33_ASAP7_75t_L g1836 ( 
.A1(n_1811),
.A2(n_1777),
.B(n_1789),
.Y(n_1836)
);

NAND3xp33_ASAP7_75t_L g1837 ( 
.A(n_1824),
.B(n_1789),
.C(n_1768),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1803),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1816),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1798),
.B(n_1763),
.Y(n_1840)
);

NAND4xp25_ASAP7_75t_L g1841 ( 
.A(n_1818),
.B(n_1763),
.C(n_1794),
.D(n_1785),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1798),
.B(n_1767),
.Y(n_1842)
);

NAND2x1_ASAP7_75t_L g1843 ( 
.A(n_1823),
.B(n_1758),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1827),
.B(n_1830),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1816),
.B(n_1758),
.Y(n_1845)
);

INVxp67_ASAP7_75t_L g1846 ( 
.A(n_1797),
.Y(n_1846)
);

AOI221xp5_ASAP7_75t_L g1847 ( 
.A1(n_1799),
.A2(n_1653),
.B1(n_1771),
.B2(n_1779),
.C(n_1732),
.Y(n_1847)
);

INVxp67_ASAP7_75t_L g1848 ( 
.A(n_1802),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1800),
.B(n_1770),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1803),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1801),
.B(n_1774),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1808),
.Y(n_1852)
);

OAI22xp5_ASAP7_75t_L g1853 ( 
.A1(n_1804),
.A2(n_1772),
.B1(n_1767),
.B2(n_1774),
.Y(n_1853)
);

AOI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1802),
.A2(n_1779),
.B(n_1771),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_SL g1855 ( 
.A1(n_1804),
.A2(n_1637),
.B1(n_1642),
.B2(n_1779),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_SL g1856 ( 
.A(n_1806),
.B(n_1787),
.Y(n_1856)
);

AOI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1812),
.A2(n_1637),
.B1(n_1787),
.B2(n_1642),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1801),
.B(n_1782),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1858),
.B(n_1782),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1845),
.B(n_1839),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1846),
.B(n_1828),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1846),
.B(n_1829),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1842),
.Y(n_1863)
);

NOR3xp33_ASAP7_75t_SL g1864 ( 
.A(n_1833),
.B(n_1825),
.C(n_1832),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1840),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1834),
.B(n_1808),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1851),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1838),
.Y(n_1868)
);

OAI22xp33_ASAP7_75t_L g1869 ( 
.A1(n_1857),
.A2(n_1772),
.B1(n_1621),
.B2(n_1826),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1841),
.B(n_1809),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1850),
.Y(n_1871)
);

OAI21xp33_ASAP7_75t_L g1872 ( 
.A1(n_1836),
.A2(n_1855),
.B(n_1835),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1844),
.B(n_1809),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1852),
.Y(n_1874)
);

OAI221xp5_ASAP7_75t_L g1875 ( 
.A1(n_1855),
.A2(n_1826),
.B1(n_1812),
.B2(n_1817),
.C(n_1813),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1848),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1837),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_SL g1878 ( 
.A(n_1847),
.B(n_1813),
.Y(n_1878)
);

AOI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1878),
.A2(n_1847),
.B(n_1854),
.Y(n_1879)
);

NAND2xp33_ASAP7_75t_L g1880 ( 
.A(n_1864),
.B(n_1856),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1860),
.B(n_1867),
.Y(n_1881)
);

INVxp67_ASAP7_75t_L g1882 ( 
.A(n_1866),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1860),
.B(n_1849),
.Y(n_1883)
);

NOR3x1_ASAP7_75t_L g1884 ( 
.A(n_1861),
.B(n_1843),
.C(n_1853),
.Y(n_1884)
);

AOI32xp33_ASAP7_75t_L g1885 ( 
.A1(n_1877),
.A2(n_1817),
.A3(n_1821),
.B1(n_1820),
.B2(n_1819),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1872),
.A2(n_1637),
.B1(n_1642),
.B2(n_1787),
.Y(n_1886)
);

OAI31xp33_ASAP7_75t_L g1887 ( 
.A1(n_1875),
.A2(n_1854),
.A3(n_1821),
.B(n_1820),
.Y(n_1887)
);

INVxp67_ASAP7_75t_L g1888 ( 
.A(n_1877),
.Y(n_1888)
);

NOR3xp33_ASAP7_75t_L g1889 ( 
.A(n_1878),
.B(n_1819),
.C(n_1815),
.Y(n_1889)
);

NOR4xp25_ASAP7_75t_L g1890 ( 
.A(n_1876),
.B(n_1815),
.C(n_1771),
.D(n_1697),
.Y(n_1890)
);

AOI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1889),
.A2(n_1886),
.B1(n_1882),
.B2(n_1879),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1883),
.B(n_1867),
.Y(n_1892)
);

AOI221xp5_ASAP7_75t_L g1893 ( 
.A1(n_1889),
.A2(n_1869),
.B1(n_1865),
.B2(n_1863),
.C(n_1870),
.Y(n_1893)
);

AOI222xp33_ASAP7_75t_L g1894 ( 
.A1(n_1888),
.A2(n_1873),
.B1(n_1874),
.B2(n_1871),
.C1(n_1868),
.C2(n_1862),
.Y(n_1894)
);

OAI211xp5_ASAP7_75t_L g1895 ( 
.A1(n_1890),
.A2(n_1870),
.B(n_1859),
.C(n_1794),
.Y(n_1895)
);

OAI221xp5_ASAP7_75t_SL g1896 ( 
.A1(n_1887),
.A2(n_1859),
.B1(n_1688),
.B2(n_1691),
.C(n_1689),
.Y(n_1896)
);

AOI221xp5_ASAP7_75t_SL g1897 ( 
.A1(n_1880),
.A2(n_1786),
.B1(n_1784),
.B2(n_1697),
.C(n_1788),
.Y(n_1897)
);

NOR3xp33_ASAP7_75t_L g1898 ( 
.A(n_1881),
.B(n_1787),
.C(n_1691),
.Y(n_1898)
);

AOI221xp5_ASAP7_75t_L g1899 ( 
.A1(n_1885),
.A2(n_1710),
.B1(n_1712),
.B2(n_1709),
.C(n_1627),
.Y(n_1899)
);

AOI211xp5_ASAP7_75t_L g1900 ( 
.A1(n_1884),
.A2(n_1691),
.B(n_1690),
.C(n_1689),
.Y(n_1900)
);

AOI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1889),
.A2(n_1637),
.B1(n_1739),
.B2(n_1724),
.Y(n_1901)
);

AOI21xp5_ASAP7_75t_L g1902 ( 
.A1(n_1892),
.A2(n_1784),
.B(n_1786),
.Y(n_1902)
);

NAND2xp33_ASAP7_75t_SL g1903 ( 
.A(n_1897),
.B(n_1788),
.Y(n_1903)
);

XNOR2xp5_ASAP7_75t_L g1904 ( 
.A(n_1891),
.B(n_1724),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1895),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1901),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_R g1907 ( 
.A(n_1894),
.B(n_1623),
.Y(n_1907)
);

XOR2xp5_ASAP7_75t_L g1908 ( 
.A(n_1893),
.B(n_1724),
.Y(n_1908)
);

NOR2x1_ASAP7_75t_L g1909 ( 
.A(n_1905),
.B(n_1908),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1902),
.Y(n_1910)
);

AOI221xp5_ASAP7_75t_L g1911 ( 
.A1(n_1906),
.A2(n_1896),
.B1(n_1900),
.B2(n_1898),
.C(n_1899),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_1907),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1904),
.B(n_1703),
.Y(n_1913)
);

NOR3xp33_ASAP7_75t_L g1914 ( 
.A(n_1903),
.B(n_1691),
.C(n_1739),
.Y(n_1914)
);

NOR4xp25_ASAP7_75t_L g1915 ( 
.A(n_1905),
.B(n_1749),
.C(n_1753),
.D(n_1737),
.Y(n_1915)
);

INVxp33_ASAP7_75t_L g1916 ( 
.A(n_1909),
.Y(n_1916)
);

AOI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1910),
.A2(n_1637),
.B1(n_1739),
.B2(n_1627),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1913),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1914),
.Y(n_1919)
);

NOR2x1_ASAP7_75t_L g1920 ( 
.A(n_1912),
.B(n_1723),
.Y(n_1920)
);

HB1xp67_ASAP7_75t_L g1921 ( 
.A(n_1916),
.Y(n_1921)
);

HB1xp67_ASAP7_75t_L g1922 ( 
.A(n_1918),
.Y(n_1922)
);

AOI221xp5_ASAP7_75t_L g1923 ( 
.A1(n_1919),
.A2(n_1915),
.B1(n_1911),
.B2(n_1712),
.C(n_1753),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1922),
.B(n_1920),
.Y(n_1924)
);

NAND3xp33_ASAP7_75t_L g1925 ( 
.A(n_1924),
.B(n_1921),
.C(n_1923),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1925),
.Y(n_1926)
);

NAND2xp33_ASAP7_75t_R g1927 ( 
.A(n_1925),
.B(n_1676),
.Y(n_1927)
);

AO22x1_ASAP7_75t_L g1928 ( 
.A1(n_1926),
.A2(n_1917),
.B1(n_1728),
.B2(n_1749),
.Y(n_1928)
);

NAND3xp33_ASAP7_75t_L g1929 ( 
.A(n_1927),
.B(n_1701),
.C(n_1702),
.Y(n_1929)
);

AOI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1928),
.A2(n_1791),
.B(n_1737),
.Y(n_1930)
);

AOI222xp33_ASAP7_75t_SL g1931 ( 
.A1(n_1929),
.A2(n_1651),
.B1(n_1736),
.B2(n_1728),
.C1(n_1623),
.C2(n_1706),
.Y(n_1931)
);

AOI22xp5_ASAP7_75t_SL g1932 ( 
.A1(n_1930),
.A2(n_1690),
.B1(n_1613),
.B2(n_1736),
.Y(n_1932)
);

OAI221xp5_ASAP7_75t_L g1933 ( 
.A1(n_1932),
.A2(n_1931),
.B1(n_1712),
.B2(n_1621),
.C(n_1713),
.Y(n_1933)
);

AOI211xp5_ASAP7_75t_L g1934 ( 
.A1(n_1933),
.A2(n_1685),
.B(n_1686),
.C(n_1575),
.Y(n_1934)
);


endmodule