module fake_jpeg_30126_n_138 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_138);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_138;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_4),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_18),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_37),
.Y(n_41)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_25),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_15),
.B1(n_14),
.B2(n_26),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_26),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_46),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_54),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_40),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_30),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_14),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_52),
.B(n_57),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_24),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_32),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_29),
.B(n_13),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_27),
.Y(n_69)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_33),
.C(n_31),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_66),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_69),
.Y(n_82)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_27),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_73),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_30),
.C(n_27),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_27),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_21),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_74),
.B(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_21),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_49),
.A2(n_30),
.B1(n_21),
.B2(n_12),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_76),
.A2(n_53),
.B1(n_17),
.B2(n_3),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_41),
.B(n_21),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_80),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_58),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_54),
.A2(n_12),
.B(n_17),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_79),
.A2(n_43),
.B(n_55),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_12),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_63),
.A2(n_48),
.B1(n_50),
.B2(n_60),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_81),
.A2(n_92),
.B1(n_71),
.B2(n_65),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_85),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_58),
.B(n_51),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_48),
.B(n_57),
.Y(n_86)
);

AOI22x1_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_53),
.B1(n_72),
.B2(n_65),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_88),
.B(n_96),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_70),
.A2(n_56),
.B1(n_49),
.B2(n_43),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_93),
.B1(n_78),
.B2(n_71),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_56),
.B1(n_43),
.B2(n_55),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_68),
.B(n_8),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_91),
.Y(n_97)
);

NOR4xp25_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_106),
.C(n_104),
.D(n_108),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_70),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_99),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_62),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_66),
.C(n_61),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_87),
.C(n_84),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_108),
.B(n_89),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_94),
.A2(n_78),
.B1(n_67),
.B2(n_79),
.Y(n_102)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_103),
.A2(n_88),
.B(n_92),
.Y(n_110)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_82),
.B(n_72),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_110),
.A2(n_111),
.B1(n_114),
.B2(n_115),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_100),
.C(n_98),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_108),
.A2(n_65),
.B1(n_86),
.B2(n_91),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_119),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_116),
.Y(n_118)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_99),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_120),
.A2(n_121),
.B(n_122),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_107),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

AOI322xp5_ASAP7_75t_L g127 ( 
.A1(n_123),
.A2(n_112),
.A3(n_85),
.B1(n_107),
.B2(n_103),
.C1(n_101),
.C2(n_102),
.Y(n_127)
);

NOR3xp33_ASAP7_75t_SL g131 ( 
.A(n_127),
.B(n_128),
.C(n_11),
.Y(n_131)
);

OAI321xp33_ASAP7_75t_L g128 ( 
.A1(n_121),
.A2(n_84),
.A3(n_8),
.B1(n_11),
.B2(n_7),
.C(n_2),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_118),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_130),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_117),
.C(n_119),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_131),
.B(n_1),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_131),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_134),
.B(n_135),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_126),
.C(n_5),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_1),
.C(n_5),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_17),
.Y(n_138)
);


endmodule