module real_aes_8408_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_241;
wire n_168;
wire n_175;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g420 ( .A(n_0), .Y(n_420) );
INVx1_ASAP7_75t_L g463 ( .A(n_1), .Y(n_463) );
INVx1_ASAP7_75t_L g238 ( .A(n_2), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_3), .A2(n_36), .B1(n_157), .B2(n_491), .Y(n_490) );
AOI21xp33_ASAP7_75t_L g145 ( .A1(n_4), .A2(n_146), .B(n_147), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_5), .B(n_144), .Y(n_440) );
AND2x6_ASAP7_75t_L g119 ( .A(n_6), .B(n_120), .Y(n_119) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_7), .A2(n_214), .B(n_215), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_8), .B(n_37), .Y(n_421) );
INVx1_ASAP7_75t_L g154 ( .A(n_9), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_10), .B(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g116 ( .A(n_11), .Y(n_116) );
INVx1_ASAP7_75t_L g459 ( .A(n_12), .Y(n_459) );
INVx1_ASAP7_75t_L g220 ( .A(n_13), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_14), .B(n_122), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_15), .B(n_112), .Y(n_468) );
AO32x2_ASAP7_75t_L g488 ( .A1(n_16), .A2(n_111), .A3(n_144), .B1(n_451), .B2(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_17), .B(n_157), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_18), .B(n_165), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_19), .B(n_112), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_20), .A2(n_48), .B1(n_157), .B2(n_491), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_21), .B(n_146), .Y(n_174) );
AOI22xp33_ASAP7_75t_SL g511 ( .A1(n_22), .A2(n_73), .B1(n_122), .B2(n_157), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_23), .B(n_157), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_24), .B(n_142), .Y(n_168) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_25), .A2(n_218), .B(n_219), .C(n_221), .Y(n_217) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_26), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_27), .B(n_159), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_28), .B(n_152), .Y(n_239) );
INVx1_ASAP7_75t_L g130 ( .A(n_29), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_30), .B(n_159), .Y(n_485) );
INVx2_ASAP7_75t_L g124 ( .A(n_31), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_32), .B(n_157), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_33), .B(n_159), .Y(n_502) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_34), .A2(n_101), .B1(n_718), .B2(n_727), .C1(n_736), .C2(n_742), .Y(n_100) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_34), .A2(n_40), .B1(n_731), .B2(n_732), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_34), .Y(n_732) );
A2O1A1Ixp33_ASAP7_75t_L g175 ( .A1(n_35), .A2(n_119), .B(n_131), .C(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g128 ( .A(n_38), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_39), .B(n_152), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_40), .Y(n_731) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_41), .B(n_157), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_42), .A2(n_84), .B1(n_182), .B2(n_491), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_43), .B(n_157), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_44), .B(n_157), .Y(n_460) );
CKINVDCx16_ASAP7_75t_R g134 ( .A(n_45), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_46), .B(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_47), .B(n_146), .Y(n_208) );
AOI22xp33_ASAP7_75t_SL g472 ( .A1(n_49), .A2(n_58), .B1(n_122), .B2(n_157), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g121 ( .A1(n_50), .A2(n_122), .B1(n_125), .B2(n_131), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_51), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_52), .B(n_157), .Y(n_450) );
CKINVDCx16_ASAP7_75t_R g235 ( .A(n_53), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_54), .B(n_157), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_L g150 ( .A1(n_55), .A2(n_151), .B(n_153), .C(n_156), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_56), .Y(n_195) );
INVx1_ASAP7_75t_L g148 ( .A(n_57), .Y(n_148) );
INVx1_ASAP7_75t_L g120 ( .A(n_59), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_60), .B(n_157), .Y(n_464) );
INVx1_ASAP7_75t_L g115 ( .A(n_61), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_62), .Y(n_723) );
AO32x2_ASAP7_75t_L g508 ( .A1(n_63), .A2(n_144), .A3(n_200), .B1(n_451), .B2(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g448 ( .A(n_64), .Y(n_448) );
INVx1_ASAP7_75t_L g480 ( .A(n_65), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_SL g164 ( .A1(n_66), .A2(n_156), .B(n_165), .C(n_166), .Y(n_164) );
INVxp67_ASAP7_75t_L g167 ( .A(n_67), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_68), .B(n_122), .Y(n_481) );
INVx1_ASAP7_75t_L g722 ( .A(n_69), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_70), .Y(n_139) );
INVx1_ASAP7_75t_L g188 ( .A(n_71), .Y(n_188) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_72), .A2(n_98), .B1(n_708), .B2(n_709), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_72), .Y(n_708) );
A2O1A1Ixp33_ASAP7_75t_L g189 ( .A1(n_74), .A2(n_119), .B(n_131), .C(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_75), .B(n_491), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_76), .B(n_122), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_77), .B(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g113 ( .A(n_78), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_79), .B(n_165), .Y(n_179) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_80), .A2(n_103), .B1(n_707), .B2(n_710), .C1(n_711), .C2(n_714), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_81), .B(n_122), .Y(n_434) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_82), .A2(n_119), .B(n_131), .C(n_237), .Y(n_236) );
OR2x2_ASAP7_75t_L g418 ( .A(n_83), .B(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g706 ( .A(n_83), .Y(n_706) );
OR2x2_ASAP7_75t_L g726 ( .A(n_83), .B(n_717), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_85), .A2(n_99), .B1(n_122), .B2(n_123), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_86), .B(n_734), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_87), .B(n_159), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_88), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_89), .A2(n_119), .B(n_131), .C(n_203), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_90), .Y(n_210) );
INVx1_ASAP7_75t_L g163 ( .A(n_91), .Y(n_163) );
CKINVDCx16_ASAP7_75t_R g216 ( .A(n_92), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_93), .B(n_178), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_94), .B(n_122), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_95), .B(n_144), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_96), .A2(n_146), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_97), .B(n_722), .Y(n_721) );
CKINVDCx16_ASAP7_75t_R g709 ( .A(n_98), .Y(n_709) );
INVxp67_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
OAI22xp5_ASAP7_75t_SL g103 ( .A1(n_104), .A2(n_416), .B1(n_422), .B2(n_703), .Y(n_103) );
INVx1_ASAP7_75t_L g712 ( .A(n_104), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_104), .A2(n_712), .B1(n_729), .B2(n_730), .Y(n_728) );
AND3x1_ASAP7_75t_L g104 ( .A(n_105), .B(n_341), .C(n_390), .Y(n_104) );
NOR3xp33_ASAP7_75t_SL g105 ( .A(n_106), .B(n_248), .C(n_286), .Y(n_105) );
OAI222xp33_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_169), .B1(n_223), .B2(n_229), .C1(n_243), .C2(n_246), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_140), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_108), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_108), .B(n_291), .Y(n_382) );
BUFx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g259 ( .A(n_109), .B(n_160), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_109), .B(n_141), .Y(n_267) );
AND2x2_ASAP7_75t_L g302 ( .A(n_109), .B(n_279), .Y(n_302) );
OR2x2_ASAP7_75t_L g326 ( .A(n_109), .B(n_141), .Y(n_326) );
OR2x2_ASAP7_75t_L g334 ( .A(n_109), .B(n_233), .Y(n_334) );
AND2x2_ASAP7_75t_L g337 ( .A(n_109), .B(n_160), .Y(n_337) );
INVx3_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g231 ( .A(n_110), .B(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g245 ( .A(n_110), .B(n_160), .Y(n_245) );
AND2x2_ASAP7_75t_L g295 ( .A(n_110), .B(n_233), .Y(n_295) );
AND2x2_ASAP7_75t_L g308 ( .A(n_110), .B(n_141), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_110), .B(n_394), .Y(n_415) );
AO21x2_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_117), .B(n_138), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_111), .B(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g183 ( .A(n_111), .Y(n_183) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_111), .A2(n_234), .B(n_241), .Y(n_233) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_112), .Y(n_144) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AND2x2_ASAP7_75t_SL g159 ( .A(n_113), .B(n_114), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
OAI22xp33_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_121), .B1(n_134), .B2(n_135), .Y(n_117) );
O2A1O1Ixp33_ASAP7_75t_L g147 ( .A1(n_118), .A2(n_148), .B(n_149), .C(n_150), .Y(n_147) );
O2A1O1Ixp33_ASAP7_75t_L g162 ( .A1(n_118), .A2(n_149), .B(n_163), .C(n_164), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_L g215 ( .A1(n_118), .A2(n_149), .B(n_216), .C(n_217), .Y(n_215) );
INVx4_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
NAND2x1p5_ASAP7_75t_L g135 ( .A(n_119), .B(n_136), .Y(n_135) );
AND2x4_ASAP7_75t_L g146 ( .A(n_119), .B(n_136), .Y(n_146) );
OAI21xp5_ASAP7_75t_L g431 ( .A1(n_119), .A2(n_432), .B(n_435), .Y(n_431) );
BUFx3_ASAP7_75t_L g451 ( .A(n_119), .Y(n_451) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_119), .A2(n_458), .B(n_462), .Y(n_457) );
OAI21xp5_ASAP7_75t_L g478 ( .A1(n_119), .A2(n_479), .B(n_482), .Y(n_478) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_119), .A2(n_495), .B(n_499), .Y(n_494) );
INVx2_ASAP7_75t_L g240 ( .A(n_122), .Y(n_240) );
INVx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g132 ( .A(n_124), .Y(n_132) );
INVx1_ASAP7_75t_L g137 ( .A(n_124), .Y(n_137) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_126), .A2(n_128), .B1(n_129), .B2(n_130), .Y(n_125) );
INVx2_ASAP7_75t_L g129 ( .A(n_126), .Y(n_129) );
INVx4_ASAP7_75t_L g218 ( .A(n_126), .Y(n_218) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g133 ( .A(n_127), .Y(n_133) );
AND2x2_ASAP7_75t_L g136 ( .A(n_127), .B(n_137), .Y(n_136) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_127), .Y(n_152) );
INVx3_ASAP7_75t_L g155 ( .A(n_127), .Y(n_155) );
INVx1_ASAP7_75t_L g165 ( .A(n_127), .Y(n_165) );
INVx5_ASAP7_75t_L g149 ( .A(n_131), .Y(n_149) );
AND2x6_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_132), .Y(n_157) );
BUFx3_ASAP7_75t_L g182 ( .A(n_132), .Y(n_182) );
INVx1_ASAP7_75t_L g491 ( .A(n_132), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g187 ( .A1(n_135), .A2(n_188), .B(n_189), .Y(n_187) );
OAI21xp5_ASAP7_75t_L g234 ( .A1(n_135), .A2(n_235), .B(n_236), .Y(n_234) );
INVx1_ASAP7_75t_L g438 ( .A(n_137), .Y(n_438) );
O2A1O1Ixp33_ASAP7_75t_L g333 ( .A1(n_140), .A2(n_334), .B(n_335), .C(n_338), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_140), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_140), .B(n_278), .Y(n_400) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_160), .Y(n_140) );
AND2x2_ASAP7_75t_SL g244 ( .A(n_141), .B(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g258 ( .A(n_141), .Y(n_258) );
AND2x2_ASAP7_75t_L g285 ( .A(n_141), .B(n_279), .Y(n_285) );
INVx1_ASAP7_75t_SL g293 ( .A(n_141), .Y(n_293) );
AND2x2_ASAP7_75t_L g316 ( .A(n_141), .B(n_317), .Y(n_316) );
BUFx2_ASAP7_75t_L g394 ( .A(n_141), .Y(n_394) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_145), .B(n_158), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NOR2xp33_ASAP7_75t_SL g184 ( .A(n_143), .B(n_185), .Y(n_184) );
NAND3xp33_ASAP7_75t_L g469 ( .A(n_143), .B(n_451), .C(n_470), .Y(n_469) );
AO21x1_ASAP7_75t_L g514 ( .A1(n_143), .A2(n_470), .B(n_515), .Y(n_514) );
INVx4_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_144), .A2(n_161), .B(n_168), .Y(n_160) );
OA21x2_ASAP7_75t_L g430 ( .A1(n_144), .A2(n_431), .B(n_440), .Y(n_430) );
BUFx2_ASAP7_75t_L g214 ( .A(n_146), .Y(n_214) );
O2A1O1Ixp5_ASAP7_75t_L g447 ( .A1(n_151), .A2(n_448), .B(n_449), .C(n_450), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_151), .A2(n_500), .B(n_501), .Y(n_499) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx4_ASAP7_75t_L g206 ( .A(n_152), .Y(n_206) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_152), .A2(n_439), .B1(n_471), .B2(n_472), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_152), .A2(n_439), .B1(n_490), .B2(n_492), .Y(n_489) );
OAI22xp5_ASAP7_75t_SL g509 ( .A1(n_152), .A2(n_155), .B1(n_510), .B2(n_511), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_155), .B(n_167), .Y(n_166) );
INVx5_ASAP7_75t_L g178 ( .A(n_155), .Y(n_178) );
O2A1O1Ixp5_ASAP7_75t_SL g479 ( .A1(n_156), .A2(n_178), .B(n_480), .C(n_481), .Y(n_479) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_157), .Y(n_207) );
INVx1_ASAP7_75t_L g196 ( .A(n_159), .Y(n_196) );
INVx2_ASAP7_75t_L g200 ( .A(n_159), .Y(n_200) );
OA21x2_ASAP7_75t_L g212 ( .A1(n_159), .A2(n_213), .B(n_222), .Y(n_212) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_159), .A2(n_478), .B(n_485), .Y(n_477) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_159), .A2(n_494), .B(n_502), .Y(n_493) );
BUFx2_ASAP7_75t_L g230 ( .A(n_160), .Y(n_230) );
INVx1_ASAP7_75t_L g292 ( .A(n_160), .Y(n_292) );
INVx3_ASAP7_75t_L g317 ( .A(n_160), .Y(n_317) );
INVx1_ASAP7_75t_L g498 ( .A(n_165), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_169), .B(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g169 ( .A(n_170), .B(n_197), .Y(n_169) );
INVx1_ASAP7_75t_L g313 ( .A(n_170), .Y(n_313) );
OAI32xp33_ASAP7_75t_L g319 ( .A1(n_170), .A2(n_258), .A3(n_320), .B1(n_321), .B2(n_322), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_170), .A2(n_324), .B1(n_327), .B2(n_332), .Y(n_323) );
INVx4_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g261 ( .A(n_171), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g339 ( .A(n_171), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g409 ( .A(n_171), .B(n_355), .Y(n_409) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_186), .Y(n_171) );
AND2x2_ASAP7_75t_L g224 ( .A(n_172), .B(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g254 ( .A(n_172), .Y(n_254) );
INVx1_ASAP7_75t_L g273 ( .A(n_172), .Y(n_273) );
OR2x2_ASAP7_75t_L g281 ( .A(n_172), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g288 ( .A(n_172), .B(n_262), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_172), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g309 ( .A(n_172), .B(n_227), .Y(n_309) );
INVx3_ASAP7_75t_L g331 ( .A(n_172), .Y(n_331) );
AND2x2_ASAP7_75t_L g356 ( .A(n_172), .B(n_228), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_172), .B(n_321), .Y(n_404) );
OR2x6_ASAP7_75t_L g172 ( .A(n_173), .B(n_184), .Y(n_172) );
AOI21xp5_ASAP7_75t_SL g173 ( .A1(n_174), .A2(n_175), .B(n_183), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_179), .B(n_180), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_L g237 ( .A1(n_178), .A2(n_238), .B(n_239), .C(n_240), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g432 ( .A1(n_178), .A2(n_433), .B(n_434), .Y(n_432) );
INVx2_ASAP7_75t_L g439 ( .A(n_178), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_178), .A2(n_445), .B(n_446), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_180), .A2(n_191), .B(n_192), .Y(n_190) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g221 ( .A(n_182), .Y(n_221) );
INVx1_ASAP7_75t_L g193 ( .A(n_183), .Y(n_193) );
OA21x2_ASAP7_75t_L g442 ( .A1(n_183), .A2(n_443), .B(n_452), .Y(n_442) );
OA21x2_ASAP7_75t_L g456 ( .A1(n_183), .A2(n_457), .B(n_465), .Y(n_456) );
INVx2_ASAP7_75t_L g228 ( .A(n_186), .Y(n_228) );
AND2x2_ASAP7_75t_L g360 ( .A(n_186), .B(n_198), .Y(n_360) );
AO21x2_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_193), .B(n_194), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_196), .B(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_196), .B(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g402 ( .A(n_197), .Y(n_402) );
OR2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_211), .Y(n_197) );
INVx1_ASAP7_75t_L g247 ( .A(n_198), .Y(n_247) );
AND2x2_ASAP7_75t_L g274 ( .A(n_198), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_198), .B(n_228), .Y(n_282) );
AND2x2_ASAP7_75t_L g340 ( .A(n_198), .B(n_263), .Y(n_340) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g226 ( .A(n_199), .Y(n_226) );
AND2x2_ASAP7_75t_L g253 ( .A(n_199), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g262 ( .A(n_199), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_199), .B(n_228), .Y(n_328) );
AO21x2_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B(n_209), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_202), .B(n_208), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_207), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_211), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g275 ( .A(n_211), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_211), .B(n_228), .Y(n_321) );
AND2x2_ASAP7_75t_L g330 ( .A(n_211), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g355 ( .A(n_211), .Y(n_355) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g227 ( .A(n_212), .B(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g263 ( .A(n_212), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_218), .B(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g461 ( .A(n_218), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_218), .A2(n_483), .B(n_484), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_223), .A2(n_233), .B1(n_392), .B2(n_395), .Y(n_391) );
INVx1_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
OAI21xp5_ASAP7_75t_SL g414 ( .A1(n_225), .A2(n_336), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_226), .B(n_331), .Y(n_348) );
INVx1_ASAP7_75t_L g373 ( .A(n_226), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_227), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g300 ( .A(n_227), .B(n_253), .Y(n_300) );
INVx2_ASAP7_75t_L g256 ( .A(n_228), .Y(n_256) );
INVx1_ASAP7_75t_L g306 ( .A(n_228), .Y(n_306) );
OAI221xp5_ASAP7_75t_L g397 ( .A1(n_229), .A2(n_381), .B1(n_398), .B2(n_401), .C(n_403), .Y(n_397) );
OR2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
INVx1_ASAP7_75t_L g268 ( .A(n_230), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_230), .B(n_279), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_231), .B(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g322 ( .A(n_231), .B(n_268), .Y(n_322) );
INVx3_ASAP7_75t_SL g363 ( .A(n_231), .Y(n_363) );
AND2x2_ASAP7_75t_L g307 ( .A(n_232), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g336 ( .A(n_232), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_232), .B(n_245), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_232), .B(n_291), .Y(n_377) );
INVx3_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx3_ASAP7_75t_L g279 ( .A(n_233), .Y(n_279) );
OAI322xp33_ASAP7_75t_L g374 ( .A1(n_233), .A2(n_305), .A3(n_327), .B1(n_375), .B2(n_377), .C1(n_378), .C2(n_379), .Y(n_374) );
O2A1O1Ixp33_ASAP7_75t_L g458 ( .A1(n_240), .A2(n_459), .B(n_460), .C(n_461), .Y(n_458) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AOI21xp33_ASAP7_75t_L g398 ( .A1(n_244), .A2(n_247), .B(n_399), .Y(n_398) );
NOR2xp33_ASAP7_75t_SL g324 ( .A(n_245), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g346 ( .A(n_245), .B(n_258), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_245), .B(n_285), .Y(n_361) );
INVxp67_ASAP7_75t_L g312 ( .A(n_247), .Y(n_312) );
AOI211xp5_ASAP7_75t_L g318 ( .A1(n_247), .A2(n_319), .B(n_323), .C(n_333), .Y(n_318) );
OAI221xp5_ASAP7_75t_SL g248 ( .A1(n_249), .A2(n_257), .B1(n_260), .B2(n_264), .C(n_269), .Y(n_248) );
INVxp67_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_255), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g272 ( .A(n_256), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g389 ( .A(n_256), .Y(n_389) );
OAI221xp5_ASAP7_75t_L g405 ( .A1(n_257), .A2(n_406), .B1(n_411), .B2(n_412), .C(n_414), .Y(n_405) );
OR2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_258), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_SL g305 ( .A(n_258), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_258), .B(n_336), .Y(n_343) );
AND2x2_ASAP7_75t_L g385 ( .A(n_258), .B(n_363), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_259), .B(n_284), .Y(n_283) );
OAI22xp33_ASAP7_75t_L g380 ( .A1(n_259), .A2(n_271), .B1(n_381), .B2(n_382), .Y(n_380) );
OR2x2_ASAP7_75t_L g411 ( .A(n_259), .B(n_279), .Y(n_411) );
CKINVDCx16_ASAP7_75t_R g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g388 ( .A(n_262), .Y(n_388) );
AND2x2_ASAP7_75t_L g413 ( .A(n_262), .B(n_356), .Y(n_413) );
INVxp67_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NOR2xp33_ASAP7_75t_SL g265 ( .A(n_266), .B(n_268), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g277 ( .A(n_267), .B(n_278), .Y(n_277) );
AOI22xp5_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_276), .B1(n_280), .B2(n_283), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
INVx1_ASAP7_75t_L g344 ( .A(n_272), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_272), .B(n_312), .Y(n_379) );
AOI322xp5_ASAP7_75t_L g303 ( .A1(n_274), .A2(n_304), .A3(n_306), .B1(n_307), .B2(n_309), .C1(n_310), .C2(n_314), .Y(n_303) );
INVxp67_ASAP7_75t_L g297 ( .A(n_275), .Y(n_297) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OAI22xp5_ASAP7_75t_L g298 ( .A1(n_277), .A2(n_282), .B1(n_299), .B2(n_301), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_278), .B(n_291), .Y(n_378) );
INVx1_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_279), .B(n_317), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_279), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g375 ( .A(n_281), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
NAND3xp33_ASAP7_75t_SL g286 ( .A(n_287), .B(n_303), .C(n_318), .Y(n_286) );
AOI221xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_289), .B1(n_294), .B2(n_296), .C(n_298), .Y(n_287) );
AND2x2_ASAP7_75t_L g294 ( .A(n_290), .B(n_295), .Y(n_294) );
INVx3_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
AND2x4_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
AND2x2_ASAP7_75t_L g304 ( .A(n_295), .B(n_305), .Y(n_304) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_297), .Y(n_376) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_302), .B(n_316), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_305), .B(n_363), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_306), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_SL g381 ( .A(n_309), .Y(n_381) );
AND2x2_ASAP7_75t_L g396 ( .A(n_309), .B(n_373), .Y(n_396) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AOI211xp5_ASAP7_75t_L g390 ( .A1(n_320), .A2(n_391), .B(n_397), .C(n_405), .Y(n_390) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g359 ( .A(n_330), .B(n_360), .Y(n_359) );
NAND2x1_ASAP7_75t_SL g401 ( .A(n_331), .B(n_402), .Y(n_401) );
CKINVDCx16_ASAP7_75t_R g371 ( .A(n_334), .Y(n_371) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g366 ( .A(n_340), .Y(n_366) );
AND2x2_ASAP7_75t_L g370 ( .A(n_340), .B(n_356), .Y(n_370) );
NOR5xp2_ASAP7_75t_L g341 ( .A(n_342), .B(n_357), .C(n_374), .D(n_380), .E(n_383), .Y(n_341) );
OAI221xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_344), .B1(n_345), .B2(n_347), .C(n_349), .Y(n_342) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_346), .B(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g372 ( .A(n_356), .B(n_373), .Y(n_372) );
OAI221xp5_ASAP7_75t_SL g357 ( .A1(n_358), .A2(n_361), .B1(n_362), .B2(n_364), .C(n_367), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_370), .B1(n_371), .B2(n_372), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g410 ( .A(n_370), .Y(n_410) );
AOI211xp5_ASAP7_75t_SL g383 ( .A1(n_384), .A2(n_386), .B(n_388), .C(n_389), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVxp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_408), .B(n_410), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
CKINVDCx14_ASAP7_75t_R g412 ( .A(n_413), .Y(n_412) );
OAI22xp5_ASAP7_75t_SL g711 ( .A1(n_416), .A2(n_423), .B1(n_712), .B2(n_713), .Y(n_711) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g705 ( .A(n_419), .B(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g717 ( .A(n_419), .Y(n_717) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NAND2x1p5_ASAP7_75t_L g423 ( .A(n_424), .B(n_627), .Y(n_423) );
AND2x2_ASAP7_75t_SL g424 ( .A(n_425), .B(n_585), .Y(n_424) );
NOR4xp25_ASAP7_75t_L g425 ( .A(n_426), .B(n_525), .C(n_561), .D(n_575), .Y(n_425) );
OAI221xp5_ASAP7_75t_SL g426 ( .A1(n_427), .A2(n_473), .B1(n_503), .B2(n_512), .C(n_516), .Y(n_426) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_427), .B(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g427 ( .A(n_428), .B(n_453), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_441), .Y(n_429) );
AND2x2_ASAP7_75t_L g522 ( .A(n_430), .B(n_442), .Y(n_522) );
INVx3_ASAP7_75t_L g530 ( .A(n_430), .Y(n_530) );
AND2x2_ASAP7_75t_L g584 ( .A(n_430), .B(n_456), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_430), .B(n_455), .Y(n_620) );
AND2x2_ASAP7_75t_L g678 ( .A(n_430), .B(n_540), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_437), .B(n_439), .Y(n_435) );
INVx2_ASAP7_75t_L g449 ( .A(n_438), .Y(n_449) );
O2A1O1Ixp33_ASAP7_75t_L g462 ( .A1(n_439), .A2(n_449), .B(n_463), .C(n_464), .Y(n_462) );
AND2x2_ASAP7_75t_L g513 ( .A(n_441), .B(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g527 ( .A(n_441), .B(n_456), .Y(n_527) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_442), .B(n_456), .Y(n_542) );
AND2x2_ASAP7_75t_L g554 ( .A(n_442), .B(n_530), .Y(n_554) );
OR2x2_ASAP7_75t_L g556 ( .A(n_442), .B(n_514), .Y(n_556) );
AND2x2_ASAP7_75t_L g591 ( .A(n_442), .B(n_514), .Y(n_591) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_442), .Y(n_636) );
INVx1_ASAP7_75t_L g644 ( .A(n_442), .Y(n_644) );
OAI21xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_447), .B(n_451), .Y(n_443) );
OAI221xp5_ASAP7_75t_L g561 ( .A1(n_453), .A2(n_562), .B1(n_566), .B2(n_570), .C(n_571), .Y(n_561) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g521 ( .A(n_454), .B(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_466), .Y(n_454) );
INVx2_ASAP7_75t_L g520 ( .A(n_455), .Y(n_520) );
AND2x2_ASAP7_75t_L g573 ( .A(n_455), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g592 ( .A(n_455), .B(n_530), .Y(n_592) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g655 ( .A(n_456), .B(n_530), .Y(n_655) );
AND2x2_ASAP7_75t_L g577 ( .A(n_466), .B(n_522), .Y(n_577) );
OAI322xp33_ASAP7_75t_L g645 ( .A1(n_466), .A2(n_601), .A3(n_646), .B1(n_648), .B2(n_651), .C1(n_653), .C2(n_657), .Y(n_645) );
INVx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NOR2x1_ASAP7_75t_L g528 ( .A(n_467), .B(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g541 ( .A(n_467), .Y(n_541) );
AND2x2_ASAP7_75t_L g650 ( .A(n_467), .B(n_530), .Y(n_650) );
AND2x2_ASAP7_75t_L g682 ( .A(n_467), .B(n_554), .Y(n_682) );
OR2x2_ASAP7_75t_L g685 ( .A(n_467), .B(n_686), .Y(n_685) );
AND2x4_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
INVx1_ASAP7_75t_L g515 ( .A(n_468), .Y(n_515) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_486), .Y(n_474) );
INVx1_ASAP7_75t_L g698 ( .A(n_475), .Y(n_698) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OR2x2_ASAP7_75t_L g505 ( .A(n_476), .B(n_493), .Y(n_505) );
INVx2_ASAP7_75t_L g538 ( .A(n_476), .Y(n_538) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g560 ( .A(n_477), .Y(n_560) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_477), .Y(n_568) );
OR2x2_ASAP7_75t_L g692 ( .A(n_477), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g517 ( .A(n_486), .B(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g557 ( .A(n_486), .B(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g609 ( .A(n_486), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_493), .Y(n_486) );
AND2x2_ASAP7_75t_L g506 ( .A(n_487), .B(n_507), .Y(n_506) );
NOR2xp67_ASAP7_75t_L g564 ( .A(n_487), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g618 ( .A(n_487), .B(n_508), .Y(n_618) );
OR2x2_ASAP7_75t_L g626 ( .A(n_487), .B(n_560), .Y(n_626) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx2_ASAP7_75t_L g535 ( .A(n_488), .Y(n_535) );
AND2x2_ASAP7_75t_L g545 ( .A(n_488), .B(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g569 ( .A(n_488), .B(n_493), .Y(n_569) );
AND2x2_ASAP7_75t_L g633 ( .A(n_488), .B(n_508), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_493), .B(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_493), .B(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g546 ( .A(n_493), .Y(n_546) );
INVx1_ASAP7_75t_L g551 ( .A(n_493), .Y(n_551) );
AND2x2_ASAP7_75t_L g563 ( .A(n_493), .B(n_564), .Y(n_563) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_493), .Y(n_641) );
INVx1_ASAP7_75t_L g693 ( .A(n_493), .Y(n_693) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_497), .B(n_498), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_506), .Y(n_503) );
AND2x2_ASAP7_75t_L g670 ( .A(n_504), .B(n_579), .Y(n_670) );
INVx2_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g597 ( .A(n_506), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g696 ( .A(n_506), .B(n_631), .Y(n_696) );
INVx1_ASAP7_75t_L g518 ( .A(n_507), .Y(n_518) );
AND2x2_ASAP7_75t_L g544 ( .A(n_507), .B(n_538), .Y(n_544) );
BUFx2_ASAP7_75t_L g603 ( .A(n_507), .Y(n_603) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_508), .Y(n_524) );
INVx1_ASAP7_75t_L g534 ( .A(n_508), .Y(n_534) );
NOR2xp67_ASAP7_75t_L g672 ( .A(n_512), .B(n_519), .Y(n_672) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AOI32xp33_ASAP7_75t_L g516 ( .A1(n_513), .A2(n_517), .A3(n_519), .B1(n_521), .B2(n_523), .Y(n_516) );
AND2x2_ASAP7_75t_L g656 ( .A(n_513), .B(n_529), .Y(n_656) );
AND2x2_ASAP7_75t_L g694 ( .A(n_513), .B(n_592), .Y(n_694) );
INVx1_ASAP7_75t_L g574 ( .A(n_514), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_518), .B(n_580), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_519), .B(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_519), .B(n_522), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g673 ( .A(n_519), .B(n_591), .Y(n_673) );
OR2x2_ASAP7_75t_L g687 ( .A(n_519), .B(n_556), .Y(n_687) );
INVx3_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g614 ( .A(n_520), .B(n_522), .Y(n_614) );
OR2x2_ASAP7_75t_L g623 ( .A(n_520), .B(n_610), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_522), .B(n_573), .Y(n_595) );
INVx2_ASAP7_75t_L g610 ( .A(n_524), .Y(n_610) );
OR2x2_ASAP7_75t_L g625 ( .A(n_524), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g640 ( .A(n_524), .B(n_641), .Y(n_640) );
A2O1A1Ixp33_ASAP7_75t_L g697 ( .A1(n_524), .A2(n_617), .B(n_698), .C(n_699), .Y(n_697) );
OAI321xp33_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_531), .A3(n_536), .B1(n_539), .B2(n_543), .C(n_547), .Y(n_525) );
INVx1_ASAP7_75t_L g638 ( .A(n_526), .Y(n_638) );
NAND2x1p5_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
AND2x2_ASAP7_75t_L g649 ( .A(n_527), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g601 ( .A(n_529), .Y(n_601) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_530), .B(n_644), .Y(n_661) );
OAI221xp5_ASAP7_75t_L g668 ( .A1(n_531), .A2(n_669), .B1(n_671), .B2(n_673), .C(n_674), .Y(n_668) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .Y(n_532) );
AND2x2_ASAP7_75t_L g606 ( .A(n_533), .B(n_580), .Y(n_606) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_534), .B(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g579 ( .A(n_535), .Y(n_579) );
A2O1A1Ixp33_ASAP7_75t_L g621 ( .A1(n_536), .A2(n_577), .B(n_622), .C(n_624), .Y(n_621) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g588 ( .A(n_538), .B(n_545), .Y(n_588) );
BUFx2_ASAP7_75t_L g598 ( .A(n_538), .Y(n_598) );
INVx1_ASAP7_75t_L g613 ( .A(n_538), .Y(n_613) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
OR2x2_ASAP7_75t_L g619 ( .A(n_541), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g702 ( .A(n_541), .Y(n_702) );
INVx1_ASAP7_75t_L g695 ( .A(n_542), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
AND2x2_ASAP7_75t_L g548 ( .A(n_544), .B(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g652 ( .A(n_544), .B(n_569), .Y(n_652) );
INVx1_ASAP7_75t_L g581 ( .A(n_545), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_552), .B1(n_555), .B2(n_557), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_549), .B(n_665), .Y(n_664) );
INVxp67_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x4_ASAP7_75t_L g617 ( .A(n_550), .B(n_618), .Y(n_617) );
BUFx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_SL g580 ( .A(n_551), .B(n_560), .Y(n_580) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g572 ( .A(n_554), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g582 ( .A(n_556), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
OAI221xp5_ASAP7_75t_L g676 ( .A1(n_559), .A2(n_677), .B1(n_679), .B2(n_680), .C(n_681), .Y(n_676) );
INVx1_ASAP7_75t_L g565 ( .A(n_560), .Y(n_565) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_560), .Y(n_631) );
INVx1_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_563), .B(n_682), .Y(n_681) );
OAI21xp5_ASAP7_75t_L g571 ( .A1(n_564), .A2(n_569), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_567), .B(n_577), .Y(n_674) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
INVx1_ASAP7_75t_L g643 ( .A(n_568), .Y(n_643) );
AND2x2_ASAP7_75t_L g602 ( .A(n_569), .B(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g691 ( .A(n_569), .Y(n_691) );
INVx1_ASAP7_75t_L g607 ( .A(n_572), .Y(n_607) );
INVx1_ASAP7_75t_L g662 ( .A(n_573), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_578), .B1(n_581), .B2(n_582), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_579), .B(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g647 ( .A(n_580), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_580), .B(n_618), .Y(n_684) );
OR2x2_ASAP7_75t_L g657 ( .A(n_581), .B(n_610), .Y(n_657) );
INVx1_ASAP7_75t_L g596 ( .A(n_582), .Y(n_596) );
INVx1_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_584), .B(n_635), .Y(n_634) );
NOR3xp33_ASAP7_75t_L g585 ( .A(n_586), .B(n_604), .C(n_615), .Y(n_585) );
OAI211xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_589), .B(n_593), .C(n_599), .Y(n_586) );
INVxp67_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_588), .A2(n_659), .B1(n_663), .B2(n_666), .C(n_668), .Y(n_658) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
AND2x2_ASAP7_75t_L g600 ( .A(n_591), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g654 ( .A(n_591), .B(n_655), .Y(n_654) );
OAI211xp5_ASAP7_75t_L g639 ( .A1(n_592), .A2(n_640), .B(n_642), .C(n_644), .Y(n_639) );
INVx2_ASAP7_75t_L g686 ( .A(n_592), .Y(n_686) );
OAI21xp5_ASAP7_75t_SL g593 ( .A1(n_594), .A2(n_596), .B(n_597), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g665 ( .A(n_598), .B(n_618), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_602), .Y(n_599) );
OAI21xp5_ASAP7_75t_SL g604 ( .A1(n_605), .A2(n_607), .B(n_608), .Y(n_604) );
INVxp67_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OAI21xp5_ASAP7_75t_SL g608 ( .A1(n_609), .A2(n_611), .B(n_614), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_609), .B(n_638), .Y(n_637) );
INVxp67_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_614), .B(n_701), .Y(n_700) );
OAI21xp33_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_619), .B(n_621), .Y(n_615) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g642 ( .A(n_618), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND4x1_ASAP7_75t_L g627 ( .A(n_628), .B(n_658), .C(n_675), .D(n_697), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_629), .B(n_645), .Y(n_628) );
OAI211xp5_ASAP7_75t_SL g629 ( .A1(n_630), .A2(n_634), .B(n_637), .C(n_639), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
INVx1_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_633), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_644), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_654), .B(n_656), .Y(n_653) );
INVx1_ASAP7_75t_L g679 ( .A(n_654), .Y(n_679) );
INVx2_ASAP7_75t_SL g667 ( .A(n_655), .Y(n_667) );
OR2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g680 ( .A(n_665), .Y(n_680) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NOR2xp33_ASAP7_75t_SL g675 ( .A(n_676), .B(n_683), .Y(n_675) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
OAI221xp5_ASAP7_75t_SL g683 ( .A1(n_684), .A2(n_685), .B1(n_687), .B2(n_688), .C(n_689), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_694), .B1(n_695), .B2(n_696), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_691), .B(n_692), .Y(n_690) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g713 ( .A(n_704), .Y(n_713) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NOR2x2_ASAP7_75t_L g716 ( .A(n_706), .B(n_717), .Y(n_716) );
CKINVDCx14_ASAP7_75t_R g710 ( .A(n_707), .Y(n_710) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
NAND2xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_724), .Y(n_719) );
NOR2xp33_ASAP7_75t_SL g720 ( .A(n_721), .B(n_723), .Y(n_720) );
INVx1_ASAP7_75t_SL g741 ( .A(n_721), .Y(n_741) );
INVx1_ASAP7_75t_L g740 ( .A(n_723), .Y(n_740) );
OA21x2_ASAP7_75t_L g743 ( .A1(n_723), .A2(n_735), .B(n_741), .Y(n_743) );
INVx1_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
OAI21xp5_ASAP7_75t_L g727 ( .A1(n_725), .A2(n_728), .B(n_733), .Y(n_727) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
BUFx2_ASAP7_75t_L g735 ( .A(n_726), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_737), .Y(n_736) );
CKINVDCx6p67_ASAP7_75t_R g737 ( .A(n_738), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_741), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
endmodule