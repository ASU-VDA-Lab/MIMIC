module real_jpeg_7553_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_1),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_1),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_1),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_1),
.B(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_2),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_3),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_3),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_3),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_3),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_3),
.B(n_221),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_3),
.B(n_243),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_3),
.B(n_188),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_4),
.B(n_178),
.Y(n_177)
);

NAND2x1p5_ASAP7_75t_L g217 ( 
.A(n_4),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_4),
.B(n_259),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_4),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_4),
.B(n_298),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_4),
.B(n_330),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_4),
.B(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_5),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_5),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_5),
.B(n_145),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_5),
.B(n_187),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_5),
.B(n_273),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_5),
.B(n_281),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_5),
.B(n_325),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_5),
.B(n_350),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_6),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_6),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_6),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_6),
.B(n_241),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_6),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_6),
.B(n_316),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_6),
.B(n_352),
.Y(n_351)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_7),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_7),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g265 ( 
.A(n_7),
.Y(n_265)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_7),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_7),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_8),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_8),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_8),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_8),
.B(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_SL g186 ( 
.A(n_8),
.B(n_187),
.Y(n_186)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_10),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_10),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_10),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_10),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_10),
.B(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_SL g235 ( 
.A(n_10),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_10),
.B(n_188),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_10),
.B(n_358),
.Y(n_357)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_11),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_11),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g344 ( 
.A(n_11),
.Y(n_344)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_12),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_13),
.Y(n_88)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_13),
.Y(n_179)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_13),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_14),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_14),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_14),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_14),
.B(n_284),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_14),
.B(n_55),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_14),
.B(n_145),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_14),
.B(n_344),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_15),
.Y(n_97)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_15),
.Y(n_238)
);

BUFx5_ASAP7_75t_L g281 ( 
.A(n_15),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_16),
.B(n_39),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_16),
.B(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_16),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_16),
.B(n_145),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_16),
.B(n_275),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_16),
.B(n_292),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_16),
.B(n_241),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_17),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_17),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_17),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_17),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_17),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_17),
.B(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_194),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_193),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_150),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_23),
.B(n_150),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_89),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_62),
.C(n_75),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_25),
.B(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_41),
.C(n_48),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_26),
.B(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_36),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_28),
.B(n_33),
.C(n_36),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_28),
.A2(n_29),
.B1(n_44),
.B2(n_172),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_42),
.C(n_44),
.Y(n_41)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_32),
.A2(n_33),
.B1(n_94),
.B2(n_115),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_33),
.B(n_92),
.C(n_94),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_35),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_35),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_38),
.Y(n_218)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_41),
.B(n_48),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_42),
.B(n_171),
.Y(n_170)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_43),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_44),
.Y(n_172)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_46),
.Y(n_273)
);

INVx8_ASAP7_75t_L g292 ( 
.A(n_46),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_47),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_53),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_49),
.B(n_54),
.C(n_57),
.Y(n_124)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_56),
.Y(n_141)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_56),
.Y(n_330)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_60),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_60),
.Y(n_241)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_61),
.Y(n_285)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_61),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_61),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_62),
.B(n_75),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_63),
.B(n_69),
.C(n_74),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_69),
.B1(n_70),
.B2(n_74),
.Y(n_64)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_69),
.A2(n_70),
.B1(n_85),
.B2(n_86),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_76),
.C(n_85),
.Y(n_75)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_77),
.B(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.C(n_82),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_78),
.B(n_82),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_79),
.B(n_159),
.Y(n_158)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_119),
.B1(n_148),
.B2(n_149),
.Y(n_89)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

BUFx24_ASAP7_75t_SL g429 ( 
.A(n_90),
.Y(n_429)
);

FAx1_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_98),
.CI(n_110),
.CON(n_90),
.SN(n_90)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_112),
.B1(n_113),
.B2(n_115),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_97),
.Y(n_190)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_97),
.Y(n_245)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_97),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.C(n_107),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_99),
.B(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_107),
.Y(n_123)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_116),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_127),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.C(n_125),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_122),
.B1(n_124),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.Y(n_131)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_142),
.B2(n_147),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_141),
.Y(n_225)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_142),
.Y(n_147)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_146),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.C(n_156),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_151),
.B(n_153),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_156),
.B(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_173),
.C(n_175),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_157),
.B(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.C(n_170),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_158),
.B(n_413),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_160),
.A2(n_161),
.B1(n_170),
.B2(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.C(n_168),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_162),
.B(n_168),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_164),
.B(n_403),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_170),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_175),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_189),
.C(n_191),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_176),
.B(n_228),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_180),
.C(n_186),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_177),
.B(n_210),
.Y(n_209)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_186),
.Y(n_210)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_184),
.Y(n_259)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_191),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_247),
.B(n_428),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_196),
.B(n_198),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.C(n_205),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_200),
.B(n_203),
.Y(n_423)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_205),
.B(n_423),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_226),
.C(n_229),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_207),
.B(n_416),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.C(n_215),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_208),
.A2(n_209),
.B1(n_394),
.B2(n_395),
.Y(n_393)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_211),
.A2(n_212),
.B(n_214),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_211),
.B(n_215),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_214),
.Y(n_211)
);

MAJx2_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.C(n_223),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_371)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx8_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_223),
.B(n_371),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_224),
.B(n_311),
.Y(n_310)
);

INVx6_ASAP7_75t_L g350 ( 
.A(n_225),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g416 ( 
.A1(n_226),
.A2(n_227),
.B1(n_229),
.B2(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_229),
.Y(n_417)
);

MAJx2_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_242),
.C(n_246),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_231),
.B(n_405),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_235),
.C(n_239),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_232),
.B(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_235),
.A2(n_239),
.B1(n_240),
.B2(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_235),
.Y(n_384)
);

INVx8_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_237),
.Y(n_262)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_238),
.Y(n_311)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_242),
.B(n_246),
.Y(n_405)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

AOI21x1_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_421),
.B(n_427),
.Y(n_247)
);

OAI21x1_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_408),
.B(n_420),
.Y(n_248)
);

AOI21x1_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_390),
.B(n_407),
.Y(n_249)
);

OAI21x1_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_364),
.B(n_389),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_334),
.B(n_363),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_303),
.B(n_333),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_287),
.B(n_302),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_267),
.B(n_286),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_263),
.B(n_266),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_261),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_261),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_264),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_260),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_269),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_277),
.B2(n_278),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_270),
.B(n_280),
.C(n_282),
.Y(n_301)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_274),
.Y(n_295)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_282),
.B2(n_283),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_301),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_301),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_296),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_295),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_295),
.C(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_293),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_293),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_296),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g430 ( 
.A(n_296),
.Y(n_430)
);

FAx1_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.CI(n_300),
.CON(n_296),
.SN(n_296)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_297),
.B(n_321),
.C(n_322),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_299),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_300),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_306),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_304),
.B(n_306),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_319),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_307),
.B(n_320),
.C(n_323),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_308),
.B(n_310),
.C(n_312),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_312),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_315),
.B2(n_318),
.Y(n_312)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_313),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_314),
.B(n_318),
.Y(n_345)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_323),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_327),
.Y(n_323)
);

MAJx2_ASAP7_75t_L g361 ( 
.A(n_324),
.B(n_329),
.C(n_331),
.Y(n_361)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_328),
.A2(n_329),
.B1(n_331),
.B2(n_332),
.Y(n_327)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_328),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_329),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_362),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_335),
.B(n_362),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_347),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_346),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_337),
.B(n_346),
.C(n_388),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_345),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_343),
.Y(n_338)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_339),
.Y(n_378)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

CKINVDCx14_ASAP7_75t_R g379 ( 
.A(n_343),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_345),
.B(n_378),
.C(n_379),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_347),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_354),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_348),
.B(n_356),
.C(n_360),
.Y(n_367)
);

BUFx24_ASAP7_75t_SL g431 ( 
.A(n_348),
.Y(n_431)
);

FAx1_ASAP7_75t_SL g348 ( 
.A(n_349),
.B(n_351),
.CI(n_353),
.CON(n_348),
.SN(n_348)
);

MAJx2_ASAP7_75t_L g375 ( 
.A(n_349),
.B(n_351),
.C(n_353),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_356),
.B1(n_360),
.B2(n_361),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_359),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_357),
.B(n_359),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_361),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_387),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_365),
.B(n_387),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_376),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_367),
.B(n_368),
.C(n_376),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_369),
.A2(n_370),
.B1(n_372),
.B2(n_373),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_369),
.B(n_399),
.C(n_400),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_374),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_375),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_377),
.B(n_380),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_377),
.B(n_381),
.C(n_386),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_382),
.B1(n_385),
.B2(n_386),
.Y(n_380)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_381),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_382),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_391),
.B(n_406),
.Y(n_390)
);

NOR2xp67_ASAP7_75t_SL g407 ( 
.A(n_391),
.B(n_406),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_392),
.B(n_397),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_396),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_393),
.B(n_396),
.C(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_394),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_397),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_398),
.B(n_401),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_398),
.B(n_402),
.C(n_404),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_404),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_409),
.B(n_418),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_409),
.B(n_418),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_410),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_415),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_412),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_415),
.B(n_425),
.C(n_426),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_422),
.B(n_424),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_422),
.B(n_424),
.Y(n_427)
);


endmodule