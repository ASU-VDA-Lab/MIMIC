module fake_netlist_6_2267_n_4424 (n_992, n_52, n_591, n_435, n_1, n_91, n_793, n_326, n_801, n_256, n_853, n_440, n_587, n_695, n_507, n_968, n_909, n_580, n_762, n_1030, n_881, n_875, n_209, n_367, n_465, n_680, n_741, n_760, n_1008, n_1027, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_828, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_1033, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_933, n_740, n_578, n_703, n_1003, n_144, n_365, n_978, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_820, n_951, n_783, n_106, n_725, n_952, n_999, n_358, n_160, n_751, n_449, n_131, n_749, n_798, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_994, n_677, n_969, n_988, n_805, n_396, n_495, n_815, n_350, n_78, n_84, n_585, n_732, n_974, n_568, n_392, n_840, n_442, n_480, n_142, n_874, n_724, n_143, n_382, n_673, n_1020, n_180, n_1009, n_62, n_628, n_883, n_557, n_823, n_349, n_643, n_233, n_617, n_698, n_898, n_1032, n_845, n_255, n_807, n_1036, n_739, n_284, n_400, n_140, n_337, n_955, n_865, n_893, n_214, n_925, n_485, n_67, n_15, n_1026, n_443, n_246, n_892, n_768, n_38, n_471, n_289, n_935, n_421, n_781, n_424, n_789, n_615, n_59, n_181, n_182, n_238, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_794, n_963, n_727, n_894, n_369, n_597, n_685, n_280, n_287, n_832, n_353, n_610, n_555, n_389, n_814, n_415, n_830, n_65, n_230, n_605, n_461, n_873, n_141, n_383, n_826, n_1024, n_669, n_200, n_447, n_176, n_872, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_1018, n_747, n_852, n_667, n_71, n_74, n_229, n_542, n_847, n_644, n_682, n_851, n_621, n_305, n_72, n_721, n_996, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_901, n_111, n_504, n_923, n_314, n_378, n_413, n_377, n_791, n_35, n_183, n_510, n_837, n_836, n_1015, n_79, n_863, n_375, n_601, n_338, n_522, n_948, n_466, n_704, n_918, n_748, n_506, n_56, n_763, n_360, n_945, n_977, n_603, n_1005, n_119, n_991, n_957, n_235, n_536, n_895, n_866, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_744, n_971, n_946, n_39, n_344, n_73, n_581, n_428, n_761, n_785, n_746, n_609, n_765, n_432, n_987, n_641, n_822, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_842, n_611, n_943, n_156, n_491, n_878, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_843, n_989, n_797, n_666, n_1016, n_371, n_795, n_770, n_940, n_567, n_899, n_189, n_738, n_405, n_213, n_538, n_1035, n_294, n_302, n_499, n_380, n_838, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_844, n_448, n_886, n_953, n_20, n_1004, n_1017, n_494, n_539, n_493, n_397, n_155, n_1022, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_930, n_888, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_910, n_37, n_486, n_911, n_381, n_82, n_947, n_27, n_236, n_653, n_887, n_752, n_908, n_112, n_172, n_944, n_713, n_648, n_657, n_576, n_1028, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_782, n_976, n_490, n_803, n_290, n_220, n_809, n_1011, n_118, n_224, n_48, n_926, n_927, n_25, n_93, n_839, n_986, n_80, n_734, n_708, n_196, n_919, n_402, n_352, n_917, n_668, n_478, n_626, n_990, n_574, n_779, n_9, n_800, n_929, n_460, n_107, n_907, n_854, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_870, n_366, n_904, n_777, n_407, n_913, n_450, n_103, n_808, n_867, n_272, n_526, n_921, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_937, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_998, n_16, n_163, n_717, n_46, n_330, n_771, n_470, n_475, n_924, n_298, n_18, n_492, n_972, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_824, n_962, n_1000, n_279, n_686, n_796, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_936, n_184, n_552, n_619, n_885, n_216, n_455, n_896, n_83, n_521, n_363, n_572, n_912, n_395, n_813, n_592, n_745, n_654, n_323, n_829, n_606, n_393, n_818, n_984, n_411, n_503, n_716, n_152, n_623, n_92, n_884, n_599, n_513, n_855, n_776, n_321, n_645, n_331, n_105, n_916, n_227, n_132, n_868, n_570, n_731, n_859, n_406, n_483, n_735, n_102, n_204, n_482, n_934, n_755, n_931, n_1021, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_958, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_942, n_792, n_880, n_476, n_981, n_714, n_2, n_291, n_219, n_543, n_889, n_357, n_150, n_264, n_263, n_985, n_589, n_860, n_481, n_788, n_819, n_939, n_997, n_821, n_325, n_938, n_767, n_804, n_329, n_464, n_600, n_831, n_802, n_964, n_982, n_561, n_33, n_477, n_549, n_980, n_533, n_954, n_408, n_932, n_806, n_864, n_879, n_959, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_979, n_548, n_905, n_94, n_282, n_436, n_833, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_993, n_345, n_409, n_231, n_354, n_689, n_40, n_799, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_810, n_635, n_95, n_787, n_311, n_10, n_403, n_723, n_253, n_634, n_583, n_596, n_123, n_136, n_966, n_546, n_562, n_249, n_201, n_386, n_764, n_556, n_159, n_1034, n_157, n_162, n_692, n_733, n_754, n_941, n_975, n_1031, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_849, n_970, n_560, n_1014, n_753, n_642, n_995, n_276, n_569, n_441, n_221, n_811, n_882, n_444, n_586, n_423, n_146, n_737, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_973, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_1029, n_418, n_113, n_618, n_790, n_582, n_4, n_199, n_138, n_266, n_296, n_861, n_674, n_857, n_871, n_967, n_775, n_922, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_902, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_914, n_759, n_1010, n_355, n_426, n_317, n_149, n_915, n_632, n_702, n_431, n_90, n_347, n_812, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_1006, n_373, n_1012, n_87, n_195, n_285, n_497, n_780, n_773, n_675, n_903, n_85, n_99, n_257, n_920, n_730, n_655, n_13, n_706, n_786, n_670, n_203, n_286, n_254, n_207, n_834, n_242, n_835, n_928, n_19, n_47, n_690, n_29, n_850, n_75, n_401, n_324, n_743, n_766, n_816, n_335, n_430, n_1002, n_463, n_545, n_489, n_877, n_205, n_604, n_848, n_120, n_251, n_1019, n_301, n_274, n_636, n_825, n_728, n_681, n_729, n_110, n_151, n_876, n_774, n_412, n_640, n_81, n_660, n_965, n_36, n_26, n_55, n_267, n_438, n_339, n_784, n_315, n_434, n_515, n_983, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_906, n_688, n_722, n_961, n_862, n_135, n_165, n_351, n_869, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_890, n_637, n_295, n_385, n_701, n_817, n_950, n_629, n_388, n_190, n_858, n_262, n_484, n_613, n_736, n_187, n_897, n_900, n_846, n_501, n_841, n_956, n_960, n_531, n_827, n_1001, n_60, n_361, n_508, n_663, n_856, n_379, n_170, n_778, n_1025, n_332, n_891, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_1013, n_1023, n_194, n_664, n_171, n_949, n_678, n_192, n_57, n_169, n_1007, n_51, n_649, n_283, n_4424);

input n_992;
input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_793;
input n_326;
input n_801;
input n_256;
input n_853;
input n_440;
input n_587;
input n_695;
input n_507;
input n_968;
input n_909;
input n_580;
input n_762;
input n_1030;
input n_881;
input n_875;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_1008;
input n_1027;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_828;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_1033;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_933;
input n_740;
input n_578;
input n_703;
input n_1003;
input n_144;
input n_365;
input n_978;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_820;
input n_951;
input n_783;
input n_106;
input n_725;
input n_952;
input n_999;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_798;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_994;
input n_677;
input n_969;
input n_988;
input n_805;
input n_396;
input n_495;
input n_815;
input n_350;
input n_78;
input n_84;
input n_585;
input n_732;
input n_974;
input n_568;
input n_392;
input n_840;
input n_442;
input n_480;
input n_142;
input n_874;
input n_724;
input n_143;
input n_382;
input n_673;
input n_1020;
input n_180;
input n_1009;
input n_62;
input n_628;
input n_883;
input n_557;
input n_823;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_898;
input n_1032;
input n_845;
input n_255;
input n_807;
input n_1036;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_955;
input n_865;
input n_893;
input n_214;
input n_925;
input n_485;
input n_67;
input n_15;
input n_1026;
input n_443;
input n_246;
input n_892;
input n_768;
input n_38;
input n_471;
input n_289;
input n_935;
input n_421;
input n_781;
input n_424;
input n_789;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_794;
input n_963;
input n_727;
input n_894;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_832;
input n_353;
input n_610;
input n_555;
input n_389;
input n_814;
input n_415;
input n_830;
input n_65;
input n_230;
input n_605;
input n_461;
input n_873;
input n_141;
input n_383;
input n_826;
input n_1024;
input n_669;
input n_200;
input n_447;
input n_176;
input n_872;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_1018;
input n_747;
input n_852;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_621;
input n_305;
input n_72;
input n_721;
input n_996;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_901;
input n_111;
input n_504;
input n_923;
input n_314;
input n_378;
input n_413;
input n_377;
input n_791;
input n_35;
input n_183;
input n_510;
input n_837;
input n_836;
input n_1015;
input n_79;
input n_863;
input n_375;
input n_601;
input n_338;
input n_522;
input n_948;
input n_466;
input n_704;
input n_918;
input n_748;
input n_506;
input n_56;
input n_763;
input n_360;
input n_945;
input n_977;
input n_603;
input n_1005;
input n_119;
input n_991;
input n_957;
input n_235;
input n_536;
input n_895;
input n_866;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_971;
input n_946;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_761;
input n_785;
input n_746;
input n_609;
input n_765;
input n_432;
input n_987;
input n_641;
input n_822;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_842;
input n_611;
input n_943;
input n_156;
input n_491;
input n_878;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_843;
input n_989;
input n_797;
input n_666;
input n_1016;
input n_371;
input n_795;
input n_770;
input n_940;
input n_567;
input n_899;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_1035;
input n_294;
input n_302;
input n_499;
input n_380;
input n_838;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_844;
input n_448;
input n_886;
input n_953;
input n_20;
input n_1004;
input n_1017;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_1022;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_930;
input n_888;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_910;
input n_37;
input n_486;
input n_911;
input n_381;
input n_82;
input n_947;
input n_27;
input n_236;
input n_653;
input n_887;
input n_752;
input n_908;
input n_112;
input n_172;
input n_944;
input n_713;
input n_648;
input n_657;
input n_576;
input n_1028;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_782;
input n_976;
input n_490;
input n_803;
input n_290;
input n_220;
input n_809;
input n_1011;
input n_118;
input n_224;
input n_48;
input n_926;
input n_927;
input n_25;
input n_93;
input n_839;
input n_986;
input n_80;
input n_734;
input n_708;
input n_196;
input n_919;
input n_402;
input n_352;
input n_917;
input n_668;
input n_478;
input n_626;
input n_990;
input n_574;
input n_779;
input n_9;
input n_800;
input n_929;
input n_460;
input n_107;
input n_907;
input n_854;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_870;
input n_366;
input n_904;
input n_777;
input n_407;
input n_913;
input n_450;
input n_103;
input n_808;
input n_867;
input n_272;
input n_526;
input n_921;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_937;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_998;
input n_16;
input n_163;
input n_717;
input n_46;
input n_330;
input n_771;
input n_470;
input n_475;
input n_924;
input n_298;
input n_18;
input n_492;
input n_972;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_824;
input n_962;
input n_1000;
input n_279;
input n_686;
input n_796;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_936;
input n_184;
input n_552;
input n_619;
input n_885;
input n_216;
input n_455;
input n_896;
input n_83;
input n_521;
input n_363;
input n_572;
input n_912;
input n_395;
input n_813;
input n_592;
input n_745;
input n_654;
input n_323;
input n_829;
input n_606;
input n_393;
input n_818;
input n_984;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_92;
input n_884;
input n_599;
input n_513;
input n_855;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_916;
input n_227;
input n_132;
input n_868;
input n_570;
input n_731;
input n_859;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_934;
input n_755;
input n_931;
input n_1021;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_958;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_942;
input n_792;
input n_880;
input n_476;
input n_981;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_889;
input n_357;
input n_150;
input n_264;
input n_263;
input n_985;
input n_589;
input n_860;
input n_481;
input n_788;
input n_819;
input n_939;
input n_997;
input n_821;
input n_325;
input n_938;
input n_767;
input n_804;
input n_329;
input n_464;
input n_600;
input n_831;
input n_802;
input n_964;
input n_982;
input n_561;
input n_33;
input n_477;
input n_549;
input n_980;
input n_533;
input n_954;
input n_408;
input n_932;
input n_806;
input n_864;
input n_879;
input n_959;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_979;
input n_548;
input n_905;
input n_94;
input n_282;
input n_436;
input n_833;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_993;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_799;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_810;
input n_635;
input n_95;
input n_787;
input n_311;
input n_10;
input n_403;
input n_723;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_966;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_764;
input n_556;
input n_159;
input n_1034;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_941;
input n_975;
input n_1031;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_849;
input n_970;
input n_560;
input n_1014;
input n_753;
input n_642;
input n_995;
input n_276;
input n_569;
input n_441;
input n_221;
input n_811;
input n_882;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_973;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_1029;
input n_418;
input n_113;
input n_618;
input n_790;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_861;
input n_674;
input n_857;
input n_871;
input n_967;
input n_775;
input n_922;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_902;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_914;
input n_759;
input n_1010;
input n_355;
input n_426;
input n_317;
input n_149;
input n_915;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_812;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_1006;
input n_373;
input n_1012;
input n_87;
input n_195;
input n_285;
input n_497;
input n_780;
input n_773;
input n_675;
input n_903;
input n_85;
input n_99;
input n_257;
input n_920;
input n_730;
input n_655;
input n_13;
input n_706;
input n_786;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_834;
input n_242;
input n_835;
input n_928;
input n_19;
input n_47;
input n_690;
input n_29;
input n_850;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_816;
input n_335;
input n_430;
input n_1002;
input n_463;
input n_545;
input n_489;
input n_877;
input n_205;
input n_604;
input n_848;
input n_120;
input n_251;
input n_1019;
input n_301;
input n_274;
input n_636;
input n_825;
input n_728;
input n_681;
input n_729;
input n_110;
input n_151;
input n_876;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_965;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_784;
input n_315;
input n_434;
input n_515;
input n_983;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_906;
input n_688;
input n_722;
input n_961;
input n_862;
input n_135;
input n_165;
input n_351;
input n_869;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_890;
input n_637;
input n_295;
input n_385;
input n_701;
input n_817;
input n_950;
input n_629;
input n_388;
input n_190;
input n_858;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_897;
input n_900;
input n_846;
input n_501;
input n_841;
input n_956;
input n_960;
input n_531;
input n_827;
input n_1001;
input n_60;
input n_361;
input n_508;
input n_663;
input n_856;
input n_379;
input n_170;
input n_778;
input n_1025;
input n_332;
input n_891;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_1013;
input n_1023;
input n_194;
input n_664;
input n_171;
input n_949;
input n_678;
input n_192;
input n_57;
input n_169;
input n_1007;
input n_51;
input n_649;
input n_283;

output n_4424;

wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_3766;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_3254;
wire n_3684;
wire n_1199;
wire n_1674;
wire n_3392;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_3152;
wire n_4154;
wire n_3579;
wire n_1212;
wire n_4251;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3773;
wire n_3783;
wire n_4177;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_4127;
wire n_1038;
wire n_1581;
wire n_3844;
wire n_4388;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_4395;
wire n_4099;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_3741;
wire n_4168;
wire n_4372;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_2324;
wire n_1854;
wire n_1575;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_2260;
wire n_1387;
wire n_3222;
wire n_1708;
wire n_1151;
wire n_2977;
wire n_3952;
wire n_1739;
wire n_2051;
wire n_4370;
wire n_2317;
wire n_1380;
wire n_3911;
wire n_2359;
wire n_2847;
wire n_2557;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_3332;
wire n_4134;
wire n_4285;
wire n_3465;
wire n_1975;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_3706;
wire n_4050;
wire n_1160;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_4092;
wire n_1724;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_4078;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_4249;
wire n_1264;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_3619;
wire n_4359;
wire n_4087;
wire n_1700;
wire n_1555;
wire n_2211;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_4302;
wire n_2291;
wire n_2299;
wire n_3340;
wire n_4179;
wire n_1371;
wire n_1285;
wire n_2886;
wire n_2974;
wire n_3946;
wire n_1985;
wire n_4213;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_2509;
wire n_4065;
wire n_4026;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_3904;
wire n_4178;
wire n_1393;
wire n_1867;
wire n_1517;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_2247;
wire n_1711;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_4273;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_4029;
wire n_3345;
wire n_2074;
wire n_4417;
wire n_2447;
wire n_2919;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_3879;
wire n_4010;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1772;
wire n_1232;
wire n_1572;
wire n_3979;
wire n_4308;
wire n_1874;
wire n_4347;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_2510;
wire n_2739;
wire n_1541;
wire n_1300;
wire n_2480;
wire n_3023;
wire n_3890;
wire n_3232;
wire n_2791;
wire n_1313;
wire n_3750;
wire n_3607;
wire n_4325;
wire n_3251;
wire n_1056;
wire n_3877;
wire n_3316;
wire n_2212;
wire n_3929;
wire n_3494;
wire n_3048;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_2729;
wire n_1163;
wire n_3063;
wire n_4311;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_1798;
wire n_4060;
wire n_1550;
wire n_2703;
wire n_3998;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_4187;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_4164;
wire n_2004;
wire n_1106;
wire n_1471;
wire n_1094;
wire n_3624;
wire n_3077;
wire n_3737;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3655;
wire n_3107;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_4117;
wire n_3948;
wire n_2836;
wire n_1421;
wire n_3664;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_1660;
wire n_4327;
wire n_1961;
wire n_3047;
wire n_4414;
wire n_1280;
wire n_3765;
wire n_2655;
wire n_4125;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_4221;
wire n_1467;
wire n_3297;
wire n_4250;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_3906;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_1088;
wire n_4262;
wire n_4392;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3963;
wire n_3368;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_2591;
wire n_3507;
wire n_4334;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_4253;
wire n_4110;
wire n_1658;
wire n_2593;
wire n_4071;
wire n_4255;
wire n_4403;
wire n_3506;
wire n_4268;
wire n_3568;
wire n_3269;
wire n_4047;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_1967;
wire n_1193;
wire n_3999;
wire n_1054;
wire n_3928;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_4139;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_1986;
wire n_3943;
wire n_4320;
wire n_4305;
wire n_2397;
wire n_3884;
wire n_3931;
wire n_4349;
wire n_4102;
wire n_4297;
wire n_2113;
wire n_1641;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_3871;
wire n_2907;
wire n_3438;
wire n_2735;
wire n_4141;
wire n_1843;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_4227;
wire n_2850;
wire n_4314;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_3822;
wire n_4163;
wire n_1441;
wire n_3373;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_1699;
wire n_3910;
wire n_3934;
wire n_2093;
wire n_4033;
wire n_4415;
wire n_4296;
wire n_4009;
wire n_2633;
wire n_3883;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_3728;
wire n_2669;
wire n_2925;
wire n_4094;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_2522;
wire n_3949;
wire n_4364;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_4354;
wire n_2616;
wire n_3912;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_3923;
wire n_2529;
wire n_3900;
wire n_4393;
wire n_1162;
wire n_1530;
wire n_3798;
wire n_3488;
wire n_1543;
wire n_2811;
wire n_1302;
wire n_1599;
wire n_1068;
wire n_3732;
wire n_4257;
wire n_2674;
wire n_2832;
wire n_4226;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_2831;
wire n_2998;
wire n_4318;
wire n_4377;
wire n_3446;
wire n_4158;
wire n_4366;
wire n_3317;
wire n_3857;
wire n_3978;
wire n_1876;
wire n_4107;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_4074;
wire n_3716;
wire n_1873;
wire n_4294;
wire n_3630;
wire n_3518;
wire n_3824;
wire n_3859;
wire n_1866;
wire n_4013;
wire n_2692;
wire n_1680;
wire n_3842;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3914;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_4032;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_2355;
wire n_3927;
wire n_4147;
wire n_3888;
wire n_2908;
wire n_3168;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_4130;
wire n_4161;
wire n_4337;
wire n_2895;
wire n_2009;
wire n_4172;
wire n_3403;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_3882;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_3055;
wire n_3092;
wire n_3492;
wire n_3895;
wire n_3966;
wire n_4369;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_3734;
wire n_4331;
wire n_3686;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_4118;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_2459;
wire n_3746;
wire n_1111;
wire n_2971;
wire n_1713;
wire n_4375;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_3935;
wire n_1265;
wire n_4277;
wire n_2711;
wire n_3490;
wire n_4291;
wire n_4199;
wire n_1950;
wire n_1726;
wire n_1912;
wire n_1563;
wire n_2434;
wire n_4319;
wire n_3369;
wire n_3419;
wire n_1982;
wire n_3872;
wire n_2878;
wire n_3012;
wire n_3772;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3875;
wire n_1167;
wire n_2818;
wire n_1359;
wire n_2428;
wire n_3581;
wire n_3794;
wire n_3247;
wire n_3069;
wire n_3921;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_2641;
wire n_1722;
wire n_1664;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_3933;
wire n_2749;
wire n_2008;
wire n_3298;
wire n_2192;
wire n_3346;
wire n_2345;
wire n_2254;
wire n_3281;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_2311;
wire n_1386;
wire n_1896;
wire n_2965;
wire n_3058;
wire n_1747;
wire n_3691;
wire n_3861;
wire n_2624;
wire n_4066;
wire n_4386;
wire n_4146;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_4340;
wire n_3891;
wire n_2193;
wire n_3961;
wire n_2676;
wire n_1655;
wire n_3940;
wire n_4072;
wire n_4220;
wire n_1801;
wire n_1214;
wire n_2347;
wire n_1886;
wire n_2092;
wire n_3917;
wire n_1654;
wire n_4371;
wire n_1157;
wire n_3453;
wire n_2994;
wire n_1750;
wire n_1462;
wire n_3410;
wire n_3153;
wire n_3428;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_4004;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_4043;
wire n_4313;
wire n_4353;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_4292;
wire n_1588;
wire n_3785;
wire n_3942;
wire n_3997;
wire n_2963;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_4381;
wire n_1124;
wire n_1624;
wire n_3873;
wire n_3983;
wire n_2096;
wire n_2980;
wire n_3968;
wire n_4418;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_3434;
wire n_1515;
wire n_4356;
wire n_3510;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_4169;
wire n_4055;
wire n_2377;
wire n_3271;
wire n_2178;
wire n_4362;
wire n_4248;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_3009;
wire n_1709;
wire n_2652;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_4361;
wire n_2393;
wire n_1796;
wire n_1757;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_3889;
wire n_2687;
wire n_3237;
wire n_1630;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_3707;
wire n_2075;
wire n_4045;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_4367;
wire n_2763;
wire n_2762;
wire n_4070;
wire n_1987;
wire n_3545;
wire n_1369;
wire n_3578;
wire n_3885;
wire n_2271;
wire n_3192;
wire n_3993;
wire n_1546;
wire n_2583;
wire n_4394;
wire n_4116;
wire n_2606;
wire n_4031;
wire n_2279;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_3073;
wire n_2431;
wire n_4018;
wire n_2987;
wire n_2938;
wire n_2150;
wire n_2943;
wire n_1294;
wire n_1420;
wire n_3696;
wire n_3780;
wire n_4082;
wire n_2078;
wire n_1634;
wire n_3252;
wire n_2932;
wire n_1767;
wire n_3253;
wire n_1779;
wire n_1465;
wire n_3337;
wire n_3431;
wire n_3450;
wire n_4002;
wire n_3209;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_4329;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_2750;
wire n_2558;
wire n_2893;
wire n_1523;
wire n_2775;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1735;
wire n_2954;
wire n_3477;
wire n_4288;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_4289;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_3953;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_3421;
wire n_2913;
wire n_3614;
wire n_1756;
wire n_3183;
wire n_2493;
wire n_1128;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_4019;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_4385;
wire n_1952;
wire n_3616;
wire n_4228;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_4044;
wire n_3436;
wire n_1932;
wire n_1101;
wire n_1880;
wire n_2535;
wire n_3366;
wire n_3442;
wire n_2631;
wire n_4191;
wire n_1364;
wire n_4322;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_3937;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_4287;
wire n_1293;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_3941;
wire n_2767;
wire n_3793;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_1514;
wire n_1863;
wire n_3385;
wire n_4350;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_1714;
wire n_1139;
wire n_3922;
wire n_3179;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_4330;
wire n_2897;
wire n_2537;
wire n_3970;
wire n_4389;
wire n_4345;
wire n_2554;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_2747;
wire n_1513;
wire n_3924;
wire n_3171;
wire n_1913;
wire n_4216;
wire n_3608;
wire n_4315;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_4156;
wire n_3491;
wire n_4240;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_2148;
wire n_4284;
wire n_4162;
wire n_2339;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_2643;
wire n_2590;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_3782;
wire n_3975;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_4011;
wire n_1835;
wire n_3470;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_4098;
wire n_4021;
wire n_1492;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_4058;
wire n_4103;
wire n_3104;
wire n_3435;
wire n_3148;
wire n_2262;
wire n_3348;
wire n_3229;
wire n_4022;
wire n_2239;
wire n_3082;
wire n_1707;
wire n_3611;
wire n_4310;
wire n_1432;
wire n_2208;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_2717;
wire n_1723;
wire n_1246;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_3580;
wire n_3775;
wire n_3537;
wire n_1176;
wire n_2134;
wire n_2335;
wire n_1529;
wire n_2473;
wire n_3887;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_4123;
wire n_1431;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_3835;
wire n_4286;
wire n_1809;
wire n_3119;
wire n_4280;
wire n_2958;
wire n_2948;
wire n_3735;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_4379;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1448;
wire n_1087;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_1049;
wire n_3223;
wire n_3996;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_4097;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_4218;
wire n_4402;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_3880;
wire n_1849;
wire n_2848;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_4100;
wire n_2231;
wire n_3609;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_4264;
wire n_2857;
wire n_3693;
wire n_3788;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_1299;
wire n_2896;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_4079;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_4175;
wire n_3200;
wire n_1665;
wire n_4306;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_4224;
wire n_3390;
wire n_3656;
wire n_4339;
wire n_1178;
wire n_2127;
wire n_2338;
wire n_1424;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_3867;
wire n_1073;
wire n_1195;
wire n_3559;
wire n_3025;
wire n_2137;
wire n_3191;
wire n_1626;
wire n_4005;
wire n_2482;
wire n_1507;
wire n_3810;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_2424;
wire n_2296;
wire n_1284;
wire n_3201;
wire n_3633;
wire n_1604;
wire n_3447;
wire n_3971;
wire n_1142;
wire n_2849;
wire n_1475;
wire n_1048;
wire n_1201;
wire n_2354;
wire n_1398;
wire n_2682;
wire n_3032;
wire n_3103;
wire n_3638;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_3393;
wire n_2442;
wire n_1207;
wire n_3627;
wire n_3451;
wire n_1791;
wire n_1368;
wire n_3480;
wire n_1418;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_4222;
wire n_2545;
wire n_3540;
wire n_3577;
wire n_4401;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_4368;
wire n_1478;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_2966;
wire n_2294;
wire n_2581;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_3591;
wire n_3641;
wire n_1837;
wire n_2218;
wire n_1314;
wire n_2788;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_4419;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_4120;
wire n_1382;
wire n_1534;
wire n_3892;
wire n_1736;
wire n_1564;
wire n_4069;
wire n_2748;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2860;
wire n_2292;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_3964;
wire n_1993;
wire n_2281;
wire n_4167;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_3944;
wire n_3909;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2323;
wire n_1220;
wire n_1893;
wire n_2784;
wire n_2301;
wire n_2209;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_4223;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_4387;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_3481;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_4299;
wire n_3033;
wire n_3724;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_1774;
wire n_1223;
wire n_3571;
wire n_3913;
wire n_4276;
wire n_2990;
wire n_3847;
wire n_1286;
wire n_1775;
wire n_2115;
wire n_1773;
wire n_2552;
wire n_2410;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_4348;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_2929;
wire n_1597;
wire n_2780;
wire n_3323;
wire n_3226;
wire n_3364;
wire n_4020;
wire n_4176;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_4404;
wire n_1153;
wire n_3407;
wire n_1618;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_2384;
wire n_3894;
wire n_4204;
wire n_4261;
wire n_1745;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_4063;
wire n_1625;
wire n_3986;
wire n_4237;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_1453;
wire n_2146;
wire n_4006;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_3646;
wire n_2920;
wire n_4015;
wire n_3547;
wire n_1901;
wire n_3869;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1892;
wire n_1459;
wire n_3188;
wire n_3742;
wire n_1614;
wire n_4410;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_4034;
wire n_1617;
wire n_4056;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_3960;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_3175;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_2732;
wire n_2928;
wire n_4206;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_3862;
wire n_4267;
wire n_1580;
wire n_2227;
wire n_4247;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_4180;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_3284;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_2720;
wire n_1520;
wire n_3126;
wire n_2159;
wire n_2289;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2863;
wire n_1390;
wire n_1419;
wire n_3299;
wire n_3663;
wire n_4132;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_3360;
wire n_2087;
wire n_1855;
wire n_3051;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_3956;
wire n_3367;
wire n_1832;
wire n_1645;
wire n_4001;
wire n_1687;
wire n_2328;
wire n_1439;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_2049;
wire n_4149;
wire n_1331;
wire n_2627;
wire n_4355;
wire n_2276;
wire n_3234;
wire n_4422;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_2993;
wire n_3016;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_4003;
wire n_4126;
wire n_1129;
wire n_3870;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_2181;
wire n_3751;
wire n_3845;
wire n_1869;
wire n_2911;
wire n_3625;
wire n_3804;
wire n_1594;
wire n_1764;
wire n_4207;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_4113;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_1202;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_2942;
wire n_1635;
wire n_4014;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_2139;
wire n_2142;
wire n_4067;
wire n_4252;
wire n_4357;
wire n_1551;
wire n_4028;
wire n_4054;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_3907;
wire n_2555;
wire n_4048;
wire n_3338;
wire n_4217;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_2327;
wire n_4374;
wire n_2201;
wire n_3919;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_2984;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_4024;
wire n_1508;
wire n_2487;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_2597;
wire n_2375;
wire n_3194;
wire n_3113;
wire n_3250;
wire n_1934;
wire n_3276;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_4214;
wire n_1728;
wire n_3973;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_4338;
wire n_3886;
wire n_2924;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_4420;
wire n_1510;
wire n_3637;
wire n_3120;
wire n_1468;
wire n_3991;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3797;
wire n_3926;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_2598;
wire n_1916;
wire n_1683;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_4405;
wire n_4234;
wire n_4304;
wire n_4413;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_4101;
wire n_3548;
wire n_3767;
wire n_3864;
wire n_4036;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_3974;
wire n_2052;
wire n_1847;
wire n_3634;
wire n_2302;
wire n_4211;
wire n_4182;
wire n_1667;
wire n_1206;
wire n_3230;
wire n_4016;
wire n_1037;
wire n_1397;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_3592;
wire n_2755;
wire n_3141;
wire n_1409;
wire n_4230;
wire n_1841;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_3967;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_4328;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_4274;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_2785;
wire n_1657;
wire n_4189;
wire n_4270;
wire n_4151;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_1818;
wire n_1108;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3730;
wire n_1298;
wire n_4124;
wire n_3659;
wire n_2559;
wire n_2595;
wire n_2177;
wire n_3399;
wire n_4397;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_4155;
wire n_2740;
wire n_4238;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_3042;
wire n_1356;
wire n_1589;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1943;
wire n_1216;
wire n_3228;
wire n_3249;
wire n_2716;
wire n_1320;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_4152;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_4406;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_3177;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_4380;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_4398;
wire n_2498;
wire n_4219;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_3238;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3529;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_4109;
wire n_4192;
wire n_1443;
wire n_2392;
wire n_1272;
wire n_2894;
wire n_3424;
wire n_3957;
wire n_4038;
wire n_2790;
wire n_4131;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_4195;
wire n_4159;
wire n_3784;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_1043;
wire n_3819;
wire n_4090;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_4144;
wire n_1870;
wire n_2964;
wire n_4174;
wire n_1692;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3501;
wire n_3475;
wire n_1840;
wire n_1152;
wire n_1705;
wire n_3905;
wire n_3262;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_4008;
wire n_2244;
wire n_4290;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_2789;
wire n_3105;
wire n_1352;
wire n_3210;
wire n_2872;
wire n_2257;
wire n_3692;
wire n_2017;
wire n_1682;
wire n_1828;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_4258;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_2376;
wire n_1405;
wire n_3826;
wire n_1406;
wire n_3790;
wire n_3878;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_4323;
wire n_1041;
wire n_2346;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_4300;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_3320;
wire n_2541;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_1974;
wire n_3988;
wire n_4122;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_1637;
wire n_2635;
wire n_3307;
wire n_3439;
wire n_3588;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_4135;
wire n_4209;
wire n_2871;
wire n_4279;
wire n_2688;
wire n_3858;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_4183;
wire n_1489;
wire n_4321;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_4128;
wire n_2229;
wire n_1964;
wire n_4133;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_4145;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_4271;
wire n_1946;
wire n_1355;
wire n_4181;
wire n_1225;
wire n_3184;
wire n_2258;
wire n_1485;
wire n_1544;
wire n_1640;
wire n_4040;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_4111;
wire n_2390;
wire n_4007;
wire n_3712;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_4239;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_4184;
wire n_2626;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_4037;
wire n_1319;
wire n_2986;
wire n_1900;
wire n_3930;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_3915;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_4343;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_4215;
wire n_1282;
wire n_2561;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2962;
wire n_2154;
wire n_2727;
wire n_3377;
wire n_2939;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_2533;
wire n_3157;
wire n_1672;
wire n_3530;
wire n_4185;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_4378;
wire n_4407;
wire n_1914;
wire n_1318;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_3893;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_3762;
wire n_3469;
wire n_3958;
wire n_2266;
wire n_2960;
wire n_3932;
wire n_3005;
wire n_3985;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_4196;
wire n_3779;
wire n_1447;
wire n_2388;
wire n_3984;
wire n_2056;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_4358;
wire n_1706;
wire n_4242;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_4232;
wire n_4190;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_2189;
wire n_2680;
wire n_4052;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_3899;
wire n_4084;
wire n_3558;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_4326;
wire n_3156;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_2668;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_3939;
wire n_1941;
wire n_1375;
wire n_3483;
wire n_3613;
wire n_3972;
wire n_4153;
wire n_2128;
wire n_1045;
wire n_1794;
wire n_1962;
wire n_1236;
wire n_1650;
wire n_1559;
wire n_2398;
wire n_1928;
wire n_1725;
wire n_3743;
wire n_3855;
wire n_1872;
wire n_3091;
wire n_4317;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_4269;
wire n_3124;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_4088;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_3524;
wire n_2671;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2888;
wire n_1804;
wire n_2923;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_1727;
wire n_2508;
wire n_4301;
wire n_3511;
wire n_2054;
wire n_4143;
wire n_4170;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_4421;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_1154;
wire n_3308;
wire n_1113;
wire n_2833;
wire n_1600;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_2261;
wire n_4423;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_1476;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_4376;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_3515;
wire n_1150;
wire n_4203;
wire n_3808;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_4365;
wire n_1826;
wire n_1882;
wire n_2951;
wire n_1118;
wire n_1076;
wire n_2949;
wire n_3726;
wire n_1807;
wire n_1929;
wire n_2369;
wire n_1378;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_3758;
wire n_1879;
wire n_3806;
wire n_4081;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_3866;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_1953;
wire n_3343;
wire n_3303;
wire n_4157;
wire n_2752;
wire n_4173;
wire n_3135;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_4229;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_3990;
wire n_3865;
wire n_1824;
wire n_3954;
wire n_1628;
wire n_4073;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_3658;
wire n_1516;
wire n_1536;
wire n_3846;
wire n_2163;
wire n_2186;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3951;
wire n_3034;
wire n_4408;
wire n_1132;
wire n_1074;
wire n_1394;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_3874;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_2969;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_3027;
wire n_1554;
wire n_3231;
wire n_4083;
wire n_1130;
wire n_3083;
wire n_4212;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_2380;
wire n_4295;
wire n_1120;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_4225;
wire n_4171;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_3541;
wire n_2565;
wire n_4023;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_1461;
wire n_3432;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_3860;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_4282;
wire n_1598;
wire n_3493;
wire n_4344;
wire n_2935;
wire n_4046;
wire n_3807;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_2385;
wire n_1283;
wire n_4112;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_3268;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3701;
wire n_3154;
wire n_4027;
wire n_2396;
wire n_2584;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_1994;
wire n_3473;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_3739;
wire n_2284;
wire n_3898;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_4352;
wire n_4391;
wire n_4416;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_1303;
wire n_2769;
wire n_4342;
wire n_3622;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_4095;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3897;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1347;
wire n_4106;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_4373;
wire n_1245;
wire n_3215;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_2952;
wire n_3068;
wire n_3853;
wire n_2117;
wire n_2234;
wire n_4256;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_3553;
wire n_1561;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_3811;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_2112;
wire n_2255;
wire n_1737;
wire n_2430;
wire n_3584;
wire n_3486;
wire n_1414;
wire n_1464;
wire n_4086;
wire n_2649;
wire n_2721;
wire n_4335;
wire n_3556;
wire n_2034;
wire n_3836;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_4068;
wire n_2032;
wire n_4409;
wire n_2744;
wire n_4309;
wire n_4363;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_2437;
wire n_2743;
wire n_3962;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_4166;
wire n_1821;
wire n_1500;
wire n_1537;
wire n_2205;
wire n_3699;
wire n_4243;
wire n_3204;
wire n_1104;
wire n_1058;
wire n_3378;
wire n_4025;
wire n_2312;
wire n_3404;
wire n_1122;
wire n_1253;
wire n_1266;
wire n_2242;
wire n_3362;
wire n_3745;
wire n_4059;
wire n_1509;
wire n_4188;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_4121;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_3256;
wire n_1276;
wire n_3802;
wire n_3868;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_4142;
wire n_2111;
wire n_2466;
wire n_3982;
wire n_4266;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_3796;
wire n_2999;
wire n_4115;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3643;
wire n_3697;
wire n_1584;
wire n_2425;
wire n_3461;
wire n_3408;
wire n_1582;
wire n_3680;
wire n_4265;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_2408;
wire n_4246;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_4383;
wire n_3098;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_2666;
wire n_4105;
wire n_1851;
wire n_1585;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_4244;
wire n_1816;
wire n_4064;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_4049;
wire n_1156;
wire n_1362;
wire n_4259;
wire n_3123;
wire n_2600;
wire n_3380;
wire n_1829;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_3038;
wire n_3086;
wire n_2033;
wire n_4104;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_3285;
wire n_4208;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_3361;
wire n_3596;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_4089;
wire n_4346;
wire n_4351;
wire n_1144;
wire n_2071;
wire n_3669;
wire n_3863;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_4316;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_3521;
wire n_3233;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_1301;
wire n_2805;
wire n_3310;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_4390;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_4061;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_4075;
wire n_3344;
wire n_2334;
wire n_3902;
wire n_4062;
wire n_3881;
wire n_3295;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_4396;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_3989;
wire n_2303;
wire n_2478;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_4233;
wire n_1606;
wire n_4332;
wire n_4108;
wire n_1133;
wire n_3374;
wire n_1194;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_2640;
wire n_3695;
wire n_4051;
wire n_1051;
wire n_3976;
wire n_4254;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_3992;
wire n_2367;
wire n_4307;
wire n_3876;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_2043;
wire n_4303;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_4293;
wire n_3552;
wire n_3206;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_2662;
wire n_3147;
wire n_3116;
wire n_3383;
wire n_3709;
wire n_3925;
wire n_4091;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_4186;
wire n_3187;
wire n_2540;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_2217;
wire n_2197;
wire n_1675;
wire n_2065;
wire n_2879;
wire n_3717;
wire n_4148;
wire n_2461;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_4341;
wire n_1884;
wire n_2040;
wire n_4057;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_1629;
wire n_1170;
wire n_2221;
wire n_4263;
wire n_1819;
wire n_2055;
wire n_1260;
wire n_3555;
wire n_3444;
wire n_4210;
wire n_2553;
wire n_1040;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_1578;
wire n_1861;
wire n_3110;
wire n_1890;
wire n_1632;
wire n_3017;
wire n_3955;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_2280;
wire n_1557;
wire n_1833;
wire n_3903;
wire n_1311;
wire n_3945;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_4205;
wire n_2162;
wire n_3908;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_4278;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3950;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_1417;
wire n_2185;
wire n_2086;
wire n_1242;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_3833;
wire n_4281;
wire n_3815;
wire n_2774;
wire n_3896;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3333;
wire n_3274;
wire n_3186;
wire n_1322;
wire n_4129;
wire n_1899;
wire n_1428;
wire n_4093;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_3965;
wire n_2632;
wire n_2579;
wire n_2105;
wire n_3079;
wire n_4360;
wire n_2098;
wire n_3085;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_4039;
wire n_3387;
wire n_2027;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_4197;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_4275;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_4283;
wire n_3504;
wire n_4194;
wire n_1449;
wire n_2912;
wire n_4272;
wire n_2659;
wire n_2930;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_1742;
wire n_4030;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g1037 ( 
.A(n_892),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_60),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_165),
.Y(n_1039)
);

INVx2_ASAP7_75t_SL g1040 ( 
.A(n_972),
.Y(n_1040)
);

CKINVDCx20_ASAP7_75t_R g1041 ( 
.A(n_742),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_197),
.Y(n_1042)
);

INVx1_ASAP7_75t_SL g1043 ( 
.A(n_940),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_529),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_858),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_898),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_869),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_991),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_698),
.Y(n_1049)
);

INVx1_ASAP7_75t_SL g1050 ( 
.A(n_159),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_392),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_284),
.Y(n_1052)
);

BUFx10_ASAP7_75t_L g1053 ( 
.A(n_101),
.Y(n_1053)
);

CKINVDCx20_ASAP7_75t_R g1054 ( 
.A(n_12),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_174),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_276),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_201),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_222),
.Y(n_1058)
);

INVx1_ASAP7_75t_SL g1059 ( 
.A(n_330),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_533),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_917),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_491),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_306),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_443),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_930),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_706),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_994),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_796),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_761),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_784),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_21),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_427),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_302),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_419),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_984),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_356),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_455),
.Y(n_1077)
);

CKINVDCx20_ASAP7_75t_R g1078 ( 
.A(n_967),
.Y(n_1078)
);

INVx1_ASAP7_75t_SL g1079 ( 
.A(n_755),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_866),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_865),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_730),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_647),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_30),
.Y(n_1084)
);

INVx3_ASAP7_75t_L g1085 ( 
.A(n_726),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_414),
.Y(n_1086)
);

CKINVDCx20_ASAP7_75t_R g1087 ( 
.A(n_655),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_17),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_459),
.Y(n_1089)
);

BUFx2_ASAP7_75t_L g1090 ( 
.A(n_175),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_964),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_18),
.Y(n_1092)
);

INVx1_ASAP7_75t_SL g1093 ( 
.A(n_551),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_725),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_331),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_314),
.Y(n_1096)
);

BUFx10_ASAP7_75t_L g1097 ( 
.A(n_296),
.Y(n_1097)
);

CKINVDCx20_ASAP7_75t_R g1098 ( 
.A(n_931),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_795),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_845),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_67),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_320),
.Y(n_1102)
);

BUFx10_ASAP7_75t_L g1103 ( 
.A(n_210),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_815),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_623),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_820),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_478),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_650),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_906),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_423),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_193),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_968),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_819),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_752),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_1033),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_927),
.Y(n_1116)
);

CKINVDCx14_ASAP7_75t_R g1117 ( 
.A(n_1011),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_981),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_999),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_579),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_439),
.Y(n_1121)
);

INVx1_ASAP7_75t_SL g1122 ( 
.A(n_850),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_585),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_1025),
.Y(n_1124)
);

INVx2_ASAP7_75t_SL g1125 ( 
.A(n_949),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_1022),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_141),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_480),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_141),
.Y(n_1129)
);

INVx1_ASAP7_75t_SL g1130 ( 
.A(n_881),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_932),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_700),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_184),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_688),
.Y(n_1134)
);

CKINVDCx20_ASAP7_75t_R g1135 ( 
.A(n_589),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_804),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_913),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_960),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_894),
.Y(n_1139)
);

CKINVDCx14_ASAP7_75t_R g1140 ( 
.A(n_339),
.Y(n_1140)
);

BUFx2_ASAP7_75t_SL g1141 ( 
.A(n_885),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_123),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_780),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_587),
.Y(n_1144)
);

CKINVDCx20_ASAP7_75t_R g1145 ( 
.A(n_268),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_674),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_52),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_938),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_823),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_91),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_737),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_829),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_765),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_966),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_502),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1023),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_369),
.Y(n_1157)
);

HB1xp67_ASAP7_75t_L g1158 ( 
.A(n_711),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_356),
.Y(n_1159)
);

INVx1_ASAP7_75t_SL g1160 ( 
.A(n_674),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_772),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_722),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_122),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_390),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_826),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_963),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_139),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_946),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_369),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_799),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_409),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_747),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_173),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_489),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_859),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_808),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_630),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_886),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_32),
.Y(n_1179)
);

CKINVDCx20_ASAP7_75t_R g1180 ( 
.A(n_36),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_740),
.Y(n_1181)
);

BUFx10_ASAP7_75t_L g1182 ( 
.A(n_658),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_503),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_21),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_668),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_308),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_777),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_471),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_952),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_401),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_187),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_699),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_136),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_209),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_350),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_187),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_934),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_178),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_297),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_800),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_910),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_614),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_458),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_196),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_776),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_988),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_53),
.Y(n_1207)
);

CKINVDCx20_ASAP7_75t_R g1208 ( 
.A(n_773),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_118),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_5),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_27),
.Y(n_1211)
);

INVx1_ASAP7_75t_SL g1212 ( 
.A(n_849),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_813),
.Y(n_1213)
);

CKINVDCx20_ASAP7_75t_R g1214 ( 
.A(n_610),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_921),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_848),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_720),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1016),
.Y(n_1218)
);

BUFx10_ASAP7_75t_L g1219 ( 
.A(n_929),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_7),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_836),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_679),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_900),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_22),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_173),
.Y(n_1225)
);

CKINVDCx12_ASAP7_75t_R g1226 ( 
.A(n_926),
.Y(n_1226)
);

CKINVDCx20_ASAP7_75t_R g1227 ( 
.A(n_571),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_52),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_944),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_264),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_883),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_947),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_980),
.Y(n_1233)
);

CKINVDCx20_ASAP7_75t_R g1234 ( 
.A(n_99),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_928),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_833),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1010),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_893),
.Y(n_1238)
);

INVx1_ASAP7_75t_SL g1239 ( 
.A(n_109),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_879),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_781),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_718),
.Y(n_1242)
);

CKINVDCx20_ASAP7_75t_R g1243 ( 
.A(n_266),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_557),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_342),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_523),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_576),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_549),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_680),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_362),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_1002),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_979),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_641),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_622),
.Y(n_1254)
);

INVx1_ASAP7_75t_SL g1255 ( 
.A(n_717),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_759),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_449),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_705),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_709),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_393),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_616),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_852),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_997),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_227),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_959),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_908),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_986),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_61),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1032),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_877),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_798),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1034),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_439),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_647),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_479),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_933),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_746),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_692),
.Y(n_1278)
);

CKINVDCx20_ASAP7_75t_R g1279 ( 
.A(n_889),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_783),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_196),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_982),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_648),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_1012),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_92),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_531),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_899),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_646),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_871),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_789),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_346),
.Y(n_1291)
);

INVx1_ASAP7_75t_SL g1292 ( 
.A(n_767),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_987),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_140),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_658),
.Y(n_1295)
);

CKINVDCx20_ASAP7_75t_R g1296 ( 
.A(n_962),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_495),
.Y(n_1297)
);

CKINVDCx16_ASAP7_75t_R g1298 ( 
.A(n_916),
.Y(n_1298)
);

BUFx8_ASAP7_75t_SL g1299 ( 
.A(n_924),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_436),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_155),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_810),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_666),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1005),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_817),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_809),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_702),
.Y(n_1307)
);

INVxp67_ASAP7_75t_L g1308 ( 
.A(n_880),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_1035),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_969),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_471),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_766),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_925),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_331),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_801),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_802),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_384),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_343),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_224),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_41),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_61),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_697),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_236),
.Y(n_1323)
);

BUFx10_ASAP7_75t_L g1324 ( 
.A(n_920),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1026),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_340),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_935),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_551),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_945),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_457),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_263),
.Y(n_1331)
);

BUFx6f_ASAP7_75t_L g1332 ( 
.A(n_722),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_863),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_970),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_282),
.Y(n_1335)
);

INVx1_ASAP7_75t_SL g1336 ( 
.A(n_714),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_78),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_328),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_210),
.Y(n_1339)
);

INVxp67_ASAP7_75t_L g1340 ( 
.A(n_479),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_123),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_1015),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_703),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_974),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_983),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_195),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_793),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_679),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1024),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_953),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_758),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_965),
.Y(n_1352)
);

BUFx5_ASAP7_75t_L g1353 ( 
.A(n_992),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_498),
.Y(n_1354)
);

CKINVDCx20_ASAP7_75t_R g1355 ( 
.A(n_846),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_217),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1013),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_26),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1014),
.Y(n_1359)
);

BUFx10_ASAP7_75t_L g1360 ( 
.A(n_234),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_680),
.Y(n_1361)
);

BUFx10_ASAP7_75t_L g1362 ( 
.A(n_601),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_1031),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_458),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_710),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_380),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_6),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_493),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_603),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_782),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_320),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_923),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_903),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_326),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_751),
.Y(n_1375)
);

INVx2_ASAP7_75t_SL g1376 ( 
.A(n_843),
.Y(n_1376)
);

CKINVDCx20_ASAP7_75t_R g1377 ( 
.A(n_1036),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_134),
.Y(n_1378)
);

CKINVDCx20_ASAP7_75t_R g1379 ( 
.A(n_453),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_870),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_595),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_943),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_257),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_895),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_830),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_657),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_283),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_668),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_995),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_712),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_710),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_428),
.Y(n_1392)
);

INVx1_ASAP7_75t_SL g1393 ( 
.A(n_650),
.Y(n_1393)
);

BUFx6f_ASAP7_75t_L g1394 ( 
.A(n_32),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_209),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_922),
.Y(n_1396)
);

INVx2_ASAP7_75t_SL g1397 ( 
.A(n_601),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_724),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_545),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_851),
.Y(n_1400)
);

INVx2_ASAP7_75t_SL g1401 ( 
.A(n_585),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_217),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_790),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_838),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_586),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_860),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_681),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_753),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_329),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_857),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_769),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_821),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_904),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_15),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_446),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_856),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1007),
.Y(n_1417)
);

BUFx10_ASAP7_75t_L g1418 ( 
.A(n_902),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_168),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_978),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_156),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_53),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_58),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_147),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_58),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_422),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_779),
.Y(n_1427)
);

BUFx10_ASAP7_75t_L g1428 ( 
.A(n_827),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_842),
.Y(n_1429)
);

CKINVDCx20_ASAP7_75t_R g1430 ( 
.A(n_1027),
.Y(n_1430)
);

BUFx10_ASAP7_75t_L g1431 ( 
.A(n_692),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_623),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1028),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_803),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_715),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_174),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_642),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_310),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_258),
.Y(n_1439)
);

INVx2_ASAP7_75t_SL g1440 ( 
.A(n_744),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_977),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_444),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_59),
.Y(n_1443)
);

CKINVDCx14_ASAP7_75t_R g1444 ( 
.A(n_825),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_432),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_25),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_794),
.Y(n_1447)
);

CKINVDCx16_ASAP7_75t_R g1448 ( 
.A(n_343),
.Y(n_1448)
);

BUFx10_ASAP7_75t_L g1449 ( 
.A(n_241),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_948),
.Y(n_1450)
);

CKINVDCx20_ASAP7_75t_R g1451 ( 
.A(n_407),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_516),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_93),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_164),
.Y(n_1454)
);

CKINVDCx20_ASAP7_75t_R g1455 ( 
.A(n_901),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_610),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_750),
.Y(n_1457)
);

CKINVDCx20_ASAP7_75t_R g1458 ( 
.A(n_589),
.Y(n_1458)
);

INVx2_ASAP7_75t_SL g1459 ( 
.A(n_1018),
.Y(n_1459)
);

CKINVDCx20_ASAP7_75t_R g1460 ( 
.A(n_690),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_313),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_1001),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_403),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_775),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_669),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_835),
.Y(n_1466)
);

CKINVDCx16_ASAP7_75t_R g1467 ( 
.A(n_985),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_536),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_354),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_424),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_664),
.Y(n_1471)
);

CKINVDCx20_ASAP7_75t_R g1472 ( 
.A(n_937),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_L g1473 ( 
.A(n_644),
.Y(n_1473)
);

CKINVDCx16_ASAP7_75t_R g1474 ( 
.A(n_257),
.Y(n_1474)
);

CKINVDCx20_ASAP7_75t_R g1475 ( 
.A(n_812),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_503),
.Y(n_1476)
);

CKINVDCx20_ASAP7_75t_R g1477 ( 
.A(n_873),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_874),
.Y(n_1478)
);

INVx1_ASAP7_75t_SL g1479 ( 
.A(n_118),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_887),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_685),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_545),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_108),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_936),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_748),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_749),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_592),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_723),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_764),
.Y(n_1489)
);

BUFx6f_ASAP7_75t_L g1490 ( 
.A(n_876),
.Y(n_1490)
);

BUFx10_ASAP7_75t_L g1491 ( 
.A(n_480),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_695),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_284),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_335),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_512),
.Y(n_1495)
);

BUFx8_ASAP7_75t_SL g1496 ( 
.A(n_40),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_708),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_572),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_380),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_560),
.Y(n_1500)
);

CKINVDCx14_ASAP7_75t_R g1501 ( 
.A(n_98),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_556),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_791),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_834),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_165),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_412),
.Y(n_1506)
);

BUFx10_ASAP7_75t_L g1507 ( 
.A(n_368),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_961),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_646),
.Y(n_1509)
);

CKINVDCx20_ASAP7_75t_R g1510 ( 
.A(n_847),
.Y(n_1510)
);

CKINVDCx14_ASAP7_75t_R g1511 ( 
.A(n_941),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_425),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_333),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_743),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_152),
.Y(n_1515)
);

CKINVDCx20_ASAP7_75t_R g1516 ( 
.A(n_300),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_608),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_884),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_875),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_79),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_768),
.Y(n_1521)
);

CKINVDCx20_ASAP7_75t_R g1522 ( 
.A(n_681),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_614),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_36),
.Y(n_1524)
);

INVxp67_ASAP7_75t_L g1525 ( 
.A(n_142),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_214),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_919),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_546),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_324),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_993),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_530),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_590),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_716),
.Y(n_1533)
);

CKINVDCx20_ASAP7_75t_R g1534 ( 
.A(n_114),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_48),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_514),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_348),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_48),
.Y(n_1538)
);

CKINVDCx20_ASAP7_75t_R g1539 ( 
.A(n_872),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_939),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_717),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_667),
.Y(n_1542)
);

INVx1_ASAP7_75t_SL g1543 ( 
.A(n_299),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_957),
.Y(n_1544)
);

INVx2_ASAP7_75t_SL g1545 ( 
.A(n_861),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_146),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_818),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_955),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_283),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_583),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_219),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_837),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_147),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_342),
.Y(n_1554)
);

BUFx3_ASAP7_75t_L g1555 ( 
.A(n_294),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_721),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_349),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_497),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_841),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_543),
.Y(n_1560)
);

CKINVDCx20_ASAP7_75t_R g1561 ( 
.A(n_472),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_184),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_446),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_270),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_745),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_1030),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_676),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_516),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_603),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_291),
.Y(n_1570)
);

INVx1_ASAP7_75t_SL g1571 ( 
.A(n_1006),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_119),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_244),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_417),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_16),
.Y(n_1575)
);

INVx1_ASAP7_75t_SL g1576 ( 
.A(n_867),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_942),
.Y(n_1577)
);

BUFx2_ASAP7_75t_L g1578 ( 
.A(n_741),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_205),
.Y(n_1579)
);

BUFx2_ASAP7_75t_L g1580 ( 
.A(n_760),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_44),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_990),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_122),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_1004),
.Y(n_1584)
);

INVx2_ASAP7_75t_SL g1585 ( 
.A(n_882),
.Y(n_1585)
);

CKINVDCx20_ASAP7_75t_R g1586 ( 
.A(n_391),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_41),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_762),
.Y(n_1588)
);

CKINVDCx20_ASAP7_75t_R g1589 ( 
.A(n_179),
.Y(n_1589)
);

INVx1_ASAP7_75t_SL g1590 ( 
.A(n_148),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_421),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_206),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_735),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_950),
.Y(n_1594)
);

BUFx3_ASAP7_75t_L g1595 ( 
.A(n_327),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_909),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_392),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_914),
.Y(n_1598)
);

BUFx3_ASAP7_75t_L g1599 ( 
.A(n_33),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_18),
.Y(n_1600)
);

INVx1_ASAP7_75t_SL g1601 ( 
.A(n_756),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_971),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_150),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_792),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_71),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_738),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_629),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_99),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_424),
.Y(n_1609)
);

BUFx5_ASAP7_75t_L g1610 ( 
.A(n_918),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_563),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_811),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_426),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_754),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_785),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_797),
.Y(n_1616)
);

CKINVDCx20_ASAP7_75t_R g1617 ( 
.A(n_976),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1009),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_5),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_989),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_313),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_890),
.Y(n_1622)
);

BUFx2_ASAP7_75t_SL g1623 ( 
.A(n_251),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_260),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_432),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_831),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_361),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_238),
.Y(n_1628)
);

INVxp33_ASAP7_75t_R g1629 ( 
.A(n_523),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_221),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_171),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_816),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_495),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_146),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_517),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_390),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_853),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_854),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_687),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_907),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_348),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_139),
.Y(n_1642)
);

CKINVDCx20_ASAP7_75t_R g1643 ( 
.A(n_778),
.Y(n_1643)
);

BUFx5_ASAP7_75t_L g1644 ( 
.A(n_805),
.Y(n_1644)
);

CKINVDCx20_ASAP7_75t_R g1645 ( 
.A(n_617),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_518),
.Y(n_1646)
);

INVx1_ASAP7_75t_SL g1647 ( 
.A(n_911),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_71),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_896),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_31),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_120),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_558),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_786),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_822),
.Y(n_1654)
);

BUFx10_ASAP7_75t_L g1655 ( 
.A(n_1000),
.Y(n_1655)
);

HB1xp67_ASAP7_75t_L g1656 ( 
.A(n_153),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_286),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_855),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1003),
.Y(n_1659)
);

BUFx6f_ASAP7_75t_L g1660 ( 
.A(n_956),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_248),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_729),
.Y(n_1662)
);

BUFx2_ASAP7_75t_L g1663 ( 
.A(n_840),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_388),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_620),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1020),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_905),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_1019),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_788),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_1029),
.Y(n_1670)
);

INVx2_ASAP7_75t_SL g1671 ( 
.A(n_74),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_727),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_371),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_878),
.Y(n_1674)
);

BUFx10_ASAP7_75t_L g1675 ( 
.A(n_599),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_832),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_862),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_951),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_450),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_669),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_537),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_245),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_975),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_412),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_719),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_548),
.Y(n_1686)
);

BUFx10_ASAP7_75t_L g1687 ( 
.A(n_958),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_739),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_771),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_470),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_SL g1691 ( 
.A(n_689),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_399),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_666),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_191),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_844),
.Y(n_1695)
);

CKINVDCx16_ASAP7_75t_R g1696 ( 
.A(n_888),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_227),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_868),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_394),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_592),
.Y(n_1700)
);

CKINVDCx20_ASAP7_75t_R g1701 ( 
.A(n_864),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_150),
.Y(n_1702)
);

CKINVDCx5p33_ASAP7_75t_R g1703 ( 
.A(n_728),
.Y(n_1703)
);

HB1xp67_ASAP7_75t_L g1704 ( 
.A(n_216),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_602),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_62),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_529),
.Y(n_1707)
);

BUFx3_ASAP7_75t_L g1708 ( 
.A(n_175),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_996),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_891),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_277),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_774),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_652),
.Y(n_1713)
);

BUFx2_ASAP7_75t_L g1714 ( 
.A(n_482),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_807),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_497),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_839),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_713),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_180),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_560),
.Y(n_1720)
);

BUFx5_ASAP7_75t_L g1721 ( 
.A(n_488),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_721),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_696),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_574),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_824),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_954),
.Y(n_1726)
);

INVxp67_ASAP7_75t_SL g1727 ( 
.A(n_763),
.Y(n_1727)
);

INVxp67_ASAP7_75t_L g1728 ( 
.A(n_501),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_734),
.Y(n_1729)
);

CKINVDCx20_ASAP7_75t_R g1730 ( 
.A(n_704),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_205),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_806),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_531),
.Y(n_1733)
);

BUFx10_ASAP7_75t_L g1734 ( 
.A(n_158),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_998),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_544),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_579),
.Y(n_1737)
);

CKINVDCx5p33_ASAP7_75t_R g1738 ( 
.A(n_452),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_180),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_188),
.Y(n_1740)
);

CKINVDCx20_ASAP7_75t_R g1741 ( 
.A(n_499),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_124),
.Y(n_1742)
);

BUFx3_ASAP7_75t_L g1743 ( 
.A(n_244),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_973),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_164),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_575),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_79),
.Y(n_1747)
);

INVx1_ASAP7_75t_SL g1748 ( 
.A(n_915),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_828),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_814),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_770),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_70),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_912),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_787),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_151),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_1017),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_1008),
.Y(n_1757)
);

BUFx3_ASAP7_75t_L g1758 ( 
.A(n_667),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_566),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_485),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_701),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_463),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_584),
.Y(n_1763)
);

BUFx10_ASAP7_75t_L g1764 ( 
.A(n_452),
.Y(n_1764)
);

BUFx3_ASAP7_75t_L g1765 ( 
.A(n_607),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_522),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_177),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1021),
.Y(n_1768)
);

BUFx2_ASAP7_75t_SL g1769 ( 
.A(n_707),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_563),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_441),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_299),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_757),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_403),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_897),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_700),
.Y(n_1776)
);

INVxp67_ASAP7_75t_SL g1777 ( 
.A(n_1048),
.Y(n_1777)
);

INVxp67_ASAP7_75t_L g1778 ( 
.A(n_1090),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1721),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1721),
.Y(n_1780)
);

BUFx3_ASAP7_75t_L g1781 ( 
.A(n_1219),
.Y(n_1781)
);

INVxp67_ASAP7_75t_L g1782 ( 
.A(n_1285),
.Y(n_1782)
);

INVxp67_ASAP7_75t_SL g1783 ( 
.A(n_1115),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1721),
.Y(n_1784)
);

INVxp67_ASAP7_75t_SL g1785 ( 
.A(n_1578),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1721),
.Y(n_1786)
);

INVxp67_ASAP7_75t_SL g1787 ( 
.A(n_1580),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1721),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1085),
.Y(n_1789)
);

CKINVDCx16_ASAP7_75t_R g1790 ( 
.A(n_1448),
.Y(n_1790)
);

CKINVDCx16_ASAP7_75t_R g1791 ( 
.A(n_1474),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1085),
.Y(n_1792)
);

BUFx3_ASAP7_75t_L g1793 ( 
.A(n_1219),
.Y(n_1793)
);

INVxp33_ASAP7_75t_SL g1794 ( 
.A(n_1147),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1042),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1042),
.Y(n_1796)
);

INVxp67_ASAP7_75t_L g1797 ( 
.A(n_1303),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1042),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1196),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1196),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1196),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1225),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1225),
.Y(n_1803)
);

CKINVDCx5p33_ASAP7_75t_R g1804 ( 
.A(n_1299),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1225),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1332),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1332),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1332),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1337),
.Y(n_1809)
);

INVxp67_ASAP7_75t_SL g1810 ( 
.A(n_1663),
.Y(n_1810)
);

INVxp67_ASAP7_75t_SL g1811 ( 
.A(n_1154),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1337),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1337),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1394),
.Y(n_1814)
);

CKINVDCx5p33_ASAP7_75t_R g1815 ( 
.A(n_1496),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1394),
.Y(n_1816)
);

CKINVDCx20_ASAP7_75t_R g1817 ( 
.A(n_1041),
.Y(n_1817)
);

INVxp67_ASAP7_75t_L g1818 ( 
.A(n_1714),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1394),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1426),
.Y(n_1820)
);

INVx3_ASAP7_75t_L g1821 ( 
.A(n_1426),
.Y(n_1821)
);

CKINVDCx20_ASAP7_75t_R g1822 ( 
.A(n_1078),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1426),
.Y(n_1823)
);

INVxp67_ASAP7_75t_SL g1824 ( 
.A(n_1154),
.Y(n_1824)
);

INVxp67_ASAP7_75t_SL g1825 ( 
.A(n_1161),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1463),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_L g1827 ( 
.A(n_1140),
.B(n_1),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_1045),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1047),
.Y(n_1829)
);

INVxp33_ASAP7_75t_L g1830 ( 
.A(n_1158),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1463),
.Y(n_1831)
);

CKINVDCx5p33_ASAP7_75t_R g1832 ( 
.A(n_1061),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1463),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1473),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1473),
.Y(n_1835)
);

INVxp67_ASAP7_75t_L g1836 ( 
.A(n_1656),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1473),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_1065),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1071),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_1070),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1074),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1253),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1300),
.Y(n_1843)
);

CKINVDCx16_ASAP7_75t_R g1844 ( 
.A(n_1298),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_1081),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1321),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_1082),
.Y(n_1847)
);

INVxp67_ASAP7_75t_SL g1848 ( 
.A(n_1406),
.Y(n_1848)
);

INVxp67_ASAP7_75t_L g1849 ( 
.A(n_1704),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1443),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1353),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1555),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1556),
.Y(n_1853)
);

INVxp67_ASAP7_75t_L g1854 ( 
.A(n_1691),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1595),
.Y(n_1855)
);

CKINVDCx5p33_ASAP7_75t_R g1856 ( 
.A(n_1091),
.Y(n_1856)
);

INVxp67_ASAP7_75t_SL g1857 ( 
.A(n_1447),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_1106),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1353),
.Y(n_1859)
);

CKINVDCx16_ASAP7_75t_R g1860 ( 
.A(n_1467),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1599),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1708),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1743),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1758),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_1114),
.Y(n_1865)
);

INVxp67_ASAP7_75t_SL g1866 ( 
.A(n_1308),
.Y(n_1866)
);

INVxp67_ASAP7_75t_SL g1867 ( 
.A(n_1765),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1044),
.Y(n_1868)
);

INVxp67_ASAP7_75t_SL g1869 ( 
.A(n_1046),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1051),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1055),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1062),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1761),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1771),
.Y(n_1874)
);

INVxp67_ASAP7_75t_SL g1875 ( 
.A(n_1067),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1772),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1073),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_1116),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1086),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1094),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_1118),
.Y(n_1881)
);

INVxp67_ASAP7_75t_SL g1882 ( 
.A(n_1068),
.Y(n_1882)
);

INVxp67_ASAP7_75t_L g1883 ( 
.A(n_1053),
.Y(n_1883)
);

INVxp67_ASAP7_75t_SL g1884 ( 
.A(n_1069),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1107),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1111),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1132),
.Y(n_1887)
);

INVxp33_ASAP7_75t_SL g1888 ( 
.A(n_1038),
.Y(n_1888)
);

INVxp67_ASAP7_75t_SL g1889 ( 
.A(n_1075),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1759),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1150),
.Y(n_1891)
);

BUFx3_ASAP7_75t_L g1892 ( 
.A(n_1839),
.Y(n_1892)
);

HB1xp67_ASAP7_75t_L g1893 ( 
.A(n_1854),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1816),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1835),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1825),
.B(n_1117),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1795),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1796),
.Y(n_1898)
);

BUFx2_ASAP7_75t_L g1899 ( 
.A(n_1781),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1798),
.Y(n_1900)
);

BUFx6f_ASAP7_75t_L g1901 ( 
.A(n_1821),
.Y(n_1901)
);

BUFx6f_ASAP7_75t_L g1902 ( 
.A(n_1821),
.Y(n_1902)
);

BUFx6f_ASAP7_75t_L g1903 ( 
.A(n_1799),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1828),
.B(n_1444),
.Y(n_1904)
);

OA22x2_ASAP7_75t_SL g1905 ( 
.A1(n_1785),
.A2(n_1629),
.B1(n_1186),
.B2(n_1190),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1800),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1801),
.Y(n_1907)
);

OA21x2_ASAP7_75t_L g1908 ( 
.A1(n_1779),
.A2(n_1099),
.B(n_1080),
.Y(n_1908)
);

OAI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1794),
.A2(n_1810),
.B1(n_1787),
.B2(n_1778),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1802),
.Y(n_1910)
);

OA21x2_ASAP7_75t_L g1911 ( 
.A1(n_1780),
.A2(n_1109),
.B(n_1100),
.Y(n_1911)
);

INVx3_ASAP7_75t_L g1912 ( 
.A(n_1803),
.Y(n_1912)
);

BUFx6f_ASAP7_75t_L g1913 ( 
.A(n_1805),
.Y(n_1913)
);

NOR2xp33_ASAP7_75t_L g1914 ( 
.A(n_1888),
.B(n_1501),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1806),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1807),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1808),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1848),
.B(n_1511),
.Y(n_1918)
);

CKINVDCx5p33_ASAP7_75t_R g1919 ( 
.A(n_1829),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1809),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1832),
.B(n_1040),
.Y(n_1921)
);

HB1xp67_ASAP7_75t_L g1922 ( 
.A(n_1790),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1812),
.Y(n_1923)
);

NOR2xp33_ASAP7_75t_L g1924 ( 
.A(n_1838),
.B(n_1696),
.Y(n_1924)
);

AOI22xp33_ASAP7_75t_SL g1925 ( 
.A1(n_1791),
.A2(n_1087),
.B1(n_1134),
.B2(n_1054),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1813),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1814),
.Y(n_1927)
);

INVx3_ASAP7_75t_L g1928 ( 
.A(n_1819),
.Y(n_1928)
);

BUFx6f_ASAP7_75t_L g1929 ( 
.A(n_1820),
.Y(n_1929)
);

AND2x4_ASAP7_75t_L g1930 ( 
.A(n_1793),
.B(n_1043),
.Y(n_1930)
);

CKINVDCx20_ASAP7_75t_R g1931 ( 
.A(n_1817),
.Y(n_1931)
);

AOI22xp5_ASAP7_75t_L g1932 ( 
.A1(n_1827),
.A2(n_1104),
.B1(n_1126),
.B2(n_1098),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1823),
.Y(n_1933)
);

OA21x2_ASAP7_75t_L g1934 ( 
.A1(n_1784),
.A2(n_1113),
.B(n_1112),
.Y(n_1934)
);

AND2x4_ASAP7_75t_L g1935 ( 
.A(n_1857),
.B(n_1079),
.Y(n_1935)
);

BUFx6f_ASAP7_75t_L g1936 ( 
.A(n_1826),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1831),
.Y(n_1937)
);

BUFx6f_ASAP7_75t_L g1938 ( 
.A(n_1833),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1834),
.Y(n_1939)
);

OAI22xp5_ASAP7_75t_SL g1940 ( 
.A1(n_1822),
.A2(n_1145),
.B1(n_1180),
.B2(n_1135),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1837),
.Y(n_1941)
);

INVx3_ASAP7_75t_L g1942 ( 
.A(n_1841),
.Y(n_1942)
);

BUFx3_ASAP7_75t_L g1943 ( 
.A(n_1842),
.Y(n_1943)
);

NOR2xp33_ASAP7_75t_L g1944 ( 
.A(n_1840),
.B(n_1845),
.Y(n_1944)
);

OAI22x1_ASAP7_75t_SL g1945 ( 
.A1(n_1815),
.A2(n_1222),
.B1(n_1227),
.B2(n_1214),
.Y(n_1945)
);

OAI21x1_ASAP7_75t_L g1946 ( 
.A1(n_1851),
.A2(n_1156),
.B(n_1037),
.Y(n_1946)
);

AND2x4_ASAP7_75t_L g1947 ( 
.A(n_1777),
.B(n_1122),
.Y(n_1947)
);

OAI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1782),
.A2(n_1525),
.B1(n_1728),
.B2(n_1340),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1786),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1788),
.Y(n_1950)
);

AND2x4_ASAP7_75t_L g1951 ( 
.A(n_1783),
.B(n_1130),
.Y(n_1951)
);

AOI22xp5_ASAP7_75t_L g1952 ( 
.A1(n_1844),
.A2(n_1860),
.B1(n_1818),
.B2(n_1797),
.Y(n_1952)
);

NOR2xp33_ASAP7_75t_L g1953 ( 
.A(n_1847),
.B(n_1212),
.Y(n_1953)
);

BUFx6f_ASAP7_75t_L g1954 ( 
.A(n_1868),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1866),
.B(n_1324),
.Y(n_1955)
);

BUFx6f_ASAP7_75t_L g1956 ( 
.A(n_1870),
.Y(n_1956)
);

BUFx12f_ASAP7_75t_L g1957 ( 
.A(n_1804),
.Y(n_1957)
);

INVxp67_ASAP7_75t_L g1958 ( 
.A(n_1867),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1789),
.Y(n_1959)
);

INVx3_ASAP7_75t_L g1960 ( 
.A(n_1843),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1792),
.Y(n_1961)
);

AOI22xp5_ASAP7_75t_L g1962 ( 
.A1(n_1836),
.A2(n_1266),
.B1(n_1279),
.B2(n_1208),
.Y(n_1962)
);

INVxp67_ASAP7_75t_L g1963 ( 
.A(n_1846),
.Y(n_1963)
);

AND2x4_ASAP7_75t_L g1964 ( 
.A(n_1849),
.B(n_1292),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1871),
.Y(n_1965)
);

BUFx6f_ASAP7_75t_L g1966 ( 
.A(n_1872),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1873),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1874),
.Y(n_1968)
);

BUFx6f_ASAP7_75t_L g1969 ( 
.A(n_1876),
.Y(n_1969)
);

INVx6_ASAP7_75t_L g1970 ( 
.A(n_1883),
.Y(n_1970)
);

OAI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1830),
.A2(n_1049),
.B1(n_1052),
.B2(n_1039),
.Y(n_1971)
);

BUFx6f_ASAP7_75t_L g1972 ( 
.A(n_1877),
.Y(n_1972)
);

BUFx12f_ASAP7_75t_L g1973 ( 
.A(n_1856),
.Y(n_1973)
);

BUFx3_ASAP7_75t_L g1974 ( 
.A(n_1850),
.Y(n_1974)
);

BUFx6f_ASAP7_75t_L g1975 ( 
.A(n_1879),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1880),
.Y(n_1976)
);

INVx3_ASAP7_75t_L g1977 ( 
.A(n_1852),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1885),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1886),
.Y(n_1979)
);

INVx3_ASAP7_75t_L g1980 ( 
.A(n_1853),
.Y(n_1980)
);

OA21x2_ASAP7_75t_L g1981 ( 
.A1(n_1811),
.A2(n_1131),
.B(n_1119),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1858),
.B(n_1324),
.Y(n_1982)
);

AND2x4_ASAP7_75t_L g1983 ( 
.A(n_1824),
.B(n_1571),
.Y(n_1983)
);

BUFx2_ASAP7_75t_L g1984 ( 
.A(n_1865),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1878),
.B(n_1125),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1887),
.Y(n_1986)
);

BUFx2_ASAP7_75t_L g1987 ( 
.A(n_1881),
.Y(n_1987)
);

BUFx3_ASAP7_75t_L g1988 ( 
.A(n_1855),
.Y(n_1988)
);

AND2x4_ASAP7_75t_L g1989 ( 
.A(n_1869),
.B(n_1576),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1890),
.Y(n_1990)
);

AND2x4_ASAP7_75t_L g1991 ( 
.A(n_1875),
.B(n_1601),
.Y(n_1991)
);

INVx4_ASAP7_75t_L g1992 ( 
.A(n_1859),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1882),
.B(n_1418),
.Y(n_1993)
);

OA21x2_ASAP7_75t_L g1994 ( 
.A1(n_1884),
.A2(n_1165),
.B(n_1143),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1889),
.B(n_1376),
.Y(n_1995)
);

INVx5_ASAP7_75t_L g1996 ( 
.A(n_1891),
.Y(n_1996)
);

AOI22x1_ASAP7_75t_SL g1997 ( 
.A1(n_1861),
.A2(n_1243),
.B1(n_1346),
.B2(n_1234),
.Y(n_1997)
);

BUFx6f_ASAP7_75t_L g1998 ( 
.A(n_1862),
.Y(n_1998)
);

AND2x4_ASAP7_75t_L g1999 ( 
.A(n_1863),
.B(n_1647),
.Y(n_1999)
);

AOI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1864),
.A2(n_1342),
.B1(n_1355),
.B2(n_1296),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1816),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1816),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1828),
.B(n_1440),
.Y(n_2003)
);

OAI22x1_ASAP7_75t_L g2004 ( 
.A1(n_1883),
.A2(n_1059),
.B1(n_1093),
.B2(n_1050),
.Y(n_2004)
);

BUFx8_ASAP7_75t_L g2005 ( 
.A(n_1781),
.Y(n_2005)
);

BUFx6f_ASAP7_75t_L g2006 ( 
.A(n_1816),
.Y(n_2006)
);

OAI21x1_ASAP7_75t_L g2007 ( 
.A1(n_1851),
.A2(n_1256),
.B(n_1238),
.Y(n_2007)
);

BUFx12f_ASAP7_75t_L g2008 ( 
.A(n_1804),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1825),
.B(n_1418),
.Y(n_2009)
);

AND2x6_ASAP7_75t_L g2010 ( 
.A(n_1827),
.B(n_1160),
.Y(n_2010)
);

AND2x4_ASAP7_75t_L g2011 ( 
.A(n_1781),
.B(n_1748),
.Y(n_2011)
);

INVx5_ASAP7_75t_L g2012 ( 
.A(n_1821),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1816),
.Y(n_2013)
);

NOR2xp33_ASAP7_75t_SL g2014 ( 
.A(n_1844),
.B(n_1428),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1828),
.B(n_1459),
.Y(n_2015)
);

HB1xp67_ASAP7_75t_L g2016 ( 
.A(n_1854),
.Y(n_2016)
);

XNOR2xp5_ASAP7_75t_L g2017 ( 
.A(n_1817),
.B(n_1379),
.Y(n_2017)
);

INVx3_ASAP7_75t_L g2018 ( 
.A(n_1821),
.Y(n_2018)
);

CKINVDCx20_ASAP7_75t_R g2019 ( 
.A(n_1817),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1816),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1828),
.B(n_1545),
.Y(n_2021)
);

BUFx6f_ASAP7_75t_L g2022 ( 
.A(n_1816),
.Y(n_2022)
);

AND2x4_ASAP7_75t_L g2023 ( 
.A(n_1781),
.B(n_1727),
.Y(n_2023)
);

INVx1_ASAP7_75t_SL g2024 ( 
.A(n_1817),
.Y(n_2024)
);

INVx3_ASAP7_75t_L g2025 ( 
.A(n_1821),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1825),
.B(n_1428),
.Y(n_2026)
);

BUFx6f_ASAP7_75t_L g2027 ( 
.A(n_1816),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1828),
.B(n_1585),
.Y(n_2028)
);

BUFx6f_ASAP7_75t_L g2029 ( 
.A(n_1816),
.Y(n_2029)
);

AND2x4_ASAP7_75t_L g2030 ( 
.A(n_1781),
.B(n_1176),
.Y(n_2030)
);

OAI21x1_ASAP7_75t_L g2031 ( 
.A1(n_1851),
.A2(n_1357),
.B(n_1325),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1816),
.Y(n_2032)
);

OA21x2_ASAP7_75t_L g2033 ( 
.A1(n_1779),
.A2(n_1187),
.B(n_1178),
.Y(n_2033)
);

BUFx6f_ASAP7_75t_L g2034 ( 
.A(n_1816),
.Y(n_2034)
);

INVx4_ASAP7_75t_L g2035 ( 
.A(n_1828),
.Y(n_2035)
);

AOI22xp5_ASAP7_75t_L g2036 ( 
.A1(n_1794),
.A2(n_1430),
.B1(n_1455),
.B2(n_1377),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1825),
.B(n_1655),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1816),
.Y(n_2038)
);

INVx3_ASAP7_75t_L g2039 ( 
.A(n_1821),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1828),
.B(n_1370),
.Y(n_2040)
);

OAI22xp5_ASAP7_75t_L g2041 ( 
.A1(n_1794),
.A2(n_1056),
.B1(n_1058),
.B2(n_1057),
.Y(n_2041)
);

NOR2xp33_ASAP7_75t_SL g2042 ( 
.A(n_1844),
.B(n_1655),
.Y(n_2042)
);

BUFx12f_ASAP7_75t_L g2043 ( 
.A(n_1804),
.Y(n_2043)
);

INVx5_ASAP7_75t_L g2044 ( 
.A(n_1821),
.Y(n_2044)
);

AOI22x1_ASAP7_75t_SL g2045 ( 
.A1(n_1817),
.A2(n_1458),
.B1(n_1460),
.B2(n_1451),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1816),
.Y(n_2046)
);

INVx4_ASAP7_75t_L g2047 ( 
.A(n_1828),
.Y(n_2047)
);

BUFx3_ASAP7_75t_L g2048 ( 
.A(n_1839),
.Y(n_2048)
);

BUFx6f_ASAP7_75t_L g2049 ( 
.A(n_1816),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1816),
.Y(n_2050)
);

BUFx6f_ASAP7_75t_L g2051 ( 
.A(n_1816),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_1816),
.Y(n_2052)
);

BUFx6f_ASAP7_75t_L g2053 ( 
.A(n_1816),
.Y(n_2053)
);

INVx4_ASAP7_75t_L g2054 ( 
.A(n_1828),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1828),
.B(n_1413),
.Y(n_2055)
);

INVxp67_ASAP7_75t_L g2056 ( 
.A(n_1781),
.Y(n_2056)
);

OAI21x1_ASAP7_75t_L g2057 ( 
.A1(n_1851),
.A2(n_1612),
.B(n_1602),
.Y(n_2057)
);

AOI22x1_ASAP7_75t_SL g2058 ( 
.A1(n_1817),
.A2(n_1522),
.B1(n_1534),
.B2(n_1516),
.Y(n_2058)
);

OAI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_1794),
.A2(n_1060),
.B1(n_1064),
.B2(n_1063),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1828),
.B(n_1654),
.Y(n_2060)
);

AND2x4_ASAP7_75t_L g2061 ( 
.A(n_1781),
.B(n_1197),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1828),
.B(n_1666),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1816),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1816),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1816),
.Y(n_2065)
);

BUFx2_ASAP7_75t_L g2066 ( 
.A(n_1854),
.Y(n_2066)
);

BUFx6f_ASAP7_75t_L g2067 ( 
.A(n_1816),
.Y(n_2067)
);

BUFx6f_ASAP7_75t_L g2068 ( 
.A(n_1816),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1816),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1816),
.Y(n_2070)
);

BUFx8_ASAP7_75t_L g2071 ( 
.A(n_1781),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1828),
.B(n_1667),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1816),
.Y(n_2073)
);

OAI22xp5_ASAP7_75t_SL g2074 ( 
.A1(n_1794),
.A2(n_1586),
.B1(n_1589),
.B2(n_1561),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1816),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1816),
.Y(n_2076)
);

XNOR2xp5_ASAP7_75t_L g2077 ( 
.A(n_1817),
.B(n_1645),
.Y(n_2077)
);

AOI22xp5_ASAP7_75t_SL g2078 ( 
.A1(n_1794),
.A2(n_1741),
.B1(n_1730),
.B2(n_1475),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1816),
.Y(n_2079)
);

INVx3_ASAP7_75t_L g2080 ( 
.A(n_1821),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1816),
.Y(n_2081)
);

OAI22xp5_ASAP7_75t_SL g2082 ( 
.A1(n_1794),
.A2(n_1255),
.B1(n_1336),
.B2(n_1239),
.Y(n_2082)
);

BUFx6f_ASAP7_75t_L g2083 ( 
.A(n_1816),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_1816),
.Y(n_2084)
);

OA21x2_ASAP7_75t_L g2085 ( 
.A1(n_1779),
.A2(n_1201),
.B(n_1200),
.Y(n_2085)
);

INVx4_ASAP7_75t_L g2086 ( 
.A(n_1828),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_1828),
.B(n_1695),
.Y(n_2087)
);

BUFx6f_ASAP7_75t_L g2088 ( 
.A(n_1816),
.Y(n_2088)
);

OAI22x1_ASAP7_75t_L g2089 ( 
.A1(n_1883),
.A2(n_1479),
.B1(n_1543),
.B2(n_1393),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_1816),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_1828),
.B(n_1206),
.Y(n_2091)
);

AND2x4_ASAP7_75t_L g2092 ( 
.A(n_1781),
.B(n_1218),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1816),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1816),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1816),
.Y(n_2095)
);

NOR2xp33_ASAP7_75t_L g2096 ( 
.A(n_1888),
.B(n_1229),
.Y(n_2096)
);

INVx4_ASAP7_75t_L g2097 ( 
.A(n_1828),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1816),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1816),
.Y(n_2099)
);

BUFx6f_ASAP7_75t_L g2100 ( 
.A(n_1816),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_1816),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1816),
.Y(n_2102)
);

CKINVDCx5p33_ASAP7_75t_R g2103 ( 
.A(n_1828),
.Y(n_2103)
);

BUFx6f_ASAP7_75t_L g2104 ( 
.A(n_1816),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1816),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1828),
.B(n_1231),
.Y(n_2106)
);

NOR2xp33_ASAP7_75t_L g2107 ( 
.A(n_1888),
.B(n_1240),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1816),
.Y(n_2108)
);

NOR2xp33_ASAP7_75t_SL g2109 ( 
.A(n_1844),
.B(n_1687),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1816),
.Y(n_2110)
);

INVx3_ASAP7_75t_L g2111 ( 
.A(n_1821),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1816),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1816),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1816),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1816),
.Y(n_2115)
);

INVx6_ASAP7_75t_L g2116 ( 
.A(n_1781),
.Y(n_2116)
);

BUFx12f_ASAP7_75t_L g2117 ( 
.A(n_1804),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_1816),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_1825),
.B(n_1687),
.Y(n_2119)
);

AND2x4_ASAP7_75t_L g2120 ( 
.A(n_1781),
.B(n_1241),
.Y(n_2120)
);

BUFx8_ASAP7_75t_L g2121 ( 
.A(n_1781),
.Y(n_2121)
);

AOI22xp5_ASAP7_75t_L g2122 ( 
.A1(n_1794),
.A2(n_1477),
.B1(n_1510),
.B2(n_1472),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_1816),
.Y(n_2123)
);

BUFx6f_ASAP7_75t_L g2124 ( 
.A(n_1816),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1816),
.Y(n_2125)
);

BUFx2_ASAP7_75t_L g2126 ( 
.A(n_1854),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_1816),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1816),
.Y(n_2128)
);

OA21x2_ASAP7_75t_L g2129 ( 
.A1(n_1779),
.A2(n_1282),
.B(n_1269),
.Y(n_2129)
);

AND2x4_ASAP7_75t_L g2130 ( 
.A(n_1781),
.B(n_1289),
.Y(n_2130)
);

CKINVDCx6p67_ASAP7_75t_R g2131 ( 
.A(n_1790),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_1825),
.B(n_1397),
.Y(n_2132)
);

INVx2_ASAP7_75t_SL g2133 ( 
.A(n_1781),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1816),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1828),
.B(n_1293),
.Y(n_2135)
);

NOR2xp33_ASAP7_75t_L g2136 ( 
.A(n_1888),
.B(n_1305),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1816),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1816),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1816),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1816),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_1816),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1816),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1816),
.Y(n_2143)
);

BUFx6f_ASAP7_75t_L g2144 ( 
.A(n_1816),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_1816),
.Y(n_2145)
);

BUFx3_ASAP7_75t_L g2146 ( 
.A(n_1839),
.Y(n_2146)
);

CKINVDCx5p33_ASAP7_75t_R g2147 ( 
.A(n_1828),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1816),
.Y(n_2148)
);

BUFx6f_ASAP7_75t_L g2149 ( 
.A(n_1816),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1828),
.B(n_1310),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_SL g2151 ( 
.A(n_1844),
.B(n_1053),
.Y(n_2151)
);

AOI22xp5_ASAP7_75t_L g2152 ( 
.A1(n_1794),
.A2(n_1617),
.B1(n_1643),
.B2(n_1539),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1816),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1816),
.Y(n_2154)
);

INVxp67_ASAP7_75t_SL g2155 ( 
.A(n_1825),
.Y(n_2155)
);

BUFx3_ASAP7_75t_L g2156 ( 
.A(n_1839),
.Y(n_2156)
);

BUFx6f_ASAP7_75t_L g2157 ( 
.A(n_1816),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1816),
.Y(n_2158)
);

AND2x4_ASAP7_75t_L g2159 ( 
.A(n_1781),
.B(n_1312),
.Y(n_2159)
);

AOI22x1_ASAP7_75t_SL g2160 ( 
.A1(n_1817),
.A2(n_1072),
.B1(n_1076),
.B2(n_1066),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1816),
.Y(n_2161)
);

HB1xp67_ASAP7_75t_L g2162 ( 
.A(n_1854),
.Y(n_2162)
);

OAI21x1_ASAP7_75t_L g2163 ( 
.A1(n_1851),
.A2(n_1327),
.B(n_1315),
.Y(n_2163)
);

CKINVDCx5p33_ASAP7_75t_R g2164 ( 
.A(n_1919),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_2103),
.Y(n_2165)
);

HB1xp67_ASAP7_75t_L g2166 ( 
.A(n_1922),
.Y(n_2166)
);

AND3x2_ASAP7_75t_L g2167 ( 
.A(n_2014),
.B(n_1144),
.C(n_1101),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2155),
.B(n_1124),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1965),
.Y(n_2169)
);

CKINVDCx5p33_ASAP7_75t_R g2170 ( 
.A(n_2147),
.Y(n_2170)
);

CKINVDCx16_ASAP7_75t_R g2171 ( 
.A(n_1931),
.Y(n_2171)
);

INVxp33_ASAP7_75t_SL g2172 ( 
.A(n_2017),
.Y(n_2172)
);

CKINVDCx20_ASAP7_75t_R g2173 ( 
.A(n_2019),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1968),
.Y(n_2174)
);

CKINVDCx5p33_ASAP7_75t_R g2175 ( 
.A(n_1973),
.Y(n_2175)
);

CKINVDCx5p33_ASAP7_75t_R g2176 ( 
.A(n_1957),
.Y(n_2176)
);

CKINVDCx5p33_ASAP7_75t_R g2177 ( 
.A(n_2008),
.Y(n_2177)
);

CKINVDCx20_ASAP7_75t_R g2178 ( 
.A(n_2131),
.Y(n_2178)
);

AO22x2_ASAP7_75t_L g2179 ( 
.A1(n_1909),
.A2(n_1623),
.B1(n_1769),
.B2(n_1671),
.Y(n_2179)
);

CKINVDCx5p33_ASAP7_75t_R g2180 ( 
.A(n_2043),
.Y(n_2180)
);

INVx1_ASAP7_75t_SL g2181 ( 
.A(n_1970),
.Y(n_2181)
);

CKINVDCx5p33_ASAP7_75t_R g2182 ( 
.A(n_2117),
.Y(n_2182)
);

CKINVDCx5p33_ASAP7_75t_R g2183 ( 
.A(n_1984),
.Y(n_2183)
);

CKINVDCx5p33_ASAP7_75t_R g2184 ( 
.A(n_1987),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_2029),
.Y(n_2185)
);

BUFx3_ASAP7_75t_L g2186 ( 
.A(n_2116),
.Y(n_2186)
);

CKINVDCx5p33_ASAP7_75t_R g2187 ( 
.A(n_2035),
.Y(n_2187)
);

INVxp67_ASAP7_75t_L g2188 ( 
.A(n_2066),
.Y(n_2188)
);

OAI21x1_ASAP7_75t_L g2189 ( 
.A1(n_1946),
.A2(n_1333),
.B(n_1329),
.Y(n_2189)
);

INVx3_ASAP7_75t_L g2190 ( 
.A(n_1992),
.Y(n_2190)
);

CKINVDCx5p33_ASAP7_75t_R g2191 ( 
.A(n_2047),
.Y(n_2191)
);

CKINVDCx5p33_ASAP7_75t_R g2192 ( 
.A(n_2054),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_2029),
.Y(n_2193)
);

CKINVDCx5p33_ASAP7_75t_R g2194 ( 
.A(n_2086),
.Y(n_2194)
);

CKINVDCx5p33_ASAP7_75t_R g2195 ( 
.A(n_2097),
.Y(n_2195)
);

CKINVDCx5p33_ASAP7_75t_R g2196 ( 
.A(n_1944),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1990),
.Y(n_2197)
);

BUFx6f_ASAP7_75t_L g2198 ( 
.A(n_1901),
.Y(n_2198)
);

CKINVDCx20_ASAP7_75t_R g2199 ( 
.A(n_2024),
.Y(n_2199)
);

CKINVDCx5p33_ASAP7_75t_R g2200 ( 
.A(n_2077),
.Y(n_2200)
);

CKINVDCx5p33_ASAP7_75t_R g2201 ( 
.A(n_1953),
.Y(n_2201)
);

INVxp67_ASAP7_75t_L g2202 ( 
.A(n_2126),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1954),
.Y(n_2203)
);

CKINVDCx5p33_ASAP7_75t_R g2204 ( 
.A(n_1924),
.Y(n_2204)
);

CKINVDCx5p33_ASAP7_75t_R g2205 ( 
.A(n_1899),
.Y(n_2205)
);

CKINVDCx5p33_ASAP7_75t_R g2206 ( 
.A(n_2036),
.Y(n_2206)
);

NOR2xp67_ASAP7_75t_L g2207 ( 
.A(n_2056),
.B(n_1136),
.Y(n_2207)
);

CKINVDCx5p33_ASAP7_75t_R g2208 ( 
.A(n_2122),
.Y(n_2208)
);

CKINVDCx16_ASAP7_75t_R g2209 ( 
.A(n_2042),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1956),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_1896),
.B(n_1137),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1966),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_2006),
.Y(n_2213)
);

CKINVDCx20_ASAP7_75t_R g2214 ( 
.A(n_2152),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1969),
.Y(n_2215)
);

BUFx10_ASAP7_75t_L g2216 ( 
.A(n_1914),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_R g2217 ( 
.A(n_2109),
.B(n_1701),
.Y(n_2217)
);

CKINVDCx16_ASAP7_75t_R g2218 ( 
.A(n_1940),
.Y(n_2218)
);

BUFx3_ASAP7_75t_L g2219 ( 
.A(n_1892),
.Y(n_2219)
);

CKINVDCx5p33_ASAP7_75t_R g2220 ( 
.A(n_1893),
.Y(n_2220)
);

CKINVDCx5p33_ASAP7_75t_R g2221 ( 
.A(n_2016),
.Y(n_2221)
);

BUFx10_ASAP7_75t_L g2222 ( 
.A(n_1930),
.Y(n_2222)
);

CKINVDCx5p33_ASAP7_75t_R g2223 ( 
.A(n_2162),
.Y(n_2223)
);

HB1xp67_ASAP7_75t_L g2224 ( 
.A(n_2011),
.Y(n_2224)
);

NOR2xp33_ASAP7_75t_R g2225 ( 
.A(n_2133),
.B(n_1138),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_2022),
.Y(n_2226)
);

AOI21x1_ASAP7_75t_L g2227 ( 
.A1(n_1950),
.A2(n_1345),
.B(n_1334),
.Y(n_2227)
);

CKINVDCx5p33_ASAP7_75t_R g2228 ( 
.A(n_1962),
.Y(n_2228)
);

OAI22xp5_ASAP7_75t_SL g2229 ( 
.A1(n_1925),
.A2(n_1590),
.B1(n_1083),
.B2(n_1084),
.Y(n_2229)
);

AND3x2_ASAP7_75t_L g2230 ( 
.A(n_2096),
.B(n_2136),
.C(n_2107),
.Y(n_2230)
);

BUFx3_ASAP7_75t_L g2231 ( 
.A(n_1943),
.Y(n_2231)
);

CKINVDCx5p33_ASAP7_75t_R g2232 ( 
.A(n_2005),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1972),
.Y(n_2233)
);

CKINVDCx5p33_ASAP7_75t_R g2234 ( 
.A(n_2071),
.Y(n_2234)
);

CKINVDCx5p33_ASAP7_75t_R g2235 ( 
.A(n_2121),
.Y(n_2235)
);

CKINVDCx5p33_ASAP7_75t_R g2236 ( 
.A(n_1932),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1975),
.Y(n_2237)
);

CKINVDCx5p33_ASAP7_75t_R g2238 ( 
.A(n_2160),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1986),
.Y(n_2239)
);

CKINVDCx5p33_ASAP7_75t_R g2240 ( 
.A(n_1982),
.Y(n_2240)
);

BUFx3_ASAP7_75t_L g2241 ( 
.A(n_1974),
.Y(n_2241)
);

BUFx10_ASAP7_75t_L g2242 ( 
.A(n_1964),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1949),
.Y(n_2243)
);

CKINVDCx5p33_ASAP7_75t_R g2244 ( 
.A(n_1921),
.Y(n_2244)
);

NOR2xp67_ASAP7_75t_L g2245 ( 
.A(n_1904),
.B(n_2000),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1988),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2048),
.Y(n_2247)
);

CKINVDCx5p33_ASAP7_75t_R g2248 ( 
.A(n_1985),
.Y(n_2248)
);

BUFx6f_ASAP7_75t_L g2249 ( 
.A(n_1902),
.Y(n_2249)
);

NOR2xp67_ASAP7_75t_L g2250 ( 
.A(n_1958),
.B(n_1139),
.Y(n_2250)
);

NOR2xp33_ASAP7_75t_L g2251 ( 
.A(n_2040),
.B(n_2055),
.Y(n_2251)
);

NAND2xp33_ASAP7_75t_R g2252 ( 
.A(n_1947),
.B(n_1077),
.Y(n_2252)
);

BUFx3_ASAP7_75t_L g2253 ( 
.A(n_2146),
.Y(n_2253)
);

INVxp33_ASAP7_75t_L g2254 ( 
.A(n_2074),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2156),
.Y(n_2255)
);

CKINVDCx5p33_ASAP7_75t_R g2256 ( 
.A(n_2003),
.Y(n_2256)
);

AOI21x1_ASAP7_75t_L g2257 ( 
.A1(n_2060),
.A2(n_1350),
.B(n_1349),
.Y(n_2257)
);

INVx3_ASAP7_75t_L g2258 ( 
.A(n_2027),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1959),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2034),
.Y(n_2260)
);

CKINVDCx5p33_ASAP7_75t_R g2261 ( 
.A(n_2015),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_1961),
.Y(n_2262)
);

INVx3_ASAP7_75t_L g2263 ( 
.A(n_2049),
.Y(n_2263)
);

INVx3_ASAP7_75t_L g2264 ( 
.A(n_2051),
.Y(n_2264)
);

AO21x2_ASAP7_75t_L g2265 ( 
.A1(n_2091),
.A2(n_1411),
.B(n_1400),
.Y(n_2265)
);

CKINVDCx5p33_ASAP7_75t_R g2266 ( 
.A(n_2021),
.Y(n_2266)
);

CKINVDCx5p33_ASAP7_75t_R g2267 ( 
.A(n_2028),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1998),
.Y(n_2268)
);

NOR2xp33_ASAP7_75t_R g2269 ( 
.A(n_2106),
.B(n_1148),
.Y(n_2269)
);

NOR2xp67_ASAP7_75t_L g2270 ( 
.A(n_1996),
.B(n_1149),
.Y(n_2270)
);

CKINVDCx5p33_ASAP7_75t_R g2271 ( 
.A(n_2062),
.Y(n_2271)
);

CKINVDCx5p33_ASAP7_75t_R g2272 ( 
.A(n_2072),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_1967),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1976),
.Y(n_2274)
);

NOR2xp33_ASAP7_75t_R g2275 ( 
.A(n_2135),
.B(n_1151),
.Y(n_2275)
);

CKINVDCx5p33_ASAP7_75t_R g2276 ( 
.A(n_2087),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_2053),
.Y(n_2277)
);

BUFx2_ASAP7_75t_L g2278 ( 
.A(n_2010),
.Y(n_2278)
);

CKINVDCx5p33_ASAP7_75t_R g2279 ( 
.A(n_2045),
.Y(n_2279)
);

CKINVDCx5p33_ASAP7_75t_R g2280 ( 
.A(n_2058),
.Y(n_2280)
);

CKINVDCx5p33_ASAP7_75t_R g2281 ( 
.A(n_2010),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_2067),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1978),
.Y(n_2283)
);

CKINVDCx5p33_ASAP7_75t_R g2284 ( 
.A(n_2150),
.Y(n_2284)
);

CKINVDCx5p33_ASAP7_75t_R g2285 ( 
.A(n_2041),
.Y(n_2285)
);

NOR2xp67_ASAP7_75t_L g2286 ( 
.A(n_1996),
.B(n_1963),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1979),
.Y(n_2287)
);

CKINVDCx20_ASAP7_75t_R g2288 ( 
.A(n_1952),
.Y(n_2288)
);

CKINVDCx5p33_ASAP7_75t_R g2289 ( 
.A(n_2059),
.Y(n_2289)
);

CKINVDCx5p33_ASAP7_75t_R g2290 ( 
.A(n_1997),
.Y(n_2290)
);

AND2x2_ASAP7_75t_L g2291 ( 
.A(n_1983),
.B(n_1097),
.Y(n_2291)
);

NOR2xp33_ASAP7_75t_R g2292 ( 
.A(n_1918),
.B(n_1152),
.Y(n_2292)
);

CKINVDCx5p33_ASAP7_75t_R g2293 ( 
.A(n_2023),
.Y(n_2293)
);

NOR2xp33_ASAP7_75t_R g2294 ( 
.A(n_1995),
.B(n_1168),
.Y(n_2294)
);

CKINVDCx5p33_ASAP7_75t_R g2295 ( 
.A(n_2078),
.Y(n_2295)
);

CKINVDCx5p33_ASAP7_75t_R g2296 ( 
.A(n_1951),
.Y(n_2296)
);

CKINVDCx5p33_ASAP7_75t_R g2297 ( 
.A(n_1971),
.Y(n_2297)
);

CKINVDCx5p33_ASAP7_75t_R g2298 ( 
.A(n_1935),
.Y(n_2298)
);

NOR2x1p5_ASAP7_75t_L g2299 ( 
.A(n_1942),
.B(n_1088),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2018),
.Y(n_2300)
);

CKINVDCx5p33_ASAP7_75t_R g2301 ( 
.A(n_2009),
.Y(n_2301)
);

CKINVDCx5p33_ASAP7_75t_R g2302 ( 
.A(n_2026),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2025),
.Y(n_2303)
);

CKINVDCx5p33_ASAP7_75t_R g2304 ( 
.A(n_2037),
.Y(n_2304)
);

CKINVDCx5p33_ASAP7_75t_R g2305 ( 
.A(n_2119),
.Y(n_2305)
);

CKINVDCx5p33_ASAP7_75t_R g2306 ( 
.A(n_1945),
.Y(n_2306)
);

XNOR2xp5_ASAP7_75t_L g2307 ( 
.A(n_2151),
.B(n_1089),
.Y(n_2307)
);

CKINVDCx5p33_ASAP7_75t_R g2308 ( 
.A(n_1955),
.Y(n_2308)
);

CKINVDCx5p33_ASAP7_75t_R g2309 ( 
.A(n_1993),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2068),
.Y(n_2310)
);

INVxp67_ASAP7_75t_L g2311 ( 
.A(n_1999),
.Y(n_2311)
);

HB1xp67_ASAP7_75t_L g2312 ( 
.A(n_2083),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2039),
.Y(n_2313)
);

NOR2xp33_ASAP7_75t_R g2314 ( 
.A(n_2132),
.B(n_1170),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2080),
.Y(n_2315)
);

NOR2xp33_ASAP7_75t_R g2316 ( 
.A(n_1960),
.B(n_1172),
.Y(n_2316)
);

CKINVDCx5p33_ASAP7_75t_R g2317 ( 
.A(n_1989),
.Y(n_2317)
);

NOR2xp67_ASAP7_75t_L g2318 ( 
.A(n_1977),
.B(n_1980),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2111),
.Y(n_2319)
);

CKINVDCx5p33_ASAP7_75t_R g2320 ( 
.A(n_1991),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_1897),
.Y(n_2321)
);

CKINVDCx5p33_ASAP7_75t_R g2322 ( 
.A(n_2030),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_1898),
.Y(n_2323)
);

CKINVDCx5p33_ASAP7_75t_R g2324 ( 
.A(n_2061),
.Y(n_2324)
);

NOR2xp33_ASAP7_75t_L g2325 ( 
.A(n_2092),
.B(n_1401),
.Y(n_2325)
);

INVx3_ASAP7_75t_L g2326 ( 
.A(n_2088),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_2100),
.Y(n_2327)
);

NOR2xp33_ASAP7_75t_R g2328 ( 
.A(n_1912),
.B(n_1175),
.Y(n_2328)
);

BUFx10_ASAP7_75t_L g2329 ( 
.A(n_2120),
.Y(n_2329)
);

CKINVDCx20_ASAP7_75t_R g2330 ( 
.A(n_2082),
.Y(n_2330)
);

BUFx6f_ASAP7_75t_L g2331 ( 
.A(n_2104),
.Y(n_2331)
);

AND2x2_ASAP7_75t_L g2332 ( 
.A(n_2130),
.B(n_1097),
.Y(n_2332)
);

CKINVDCx20_ASAP7_75t_R g2333 ( 
.A(n_1948),
.Y(n_2333)
);

NOR2xp33_ASAP7_75t_R g2334 ( 
.A(n_1928),
.B(n_1181),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_1900),
.Y(n_2335)
);

NOR2xp33_ASAP7_75t_R g2336 ( 
.A(n_1907),
.B(n_1189),
.Y(n_2336)
);

NOR2xp33_ASAP7_75t_L g2337 ( 
.A(n_2159),
.B(n_1092),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_1916),
.Y(n_2338)
);

HB1xp67_ASAP7_75t_L g2339 ( 
.A(n_2124),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_2144),
.Y(n_2340)
);

CKINVDCx5p33_ASAP7_75t_R g2341 ( 
.A(n_2004),
.Y(n_2341)
);

INVxp67_ASAP7_75t_SL g2342 ( 
.A(n_2149),
.Y(n_2342)
);

CKINVDCx5p33_ASAP7_75t_R g2343 ( 
.A(n_2089),
.Y(n_2343)
);

CKINVDCx5p33_ASAP7_75t_R g2344 ( 
.A(n_2157),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_2001),
.Y(n_2345)
);

CKINVDCx5p33_ASAP7_75t_R g2346 ( 
.A(n_1903),
.Y(n_2346)
);

NOR2xp67_ASAP7_75t_L g2347 ( 
.A(n_2012),
.B(n_1205),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_1923),
.Y(n_2348)
);

CKINVDCx5p33_ASAP7_75t_R g2349 ( 
.A(n_1913),
.Y(n_2349)
);

CKINVDCx5p33_ASAP7_75t_R g2350 ( 
.A(n_1929),
.Y(n_2350)
);

CKINVDCx20_ASAP7_75t_R g2351 ( 
.A(n_1994),
.Y(n_2351)
);

CKINVDCx5p33_ASAP7_75t_R g2352 ( 
.A(n_1936),
.Y(n_2352)
);

CKINVDCx5p33_ASAP7_75t_R g2353 ( 
.A(n_1938),
.Y(n_2353)
);

CKINVDCx5p33_ASAP7_75t_R g2354 ( 
.A(n_2002),
.Y(n_2354)
);

CKINVDCx20_ASAP7_75t_R g2355 ( 
.A(n_1981),
.Y(n_2355)
);

CKINVDCx20_ASAP7_75t_R g2356 ( 
.A(n_1908),
.Y(n_2356)
);

CKINVDCx5p33_ASAP7_75t_R g2357 ( 
.A(n_2013),
.Y(n_2357)
);

CKINVDCx5p33_ASAP7_75t_R g2358 ( 
.A(n_2020),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_1926),
.Y(n_2359)
);

AOI21x1_ASAP7_75t_L g2360 ( 
.A1(n_1911),
.A2(n_1427),
.B(n_1417),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_1927),
.Y(n_2361)
);

CKINVDCx5p33_ASAP7_75t_R g2362 ( 
.A(n_2032),
.Y(n_2362)
);

INVx3_ASAP7_75t_L g2363 ( 
.A(n_2046),
.Y(n_2363)
);

CKINVDCx5p33_ASAP7_75t_R g2364 ( 
.A(n_2050),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_1933),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_2052),
.Y(n_2366)
);

NOR2xp33_ASAP7_75t_L g2367 ( 
.A(n_2063),
.B(n_1095),
.Y(n_2367)
);

CKINVDCx5p33_ASAP7_75t_R g2368 ( 
.A(n_2064),
.Y(n_2368)
);

CKINVDCx5p33_ASAP7_75t_R g2369 ( 
.A(n_2069),
.Y(n_2369)
);

BUFx2_ASAP7_75t_L g2370 ( 
.A(n_2070),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_1941),
.Y(n_2371)
);

AND2x4_ASAP7_75t_L g2372 ( 
.A(n_2073),
.B(n_1177),
.Y(n_2372)
);

OR2x2_ASAP7_75t_L g2373 ( 
.A(n_2084),
.B(n_1096),
.Y(n_2373)
);

INVxp67_ASAP7_75t_L g2374 ( 
.A(n_1906),
.Y(n_2374)
);

CKINVDCx20_ASAP7_75t_R g2375 ( 
.A(n_1934),
.Y(n_2375)
);

CKINVDCx5p33_ASAP7_75t_R g2376 ( 
.A(n_2090),
.Y(n_2376)
);

NOR2xp67_ASAP7_75t_L g2377 ( 
.A(n_2012),
.B(n_1213),
.Y(n_2377)
);

CKINVDCx16_ASAP7_75t_R g2378 ( 
.A(n_1905),
.Y(n_2378)
);

BUFx2_ASAP7_75t_L g2379 ( 
.A(n_2093),
.Y(n_2379)
);

CKINVDCx5p33_ASAP7_75t_R g2380 ( 
.A(n_2095),
.Y(n_2380)
);

CKINVDCx20_ASAP7_75t_R g2381 ( 
.A(n_2033),
.Y(n_2381)
);

AND2x2_ASAP7_75t_L g2382 ( 
.A(n_2098),
.B(n_1103),
.Y(n_2382)
);

CKINVDCx20_ASAP7_75t_R g2383 ( 
.A(n_2085),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2099),
.Y(n_2384)
);

CKINVDCx5p33_ASAP7_75t_R g2385 ( 
.A(n_2101),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_2108),
.Y(n_2386)
);

CKINVDCx5p33_ASAP7_75t_R g2387 ( 
.A(n_2110),
.Y(n_2387)
);

CKINVDCx5p33_ASAP7_75t_R g2388 ( 
.A(n_2112),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_2113),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2118),
.Y(n_2390)
);

BUFx10_ASAP7_75t_L g2391 ( 
.A(n_1894),
.Y(n_2391)
);

BUFx3_ASAP7_75t_L g2392 ( 
.A(n_2044),
.Y(n_2392)
);

CKINVDCx20_ASAP7_75t_R g2393 ( 
.A(n_2129),
.Y(n_2393)
);

BUFx6f_ASAP7_75t_L g2394 ( 
.A(n_2163),
.Y(n_2394)
);

CKINVDCx5p33_ASAP7_75t_R g2395 ( 
.A(n_2123),
.Y(n_2395)
);

CKINVDCx5p33_ASAP7_75t_R g2396 ( 
.A(n_2127),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2138),
.Y(n_2397)
);

AOI21x1_ASAP7_75t_L g2398 ( 
.A1(n_2007),
.A2(n_1434),
.B(n_1433),
.Y(n_2398)
);

BUFx10_ASAP7_75t_L g2399 ( 
.A(n_1895),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_2141),
.Y(n_2400)
);

CKINVDCx5p33_ASAP7_75t_R g2401 ( 
.A(n_2145),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2154),
.Y(n_2402)
);

CKINVDCx5p33_ASAP7_75t_R g2403 ( 
.A(n_2158),
.Y(n_2403)
);

BUFx10_ASAP7_75t_L g2404 ( 
.A(n_2038),
.Y(n_2404)
);

NAND2xp33_ASAP7_75t_L g2405 ( 
.A(n_2201),
.B(n_1215),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_SL g2406 ( 
.A(n_2284),
.B(n_1216),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2370),
.Y(n_2407)
);

INVx2_ASAP7_75t_L g2408 ( 
.A(n_2345),
.Y(n_2408)
);

INVx3_ASAP7_75t_L g2409 ( 
.A(n_2198),
.Y(n_2409)
);

BUFx6f_ASAP7_75t_L g2410 ( 
.A(n_2198),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2379),
.Y(n_2411)
);

BUFx2_ASAP7_75t_L g2412 ( 
.A(n_2199),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2366),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2169),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2174),
.Y(n_2415)
);

BUFx6f_ASAP7_75t_L g2416 ( 
.A(n_2198),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2251),
.B(n_2271),
.Y(n_2417)
);

AND2x2_ASAP7_75t_L g2418 ( 
.A(n_2291),
.B(n_2065),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2197),
.Y(n_2419)
);

AND2x6_ASAP7_75t_L g2420 ( 
.A(n_2332),
.B(n_1193),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2259),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2224),
.B(n_2075),
.Y(n_2422)
);

BUFx3_ASAP7_75t_L g2423 ( 
.A(n_2186),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2262),
.Y(n_2424)
);

BUFx3_ASAP7_75t_L g2425 ( 
.A(n_2346),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2321),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2323),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_2272),
.B(n_1450),
.Y(n_2428)
);

CKINVDCx5p33_ASAP7_75t_R g2429 ( 
.A(n_2164),
.Y(n_2429)
);

AND2x2_ASAP7_75t_L g2430 ( 
.A(n_2317),
.B(n_2076),
.Y(n_2430)
);

NAND2x1p5_ASAP7_75t_L g2431 ( 
.A(n_2219),
.B(n_2044),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2335),
.Y(n_2432)
);

AND2x2_ASAP7_75t_L g2433 ( 
.A(n_2320),
.B(n_2079),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2276),
.B(n_1466),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2386),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2244),
.B(n_1478),
.Y(n_2436)
);

AND2x6_ASAP7_75t_L g2437 ( 
.A(n_2382),
.B(n_1198),
.Y(n_2437)
);

HB1xp67_ASAP7_75t_L g2438 ( 
.A(n_2181),
.Y(n_2438)
);

INVx5_ASAP7_75t_L g2439 ( 
.A(n_2242),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2338),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2348),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2359),
.Y(n_2442)
);

BUFx6f_ASAP7_75t_L g2443 ( 
.A(n_2249),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2361),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2365),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_SL g2446 ( 
.A(n_2248),
.B(n_1221),
.Y(n_2446)
);

INVx3_ASAP7_75t_L g2447 ( 
.A(n_2249),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_SL g2448 ( 
.A(n_2256),
.B(n_1223),
.Y(n_2448)
);

AND2x2_ASAP7_75t_L g2449 ( 
.A(n_2311),
.B(n_2081),
.Y(n_2449)
);

BUFx2_ASAP7_75t_L g2450 ( 
.A(n_2296),
.Y(n_2450)
);

AND2x6_ASAP7_75t_L g2451 ( 
.A(n_2337),
.B(n_1199),
.Y(n_2451)
);

OR2x6_ASAP7_75t_L g2452 ( 
.A(n_2278),
.B(n_1141),
.Y(n_2452)
);

INVx4_ASAP7_75t_SL g2453 ( 
.A(n_2249),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_SL g2454 ( 
.A(n_2261),
.B(n_1232),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2371),
.Y(n_2455)
);

AND2x4_ASAP7_75t_L g2456 ( 
.A(n_2231),
.B(n_1910),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2389),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2400),
.Y(n_2458)
);

BUFx2_ASAP7_75t_L g2459 ( 
.A(n_2298),
.Y(n_2459)
);

BUFx2_ASAP7_75t_L g2460 ( 
.A(n_2166),
.Y(n_2460)
);

OR2x6_ASAP7_75t_L g2461 ( 
.A(n_2241),
.B(n_1157),
.Y(n_2461)
);

INVx5_ASAP7_75t_L g2462 ( 
.A(n_2242),
.Y(n_2462)
);

INVx3_ASAP7_75t_L g2463 ( 
.A(n_2331),
.Y(n_2463)
);

CKINVDCx5p33_ASAP7_75t_R g2464 ( 
.A(n_2165),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2384),
.Y(n_2465)
);

INVx2_ASAP7_75t_SL g2466 ( 
.A(n_2222),
.Y(n_2466)
);

INVxp67_ASAP7_75t_L g2467 ( 
.A(n_2252),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_SL g2468 ( 
.A(n_2266),
.B(n_1233),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2390),
.Y(n_2469)
);

INVx2_ASAP7_75t_L g2470 ( 
.A(n_2363),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2397),
.Y(n_2471)
);

NOR2xp33_ASAP7_75t_L g2472 ( 
.A(n_2267),
.B(n_1102),
.Y(n_2472)
);

INVx2_ASAP7_75t_L g2473 ( 
.A(n_2363),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_L g2474 ( 
.A(n_2265),
.B(n_1508),
.Y(n_2474)
);

BUFx6f_ASAP7_75t_L g2475 ( 
.A(n_2331),
.Y(n_2475)
);

CKINVDCx8_ASAP7_75t_R g2476 ( 
.A(n_2171),
.Y(n_2476)
);

AND2x6_ASAP7_75t_L g2477 ( 
.A(n_2246),
.B(n_1203),
.Y(n_2477)
);

AND2x2_ASAP7_75t_L g2478 ( 
.A(n_2222),
.B(n_2094),
.Y(n_2478)
);

AND2x4_ASAP7_75t_L g2479 ( 
.A(n_2253),
.B(n_1915),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2402),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_SL g2481 ( 
.A(n_2309),
.B(n_1235),
.Y(n_2481)
);

NOR2xp33_ASAP7_75t_SL g2482 ( 
.A(n_2170),
.B(n_1103),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2273),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2274),
.Y(n_2484)
);

AND2x6_ASAP7_75t_L g2485 ( 
.A(n_2247),
.B(n_1204),
.Y(n_2485)
);

INVxp67_ASAP7_75t_SL g2486 ( 
.A(n_2374),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2283),
.Y(n_2487)
);

INVx1_ASAP7_75t_SL g2488 ( 
.A(n_2205),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2287),
.Y(n_2489)
);

NOR2xp33_ASAP7_75t_L g2490 ( 
.A(n_2204),
.B(n_1105),
.Y(n_2490)
);

INVx2_ASAP7_75t_L g2491 ( 
.A(n_2243),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2372),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2308),
.B(n_2102),
.Y(n_2493)
);

INVx3_ASAP7_75t_L g2494 ( 
.A(n_2331),
.Y(n_2494)
);

HB1xp67_ASAP7_75t_L g2495 ( 
.A(n_2188),
.Y(n_2495)
);

NOR2xp33_ASAP7_75t_L g2496 ( 
.A(n_2230),
.B(n_1108),
.Y(n_2496)
);

INVx2_ASAP7_75t_SL g2497 ( 
.A(n_2373),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2265),
.B(n_1518),
.Y(n_2498)
);

BUFx3_ASAP7_75t_L g2499 ( 
.A(n_2349),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2372),
.Y(n_2500)
);

INVx3_ASAP7_75t_L g2501 ( 
.A(n_2258),
.Y(n_2501)
);

INVx3_ASAP7_75t_L g2502 ( 
.A(n_2258),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2300),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2190),
.B(n_1530),
.Y(n_2504)
);

AND2x4_ASAP7_75t_L g2505 ( 
.A(n_2263),
.B(n_1917),
.Y(n_2505)
);

BUFx6f_ASAP7_75t_L g2506 ( 
.A(n_2392),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2190),
.B(n_2211),
.Y(n_2507)
);

INVxp67_ASAP7_75t_SL g2508 ( 
.A(n_2318),
.Y(n_2508)
);

AND2x2_ASAP7_75t_L g2509 ( 
.A(n_2301),
.B(n_2302),
.Y(n_2509)
);

AND2x2_ASAP7_75t_L g2510 ( 
.A(n_2304),
.B(n_2305),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2303),
.Y(n_2511)
);

AND2x4_ASAP7_75t_L g2512 ( 
.A(n_2263),
.B(n_1920),
.Y(n_2512)
);

BUFx3_ASAP7_75t_L g2513 ( 
.A(n_2350),
.Y(n_2513)
);

INVx4_ASAP7_75t_L g2514 ( 
.A(n_2352),
.Y(n_2514)
);

OR2x2_ASAP7_75t_L g2515 ( 
.A(n_2202),
.B(n_2105),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_SL g2516 ( 
.A(n_2245),
.B(n_1236),
.Y(n_2516)
);

CKINVDCx5p33_ASAP7_75t_R g2517 ( 
.A(n_2196),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2313),
.Y(n_2518)
);

OR2x2_ASAP7_75t_SL g2519 ( 
.A(n_2209),
.B(n_1224),
.Y(n_2519)
);

AND2x2_ASAP7_75t_L g2520 ( 
.A(n_2240),
.B(n_2114),
.Y(n_2520)
);

NAND3x1_ASAP7_75t_L g2521 ( 
.A(n_2254),
.B(n_1244),
.C(n_1207),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2315),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2319),
.Y(n_2523)
);

BUFx2_ASAP7_75t_L g2524 ( 
.A(n_2173),
.Y(n_2524)
);

INVxp67_ASAP7_75t_L g2525 ( 
.A(n_2325),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2354),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2185),
.Y(n_2527)
);

AND2x4_ASAP7_75t_L g2528 ( 
.A(n_2264),
.B(n_1937),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2357),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2168),
.B(n_1548),
.Y(n_2530)
);

AND2x4_ASAP7_75t_L g2531 ( 
.A(n_2264),
.B(n_1939),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2358),
.Y(n_2532)
);

INVx3_ASAP7_75t_L g2533 ( 
.A(n_2326),
.Y(n_2533)
);

INVx3_ASAP7_75t_L g2534 ( 
.A(n_2326),
.Y(n_2534)
);

AND2x4_ASAP7_75t_L g2535 ( 
.A(n_2213),
.B(n_2115),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2362),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_SL g2537 ( 
.A(n_2269),
.B(n_2275),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_L g2538 ( 
.A(n_2250),
.B(n_2294),
.Y(n_2538)
);

CKINVDCx20_ASAP7_75t_R g2539 ( 
.A(n_2178),
.Y(n_2539)
);

NOR2xp33_ASAP7_75t_R g2540 ( 
.A(n_2200),
.B(n_1237),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2364),
.Y(n_2541)
);

BUFx3_ASAP7_75t_L g2542 ( 
.A(n_2353),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_2193),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2368),
.Y(n_2544)
);

INVxp67_ASAP7_75t_L g2545 ( 
.A(n_2220),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2369),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_2314),
.B(n_1559),
.Y(n_2547)
);

BUFx6f_ASAP7_75t_L g2548 ( 
.A(n_2329),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2376),
.Y(n_2549)
);

INVx5_ASAP7_75t_L g2550 ( 
.A(n_2329),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2380),
.Y(n_2551)
);

HB1xp67_ASAP7_75t_L g2552 ( 
.A(n_2221),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2385),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_2387),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2388),
.Y(n_2555)
);

INVx4_ASAP7_75t_SL g2556 ( 
.A(n_2307),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_L g2557 ( 
.A(n_2292),
.B(n_1565),
.Y(n_2557)
);

AND2x2_ASAP7_75t_L g2558 ( 
.A(n_2223),
.B(n_2125),
.Y(n_2558)
);

INVx2_ASAP7_75t_SL g2559 ( 
.A(n_2299),
.Y(n_2559)
);

INVxp67_ASAP7_75t_SL g2560 ( 
.A(n_2312),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_SL g2561 ( 
.A(n_2187),
.B(n_1251),
.Y(n_2561)
);

INVx3_ASAP7_75t_L g2562 ( 
.A(n_2226),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_SL g2563 ( 
.A(n_2191),
.B(n_1252),
.Y(n_2563)
);

NOR2xp33_ASAP7_75t_SL g2564 ( 
.A(n_2175),
.B(n_1182),
.Y(n_2564)
);

INVx5_ASAP7_75t_L g2565 ( 
.A(n_2391),
.Y(n_2565)
);

AND2x4_ASAP7_75t_L g2566 ( 
.A(n_2260),
.B(n_2128),
.Y(n_2566)
);

CKINVDCx5p33_ASAP7_75t_R g2567 ( 
.A(n_2192),
.Y(n_2567)
);

INVx2_ASAP7_75t_SL g2568 ( 
.A(n_2391),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2395),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2396),
.B(n_1582),
.Y(n_2570)
);

AOI22xp5_ASAP7_75t_L g2571 ( 
.A1(n_2417),
.A2(n_2351),
.B1(n_2375),
.B2(n_2356),
.Y(n_2571)
);

OAI221xp5_ASAP7_75t_L g2572 ( 
.A1(n_2428),
.A2(n_2229),
.B1(n_2297),
.B2(n_2236),
.C(n_2228),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_2408),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2414),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2415),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_2507),
.B(n_2194),
.Y(n_2576)
);

BUFx6f_ASAP7_75t_L g2577 ( 
.A(n_2475),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2434),
.B(n_2195),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_SL g2579 ( 
.A(n_2467),
.B(n_2183),
.Y(n_2579)
);

INVx4_ASAP7_75t_L g2580 ( 
.A(n_2548),
.Y(n_2580)
);

AOI22x1_ASAP7_75t_L g2581 ( 
.A1(n_2503),
.A2(n_2285),
.B1(n_2289),
.B2(n_2179),
.Y(n_2581)
);

INVx3_ASAP7_75t_L g2582 ( 
.A(n_2475),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2419),
.Y(n_2583)
);

OR2x6_ASAP7_75t_L g2584 ( 
.A(n_2425),
.B(n_2277),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2413),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2421),
.Y(n_2586)
);

AOI22xp33_ASAP7_75t_L g2587 ( 
.A1(n_2474),
.A2(n_2355),
.B1(n_2383),
.B2(n_2381),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_L g2588 ( 
.A(n_2436),
.B(n_2207),
.Y(n_2588)
);

CKINVDCx5p33_ASAP7_75t_R g2589 ( 
.A(n_2429),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2424),
.Y(n_2590)
);

NOR2xp33_ASAP7_75t_L g2591 ( 
.A(n_2490),
.B(n_2206),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2426),
.Y(n_2592)
);

AOI22xp5_ASAP7_75t_L g2593 ( 
.A1(n_2472),
.A2(n_2393),
.B1(n_2208),
.B2(n_2214),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_2435),
.Y(n_2594)
);

HB1xp67_ASAP7_75t_L g2595 ( 
.A(n_2438),
.Y(n_2595)
);

OAI22xp5_ASAP7_75t_L g2596 ( 
.A1(n_2525),
.A2(n_2293),
.B1(n_2184),
.B2(n_2281),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2427),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2432),
.Y(n_2598)
);

INVx2_ASAP7_75t_L g2599 ( 
.A(n_2440),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2441),
.Y(n_2600)
);

INVxp67_ASAP7_75t_L g2601 ( 
.A(n_2460),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2442),
.Y(n_2602)
);

INVxp67_ASAP7_75t_L g2603 ( 
.A(n_2495),
.Y(n_2603)
);

OAI22xp5_ASAP7_75t_SL g2604 ( 
.A1(n_2517),
.A2(n_2218),
.B1(n_2330),
.B2(n_2288),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2444),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2445),
.Y(n_2606)
);

BUFx2_ASAP7_75t_L g2607 ( 
.A(n_2412),
.Y(n_2607)
);

OAI221xp5_ASAP7_75t_L g2608 ( 
.A1(n_2570),
.A2(n_2341),
.B1(n_2343),
.B2(n_2367),
.C(n_2255),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2455),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_2530),
.B(n_2401),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2509),
.B(n_2217),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2492),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2457),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_SL g2614 ( 
.A(n_2565),
.B(n_2216),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2500),
.Y(n_2615)
);

AND2x4_ASAP7_75t_L g2616 ( 
.A(n_2423),
.B(n_2339),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2458),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_SL g2618 ( 
.A(n_2565),
.B(n_2216),
.Y(n_2618)
);

INVx2_ASAP7_75t_L g2619 ( 
.A(n_2491),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2465),
.Y(n_2620)
);

INVx2_ASAP7_75t_L g2621 ( 
.A(n_2469),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2471),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2480),
.Y(n_2623)
);

NAND2x1p5_ASAP7_75t_L g2624 ( 
.A(n_2514),
.B(n_2268),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2483),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2484),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2486),
.B(n_2403),
.Y(n_2627)
);

BUFx2_ASAP7_75t_L g2628 ( 
.A(n_2552),
.Y(n_2628)
);

A2O1A1Ixp33_ASAP7_75t_L g2629 ( 
.A1(n_2498),
.A2(n_2189),
.B(n_1615),
.C(n_1616),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_SL g2630 ( 
.A(n_2546),
.B(n_2225),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_L g2631 ( 
.A(n_2538),
.B(n_2179),
.Y(n_2631)
);

A2O1A1Ixp33_ASAP7_75t_L g2632 ( 
.A1(n_2496),
.A2(n_1620),
.B(n_1632),
.C(n_1598),
.Y(n_2632)
);

AOI22xp33_ASAP7_75t_L g2633 ( 
.A1(n_2451),
.A2(n_2394),
.B1(n_1638),
.B2(n_1653),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2487),
.Y(n_2634)
);

INVxp67_ASAP7_75t_L g2635 ( 
.A(n_2558),
.Y(n_2635)
);

OR2x6_ASAP7_75t_SL g2636 ( 
.A(n_2567),
.B(n_2232),
.Y(n_2636)
);

AND2x4_ASAP7_75t_L g2637 ( 
.A(n_2499),
.B(n_2344),
.Y(n_2637)
);

INVxp67_ASAP7_75t_L g2638 ( 
.A(n_2493),
.Y(n_2638)
);

NOR2xp33_ASAP7_75t_L g2639 ( 
.A(n_2551),
.B(n_2172),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2489),
.Y(n_2640)
);

NAND2xp33_ASAP7_75t_L g2641 ( 
.A(n_2451),
.B(n_2394),
.Y(n_2641)
);

AO22x2_ASAP7_75t_L g2642 ( 
.A1(n_2556),
.A2(n_1249),
.B1(n_1258),
.B2(n_1257),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2449),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2518),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2523),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_2508),
.B(n_2167),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2470),
.Y(n_2647)
);

BUFx6f_ASAP7_75t_L g2648 ( 
.A(n_2410),
.Y(n_2648)
);

HB1xp67_ASAP7_75t_L g2649 ( 
.A(n_2407),
.Y(n_2649)
);

AND2x4_ASAP7_75t_L g2650 ( 
.A(n_2513),
.B(n_2282),
.Y(n_2650)
);

OR2x2_ASAP7_75t_L g2651 ( 
.A(n_2488),
.B(n_2378),
.Y(n_2651)
);

CKINVDCx20_ASAP7_75t_R g2652 ( 
.A(n_2539),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2547),
.B(n_2316),
.Y(n_2653)
);

AOI22xp33_ASAP7_75t_L g2654 ( 
.A1(n_2437),
.A2(n_2394),
.B1(n_1658),
.B2(n_1659),
.Y(n_2654)
);

AOI22xp33_ASAP7_75t_L g2655 ( 
.A1(n_2437),
.A2(n_1677),
.B1(n_1688),
.B2(n_1637),
.Y(n_2655)
);

CKINVDCx5p33_ASAP7_75t_R g2656 ( 
.A(n_2464),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2473),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2511),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2522),
.Y(n_2659)
);

AOI22xp33_ASAP7_75t_L g2660 ( 
.A1(n_2504),
.A2(n_1698),
.B1(n_1710),
.B2(n_1689),
.Y(n_2660)
);

AND2x4_ASAP7_75t_L g2661 ( 
.A(n_2542),
.B(n_2453),
.Y(n_2661)
);

NOR2xp33_ASAP7_75t_L g2662 ( 
.A(n_2554),
.B(n_2333),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2535),
.Y(n_2663)
);

AND2x4_ASAP7_75t_L g2664 ( 
.A(n_2550),
.B(n_2310),
.Y(n_2664)
);

AND2x4_ASAP7_75t_L g2665 ( 
.A(n_2550),
.B(n_2327),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2566),
.Y(n_2666)
);

AO22x2_ASAP7_75t_L g2667 ( 
.A1(n_2510),
.A2(n_1291),
.B1(n_1295),
.B2(n_1259),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2422),
.Y(n_2668)
);

INVx2_ASAP7_75t_SL g2669 ( 
.A(n_2430),
.Y(n_2669)
);

AOI21xp5_ASAP7_75t_L g2670 ( 
.A1(n_2588),
.A2(n_2537),
.B(n_2516),
.Y(n_2670)
);

AOI22xp5_ASAP7_75t_L g2671 ( 
.A1(n_2591),
.A2(n_2405),
.B1(n_2497),
.B2(n_2406),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_L g2672 ( 
.A(n_2576),
.B(n_2526),
.Y(n_2672)
);

AOI21xp5_ASAP7_75t_L g2673 ( 
.A1(n_2641),
.A2(n_2557),
.B(n_2559),
.Y(n_2673)
);

OAI21xp5_ASAP7_75t_L g2674 ( 
.A1(n_2631),
.A2(n_2448),
.B(n_2446),
.Y(n_2674)
);

AOI21xp5_ASAP7_75t_L g2675 ( 
.A1(n_2653),
.A2(n_2468),
.B(n_2454),
.Y(n_2675)
);

AOI21xp5_ASAP7_75t_L g2676 ( 
.A1(n_2610),
.A2(n_2418),
.B(n_2560),
.Y(n_2676)
);

AOI21xp5_ASAP7_75t_L g2677 ( 
.A1(n_2629),
.A2(n_2478),
.B(n_2481),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2574),
.Y(n_2678)
);

CKINVDCx20_ASAP7_75t_R g2679 ( 
.A(n_2652),
.Y(n_2679)
);

AOI21xp5_ASAP7_75t_L g2680 ( 
.A1(n_2578),
.A2(n_2563),
.B(n_2561),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2599),
.Y(n_2681)
);

OAI21x1_ASAP7_75t_L g2682 ( 
.A1(n_2613),
.A2(n_2398),
.B(n_2360),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2575),
.Y(n_2683)
);

AOI21xp5_ASAP7_75t_L g2684 ( 
.A1(n_2646),
.A2(n_2627),
.B(n_2630),
.Y(n_2684)
);

AOI33xp33_ASAP7_75t_L g2685 ( 
.A1(n_2668),
.A2(n_2643),
.A3(n_2529),
.B1(n_2532),
.B2(n_2544),
.B3(n_2541),
.Y(n_2685)
);

AND2x4_ASAP7_75t_L g2686 ( 
.A(n_2661),
.B(n_2456),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_L g2687 ( 
.A(n_2583),
.B(n_2536),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2609),
.Y(n_2688)
);

OAI22xp5_ASAP7_75t_L g2689 ( 
.A1(n_2587),
.A2(n_2553),
.B1(n_2555),
.B2(n_2549),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2621),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_SL g2691 ( 
.A(n_2669),
.B(n_2569),
.Y(n_2691)
);

HB1xp67_ASAP7_75t_L g2692 ( 
.A(n_2595),
.Y(n_2692)
);

OAI22xp5_ASAP7_75t_L g2693 ( 
.A1(n_2571),
.A2(n_2545),
.B1(n_2568),
.B2(n_2519),
.Y(n_2693)
);

AOI21x1_ASAP7_75t_L g2694 ( 
.A1(n_2647),
.A2(n_2257),
.B(n_2227),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2586),
.Y(n_2695)
);

AOI21x1_ASAP7_75t_L g2696 ( 
.A1(n_2657),
.A2(n_2543),
.B(n_2527),
.Y(n_2696)
);

AOI21xp5_ASAP7_75t_L g2697 ( 
.A1(n_2573),
.A2(n_2433),
.B(n_2411),
.Y(n_2697)
);

OAI21xp5_ASAP7_75t_L g2698 ( 
.A1(n_2590),
.A2(n_2521),
.B(n_2520),
.Y(n_2698)
);

AOI21x1_ASAP7_75t_L g2699 ( 
.A1(n_2617),
.A2(n_2057),
.B(n_2031),
.Y(n_2699)
);

INVx2_ASAP7_75t_SL g2700 ( 
.A(n_2577),
.Y(n_2700)
);

AO32x1_ASAP7_75t_L g2701 ( 
.A1(n_2612),
.A2(n_1311),
.A3(n_1314),
.B1(n_1301),
.B2(n_1297),
.Y(n_2701)
);

OAI22xp5_ASAP7_75t_L g2702 ( 
.A1(n_2638),
.A2(n_2459),
.B1(n_2450),
.B2(n_2466),
.Y(n_2702)
);

INVx2_ASAP7_75t_SL g2703 ( 
.A(n_2577),
.Y(n_2703)
);

AND2x4_ASAP7_75t_L g2704 ( 
.A(n_2580),
.B(n_2479),
.Y(n_2704)
);

NOR2x1_ASAP7_75t_L g2705 ( 
.A(n_2611),
.B(n_2637),
.Y(n_2705)
);

NOR2xp33_ASAP7_75t_SL g2706 ( 
.A(n_2589),
.B(n_2176),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2592),
.B(n_2420),
.Y(n_2707)
);

OAI21xp5_ASAP7_75t_L g2708 ( 
.A1(n_2597),
.A2(n_2515),
.B(n_2420),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2598),
.Y(n_2709)
);

O2A1O1Ixp33_ASAP7_75t_L g2710 ( 
.A1(n_2572),
.A2(n_2482),
.B(n_2452),
.C(n_2501),
.Y(n_2710)
);

OAI21xp5_ASAP7_75t_L g2711 ( 
.A1(n_2600),
.A2(n_1715),
.B(n_1712),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2585),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_2594),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2620),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2602),
.B(n_2477),
.Y(n_2715)
);

BUFx2_ASAP7_75t_L g2716 ( 
.A(n_2607),
.Y(n_2716)
);

AOI22xp33_ASAP7_75t_L g2717 ( 
.A1(n_2581),
.A2(n_2295),
.B1(n_2485),
.B2(n_2477),
.Y(n_2717)
);

OAI22xp5_ASAP7_75t_L g2718 ( 
.A1(n_2635),
.A2(n_2462),
.B1(n_2439),
.B2(n_2548),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2622),
.Y(n_2719)
);

BUFx2_ASAP7_75t_L g2720 ( 
.A(n_2628),
.Y(n_2720)
);

NOR2xp67_ASAP7_75t_L g2721 ( 
.A(n_2656),
.B(n_2439),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_SL g2722 ( 
.A(n_2662),
.B(n_2462),
.Y(n_2722)
);

AOI21xp5_ASAP7_75t_L g2723 ( 
.A1(n_2619),
.A2(n_2324),
.B(n_2322),
.Y(n_2723)
);

AOI22xp33_ASAP7_75t_L g2724 ( 
.A1(n_2605),
.A2(n_2485),
.B1(n_1732),
.B2(n_1749),
.Y(n_2724)
);

NOR2xp33_ASAP7_75t_L g2725 ( 
.A(n_2593),
.B(n_2524),
.Y(n_2725)
);

OAI21xp5_ASAP7_75t_L g2726 ( 
.A1(n_2606),
.A2(n_1751),
.B(n_1725),
.Y(n_2726)
);

CKINVDCx20_ASAP7_75t_R g2727 ( 
.A(n_2604),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2623),
.B(n_2540),
.Y(n_2728)
);

NOR3xp33_ASAP7_75t_L g2729 ( 
.A(n_2639),
.B(n_2290),
.C(n_2238),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_L g2730 ( 
.A(n_2625),
.B(n_2463),
.Y(n_2730)
);

AOI21xp5_ASAP7_75t_L g2731 ( 
.A1(n_2633),
.A2(n_2533),
.B(n_2502),
.Y(n_2731)
);

HB1xp67_ASAP7_75t_L g2732 ( 
.A(n_2649),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2626),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2634),
.B(n_2494),
.Y(n_2734)
);

OAI21xp5_ASAP7_75t_L g2735 ( 
.A1(n_2640),
.A2(n_2645),
.B(n_2644),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2615),
.B(n_2534),
.Y(n_2736)
);

OAI21xp5_ASAP7_75t_L g2737 ( 
.A1(n_2658),
.A2(n_1768),
.B(n_2505),
.Y(n_2737)
);

O2A1O1Ixp5_ASAP7_75t_L g2738 ( 
.A1(n_2632),
.A2(n_2409),
.B(n_2447),
.C(n_2562),
.Y(n_2738)
);

OAI22xp5_ASAP7_75t_L g2739 ( 
.A1(n_2654),
.A2(n_2476),
.B1(n_2416),
.B2(n_2443),
.Y(n_2739)
);

AND2x4_ASAP7_75t_L g2740 ( 
.A(n_2650),
.B(n_2506),
.Y(n_2740)
);

O2A1O1Ixp33_ASAP7_75t_L g2741 ( 
.A1(n_2608),
.A2(n_2461),
.B(n_1331),
.C(n_1338),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_L g2742 ( 
.A(n_2659),
.B(n_2512),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2660),
.B(n_2528),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2655),
.B(n_2531),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_2663),
.Y(n_2745)
);

A2O1A1Ixp33_ASAP7_75t_L g2746 ( 
.A1(n_2666),
.A2(n_2579),
.B(n_2651),
.C(n_2603),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_L g2747 ( 
.A(n_2582),
.B(n_2410),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2648),
.B(n_2416),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2648),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_SL g2750 ( 
.A(n_2601),
.B(n_2596),
.Y(n_2750)
);

AOI21xp5_ASAP7_75t_L g2751 ( 
.A1(n_2616),
.A2(n_2342),
.B(n_2443),
.Y(n_2751)
);

AOI21xp5_ASAP7_75t_L g2752 ( 
.A1(n_2664),
.A2(n_1166),
.B(n_1153),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2667),
.B(n_2336),
.Y(n_2753)
);

INVxp67_ASAP7_75t_L g2754 ( 
.A(n_2692),
.Y(n_2754)
);

INVx2_ASAP7_75t_L g2755 ( 
.A(n_2714),
.Y(n_2755)
);

AND2x2_ASAP7_75t_L g2756 ( 
.A(n_2705),
.B(n_2667),
.Y(n_2756)
);

O2A1O1Ixp33_ASAP7_75t_L g2757 ( 
.A1(n_2689),
.A2(n_2614),
.B(n_2618),
.C(n_2564),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2678),
.Y(n_2758)
);

AOI21xp5_ASAP7_75t_L g2759 ( 
.A1(n_2677),
.A2(n_2624),
.B(n_2584),
.Y(n_2759)
);

AOI21xp5_ASAP7_75t_L g2760 ( 
.A1(n_2670),
.A2(n_2584),
.B(n_2665),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2672),
.B(n_2399),
.Y(n_2761)
);

AND2x2_ASAP7_75t_L g2762 ( 
.A(n_2698),
.B(n_2732),
.Y(n_2762)
);

NAND3xp33_ASAP7_75t_SL g2763 ( 
.A(n_2671),
.B(n_2180),
.C(n_2177),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2676),
.B(n_2399),
.Y(n_2764)
);

OAI22xp5_ASAP7_75t_L g2765 ( 
.A1(n_2687),
.A2(n_2642),
.B1(n_2636),
.B2(n_2280),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_2684),
.B(n_2404),
.Y(n_2766)
);

BUFx2_ASAP7_75t_L g2767 ( 
.A(n_2720),
.Y(n_2767)
);

A2O1A1Ixp33_ASAP7_75t_L g2768 ( 
.A1(n_2674),
.A2(n_2210),
.B(n_2212),
.C(n_2203),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2719),
.B(n_2404),
.Y(n_2769)
);

AOI21xp5_ASAP7_75t_L g2770 ( 
.A1(n_2675),
.A2(n_1166),
.B(n_1153),
.Y(n_2770)
);

BUFx12f_ASAP7_75t_L g2771 ( 
.A(n_2716),
.Y(n_2771)
);

O2A1O1Ixp33_ASAP7_75t_L g2772 ( 
.A1(n_2741),
.A2(n_2233),
.B(n_2237),
.C(n_2215),
.Y(n_2772)
);

OAI21xp33_ASAP7_75t_SL g2773 ( 
.A1(n_2685),
.A2(n_1341),
.B(n_1330),
.Y(n_2773)
);

AOI21xp5_ASAP7_75t_L g2774 ( 
.A1(n_2680),
.A2(n_1166),
.B(n_1153),
.Y(n_2774)
);

INVxp67_ASAP7_75t_SL g2775 ( 
.A(n_2748),
.Y(n_2775)
);

INVx3_ASAP7_75t_L g2776 ( 
.A(n_2704),
.Y(n_2776)
);

A2O1A1Ixp33_ASAP7_75t_L g2777 ( 
.A1(n_2708),
.A2(n_2239),
.B(n_2340),
.C(n_1356),
.Y(n_2777)
);

O2A1O1Ixp33_ASAP7_75t_L g2778 ( 
.A1(n_2746),
.A2(n_1358),
.B(n_1371),
.C(n_1343),
.Y(n_2778)
);

O2A1O1Ixp33_ASAP7_75t_L g2779 ( 
.A1(n_2753),
.A2(n_1383),
.B(n_1386),
.C(n_1374),
.Y(n_2779)
);

OAI22xp5_ASAP7_75t_L g2780 ( 
.A1(n_2735),
.A2(n_2642),
.B1(n_2279),
.B2(n_1263),
.Y(n_2780)
);

AOI22xp33_ASAP7_75t_L g2781 ( 
.A1(n_2725),
.A2(n_2334),
.B1(n_2328),
.B2(n_2506),
.Y(n_2781)
);

AND2x4_ASAP7_75t_L g2782 ( 
.A(n_2740),
.B(n_2182),
.Y(n_2782)
);

O2A1O1Ixp33_ASAP7_75t_L g2783 ( 
.A1(n_2693),
.A2(n_1398),
.B(n_1405),
.C(n_1392),
.Y(n_2783)
);

NOR2xp33_ASAP7_75t_R g2784 ( 
.A(n_2679),
.B(n_2234),
.Y(n_2784)
);

AND2x4_ASAP7_75t_L g2785 ( 
.A(n_2686),
.B(n_2704),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_SL g2786 ( 
.A(n_2728),
.B(n_2431),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2683),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_SL g2788 ( 
.A(n_2721),
.B(n_2306),
.Y(n_2788)
);

NOR2xp33_ASAP7_75t_L g2789 ( 
.A(n_2750),
.B(n_2235),
.Y(n_2789)
);

AOI21xp5_ASAP7_75t_L g2790 ( 
.A1(n_2673),
.A2(n_1363),
.B(n_1351),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_L g2791 ( 
.A(n_2695),
.B(n_2709),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2733),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_SL g2793 ( 
.A(n_2706),
.B(n_2286),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2681),
.B(n_2134),
.Y(n_2794)
);

AND2x2_ASAP7_75t_L g2795 ( 
.A(n_2745),
.B(n_2137),
.Y(n_2795)
);

A2O1A1Ixp33_ASAP7_75t_L g2796 ( 
.A1(n_2697),
.A2(n_1423),
.B(n_1432),
.C(n_1415),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_SL g2797 ( 
.A(n_2702),
.B(n_2270),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_SL g2798 ( 
.A(n_2710),
.B(n_2347),
.Y(n_2798)
);

BUFx3_ASAP7_75t_L g2799 ( 
.A(n_2740),
.Y(n_2799)
);

BUFx12f_ASAP7_75t_L g2800 ( 
.A(n_2686),
.Y(n_2800)
);

INVx2_ASAP7_75t_L g2801 ( 
.A(n_2688),
.Y(n_2801)
);

INVx2_ASAP7_75t_L g2802 ( 
.A(n_2690),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2712),
.B(n_2139),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2713),
.Y(n_2804)
);

AND2x4_ASAP7_75t_L g2805 ( 
.A(n_2749),
.B(n_2140),
.Y(n_2805)
);

OAI22xp5_ASAP7_75t_L g2806 ( 
.A1(n_2744),
.A2(n_1265),
.B1(n_1267),
.B2(n_1262),
.Y(n_2806)
);

O2A1O1Ixp33_ASAP7_75t_L g2807 ( 
.A1(n_2722),
.A2(n_1461),
.B(n_1482),
.C(n_1435),
.Y(n_2807)
);

AOI21xp5_ASAP7_75t_L g2808 ( 
.A1(n_2731),
.A2(n_1363),
.B(n_1351),
.Y(n_2808)
);

A2O1A1Ixp33_ASAP7_75t_L g2809 ( 
.A1(n_2711),
.A2(n_1487),
.B(n_1495),
.C(n_1483),
.Y(n_2809)
);

CKINVDCx16_ASAP7_75t_R g2810 ( 
.A(n_2727),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2730),
.Y(n_2811)
);

OAI22xp5_ASAP7_75t_L g2812 ( 
.A1(n_2736),
.A2(n_1271),
.B1(n_1272),
.B2(n_1270),
.Y(n_2812)
);

AND2x2_ASAP7_75t_L g2813 ( 
.A(n_2717),
.B(n_2142),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2734),
.Y(n_2814)
);

AOI21x1_ASAP7_75t_L g2815 ( 
.A1(n_2696),
.A2(n_2148),
.B(n_2143),
.Y(n_2815)
);

O2A1O1Ixp5_ASAP7_75t_L g2816 ( 
.A1(n_2726),
.A2(n_1500),
.B(n_1502),
.C(n_1497),
.Y(n_2816)
);

O2A1O1Ixp33_ASAP7_75t_SL g2817 ( 
.A1(n_2715),
.A2(n_1524),
.B(n_1532),
.C(n_1520),
.Y(n_2817)
);

O2A1O1Ixp5_ASAP7_75t_L g2818 ( 
.A1(n_2737),
.A2(n_1541),
.B(n_1549),
.C(n_1537),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2791),
.Y(n_2819)
);

OAI22xp5_ASAP7_75t_L g2820 ( 
.A1(n_2761),
.A2(n_2781),
.B1(n_2789),
.B2(n_2775),
.Y(n_2820)
);

BUFx3_ASAP7_75t_L g2821 ( 
.A(n_2771),
.Y(n_2821)
);

INVx2_ASAP7_75t_SL g2822 ( 
.A(n_2782),
.Y(n_2822)
);

OAI22xp5_ASAP7_75t_L g2823 ( 
.A1(n_2762),
.A2(n_2707),
.B1(n_2739),
.B2(n_2691),
.Y(n_2823)
);

BUFx4f_ASAP7_75t_L g2824 ( 
.A(n_2800),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2792),
.Y(n_2825)
);

BUFx8_ASAP7_75t_L g2826 ( 
.A(n_2767),
.Y(n_2826)
);

BUFx6f_ASAP7_75t_L g2827 ( 
.A(n_2799),
.Y(n_2827)
);

CKINVDCx6p67_ASAP7_75t_R g2828 ( 
.A(n_2810),
.Y(n_2828)
);

BUFx2_ASAP7_75t_SL g2829 ( 
.A(n_2785),
.Y(n_2829)
);

BUFx3_ASAP7_75t_L g2830 ( 
.A(n_2785),
.Y(n_2830)
);

BUFx3_ASAP7_75t_L g2831 ( 
.A(n_2776),
.Y(n_2831)
);

AND2x2_ASAP7_75t_L g2832 ( 
.A(n_2756),
.B(n_2742),
.Y(n_2832)
);

INVxp33_ASAP7_75t_L g2833 ( 
.A(n_2784),
.Y(n_2833)
);

INVx3_ASAP7_75t_SL g2834 ( 
.A(n_2788),
.Y(n_2834)
);

BUFx3_ASAP7_75t_L g2835 ( 
.A(n_2805),
.Y(n_2835)
);

INVx8_ASAP7_75t_L g2836 ( 
.A(n_2805),
.Y(n_2836)
);

INVx2_ASAP7_75t_L g2837 ( 
.A(n_2755),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2758),
.Y(n_2838)
);

BUFx4f_ASAP7_75t_SL g2839 ( 
.A(n_2786),
.Y(n_2839)
);

INVx2_ASAP7_75t_L g2840 ( 
.A(n_2801),
.Y(n_2840)
);

INVx2_ASAP7_75t_L g2841 ( 
.A(n_2802),
.Y(n_2841)
);

BUFx10_ASAP7_75t_L g2842 ( 
.A(n_2804),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2811),
.B(n_2729),
.Y(n_2843)
);

BUFx8_ASAP7_75t_SL g2844 ( 
.A(n_2769),
.Y(n_2844)
);

CKINVDCx5p33_ASAP7_75t_R g2845 ( 
.A(n_2754),
.Y(n_2845)
);

AND2x2_ASAP7_75t_L g2846 ( 
.A(n_2795),
.B(n_2747),
.Y(n_2846)
);

NOR2xp33_ASAP7_75t_L g2847 ( 
.A(n_2780),
.B(n_2814),
.Y(n_2847)
);

INVx5_ASAP7_75t_L g2848 ( 
.A(n_2813),
.Y(n_2848)
);

INVx1_ASAP7_75t_SL g2849 ( 
.A(n_2787),
.Y(n_2849)
);

INVx3_ASAP7_75t_SL g2850 ( 
.A(n_2793),
.Y(n_2850)
);

INVx2_ASAP7_75t_SL g2851 ( 
.A(n_2765),
.Y(n_2851)
);

INVx2_ASAP7_75t_SL g2852 ( 
.A(n_2794),
.Y(n_2852)
);

BUFx3_ASAP7_75t_L g2853 ( 
.A(n_2803),
.Y(n_2853)
);

INVx4_ASAP7_75t_L g2854 ( 
.A(n_2760),
.Y(n_2854)
);

INVx1_ASAP7_75t_SL g2855 ( 
.A(n_2766),
.Y(n_2855)
);

BUFx3_ASAP7_75t_L g2856 ( 
.A(n_2764),
.Y(n_2856)
);

BUFx3_ASAP7_75t_L g2857 ( 
.A(n_2812),
.Y(n_2857)
);

BUFx3_ASAP7_75t_L g2858 ( 
.A(n_2806),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2796),
.Y(n_2859)
);

AND2x4_ASAP7_75t_L g2860 ( 
.A(n_2759),
.B(n_2700),
.Y(n_2860)
);

BUFx2_ASAP7_75t_SL g2861 ( 
.A(n_2797),
.Y(n_2861)
);

BUFx12f_ASAP7_75t_L g2862 ( 
.A(n_2763),
.Y(n_2862)
);

INVx6_ASAP7_75t_SL g2863 ( 
.A(n_2773),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2778),
.Y(n_2864)
);

AND2x2_ASAP7_75t_L g2865 ( 
.A(n_2809),
.B(n_2703),
.Y(n_2865)
);

NOR2x1_ASAP7_75t_L g2866 ( 
.A(n_2757),
.B(n_2718),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2817),
.Y(n_2867)
);

INVx8_ASAP7_75t_L g2868 ( 
.A(n_2783),
.Y(n_2868)
);

INVx4_ASAP7_75t_L g2869 ( 
.A(n_2772),
.Y(n_2869)
);

AND2x4_ASAP7_75t_L g2870 ( 
.A(n_2768),
.B(n_2751),
.Y(n_2870)
);

BUFx3_ASAP7_75t_L g2871 ( 
.A(n_2807),
.Y(n_2871)
);

INVx2_ASAP7_75t_L g2872 ( 
.A(n_2815),
.Y(n_2872)
);

BUFx3_ASAP7_75t_L g2873 ( 
.A(n_2779),
.Y(n_2873)
);

CKINVDCx20_ASAP7_75t_R g2874 ( 
.A(n_2798),
.Y(n_2874)
);

BUFx3_ASAP7_75t_L g2875 ( 
.A(n_2777),
.Y(n_2875)
);

INVx3_ASAP7_75t_L g2876 ( 
.A(n_2818),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2816),
.Y(n_2877)
);

INVx2_ASAP7_75t_SL g2878 ( 
.A(n_2774),
.Y(n_2878)
);

INVx3_ASAP7_75t_L g2879 ( 
.A(n_2770),
.Y(n_2879)
);

INVx2_ASAP7_75t_L g2880 ( 
.A(n_2825),
.Y(n_2880)
);

OR2x6_ASAP7_75t_L g2881 ( 
.A(n_2829),
.B(n_2723),
.Y(n_2881)
);

AOI22xp33_ASAP7_75t_SL g2882 ( 
.A1(n_2868),
.A2(n_1360),
.B1(n_1362),
.B2(n_1182),
.Y(n_2882)
);

AO21x1_ASAP7_75t_L g2883 ( 
.A1(n_2847),
.A2(n_2808),
.B(n_2790),
.Y(n_2883)
);

AND2x2_ASAP7_75t_L g2884 ( 
.A(n_2832),
.B(n_1353),
.Y(n_2884)
);

AOI21xp5_ASAP7_75t_L g2885 ( 
.A1(n_2854),
.A2(n_2743),
.B(n_2701),
.Y(n_2885)
);

OR2x2_ASAP7_75t_L g2886 ( 
.A(n_2855),
.B(n_2153),
.Y(n_2886)
);

OAI22xp5_ASAP7_75t_L g2887 ( 
.A1(n_2874),
.A2(n_2724),
.B1(n_2752),
.B2(n_1120),
.Y(n_2887)
);

OA21x2_ASAP7_75t_L g2888 ( 
.A1(n_2877),
.A2(n_2738),
.B(n_2682),
.Y(n_2888)
);

AND2x2_ASAP7_75t_L g2889 ( 
.A(n_2846),
.B(n_1353),
.Y(n_2889)
);

AOI221xp5_ASAP7_75t_L g2890 ( 
.A1(n_2873),
.A2(n_1123),
.B1(n_1127),
.B2(n_1121),
.C(n_1110),
.Y(n_2890)
);

OAI22xp5_ASAP7_75t_L g2891 ( 
.A1(n_2851),
.A2(n_1129),
.B1(n_1133),
.B2(n_1128),
.Y(n_2891)
);

OA21x2_ASAP7_75t_L g2892 ( 
.A1(n_2872),
.A2(n_2694),
.B(n_2699),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2838),
.Y(n_2893)
);

NOR2xp33_ASAP7_75t_L g2894 ( 
.A(n_2820),
.B(n_1276),
.Y(n_2894)
);

CKINVDCx16_ASAP7_75t_R g2895 ( 
.A(n_2821),
.Y(n_2895)
);

OAI21xp5_ASAP7_75t_L g2896 ( 
.A1(n_2843),
.A2(n_2377),
.B(n_2161),
.Y(n_2896)
);

BUFx2_ASAP7_75t_L g2897 ( 
.A(n_2826),
.Y(n_2897)
);

O2A1O1Ixp33_ASAP7_75t_L g2898 ( 
.A1(n_2823),
.A2(n_1557),
.B(n_1563),
.C(n_1554),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2849),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2819),
.Y(n_2900)
);

AOI22xp33_ASAP7_75t_L g2901 ( 
.A1(n_2871),
.A2(n_1360),
.B1(n_1431),
.B2(n_1362),
.Y(n_2901)
);

OAI21x1_ASAP7_75t_L g2902 ( 
.A1(n_2879),
.A2(n_2701),
.B(n_1572),
.Y(n_2902)
);

AND2x4_ASAP7_75t_L g2903 ( 
.A(n_2830),
.B(n_731),
.Y(n_2903)
);

AND2x4_ASAP7_75t_L g2904 ( 
.A(n_2835),
.B(n_732),
.Y(n_2904)
);

OAI21x1_ASAP7_75t_L g2905 ( 
.A1(n_2876),
.A2(n_1579),
.B(n_1569),
.Y(n_2905)
);

AOI21xp5_ASAP7_75t_L g2906 ( 
.A1(n_2878),
.A2(n_1363),
.B(n_1351),
.Y(n_2906)
);

NAND2xp33_ASAP7_75t_SL g2907 ( 
.A(n_2833),
.B(n_1142),
.Y(n_2907)
);

NAND2x1p5_ASAP7_75t_L g2908 ( 
.A(n_2848),
.B(n_1490),
.Y(n_2908)
);

INVx2_ASAP7_75t_L g2909 ( 
.A(n_2837),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_L g2910 ( 
.A(n_2856),
.B(n_1762),
.Y(n_2910)
);

INVx2_ASAP7_75t_L g2911 ( 
.A(n_2840),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2841),
.Y(n_2912)
);

OAI21x1_ASAP7_75t_L g2913 ( 
.A1(n_2867),
.A2(n_1592),
.B(n_1591),
.Y(n_2913)
);

NAND3xp33_ASAP7_75t_L g2914 ( 
.A(n_2866),
.B(n_1155),
.C(n_1146),
.Y(n_2914)
);

OR2x2_ASAP7_75t_L g2915 ( 
.A(n_2853),
.B(n_1613),
.Y(n_2915)
);

AOI221xp5_ASAP7_75t_L g2916 ( 
.A1(n_2864),
.A2(n_1163),
.B1(n_1164),
.B2(n_1162),
.C(n_1159),
.Y(n_2916)
);

OAI22xp5_ASAP7_75t_L g2917 ( 
.A1(n_2839),
.A2(n_1169),
.B1(n_1171),
.B2(n_1167),
.Y(n_2917)
);

OAI21x1_ASAP7_75t_SL g2918 ( 
.A1(n_2869),
.A2(n_2859),
.B(n_2852),
.Y(n_2918)
);

AO21x2_ASAP7_75t_L g2919 ( 
.A1(n_2870),
.A2(n_1625),
.B(n_1619),
.Y(n_2919)
);

AND2x2_ASAP7_75t_L g2920 ( 
.A(n_2848),
.B(n_1353),
.Y(n_2920)
);

OA21x2_ASAP7_75t_L g2921 ( 
.A1(n_2860),
.A2(n_1631),
.B(n_1627),
.Y(n_2921)
);

CKINVDCx5p33_ASAP7_75t_R g2922 ( 
.A(n_2828),
.Y(n_2922)
);

OAI22xp5_ASAP7_75t_SL g2923 ( 
.A1(n_2834),
.A2(n_1174),
.B1(n_1179),
.B2(n_1173),
.Y(n_2923)
);

NOR3xp33_ASAP7_75t_L g2924 ( 
.A(n_2858),
.B(n_1646),
.C(n_1641),
.Y(n_2924)
);

NOR2xp33_ASAP7_75t_R g2925 ( 
.A(n_2845),
.B(n_1226),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2842),
.Y(n_2926)
);

BUFx12f_ASAP7_75t_L g2927 ( 
.A(n_2827),
.Y(n_2927)
);

AO21x2_ASAP7_75t_L g2928 ( 
.A1(n_2865),
.A2(n_1651),
.B(n_1648),
.Y(n_2928)
);

CKINVDCx12_ASAP7_75t_R g2929 ( 
.A(n_2824),
.Y(n_2929)
);

OAI21x1_ASAP7_75t_L g2930 ( 
.A1(n_2863),
.A2(n_2861),
.B(n_1662),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_L g2931 ( 
.A(n_2850),
.B(n_1755),
.Y(n_2931)
);

BUFx4f_ASAP7_75t_SL g2932 ( 
.A(n_2827),
.Y(n_2932)
);

CKINVDCx5p33_ASAP7_75t_R g2933 ( 
.A(n_2844),
.Y(n_2933)
);

NOR2xp67_ASAP7_75t_SL g2934 ( 
.A(n_2862),
.B(n_1490),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2893),
.Y(n_2935)
);

BUFx2_ASAP7_75t_L g2936 ( 
.A(n_2899),
.Y(n_2936)
);

OR2x2_ASAP7_75t_L g2937 ( 
.A(n_2884),
.B(n_2822),
.Y(n_2937)
);

INVx2_ASAP7_75t_L g2938 ( 
.A(n_2900),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2912),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2880),
.Y(n_2940)
);

INVx2_ASAP7_75t_L g2941 ( 
.A(n_2909),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2911),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2889),
.Y(n_2943)
);

INVx2_ASAP7_75t_L g2944 ( 
.A(n_2918),
.Y(n_2944)
);

AOI22xp33_ASAP7_75t_SL g2945 ( 
.A1(n_2894),
.A2(n_2857),
.B1(n_2875),
.B2(n_2836),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2920),
.Y(n_2946)
);

OA21x2_ASAP7_75t_L g2947 ( 
.A1(n_2885),
.A2(n_2905),
.B(n_2896),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2886),
.Y(n_2948)
);

AND2x2_ASAP7_75t_L g2949 ( 
.A(n_2926),
.B(n_2831),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2921),
.Y(n_2950)
);

AND2x2_ASAP7_75t_L g2951 ( 
.A(n_2928),
.B(n_1610),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2915),
.Y(n_2952)
);

INVx2_ASAP7_75t_L g2953 ( 
.A(n_2888),
.Y(n_2953)
);

OAI21xp5_ASAP7_75t_L g2954 ( 
.A1(n_2914),
.A2(n_1665),
.B(n_1661),
.Y(n_2954)
);

AOI22xp33_ASAP7_75t_L g2955 ( 
.A1(n_2924),
.A2(n_1610),
.B1(n_1644),
.B2(n_1679),
.Y(n_2955)
);

OAI21x1_ASAP7_75t_L g2956 ( 
.A1(n_2906),
.A2(n_1684),
.B(n_1680),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2892),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2919),
.Y(n_2958)
);

AND2x2_ASAP7_75t_L g2959 ( 
.A(n_2895),
.B(n_1610),
.Y(n_2959)
);

AOI22xp33_ASAP7_75t_L g2960 ( 
.A1(n_2882),
.A2(n_1610),
.B1(n_1644),
.B2(n_1685),
.Y(n_2960)
);

BUFx12f_ASAP7_75t_L g2961 ( 
.A(n_2922),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2898),
.Y(n_2962)
);

BUFx6f_ASAP7_75t_L g2963 ( 
.A(n_2927),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2913),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_2881),
.Y(n_2965)
);

AND2x2_ASAP7_75t_L g2966 ( 
.A(n_2930),
.B(n_1610),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_L g2967 ( 
.A(n_2910),
.B(n_1644),
.Y(n_2967)
);

OA21x2_ASAP7_75t_L g2968 ( 
.A1(n_2902),
.A2(n_1693),
.B(n_1686),
.Y(n_2968)
);

INVxp33_ASAP7_75t_L g2969 ( 
.A(n_2931),
.Y(n_2969)
);

BUFx2_ASAP7_75t_L g2970 ( 
.A(n_2908),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_L g2971 ( 
.A(n_2881),
.B(n_1644),
.Y(n_2971)
);

INVx2_ASAP7_75t_SL g2972 ( 
.A(n_2932),
.Y(n_2972)
);

AOI21xp33_ASAP7_75t_L g2973 ( 
.A1(n_2887),
.A2(n_2891),
.B(n_2883),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2904),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2903),
.Y(n_2975)
);

HB1xp67_ASAP7_75t_L g2976 ( 
.A(n_2929),
.Y(n_2976)
);

INVx2_ASAP7_75t_L g2977 ( 
.A(n_2897),
.Y(n_2977)
);

AO21x2_ASAP7_75t_L g2978 ( 
.A1(n_2925),
.A2(n_1711),
.B(n_1706),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2934),
.Y(n_2979)
);

AND2x2_ASAP7_75t_L g2980 ( 
.A(n_2933),
.B(n_1644),
.Y(n_2980)
);

INVx5_ASAP7_75t_L g2981 ( 
.A(n_2907),
.Y(n_2981)
);

NOR2xp33_ASAP7_75t_R g2982 ( 
.A(n_2961),
.B(n_0),
.Y(n_2982)
);

AOI22xp5_ASAP7_75t_L g2983 ( 
.A1(n_2962),
.A2(n_2901),
.B1(n_2923),
.B2(n_2916),
.Y(n_2983)
);

CKINVDCx20_ASAP7_75t_R g2984 ( 
.A(n_2976),
.Y(n_2984)
);

CKINVDCx5p33_ASAP7_75t_R g2985 ( 
.A(n_2972),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2935),
.Y(n_2986)
);

OR2x2_ASAP7_75t_L g2987 ( 
.A(n_2936),
.B(n_1719),
.Y(n_2987)
);

NOR2xp33_ASAP7_75t_R g2988 ( 
.A(n_2963),
.B(n_0),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2938),
.Y(n_2989)
);

NAND2xp33_ASAP7_75t_R g2990 ( 
.A(n_2959),
.B(n_1),
.Y(n_2990)
);

INVx2_ASAP7_75t_L g2991 ( 
.A(n_2939),
.Y(n_2991)
);

AND2x2_ASAP7_75t_L g2992 ( 
.A(n_2977),
.B(n_1720),
.Y(n_2992)
);

INVx3_ASAP7_75t_L g2993 ( 
.A(n_2937),
.Y(n_2993)
);

O2A1O1Ixp33_ASAP7_75t_SL g2994 ( 
.A1(n_2979),
.A2(n_1731),
.B(n_1733),
.C(n_1722),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2940),
.Y(n_2995)
);

AO31x2_ASAP7_75t_L g2996 ( 
.A1(n_2958),
.A2(n_1742),
.A3(n_1737),
.B(n_1275),
.Y(n_2996)
);

AND2x4_ASAP7_75t_L g2997 ( 
.A(n_2965),
.B(n_733),
.Y(n_2997)
);

BUFx6f_ASAP7_75t_L g2998 ( 
.A(n_2963),
.Y(n_2998)
);

CKINVDCx5p33_ASAP7_75t_R g2999 ( 
.A(n_2949),
.Y(n_2999)
);

AND2x2_ASAP7_75t_L g3000 ( 
.A(n_2948),
.B(n_2943),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2942),
.Y(n_3001)
);

INVx5_ASAP7_75t_L g3002 ( 
.A(n_2981),
.Y(n_3002)
);

NOR3xp33_ASAP7_75t_SL g3003 ( 
.A(n_2971),
.B(n_2917),
.C(n_2890),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_L g3004 ( 
.A(n_2952),
.B(n_1250),
.Y(n_3004)
);

AO31x2_ASAP7_75t_L g3005 ( 
.A1(n_2953),
.A2(n_1354),
.A3(n_1364),
.B(n_1335),
.Y(n_3005)
);

NAND2xp33_ASAP7_75t_SL g3006 ( 
.A(n_2969),
.B(n_1183),
.Y(n_3006)
);

INVx2_ASAP7_75t_L g3007 ( 
.A(n_2941),
.Y(n_3007)
);

AND2x2_ASAP7_75t_L g3008 ( 
.A(n_2946),
.B(n_1378),
.Y(n_3008)
);

OAI22xp5_ASAP7_75t_L g3009 ( 
.A1(n_2945),
.A2(n_1185),
.B1(n_1188),
.B2(n_1184),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2957),
.Y(n_3010)
);

CKINVDCx14_ASAP7_75t_R g3011 ( 
.A(n_2980),
.Y(n_3011)
);

AND2x4_ASAP7_75t_L g3012 ( 
.A(n_2944),
.B(n_736),
.Y(n_3012)
);

HB1xp67_ASAP7_75t_L g3013 ( 
.A(n_2950),
.Y(n_3013)
);

HB1xp67_ASAP7_75t_L g3014 ( 
.A(n_2964),
.Y(n_3014)
);

NAND3xp33_ASAP7_75t_SL g3015 ( 
.A(n_2960),
.B(n_1192),
.C(n_1191),
.Y(n_3015)
);

AND2x4_ASAP7_75t_L g3016 ( 
.A(n_2974),
.B(n_2975),
.Y(n_3016)
);

OAI22xp5_ASAP7_75t_L g3017 ( 
.A1(n_2981),
.A2(n_1195),
.B1(n_1202),
.B2(n_1194),
.Y(n_3017)
);

INVx2_ASAP7_75t_L g3018 ( 
.A(n_2951),
.Y(n_3018)
);

NAND2xp33_ASAP7_75t_R g3019 ( 
.A(n_2970),
.B(n_2),
.Y(n_3019)
);

OR2x2_ASAP7_75t_L g3020 ( 
.A(n_2967),
.B(n_1388),
.Y(n_3020)
);

NOR2xp33_ASAP7_75t_R g3021 ( 
.A(n_2966),
.B(n_2),
.Y(n_3021)
);

AND2x2_ASAP7_75t_L g3022 ( 
.A(n_2978),
.B(n_1476),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2973),
.B(n_1523),
.Y(n_3023)
);

AOI22xp33_ASAP7_75t_L g3024 ( 
.A1(n_2955),
.A2(n_1608),
.B1(n_1621),
.B2(n_1573),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2947),
.Y(n_3025)
);

NOR2xp33_ASAP7_75t_L g3026 ( 
.A(n_2954),
.B(n_1673),
.Y(n_3026)
);

OAI22xp5_ASAP7_75t_L g3027 ( 
.A1(n_2968),
.A2(n_1210),
.B1(n_1211),
.B2(n_1209),
.Y(n_3027)
);

INVx2_ASAP7_75t_L g3028 ( 
.A(n_2956),
.Y(n_3028)
);

NOR2xp33_ASAP7_75t_R g3029 ( 
.A(n_2961),
.B(n_3),
.Y(n_3029)
);

AND2x2_ASAP7_75t_L g3030 ( 
.A(n_2936),
.B(n_1723),
.Y(n_3030)
);

AO31x2_ASAP7_75t_L g3031 ( 
.A1(n_2958),
.A2(n_1736),
.A3(n_1449),
.B(n_1491),
.Y(n_3031)
);

OR2x6_ASAP7_75t_L g3032 ( 
.A(n_2961),
.B(n_1490),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2936),
.B(n_1217),
.Y(n_3033)
);

AOI22xp33_ASAP7_75t_L g3034 ( 
.A1(n_2973),
.A2(n_1449),
.B1(n_1491),
.B2(n_1431),
.Y(n_3034)
);

CKINVDCx16_ASAP7_75t_R g3035 ( 
.A(n_2961),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2936),
.B(n_1220),
.Y(n_3036)
);

OR2x2_ASAP7_75t_SL g3037 ( 
.A(n_2977),
.B(n_1660),
.Y(n_3037)
);

OR2x2_ASAP7_75t_L g3038 ( 
.A(n_2936),
.B(n_1660),
.Y(n_3038)
);

INVx2_ASAP7_75t_L g3039 ( 
.A(n_2938),
.Y(n_3039)
);

AND2x2_ASAP7_75t_L g3040 ( 
.A(n_2993),
.B(n_3),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_3010),
.Y(n_3041)
);

AND2x2_ASAP7_75t_L g3042 ( 
.A(n_3011),
.B(n_4),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_3000),
.B(n_1228),
.Y(n_3043)
);

INVxp67_ASAP7_75t_SL g3044 ( 
.A(n_3013),
.Y(n_3044)
);

AND2x4_ASAP7_75t_L g3045 ( 
.A(n_3016),
.B(n_1660),
.Y(n_3045)
);

AND2x2_ASAP7_75t_L g3046 ( 
.A(n_3018),
.B(n_4),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2986),
.Y(n_3047)
);

AO21x2_ASAP7_75t_L g3048 ( 
.A1(n_3025),
.A2(n_3023),
.B(n_3014),
.Y(n_3048)
);

OAI221xp5_ASAP7_75t_L g3049 ( 
.A1(n_3034),
.A2(n_1245),
.B1(n_1246),
.B2(n_1242),
.C(n_1230),
.Y(n_3049)
);

AND2x2_ASAP7_75t_L g3050 ( 
.A(n_3039),
.B(n_6),
.Y(n_3050)
);

AND2x2_ASAP7_75t_L g3051 ( 
.A(n_2989),
.B(n_7),
.Y(n_3051)
);

INVx2_ASAP7_75t_L g3052 ( 
.A(n_2991),
.Y(n_3052)
);

INVx2_ASAP7_75t_L g3053 ( 
.A(n_3007),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2995),
.Y(n_3054)
);

BUFx2_ASAP7_75t_L g3055 ( 
.A(n_3038),
.Y(n_3055)
);

AND2x2_ASAP7_75t_L g3056 ( 
.A(n_3001),
.B(n_8),
.Y(n_3056)
);

OAI22xp33_ASAP7_75t_L g3057 ( 
.A1(n_3002),
.A2(n_1248),
.B1(n_1254),
.B2(n_1247),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_3008),
.Y(n_3058)
);

INVx2_ASAP7_75t_L g3059 ( 
.A(n_2987),
.Y(n_3059)
);

AND2x2_ASAP7_75t_L g3060 ( 
.A(n_2999),
.B(n_8),
.Y(n_3060)
);

OR2x2_ASAP7_75t_L g3061 ( 
.A(n_3030),
.B(n_9),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_3004),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2996),
.Y(n_3063)
);

INVx2_ASAP7_75t_L g3064 ( 
.A(n_3005),
.Y(n_3064)
);

OR2x2_ASAP7_75t_L g3065 ( 
.A(n_3020),
.B(n_9),
.Y(n_3065)
);

AND2x2_ASAP7_75t_L g3066 ( 
.A(n_3002),
.B(n_10),
.Y(n_3066)
);

INVx2_ASAP7_75t_L g3067 ( 
.A(n_3005),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2996),
.Y(n_3068)
);

INVx3_ASAP7_75t_L g3069 ( 
.A(n_2998),
.Y(n_3069)
);

INVx3_ASAP7_75t_L g3070 ( 
.A(n_2998),
.Y(n_3070)
);

OR2x2_ASAP7_75t_L g3071 ( 
.A(n_3033),
.B(n_10),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_3031),
.Y(n_3072)
);

AND2x2_ASAP7_75t_L g3073 ( 
.A(n_3035),
.B(n_11),
.Y(n_3073)
);

AND2x2_ASAP7_75t_L g3074 ( 
.A(n_2984),
.B(n_11),
.Y(n_3074)
);

BUFx3_ASAP7_75t_L g3075 ( 
.A(n_2985),
.Y(n_3075)
);

OAI21x1_ASAP7_75t_L g3076 ( 
.A1(n_3028),
.A2(n_12),
.B(n_13),
.Y(n_3076)
);

INVx2_ASAP7_75t_L g3077 ( 
.A(n_2992),
.Y(n_3077)
);

OAI21x1_ASAP7_75t_L g3078 ( 
.A1(n_3027),
.A2(n_13),
.B(n_14),
.Y(n_3078)
);

INVx2_ASAP7_75t_L g3079 ( 
.A(n_3031),
.Y(n_3079)
);

AND2x2_ASAP7_75t_L g3080 ( 
.A(n_3021),
.B(n_14),
.Y(n_3080)
);

INVx2_ASAP7_75t_SL g3081 ( 
.A(n_3036),
.Y(n_3081)
);

HB1xp67_ASAP7_75t_L g3082 ( 
.A(n_3022),
.Y(n_3082)
);

INVxp67_ASAP7_75t_SL g3083 ( 
.A(n_3019),
.Y(n_3083)
);

HB1xp67_ASAP7_75t_L g3084 ( 
.A(n_3037),
.Y(n_3084)
);

BUFx2_ASAP7_75t_L g3085 ( 
.A(n_3032),
.Y(n_3085)
);

AND2x2_ASAP7_75t_L g3086 ( 
.A(n_2997),
.B(n_15),
.Y(n_3086)
);

AND2x2_ASAP7_75t_L g3087 ( 
.A(n_3012),
.B(n_16),
.Y(n_3087)
);

AND2x2_ASAP7_75t_L g3088 ( 
.A(n_2982),
.B(n_17),
.Y(n_3088)
);

OR2x2_ASAP7_75t_L g3089 ( 
.A(n_2983),
.B(n_3006),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2994),
.Y(n_3090)
);

INVxp67_ASAP7_75t_SL g3091 ( 
.A(n_2990),
.Y(n_3091)
);

BUFx3_ASAP7_75t_L g3092 ( 
.A(n_3029),
.Y(n_3092)
);

OAI221xp5_ASAP7_75t_L g3093 ( 
.A1(n_3026),
.A2(n_3003),
.B1(n_3009),
.B2(n_3017),
.C(n_3024),
.Y(n_3093)
);

NOR2xp33_ASAP7_75t_L g3094 ( 
.A(n_3015),
.B(n_1260),
.Y(n_3094)
);

OAI21x1_ASAP7_75t_L g3095 ( 
.A1(n_2988),
.A2(n_19),
.B(n_20),
.Y(n_3095)
);

AND2x2_ASAP7_75t_L g3096 ( 
.A(n_2993),
.B(n_19),
.Y(n_3096)
);

INVx2_ASAP7_75t_L g3097 ( 
.A(n_3041),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_3047),
.Y(n_3098)
);

NOR2xp33_ASAP7_75t_L g3099 ( 
.A(n_3089),
.B(n_3062),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_3054),
.Y(n_3100)
);

AOI221x1_ASAP7_75t_L g3101 ( 
.A1(n_3066),
.A2(n_1734),
.B1(n_1764),
.B2(n_1675),
.C(n_1507),
.Y(n_3101)
);

HB1xp67_ASAP7_75t_L g3102 ( 
.A(n_3082),
.Y(n_3102)
);

NAND3xp33_ASAP7_75t_L g3103 ( 
.A(n_3072),
.B(n_1264),
.C(n_1261),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_3052),
.Y(n_3104)
);

OAI21x1_ASAP7_75t_L g3105 ( 
.A1(n_3079),
.A2(n_20),
.B(n_22),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_3055),
.B(n_3059),
.Y(n_3106)
);

INVx3_ASAP7_75t_L g3107 ( 
.A(n_3075),
.Y(n_3107)
);

HB1xp67_ASAP7_75t_L g3108 ( 
.A(n_3048),
.Y(n_3108)
);

OA21x2_ASAP7_75t_L g3109 ( 
.A1(n_3083),
.A2(n_1273),
.B(n_1268),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_3055),
.B(n_1274),
.Y(n_3110)
);

HB1xp67_ASAP7_75t_L g3111 ( 
.A(n_3044),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_3053),
.Y(n_3112)
);

OA21x2_ASAP7_75t_L g3113 ( 
.A1(n_3091),
.A2(n_1281),
.B(n_1278),
.Y(n_3113)
);

BUFx3_ASAP7_75t_L g3114 ( 
.A(n_3069),
.Y(n_3114)
);

OA21x2_ASAP7_75t_L g3115 ( 
.A1(n_3063),
.A2(n_1286),
.B(n_1283),
.Y(n_3115)
);

AND2x2_ASAP7_75t_L g3116 ( 
.A(n_3077),
.B(n_23),
.Y(n_3116)
);

AOI22xp33_ASAP7_75t_L g3117 ( 
.A1(n_3093),
.A2(n_1675),
.B1(n_1734),
.B2(n_1507),
.Y(n_3117)
);

HB1xp67_ASAP7_75t_L g3118 ( 
.A(n_3058),
.Y(n_3118)
);

HB1xp67_ASAP7_75t_L g3119 ( 
.A(n_3068),
.Y(n_3119)
);

OAI21xp33_ASAP7_75t_L g3120 ( 
.A1(n_3094),
.A2(n_1294),
.B(n_1288),
.Y(n_3120)
);

INVx2_ASAP7_75t_L g3121 ( 
.A(n_3045),
.Y(n_3121)
);

HB1xp67_ASAP7_75t_L g3122 ( 
.A(n_3056),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_3051),
.Y(n_3123)
);

AOI21xp5_ASAP7_75t_L g3124 ( 
.A1(n_3090),
.A2(n_1367),
.B(n_1318),
.Y(n_3124)
);

AOI21xp5_ASAP7_75t_L g3125 ( 
.A1(n_3081),
.A2(n_1369),
.B(n_1319),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_3050),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_3064),
.Y(n_3127)
);

HB1xp67_ASAP7_75t_L g3128 ( 
.A(n_3040),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_3067),
.Y(n_3129)
);

NAND4xp25_ASAP7_75t_L g3130 ( 
.A(n_3080),
.B(n_3071),
.C(n_3049),
.D(n_3061),
.Y(n_3130)
);

INVx3_ASAP7_75t_L g3131 ( 
.A(n_3070),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_3046),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_3096),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_3084),
.Y(n_3134)
);

OA21x2_ASAP7_75t_L g3135 ( 
.A1(n_3043),
.A2(n_1317),
.B(n_1307),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_3065),
.B(n_1320),
.Y(n_3136)
);

AOI22xp33_ASAP7_75t_L g3137 ( 
.A1(n_3073),
.A2(n_1764),
.B1(n_1323),
.B2(n_1326),
.Y(n_3137)
);

BUFx3_ASAP7_75t_L g3138 ( 
.A(n_3092),
.Y(n_3138)
);

INVx2_ASAP7_75t_L g3139 ( 
.A(n_3085),
.Y(n_3139)
);

INVxp67_ASAP7_75t_SL g3140 ( 
.A(n_3085),
.Y(n_3140)
);

INVx2_ASAP7_75t_L g3141 ( 
.A(n_3076),
.Y(n_3141)
);

OAI21x1_ASAP7_75t_L g3142 ( 
.A1(n_3078),
.A2(n_23),
.B(n_24),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_3087),
.Y(n_3143)
);

AND2x2_ASAP7_75t_L g3144 ( 
.A(n_3042),
.B(n_24),
.Y(n_3144)
);

AOI21xp5_ASAP7_75t_L g3145 ( 
.A1(n_3057),
.A2(n_1436),
.B(n_1387),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_SL g3146 ( 
.A(n_3088),
.B(n_1322),
.Y(n_3146)
);

INVx2_ASAP7_75t_L g3147 ( 
.A(n_3060),
.Y(n_3147)
);

AOI22xp33_ASAP7_75t_SL g3148 ( 
.A1(n_3074),
.A2(n_1339),
.B1(n_1348),
.B2(n_1328),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_3095),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_3086),
.Y(n_3150)
);

AOI22xp5_ASAP7_75t_L g3151 ( 
.A1(n_3083),
.A2(n_1365),
.B1(n_1366),
.B2(n_1361),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_3041),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_3041),
.Y(n_3153)
);

HB1xp67_ASAP7_75t_L g3154 ( 
.A(n_3082),
.Y(n_3154)
);

INVx3_ASAP7_75t_L g3155 ( 
.A(n_3075),
.Y(n_3155)
);

INVx4_ASAP7_75t_SL g3156 ( 
.A(n_3092),
.Y(n_3156)
);

INVx2_ASAP7_75t_L g3157 ( 
.A(n_3041),
.Y(n_3157)
);

AND2x2_ASAP7_75t_L g3158 ( 
.A(n_3055),
.B(n_25),
.Y(n_3158)
);

AOI222xp33_ASAP7_75t_L g3159 ( 
.A1(n_3091),
.A2(n_1391),
.B1(n_1381),
.B2(n_1395),
.C1(n_1390),
.C2(n_1368),
.Y(n_3159)
);

INVx2_ASAP7_75t_L g3160 ( 
.A(n_3041),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_3041),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_3041),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_L g3163 ( 
.A(n_3082),
.B(n_1399),
.Y(n_3163)
);

OAI22xp33_ASAP7_75t_L g3164 ( 
.A1(n_3083),
.A2(n_1407),
.B1(n_1409),
.B2(n_1402),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_3082),
.B(n_1414),
.Y(n_3165)
);

INVx3_ASAP7_75t_L g3166 ( 
.A(n_3075),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_3041),
.Y(n_3167)
);

NAND3xp33_ASAP7_75t_L g3168 ( 
.A(n_3072),
.B(n_1421),
.C(n_1419),
.Y(n_3168)
);

AOI21xp5_ASAP7_75t_L g3169 ( 
.A1(n_3093),
.A2(n_1445),
.B(n_1424),
.Y(n_3169)
);

INVx2_ASAP7_75t_L g3170 ( 
.A(n_3041),
.Y(n_3170)
);

INVx4_ASAP7_75t_R g3171 ( 
.A(n_3075),
.Y(n_3171)
);

NAND4xp25_ASAP7_75t_L g3172 ( 
.A(n_3093),
.B(n_28),
.C(n_26),
.D(n_27),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_3041),
.Y(n_3173)
);

AOI22xp33_ASAP7_75t_L g3174 ( 
.A1(n_3089),
.A2(n_1425),
.B1(n_1437),
.B2(n_1422),
.Y(n_3174)
);

INVx2_ASAP7_75t_L g3175 ( 
.A(n_3041),
.Y(n_3175)
);

OR2x2_ASAP7_75t_L g3176 ( 
.A(n_3082),
.B(n_28),
.Y(n_3176)
);

OAI21x1_ASAP7_75t_L g3177 ( 
.A1(n_3079),
.A2(n_29),
.B(n_30),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_3041),
.Y(n_3178)
);

OAI22xp33_ASAP7_75t_L g3179 ( 
.A1(n_3083),
.A2(n_1439),
.B1(n_1442),
.B2(n_1438),
.Y(n_3179)
);

INVx2_ASAP7_75t_L g3180 ( 
.A(n_3041),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_L g3181 ( 
.A(n_3082),
.B(n_1446),
.Y(n_3181)
);

BUFx3_ASAP7_75t_L g3182 ( 
.A(n_3075),
.Y(n_3182)
);

AO21x2_ASAP7_75t_L g3183 ( 
.A1(n_3072),
.A2(n_29),
.B(n_31),
.Y(n_3183)
);

AOI22xp33_ASAP7_75t_SL g3184 ( 
.A1(n_3083),
.A2(n_1453),
.B1(n_1454),
.B2(n_1452),
.Y(n_3184)
);

HB1xp67_ASAP7_75t_L g3185 ( 
.A(n_3082),
.Y(n_3185)
);

AO31x2_ASAP7_75t_L g3186 ( 
.A1(n_3079),
.A2(n_35),
.A3(n_33),
.B(n_34),
.Y(n_3186)
);

AO21x2_ASAP7_75t_L g3187 ( 
.A1(n_3072),
.A2(n_34),
.B(n_35),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_3041),
.Y(n_3188)
);

OAI221xp5_ASAP7_75t_L g3189 ( 
.A1(n_3083),
.A2(n_1468),
.B1(n_1469),
.B2(n_1465),
.C(n_1456),
.Y(n_3189)
);

OAI211xp5_ASAP7_75t_L g3190 ( 
.A1(n_3091),
.A2(n_1471),
.B(n_1481),
.C(n_1470),
.Y(n_3190)
);

INVx2_ASAP7_75t_L g3191 ( 
.A(n_3041),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_3041),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_3041),
.Y(n_3193)
);

OAI21xp5_ASAP7_75t_L g3194 ( 
.A1(n_3091),
.A2(n_1492),
.B(n_1488),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_3082),
.B(n_1493),
.Y(n_3195)
);

INVxp67_ASAP7_75t_SL g3196 ( 
.A(n_3082),
.Y(n_3196)
);

OAI21xp5_ASAP7_75t_L g3197 ( 
.A1(n_3091),
.A2(n_1498),
.B(n_1494),
.Y(n_3197)
);

HB1xp67_ASAP7_75t_L g3198 ( 
.A(n_3082),
.Y(n_3198)
);

AOI21xp5_ASAP7_75t_L g3199 ( 
.A1(n_3093),
.A2(n_1529),
.B(n_1499),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_3041),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_3041),
.Y(n_3201)
);

INVx2_ASAP7_75t_SL g3202 ( 
.A(n_3075),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_3082),
.B(n_1505),
.Y(n_3203)
);

AND2x2_ASAP7_75t_L g3204 ( 
.A(n_3055),
.B(n_37),
.Y(n_3204)
);

AOI21xp5_ASAP7_75t_L g3205 ( 
.A1(n_3093),
.A2(n_1535),
.B(n_1517),
.Y(n_3205)
);

OAI21xp33_ASAP7_75t_SL g3206 ( 
.A1(n_3083),
.A2(n_37),
.B(n_38),
.Y(n_3206)
);

NOR2xp33_ASAP7_75t_L g3207 ( 
.A(n_3089),
.B(n_1506),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_3098),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_3100),
.Y(n_3209)
);

AND2x2_ASAP7_75t_L g3210 ( 
.A(n_3139),
.B(n_38),
.Y(n_3210)
);

INVxp67_ASAP7_75t_SL g3211 ( 
.A(n_3108),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_3152),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_L g3213 ( 
.A(n_3099),
.B(n_1509),
.Y(n_3213)
);

AND2x2_ASAP7_75t_L g3214 ( 
.A(n_3140),
.B(n_39),
.Y(n_3214)
);

BUFx2_ASAP7_75t_L g3215 ( 
.A(n_3111),
.Y(n_3215)
);

OAI22xp5_ASAP7_75t_L g3216 ( 
.A1(n_3134),
.A2(n_1513),
.B1(n_1515),
.B2(n_1512),
.Y(n_3216)
);

AND2x2_ASAP7_75t_L g3217 ( 
.A(n_3122),
.B(n_39),
.Y(n_3217)
);

OR2x2_ASAP7_75t_L g3218 ( 
.A(n_3106),
.B(n_3102),
.Y(n_3218)
);

AOI221xp5_ASAP7_75t_L g3219 ( 
.A1(n_3172),
.A2(n_3117),
.B1(n_3205),
.B2(n_3199),
.C(n_3169),
.Y(n_3219)
);

INVx2_ASAP7_75t_L g3220 ( 
.A(n_3097),
.Y(n_3220)
);

AND2x2_ASAP7_75t_L g3221 ( 
.A(n_3128),
.B(n_40),
.Y(n_3221)
);

AND2x2_ASAP7_75t_L g3222 ( 
.A(n_3131),
.B(n_42),
.Y(n_3222)
);

AND2x2_ASAP7_75t_L g3223 ( 
.A(n_3149),
.B(n_42),
.Y(n_3223)
);

INVx2_ASAP7_75t_SL g3224 ( 
.A(n_3171),
.Y(n_3224)
);

OR2x2_ASAP7_75t_L g3225 ( 
.A(n_3154),
.B(n_43),
.Y(n_3225)
);

OAI321xp33_ASAP7_75t_L g3226 ( 
.A1(n_3194),
.A2(n_45),
.A3(n_47),
.B1(n_43),
.B2(n_44),
.C(n_46),
.Y(n_3226)
);

OR2x2_ASAP7_75t_L g3227 ( 
.A(n_3185),
.B(n_45),
.Y(n_3227)
);

OAI221xp5_ASAP7_75t_L g3228 ( 
.A1(n_3206),
.A2(n_1774),
.B1(n_1776),
.B2(n_1770),
.C(n_1767),
.Y(n_3228)
);

NOR2xp33_ASAP7_75t_L g3229 ( 
.A(n_3207),
.B(n_1526),
.Y(n_3229)
);

OAI31xp33_ASAP7_75t_SL g3230 ( 
.A1(n_3197),
.A2(n_49),
.A3(n_46),
.B(n_47),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_3157),
.Y(n_3231)
);

NAND2xp5_ASAP7_75t_L g3232 ( 
.A(n_3118),
.B(n_3141),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_3153),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_L g3234 ( 
.A(n_3196),
.B(n_1528),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_3161),
.Y(n_3235)
);

INVx3_ASAP7_75t_L g3236 ( 
.A(n_3138),
.Y(n_3236)
);

AO21x2_ASAP7_75t_L g3237 ( 
.A1(n_3110),
.A2(n_49),
.B(n_50),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_3198),
.B(n_3126),
.Y(n_3238)
);

BUFx3_ASAP7_75t_L g3239 ( 
.A(n_3182),
.Y(n_3239)
);

INVx1_ASAP7_75t_SL g3240 ( 
.A(n_3156),
.Y(n_3240)
);

INVx3_ASAP7_75t_L g3241 ( 
.A(n_3114),
.Y(n_3241)
);

AND2x2_ASAP7_75t_L g3242 ( 
.A(n_3121),
.B(n_3147),
.Y(n_3242)
);

INVx3_ASAP7_75t_L g3243 ( 
.A(n_3107),
.Y(n_3243)
);

INVx2_ASAP7_75t_L g3244 ( 
.A(n_3160),
.Y(n_3244)
);

AOI22xp33_ASAP7_75t_L g3245 ( 
.A1(n_3115),
.A2(n_1533),
.B1(n_1536),
.B2(n_1531),
.Y(n_3245)
);

HB1xp67_ASAP7_75t_L g3246 ( 
.A(n_3119),
.Y(n_3246)
);

BUFx3_ASAP7_75t_L g3247 ( 
.A(n_3155),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_3162),
.Y(n_3248)
);

AND2x2_ASAP7_75t_L g3249 ( 
.A(n_3133),
.B(n_50),
.Y(n_3249)
);

AND2x4_ASAP7_75t_L g3250 ( 
.A(n_3166),
.B(n_51),
.Y(n_3250)
);

BUFx3_ASAP7_75t_L g3251 ( 
.A(n_3202),
.Y(n_3251)
);

AND2x2_ASAP7_75t_L g3252 ( 
.A(n_3123),
.B(n_51),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_3173),
.Y(n_3253)
);

INVxp67_ASAP7_75t_SL g3254 ( 
.A(n_3113),
.Y(n_3254)
);

OAI221xp5_ASAP7_75t_L g3255 ( 
.A1(n_3184),
.A2(n_1766),
.B1(n_1763),
.B2(n_1760),
.C(n_1546),
.Y(n_3255)
);

INVx2_ASAP7_75t_SL g3256 ( 
.A(n_3156),
.Y(n_3256)
);

BUFx3_ASAP7_75t_L g3257 ( 
.A(n_3144),
.Y(n_3257)
);

AND2x2_ASAP7_75t_L g3258 ( 
.A(n_3143),
.B(n_54),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_3167),
.Y(n_3259)
);

OAI31xp33_ASAP7_75t_L g3260 ( 
.A1(n_3190),
.A2(n_56),
.A3(n_54),
.B(n_55),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_L g3261 ( 
.A(n_3204),
.B(n_1538),
.Y(n_3261)
);

AOI221xp5_ASAP7_75t_L g3262 ( 
.A1(n_3164),
.A2(n_1551),
.B1(n_1553),
.B2(n_1550),
.C(n_1542),
.Y(n_3262)
);

AND2x2_ASAP7_75t_L g3263 ( 
.A(n_3150),
.B(n_55),
.Y(n_3263)
);

AND2x4_ASAP7_75t_L g3264 ( 
.A(n_3132),
.B(n_56),
.Y(n_3264)
);

AOI22xp33_ASAP7_75t_L g3265 ( 
.A1(n_3103),
.A2(n_1560),
.B1(n_1562),
.B2(n_1558),
.Y(n_3265)
);

AND2x2_ASAP7_75t_SL g3266 ( 
.A(n_3109),
.B(n_57),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_3178),
.Y(n_3267)
);

INVx3_ASAP7_75t_L g3268 ( 
.A(n_3170),
.Y(n_3268)
);

AND2x2_ASAP7_75t_L g3269 ( 
.A(n_3175),
.B(n_57),
.Y(n_3269)
);

OR2x2_ASAP7_75t_L g3270 ( 
.A(n_3104),
.B(n_59),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_3188),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_3193),
.Y(n_3272)
);

BUFx3_ASAP7_75t_L g3273 ( 
.A(n_3116),
.Y(n_3273)
);

AND2x4_ASAP7_75t_L g3274 ( 
.A(n_3200),
.B(n_60),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_SL g3275 ( 
.A(n_3163),
.B(n_1564),
.Y(n_3275)
);

HB1xp67_ASAP7_75t_L g3276 ( 
.A(n_3180),
.Y(n_3276)
);

HB1xp67_ASAP7_75t_L g3277 ( 
.A(n_3191),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_3201),
.Y(n_3278)
);

AOI221x1_ASAP7_75t_L g3279 ( 
.A1(n_3130),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.C(n_65),
.Y(n_3279)
);

INVx2_ASAP7_75t_L g3280 ( 
.A(n_3192),
.Y(n_3280)
);

AOI31xp33_ASAP7_75t_L g3281 ( 
.A1(n_3159),
.A2(n_1568),
.A3(n_1570),
.B(n_1567),
.Y(n_3281)
);

OR2x2_ASAP7_75t_L g3282 ( 
.A(n_3112),
.B(n_63),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_L g3283 ( 
.A(n_3158),
.B(n_1574),
.Y(n_3283)
);

HB1xp67_ASAP7_75t_L g3284 ( 
.A(n_3127),
.Y(n_3284)
);

AND2x4_ASAP7_75t_L g3285 ( 
.A(n_3176),
.B(n_64),
.Y(n_3285)
);

NAND3xp33_ASAP7_75t_L g3286 ( 
.A(n_3101),
.B(n_1581),
.C(n_1575),
.Y(n_3286)
);

OAI221xp5_ASAP7_75t_SL g3287 ( 
.A1(n_3174),
.A2(n_1597),
.B1(n_1600),
.B2(n_1587),
.C(n_1583),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_3129),
.Y(n_3288)
);

AND2x4_ASAP7_75t_L g3289 ( 
.A(n_3142),
.B(n_65),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_3186),
.Y(n_3290)
);

AOI22xp5_ASAP7_75t_L g3291 ( 
.A1(n_3168),
.A2(n_3183),
.B1(n_3187),
.B2(n_3135),
.Y(n_3291)
);

OAI22xp5_ASAP7_75t_L g3292 ( 
.A1(n_3165),
.A2(n_1605),
.B1(n_1607),
.B2(n_1603),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_3186),
.Y(n_3293)
);

HB1xp67_ASAP7_75t_L g3294 ( 
.A(n_3181),
.Y(n_3294)
);

INVx2_ASAP7_75t_L g3295 ( 
.A(n_3105),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_L g3296 ( 
.A(n_3195),
.B(n_1609),
.Y(n_3296)
);

INVx2_ASAP7_75t_L g3297 ( 
.A(n_3177),
.Y(n_3297)
);

INVx2_ASAP7_75t_L g3298 ( 
.A(n_3203),
.Y(n_3298)
);

AND2x2_ASAP7_75t_SL g3299 ( 
.A(n_3137),
.B(n_3151),
.Y(n_3299)
);

AND2x2_ASAP7_75t_L g3300 ( 
.A(n_3136),
.B(n_3146),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_3189),
.Y(n_3301)
);

INVx2_ASAP7_75t_L g3302 ( 
.A(n_3179),
.Y(n_3302)
);

AND2x2_ASAP7_75t_L g3303 ( 
.A(n_3148),
.B(n_66),
.Y(n_3303)
);

BUFx3_ASAP7_75t_L g3304 ( 
.A(n_3125),
.Y(n_3304)
);

AND2x2_ASAP7_75t_L g3305 ( 
.A(n_3124),
.B(n_66),
.Y(n_3305)
);

INVx2_ASAP7_75t_L g3306 ( 
.A(n_3120),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_3145),
.Y(n_3307)
);

NOR2xp33_ASAP7_75t_L g3308 ( 
.A(n_3207),
.B(n_1611),
.Y(n_3308)
);

INVx2_ASAP7_75t_L g3309 ( 
.A(n_3139),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_3098),
.Y(n_3310)
);

HB1xp67_ASAP7_75t_L g3311 ( 
.A(n_3111),
.Y(n_3311)
);

AND2x2_ASAP7_75t_L g3312 ( 
.A(n_3139),
.B(n_67),
.Y(n_3312)
);

AO21x2_ASAP7_75t_L g3313 ( 
.A1(n_3108),
.A2(n_68),
.B(n_69),
.Y(n_3313)
);

AOI33xp33_ASAP7_75t_L g3314 ( 
.A1(n_3117),
.A2(n_1633),
.A3(n_1628),
.B1(n_1634),
.B2(n_1630),
.B3(n_1624),
.Y(n_3314)
);

AOI22xp5_ASAP7_75t_L g3315 ( 
.A1(n_3172),
.A2(n_1636),
.B1(n_1639),
.B2(n_1635),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_3098),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_L g3317 ( 
.A(n_3099),
.B(n_1642),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3098),
.Y(n_3318)
);

INVx2_ASAP7_75t_L g3319 ( 
.A(n_3139),
.Y(n_3319)
);

OR2x2_ASAP7_75t_L g3320 ( 
.A(n_3106),
.B(n_68),
.Y(n_3320)
);

INVx4_ASAP7_75t_L g3321 ( 
.A(n_3156),
.Y(n_3321)
);

NAND4xp25_ASAP7_75t_SL g3322 ( 
.A(n_3101),
.B(n_72),
.C(n_69),
.D(n_70),
.Y(n_3322)
);

INVx2_ASAP7_75t_SL g3323 ( 
.A(n_3171),
.Y(n_3323)
);

INVx2_ASAP7_75t_L g3324 ( 
.A(n_3139),
.Y(n_3324)
);

AND2x2_ASAP7_75t_L g3325 ( 
.A(n_3139),
.B(n_72),
.Y(n_3325)
);

AND2x2_ASAP7_75t_L g3326 ( 
.A(n_3139),
.B(n_73),
.Y(n_3326)
);

AO22x1_ASAP7_75t_L g3327 ( 
.A1(n_3140),
.A2(n_1652),
.B1(n_1657),
.B2(n_1650),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_3099),
.B(n_1664),
.Y(n_3328)
);

HB1xp67_ASAP7_75t_L g3329 ( 
.A(n_3111),
.Y(n_3329)
);

NAND3xp33_ASAP7_75t_L g3330 ( 
.A(n_3172),
.B(n_1681),
.C(n_1672),
.Y(n_3330)
);

INVx3_ASAP7_75t_L g3331 ( 
.A(n_3138),
.Y(n_3331)
);

BUFx3_ASAP7_75t_L g3332 ( 
.A(n_3182),
.Y(n_3332)
);

AND2x4_ASAP7_75t_L g3333 ( 
.A(n_3140),
.B(n_73),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3098),
.Y(n_3334)
);

HB1xp67_ASAP7_75t_L g3335 ( 
.A(n_3111),
.Y(n_3335)
);

AOI221xp5_ASAP7_75t_L g3336 ( 
.A1(n_3172),
.A2(n_1692),
.B1(n_1694),
.B2(n_1690),
.C(n_1682),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_L g3337 ( 
.A(n_3099),
.B(n_1697),
.Y(n_3337)
);

AND2x2_ASAP7_75t_L g3338 ( 
.A(n_3139),
.B(n_74),
.Y(n_3338)
);

OAI22xp5_ASAP7_75t_L g3339 ( 
.A1(n_3140),
.A2(n_1700),
.B1(n_1702),
.B2(n_1699),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_3098),
.Y(n_3340)
);

AND2x2_ASAP7_75t_L g3341 ( 
.A(n_3139),
.B(n_75),
.Y(n_3341)
);

OR2x2_ASAP7_75t_L g3342 ( 
.A(n_3106),
.B(n_75),
.Y(n_3342)
);

AND2x2_ASAP7_75t_L g3343 ( 
.A(n_3139),
.B(n_76),
.Y(n_3343)
);

AND2x4_ASAP7_75t_L g3344 ( 
.A(n_3140),
.B(n_76),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_3098),
.Y(n_3345)
);

OAI22xp5_ASAP7_75t_L g3346 ( 
.A1(n_3140),
.A2(n_1705),
.B1(n_1707),
.B2(n_1703),
.Y(n_3346)
);

INVx1_ASAP7_75t_SL g3347 ( 
.A(n_3156),
.Y(n_3347)
);

AND2x2_ASAP7_75t_L g3348 ( 
.A(n_3139),
.B(n_77),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_3098),
.Y(n_3349)
);

INVx4_ASAP7_75t_SL g3350 ( 
.A(n_3186),
.Y(n_3350)
);

AND2x2_ASAP7_75t_L g3351 ( 
.A(n_3139),
.B(n_77),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3098),
.Y(n_3352)
);

NOR3xp33_ASAP7_75t_SL g3353 ( 
.A(n_3206),
.B(n_1716),
.C(n_1713),
.Y(n_3353)
);

INVx2_ASAP7_75t_L g3354 ( 
.A(n_3139),
.Y(n_3354)
);

NAND3xp33_ASAP7_75t_L g3355 ( 
.A(n_3172),
.B(n_1724),
.C(n_1718),
.Y(n_3355)
);

AND2x2_ASAP7_75t_L g3356 ( 
.A(n_3139),
.B(n_78),
.Y(n_3356)
);

INVx2_ASAP7_75t_L g3357 ( 
.A(n_3139),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_3098),
.Y(n_3358)
);

OR2x2_ASAP7_75t_L g3359 ( 
.A(n_3106),
.B(n_80),
.Y(n_3359)
);

HB1xp67_ASAP7_75t_L g3360 ( 
.A(n_3111),
.Y(n_3360)
);

HB1xp67_ASAP7_75t_L g3361 ( 
.A(n_3111),
.Y(n_3361)
);

BUFx2_ASAP7_75t_L g3362 ( 
.A(n_3140),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_L g3363 ( 
.A(n_3294),
.B(n_1738),
.Y(n_3363)
);

INVxp67_ASAP7_75t_SL g3364 ( 
.A(n_3362),
.Y(n_3364)
);

AND2x2_ASAP7_75t_L g3365 ( 
.A(n_3243),
.B(n_80),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_L g3366 ( 
.A(n_3242),
.B(n_1739),
.Y(n_3366)
);

INVx2_ASAP7_75t_L g3367 ( 
.A(n_3256),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_3208),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_3298),
.B(n_1740),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_3209),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_3295),
.B(n_1745),
.Y(n_3371)
);

INVx2_ASAP7_75t_L g3372 ( 
.A(n_3240),
.Y(n_3372)
);

OR2x2_ASAP7_75t_L g3373 ( 
.A(n_3218),
.B(n_81),
.Y(n_3373)
);

AND2x2_ASAP7_75t_L g3374 ( 
.A(n_3224),
.B(n_81),
.Y(n_3374)
);

INVx2_ASAP7_75t_L g3375 ( 
.A(n_3347),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_3212),
.Y(n_3376)
);

OAI321xp33_ASAP7_75t_L g3377 ( 
.A1(n_3315),
.A2(n_84),
.A3(n_86),
.B1(n_82),
.B2(n_83),
.C(n_85),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_L g3378 ( 
.A(n_3297),
.B(n_1746),
.Y(n_3378)
);

NOR2xp33_ASAP7_75t_L g3379 ( 
.A(n_3321),
.B(n_1747),
.Y(n_3379)
);

INVx3_ASAP7_75t_L g3380 ( 
.A(n_3251),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_3233),
.Y(n_3381)
);

INVx4_ASAP7_75t_L g3382 ( 
.A(n_3250),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_3235),
.Y(n_3383)
);

AND2x2_ASAP7_75t_L g3384 ( 
.A(n_3323),
.B(n_82),
.Y(n_3384)
);

AOI22xp33_ASAP7_75t_L g3385 ( 
.A1(n_3299),
.A2(n_1752),
.B1(n_1280),
.B2(n_1284),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_3248),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3253),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_SL g3388 ( 
.A(n_3291),
.B(n_1277),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_3267),
.Y(n_3389)
);

AND2x2_ASAP7_75t_L g3390 ( 
.A(n_3241),
.B(n_83),
.Y(n_3390)
);

AND2x2_ASAP7_75t_L g3391 ( 
.A(n_3247),
.B(n_84),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3271),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_3272),
.Y(n_3393)
);

NOR2x1_ASAP7_75t_R g3394 ( 
.A(n_3304),
.B(n_1729),
.Y(n_3394)
);

INVx2_ASAP7_75t_L g3395 ( 
.A(n_3236),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_3278),
.Y(n_3396)
);

AND2x2_ASAP7_75t_L g3397 ( 
.A(n_3331),
.B(n_85),
.Y(n_3397)
);

OR2x2_ASAP7_75t_L g3398 ( 
.A(n_3238),
.B(n_3215),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_3310),
.Y(n_3399)
);

AND2x4_ASAP7_75t_L g3400 ( 
.A(n_3239),
.B(n_3332),
.Y(n_3400)
);

AND2x4_ASAP7_75t_SL g3401 ( 
.A(n_3333),
.B(n_86),
.Y(n_3401)
);

NAND2xp33_ASAP7_75t_L g3402 ( 
.A(n_3286),
.B(n_1287),
.Y(n_3402)
);

NAND2x1_ASAP7_75t_L g3403 ( 
.A(n_3268),
.B(n_3309),
.Y(n_3403)
);

INVx4_ASAP7_75t_L g3404 ( 
.A(n_3344),
.Y(n_3404)
);

INVx2_ASAP7_75t_SL g3405 ( 
.A(n_3257),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3316),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_3318),
.Y(n_3407)
);

NOR2xp33_ASAP7_75t_L g3408 ( 
.A(n_3307),
.B(n_87),
.Y(n_3408)
);

HB1xp67_ASAP7_75t_L g3409 ( 
.A(n_3311),
.Y(n_3409)
);

OR2x2_ASAP7_75t_L g3410 ( 
.A(n_3329),
.B(n_3335),
.Y(n_3410)
);

INVx3_ASAP7_75t_L g3411 ( 
.A(n_3273),
.Y(n_3411)
);

OR2x2_ASAP7_75t_SL g3412 ( 
.A(n_3330),
.B(n_87),
.Y(n_3412)
);

AND2x2_ASAP7_75t_L g3413 ( 
.A(n_3319),
.B(n_88),
.Y(n_3413)
);

INVx2_ASAP7_75t_L g3414 ( 
.A(n_3324),
.Y(n_3414)
);

HB1xp67_ASAP7_75t_L g3415 ( 
.A(n_3360),
.Y(n_3415)
);

BUFx3_ASAP7_75t_L g3416 ( 
.A(n_3264),
.Y(n_3416)
);

AND2x4_ASAP7_75t_L g3417 ( 
.A(n_3222),
.B(n_88),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_3334),
.Y(n_3418)
);

AND2x2_ASAP7_75t_L g3419 ( 
.A(n_3354),
.B(n_89),
.Y(n_3419)
);

AND2x4_ASAP7_75t_L g3420 ( 
.A(n_3357),
.B(n_89),
.Y(n_3420)
);

INVx2_ASAP7_75t_L g3421 ( 
.A(n_3220),
.Y(n_3421)
);

INVx3_ASAP7_75t_L g3422 ( 
.A(n_3274),
.Y(n_3422)
);

BUFx2_ASAP7_75t_SL g3423 ( 
.A(n_3214),
.Y(n_3423)
);

HB1xp67_ASAP7_75t_L g3424 ( 
.A(n_3361),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_3223),
.B(n_90),
.Y(n_3425)
);

INVx3_ASAP7_75t_L g3426 ( 
.A(n_3225),
.Y(n_3426)
);

AND2x2_ASAP7_75t_L g3427 ( 
.A(n_3258),
.B(n_90),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_3340),
.Y(n_3428)
);

AND2x2_ASAP7_75t_L g3429 ( 
.A(n_3263),
.B(n_91),
.Y(n_3429)
);

AND2x2_ASAP7_75t_L g3430 ( 
.A(n_3249),
.B(n_92),
.Y(n_3430)
);

AND2x2_ASAP7_75t_L g3431 ( 
.A(n_3252),
.B(n_93),
.Y(n_3431)
);

AND2x2_ASAP7_75t_L g3432 ( 
.A(n_3276),
.B(n_94),
.Y(n_3432)
);

INVx2_ASAP7_75t_L g3433 ( 
.A(n_3231),
.Y(n_3433)
);

AND2x2_ASAP7_75t_L g3434 ( 
.A(n_3277),
.B(n_3217),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_3345),
.Y(n_3435)
);

HB1xp67_ASAP7_75t_L g3436 ( 
.A(n_3350),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_3254),
.B(n_94),
.Y(n_3437)
);

INVx1_ASAP7_75t_L g3438 ( 
.A(n_3349),
.Y(n_3438)
);

NOR2xp33_ASAP7_75t_SL g3439 ( 
.A(n_3266),
.B(n_1678),
.Y(n_3439)
);

AND2x4_ASAP7_75t_L g3440 ( 
.A(n_3210),
.B(n_95),
.Y(n_3440)
);

AND2x2_ASAP7_75t_L g3441 ( 
.A(n_3221),
.B(n_95),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_3352),
.Y(n_3442)
);

INVx2_ASAP7_75t_L g3443 ( 
.A(n_3244),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_3237),
.B(n_96),
.Y(n_3444)
);

INVx4_ASAP7_75t_L g3445 ( 
.A(n_3285),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_3312),
.B(n_3325),
.Y(n_3446)
);

AND2x2_ASAP7_75t_L g3447 ( 
.A(n_3326),
.B(n_96),
.Y(n_3447)
);

AND2x2_ASAP7_75t_L g3448 ( 
.A(n_3338),
.B(n_97),
.Y(n_3448)
);

INVx2_ASAP7_75t_L g3449 ( 
.A(n_3259),
.Y(n_3449)
);

AND2x4_ASAP7_75t_L g3450 ( 
.A(n_3341),
.B(n_97),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_3358),
.Y(n_3451)
);

AND2x4_ASAP7_75t_L g3452 ( 
.A(n_3343),
.B(n_98),
.Y(n_3452)
);

AND2x2_ASAP7_75t_L g3453 ( 
.A(n_3348),
.B(n_100),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3246),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_3288),
.Y(n_3455)
);

AND2x4_ASAP7_75t_L g3456 ( 
.A(n_3351),
.B(n_100),
.Y(n_3456)
);

INVx2_ASAP7_75t_L g3457 ( 
.A(n_3280),
.Y(n_3457)
);

AND2x2_ASAP7_75t_L g3458 ( 
.A(n_3356),
.B(n_101),
.Y(n_3458)
);

AND2x2_ASAP7_75t_L g3459 ( 
.A(n_3320),
.B(n_102),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_3284),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_3290),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_3293),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_3270),
.Y(n_3463)
);

OR2x2_ASAP7_75t_L g3464 ( 
.A(n_3342),
.B(n_102),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_3282),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_3350),
.Y(n_3466)
);

AND2x2_ASAP7_75t_L g3467 ( 
.A(n_3359),
.B(n_103),
.Y(n_3467)
);

AND2x2_ASAP7_75t_L g3468 ( 
.A(n_3269),
.B(n_103),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_L g3469 ( 
.A(n_3313),
.B(n_104),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_L g3470 ( 
.A(n_3289),
.B(n_3234),
.Y(n_3470)
);

NOR2xp33_ASAP7_75t_L g3471 ( 
.A(n_3301),
.B(n_104),
.Y(n_3471)
);

AND2x2_ASAP7_75t_L g3472 ( 
.A(n_3232),
.B(n_105),
.Y(n_3472)
);

AND2x2_ASAP7_75t_L g3473 ( 
.A(n_3302),
.B(n_105),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_3213),
.B(n_106),
.Y(n_3474)
);

INVx2_ASAP7_75t_L g3475 ( 
.A(n_3227),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_3317),
.B(n_106),
.Y(n_3476)
);

AND2x2_ASAP7_75t_L g3477 ( 
.A(n_3300),
.B(n_107),
.Y(n_3477)
);

HB1xp67_ASAP7_75t_L g3478 ( 
.A(n_3211),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_3261),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3283),
.Y(n_3480)
);

INVx2_ASAP7_75t_L g3481 ( 
.A(n_3327),
.Y(n_3481)
);

AND2x2_ASAP7_75t_L g3482 ( 
.A(n_3306),
.B(n_107),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_3328),
.Y(n_3483)
);

INVx2_ASAP7_75t_L g3484 ( 
.A(n_3305),
.Y(n_3484)
);

AND2x2_ASAP7_75t_L g3485 ( 
.A(n_3337),
.B(n_108),
.Y(n_3485)
);

OR2x2_ASAP7_75t_L g3486 ( 
.A(n_3339),
.B(n_109),
.Y(n_3486)
);

INVx3_ASAP7_75t_L g3487 ( 
.A(n_3303),
.Y(n_3487)
);

HB1xp67_ASAP7_75t_L g3488 ( 
.A(n_3346),
.Y(n_3488)
);

NOR2x1_ASAP7_75t_L g3489 ( 
.A(n_3322),
.B(n_110),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_3216),
.Y(n_3490)
);

INVx2_ASAP7_75t_L g3491 ( 
.A(n_3296),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_3279),
.Y(n_3492)
);

AND2x4_ASAP7_75t_SL g3493 ( 
.A(n_3353),
.B(n_110),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3228),
.Y(n_3494)
);

NOR2x1_ASAP7_75t_L g3495 ( 
.A(n_3355),
.B(n_3275),
.Y(n_3495)
);

AND2x2_ASAP7_75t_L g3496 ( 
.A(n_3230),
.B(n_111),
.Y(n_3496)
);

AND2x4_ASAP7_75t_L g3497 ( 
.A(n_3245),
.B(n_111),
.Y(n_3497)
);

AND2x2_ASAP7_75t_L g3498 ( 
.A(n_3219),
.B(n_3229),
.Y(n_3498)
);

AND2x4_ASAP7_75t_SL g3499 ( 
.A(n_3308),
.B(n_112),
.Y(n_3499)
);

AND2x2_ASAP7_75t_L g3500 ( 
.A(n_3292),
.B(n_112),
.Y(n_3500)
);

OR2x2_ASAP7_75t_L g3501 ( 
.A(n_3260),
.B(n_113),
.Y(n_3501)
);

INVx2_ASAP7_75t_L g3502 ( 
.A(n_3255),
.Y(n_3502)
);

INVx2_ASAP7_75t_L g3503 ( 
.A(n_3226),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3314),
.Y(n_3504)
);

HB1xp67_ASAP7_75t_L g3505 ( 
.A(n_3336),
.Y(n_3505)
);

AND2x2_ASAP7_75t_L g3506 ( 
.A(n_3265),
.B(n_113),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3281),
.Y(n_3507)
);

AND2x2_ASAP7_75t_L g3508 ( 
.A(n_3262),
.B(n_114),
.Y(n_3508)
);

INVx2_ASAP7_75t_L g3509 ( 
.A(n_3287),
.Y(n_3509)
);

INVx2_ASAP7_75t_L g3510 ( 
.A(n_3256),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_3208),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_3208),
.Y(n_3512)
);

AND2x2_ASAP7_75t_L g3513 ( 
.A(n_3243),
.B(n_115),
.Y(n_3513)
);

AND2x2_ASAP7_75t_L g3514 ( 
.A(n_3243),
.B(n_115),
.Y(n_3514)
);

AND2x2_ASAP7_75t_L g3515 ( 
.A(n_3243),
.B(n_116),
.Y(n_3515)
);

INVx3_ASAP7_75t_L g3516 ( 
.A(n_3321),
.Y(n_3516)
);

INVxp67_ASAP7_75t_L g3517 ( 
.A(n_3362),
.Y(n_3517)
);

INVx2_ASAP7_75t_L g3518 ( 
.A(n_3256),
.Y(n_3518)
);

OR2x2_ASAP7_75t_L g3519 ( 
.A(n_3218),
.B(n_116),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_3208),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_3294),
.B(n_117),
.Y(n_3521)
);

AND2x2_ASAP7_75t_L g3522 ( 
.A(n_3243),
.B(n_117),
.Y(n_3522)
);

INVx2_ASAP7_75t_L g3523 ( 
.A(n_3256),
.Y(n_3523)
);

INVx2_ASAP7_75t_L g3524 ( 
.A(n_3256),
.Y(n_3524)
);

AND2x2_ASAP7_75t_L g3525 ( 
.A(n_3243),
.B(n_119),
.Y(n_3525)
);

AND2x2_ASAP7_75t_L g3526 ( 
.A(n_3243),
.B(n_120),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_L g3527 ( 
.A(n_3294),
.B(n_121),
.Y(n_3527)
);

AND2x2_ASAP7_75t_L g3528 ( 
.A(n_3243),
.B(n_121),
.Y(n_3528)
);

AND2x2_ASAP7_75t_L g3529 ( 
.A(n_3243),
.B(n_124),
.Y(n_3529)
);

INVx1_ASAP7_75t_SL g3530 ( 
.A(n_3240),
.Y(n_3530)
);

HB1xp67_ASAP7_75t_L g3531 ( 
.A(n_3362),
.Y(n_3531)
);

INVx2_ASAP7_75t_L g3532 ( 
.A(n_3256),
.Y(n_3532)
);

AND2x4_ASAP7_75t_L g3533 ( 
.A(n_3224),
.B(n_125),
.Y(n_3533)
);

OR2x2_ASAP7_75t_L g3534 ( 
.A(n_3218),
.B(n_125),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3208),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_3294),
.B(n_126),
.Y(n_3536)
);

OR2x2_ASAP7_75t_L g3537 ( 
.A(n_3218),
.B(n_126),
.Y(n_3537)
);

INVx4_ASAP7_75t_L g3538 ( 
.A(n_3321),
.Y(n_3538)
);

AND2x2_ASAP7_75t_L g3539 ( 
.A(n_3243),
.B(n_127),
.Y(n_3539)
);

INVx2_ASAP7_75t_L g3540 ( 
.A(n_3256),
.Y(n_3540)
);

NOR2xp33_ASAP7_75t_L g3541 ( 
.A(n_3321),
.B(n_127),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_3256),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_L g3543 ( 
.A(n_3294),
.B(n_128),
.Y(n_3543)
);

INVx2_ASAP7_75t_L g3544 ( 
.A(n_3256),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3208),
.Y(n_3545)
);

AND2x2_ASAP7_75t_L g3546 ( 
.A(n_3243),
.B(n_128),
.Y(n_3546)
);

INVx2_ASAP7_75t_L g3547 ( 
.A(n_3256),
.Y(n_3547)
);

INVx1_ASAP7_75t_L g3548 ( 
.A(n_3208),
.Y(n_3548)
);

AND2x2_ASAP7_75t_L g3549 ( 
.A(n_3243),
.B(n_129),
.Y(n_3549)
);

AND2x2_ASAP7_75t_L g3550 ( 
.A(n_3243),
.B(n_129),
.Y(n_3550)
);

AND2x2_ASAP7_75t_L g3551 ( 
.A(n_3243),
.B(n_130),
.Y(n_3551)
);

OR2x2_ASAP7_75t_L g3552 ( 
.A(n_3218),
.B(n_130),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_3492),
.B(n_131),
.Y(n_3553)
);

OAI31xp33_ASAP7_75t_L g3554 ( 
.A1(n_3496),
.A2(n_3501),
.A3(n_3439),
.B(n_3503),
.Y(n_3554)
);

INVxp67_ASAP7_75t_L g3555 ( 
.A(n_3423),
.Y(n_3555)
);

BUFx2_ASAP7_75t_L g3556 ( 
.A(n_3538),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3409),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3415),
.Y(n_3558)
);

INVxp67_ASAP7_75t_SL g3559 ( 
.A(n_3380),
.Y(n_3559)
);

INVx2_ASAP7_75t_L g3560 ( 
.A(n_3400),
.Y(n_3560)
);

NAND2xp67_ASAP7_75t_L g3561 ( 
.A(n_3372),
.B(n_131),
.Y(n_3561)
);

HB1xp67_ASAP7_75t_L g3562 ( 
.A(n_3531),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3424),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3461),
.Y(n_3564)
);

AND2x2_ASAP7_75t_L g3565 ( 
.A(n_3530),
.B(n_132),
.Y(n_3565)
);

OR2x2_ASAP7_75t_L g3566 ( 
.A(n_3410),
.B(n_132),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_3375),
.B(n_133),
.Y(n_3567)
);

OAI31xp33_ASAP7_75t_L g3568 ( 
.A1(n_3388),
.A2(n_135),
.A3(n_133),
.B(n_134),
.Y(n_3568)
);

A2O1A1Ixp33_ASAP7_75t_L g3569 ( 
.A1(n_3489),
.A2(n_1302),
.B(n_1304),
.C(n_1290),
.Y(n_3569)
);

AND2x2_ASAP7_75t_L g3570 ( 
.A(n_3516),
.B(n_135),
.Y(n_3570)
);

AND2x4_ASAP7_75t_L g3571 ( 
.A(n_3367),
.B(n_136),
.Y(n_3571)
);

NOR2xp33_ASAP7_75t_L g3572 ( 
.A(n_3382),
.B(n_137),
.Y(n_3572)
);

INVx1_ASAP7_75t_SL g3573 ( 
.A(n_3401),
.Y(n_3573)
);

INVx1_ASAP7_75t_SL g3574 ( 
.A(n_3533),
.Y(n_3574)
);

AOI22xp5_ASAP7_75t_L g3575 ( 
.A1(n_3498),
.A2(n_1309),
.B1(n_1313),
.B2(n_1306),
.Y(n_3575)
);

AND2x2_ASAP7_75t_L g3576 ( 
.A(n_3510),
.B(n_3518),
.Y(n_3576)
);

NAND3xp33_ASAP7_75t_L g3577 ( 
.A(n_3517),
.B(n_1344),
.C(n_1316),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3462),
.Y(n_3578)
);

INVx2_ASAP7_75t_L g3579 ( 
.A(n_3404),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3487),
.B(n_137),
.Y(n_3580)
);

NAND2x1_ASAP7_75t_L g3581 ( 
.A(n_3411),
.B(n_138),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3478),
.Y(n_3582)
);

AND2x2_ASAP7_75t_L g3583 ( 
.A(n_3523),
.B(n_138),
.Y(n_3583)
);

AND2x2_ASAP7_75t_L g3584 ( 
.A(n_3524),
.B(n_140),
.Y(n_3584)
);

INVx3_ASAP7_75t_L g3585 ( 
.A(n_3445),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3364),
.B(n_142),
.Y(n_3586)
);

NAND2x2_ASAP7_75t_L g3587 ( 
.A(n_3405),
.B(n_143),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3463),
.Y(n_3588)
);

OR2x2_ASAP7_75t_L g3589 ( 
.A(n_3426),
.B(n_143),
.Y(n_3589)
);

OR2x2_ASAP7_75t_L g3590 ( 
.A(n_3475),
.B(n_144),
.Y(n_3590)
);

INVx1_ASAP7_75t_L g3591 ( 
.A(n_3465),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_3434),
.B(n_144),
.Y(n_3592)
);

NOR2xp33_ASAP7_75t_L g3593 ( 
.A(n_3481),
.B(n_145),
.Y(n_3593)
);

INVx3_ASAP7_75t_L g3594 ( 
.A(n_3416),
.Y(n_3594)
);

NOR2xp67_ASAP7_75t_SL g3595 ( 
.A(n_3507),
.B(n_1347),
.Y(n_3595)
);

AND2x2_ASAP7_75t_L g3596 ( 
.A(n_3532),
.B(n_145),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_3368),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3484),
.B(n_3540),
.Y(n_3598)
);

AND2x2_ASAP7_75t_L g3599 ( 
.A(n_3542),
.B(n_3544),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_3370),
.Y(n_3600)
);

AND2x2_ASAP7_75t_L g3601 ( 
.A(n_3547),
.B(n_3395),
.Y(n_3601)
);

INVxp67_ASAP7_75t_SL g3602 ( 
.A(n_3436),
.Y(n_3602)
);

AND2x2_ASAP7_75t_L g3603 ( 
.A(n_3422),
.B(n_148),
.Y(n_3603)
);

INVx1_ASAP7_75t_L g3604 ( 
.A(n_3376),
.Y(n_3604)
);

AND2x2_ASAP7_75t_L g3605 ( 
.A(n_3491),
.B(n_149),
.Y(n_3605)
);

NAND2x1p5_ASAP7_75t_L g3606 ( 
.A(n_3403),
.B(n_3365),
.Y(n_3606)
);

INVx2_ASAP7_75t_L g3607 ( 
.A(n_3466),
.Y(n_3607)
);

AOI21xp33_ASAP7_75t_L g3608 ( 
.A1(n_3505),
.A2(n_149),
.B(n_151),
.Y(n_3608)
);

NAND2xp67_ASAP7_75t_SL g3609 ( 
.A(n_3472),
.B(n_152),
.Y(n_3609)
);

INVx3_ASAP7_75t_L g3610 ( 
.A(n_3420),
.Y(n_3610)
);

AND2x2_ASAP7_75t_L g3611 ( 
.A(n_3479),
.B(n_153),
.Y(n_3611)
);

INVx4_ASAP7_75t_L g3612 ( 
.A(n_3391),
.Y(n_3612)
);

NOR2xp67_ASAP7_75t_L g3613 ( 
.A(n_3398),
.B(n_154),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3381),
.Y(n_3614)
);

AOI21xp33_ASAP7_75t_L g3615 ( 
.A1(n_3394),
.A2(n_154),
.B(n_155),
.Y(n_3615)
);

INVx1_ASAP7_75t_SL g3616 ( 
.A(n_3374),
.Y(n_3616)
);

A2O1A1Ixp33_ASAP7_75t_L g3617 ( 
.A1(n_3469),
.A2(n_1359),
.B(n_1372),
.C(n_1352),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_3383),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_3386),
.Y(n_3619)
);

AND2x2_ASAP7_75t_L g3620 ( 
.A(n_3480),
.B(n_156),
.Y(n_3620)
);

AOI22xp5_ASAP7_75t_L g3621 ( 
.A1(n_3408),
.A2(n_1375),
.B1(n_1380),
.B2(n_1373),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_L g3622 ( 
.A(n_3483),
.B(n_157),
.Y(n_3622)
);

AND2x2_ASAP7_75t_L g3623 ( 
.A(n_3473),
.B(n_157),
.Y(n_3623)
);

AND2x2_ASAP7_75t_L g3624 ( 
.A(n_3477),
.B(n_158),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_L g3625 ( 
.A(n_3488),
.B(n_159),
.Y(n_3625)
);

AND2x2_ASAP7_75t_L g3626 ( 
.A(n_3454),
.B(n_160),
.Y(n_3626)
);

AND2x2_ASAP7_75t_L g3627 ( 
.A(n_3373),
.B(n_160),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_3387),
.Y(n_3628)
);

INVx1_ASAP7_75t_SL g3629 ( 
.A(n_3384),
.Y(n_3629)
);

NOR2xp33_ASAP7_75t_L g3630 ( 
.A(n_3446),
.B(n_161),
.Y(n_3630)
);

NAND2xp5_ASAP7_75t_L g3631 ( 
.A(n_3490),
.B(n_161),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3389),
.Y(n_3632)
);

AND2x2_ASAP7_75t_L g3633 ( 
.A(n_3519),
.B(n_3534),
.Y(n_3633)
);

INVxp67_ASAP7_75t_SL g3634 ( 
.A(n_3437),
.Y(n_3634)
);

INVx2_ASAP7_75t_L g3635 ( 
.A(n_3414),
.Y(n_3635)
);

INVx2_ASAP7_75t_SL g3636 ( 
.A(n_3390),
.Y(n_3636)
);

INVx1_ASAP7_75t_SL g3637 ( 
.A(n_3499),
.Y(n_3637)
);

NOR2x1_ASAP7_75t_SL g3638 ( 
.A(n_3537),
.B(n_163),
.Y(n_3638)
);

INVx1_ASAP7_75t_SL g3639 ( 
.A(n_3397),
.Y(n_3639)
);

INVx2_ASAP7_75t_L g3640 ( 
.A(n_3413),
.Y(n_3640)
);

AOI21xp33_ASAP7_75t_SL g3641 ( 
.A1(n_3552),
.A2(n_162),
.B(n_163),
.Y(n_3641)
);

NOR2x1_ASAP7_75t_R g3642 ( 
.A(n_3497),
.B(n_1382),
.Y(n_3642)
);

OR2x2_ASAP7_75t_L g3643 ( 
.A(n_3460),
.B(n_162),
.Y(n_3643)
);

OR2x2_ASAP7_75t_L g3644 ( 
.A(n_3421),
.B(n_166),
.Y(n_3644)
);

NAND2x1p5_ASAP7_75t_L g3645 ( 
.A(n_3513),
.B(n_166),
.Y(n_3645)
);

INVx2_ASAP7_75t_L g3646 ( 
.A(n_3419),
.Y(n_3646)
);

AND2x2_ASAP7_75t_L g3647 ( 
.A(n_3470),
.B(n_167),
.Y(n_3647)
);

AND2x2_ASAP7_75t_L g3648 ( 
.A(n_3459),
.B(n_167),
.Y(n_3648)
);

AOI21xp33_ASAP7_75t_L g3649 ( 
.A1(n_3371),
.A2(n_168),
.B(n_169),
.Y(n_3649)
);

OAI32xp33_ASAP7_75t_L g3650 ( 
.A1(n_3444),
.A2(n_191),
.A3(n_200),
.B1(n_181),
.B2(n_169),
.Y(n_3650)
);

INVx1_ASAP7_75t_SL g3651 ( 
.A(n_3441),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_3392),
.Y(n_3652)
);

AND2x2_ASAP7_75t_L g3653 ( 
.A(n_3467),
.B(n_170),
.Y(n_3653)
);

AND2x2_ASAP7_75t_L g3654 ( 
.A(n_3433),
.B(n_170),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3393),
.Y(n_3655)
);

INVx1_ASAP7_75t_L g3656 ( 
.A(n_3396),
.Y(n_3656)
);

AND2x2_ASAP7_75t_L g3657 ( 
.A(n_3443),
.B(n_3449),
.Y(n_3657)
);

INVxp67_ASAP7_75t_SL g3658 ( 
.A(n_3541),
.Y(n_3658)
);

INVxp67_ASAP7_75t_L g3659 ( 
.A(n_3379),
.Y(n_3659)
);

INVxp67_ASAP7_75t_L g3660 ( 
.A(n_3366),
.Y(n_3660)
);

AND2x2_ASAP7_75t_L g3661 ( 
.A(n_3457),
.B(n_171),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3399),
.Y(n_3662)
);

NAND2x1_ASAP7_75t_L g3663 ( 
.A(n_3432),
.B(n_3406),
.Y(n_3663)
);

OR2x2_ASAP7_75t_L g3664 ( 
.A(n_3378),
.B(n_172),
.Y(n_3664)
);

INVx2_ASAP7_75t_L g3665 ( 
.A(n_3514),
.Y(n_3665)
);

INVx2_ASAP7_75t_L g3666 ( 
.A(n_3515),
.Y(n_3666)
);

INVxp67_ASAP7_75t_L g3667 ( 
.A(n_3494),
.Y(n_3667)
);

OAI22xp5_ASAP7_75t_L g3668 ( 
.A1(n_3385),
.A2(n_1385),
.B1(n_1389),
.B2(n_1384),
.Y(n_3668)
);

AND2x2_ASAP7_75t_L g3669 ( 
.A(n_3447),
.B(n_3448),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_L g3670 ( 
.A(n_3471),
.B(n_172),
.Y(n_3670)
);

OR2x2_ASAP7_75t_L g3671 ( 
.A(n_3455),
.B(n_176),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_3522),
.B(n_176),
.Y(n_3672)
);

INVxp67_ASAP7_75t_SL g3673 ( 
.A(n_3495),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_3407),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3418),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_3525),
.B(n_177),
.Y(n_3676)
);

NOR2x1_ASAP7_75t_L g3677 ( 
.A(n_3521),
.B(n_178),
.Y(n_3677)
);

INVx2_ASAP7_75t_L g3678 ( 
.A(n_3526),
.Y(n_3678)
);

INVx3_ASAP7_75t_L g3679 ( 
.A(n_3417),
.Y(n_3679)
);

INVx2_ASAP7_75t_SL g3680 ( 
.A(n_3528),
.Y(n_3680)
);

OR2x2_ASAP7_75t_L g3681 ( 
.A(n_3428),
.B(n_179),
.Y(n_3681)
);

OAI21xp33_ASAP7_75t_L g3682 ( 
.A1(n_3509),
.A2(n_1403),
.B(n_1396),
.Y(n_3682)
);

AND2x4_ASAP7_75t_L g3683 ( 
.A(n_3529),
.B(n_181),
.Y(n_3683)
);

INVx1_ASAP7_75t_L g3684 ( 
.A(n_3435),
.Y(n_3684)
);

INVx2_ASAP7_75t_L g3685 ( 
.A(n_3539),
.Y(n_3685)
);

AND2x2_ASAP7_75t_L g3686 ( 
.A(n_3453),
.B(n_182),
.Y(n_3686)
);

NOR2xp33_ASAP7_75t_L g3687 ( 
.A(n_3612),
.B(n_3502),
.Y(n_3687)
);

HB1xp67_ASAP7_75t_L g3688 ( 
.A(n_3613),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_3562),
.Y(n_3689)
);

NAND2xp5_ASAP7_75t_L g3690 ( 
.A(n_3574),
.B(n_3504),
.Y(n_3690)
);

NOR2xp33_ASAP7_75t_L g3691 ( 
.A(n_3556),
.B(n_3363),
.Y(n_3691)
);

BUFx2_ASAP7_75t_L g3692 ( 
.A(n_3559),
.Y(n_3692)
);

AND2x2_ASAP7_75t_L g3693 ( 
.A(n_3560),
.B(n_3546),
.Y(n_3693)
);

OR2x2_ASAP7_75t_L g3694 ( 
.A(n_3651),
.B(n_3527),
.Y(n_3694)
);

AND2x2_ASAP7_75t_L g3695 ( 
.A(n_3585),
.B(n_3549),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3582),
.Y(n_3696)
);

AND2x4_ASAP7_75t_L g3697 ( 
.A(n_3579),
.B(n_3550),
.Y(n_3697)
);

NOR2xp33_ASAP7_75t_L g3698 ( 
.A(n_3637),
.B(n_3536),
.Y(n_3698)
);

AND2x2_ASAP7_75t_L g3699 ( 
.A(n_3594),
.B(n_3551),
.Y(n_3699)
);

NAND2x1_ASAP7_75t_L g3700 ( 
.A(n_3610),
.B(n_3438),
.Y(n_3700)
);

HB1xp67_ASAP7_75t_L g3701 ( 
.A(n_3555),
.Y(n_3701)
);

NAND2x1p5_ASAP7_75t_L g3702 ( 
.A(n_3581),
.B(n_3440),
.Y(n_3702)
);

INVx2_ASAP7_75t_L g3703 ( 
.A(n_3606),
.Y(n_3703)
);

OR2x2_ASAP7_75t_L g3704 ( 
.A(n_3616),
.B(n_3543),
.Y(n_3704)
);

INVx2_ASAP7_75t_L g3705 ( 
.A(n_3576),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3557),
.Y(n_3706)
);

INVx2_ASAP7_75t_SL g3707 ( 
.A(n_3599),
.Y(n_3707)
);

AOI22xp33_ASAP7_75t_L g3708 ( 
.A1(n_3673),
.A2(n_3508),
.B1(n_3451),
.B2(n_3442),
.Y(n_3708)
);

AND2x2_ASAP7_75t_L g3709 ( 
.A(n_3669),
.B(n_3485),
.Y(n_3709)
);

BUFx2_ASAP7_75t_L g3710 ( 
.A(n_3602),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3558),
.Y(n_3711)
);

HB1xp67_ASAP7_75t_L g3712 ( 
.A(n_3663),
.Y(n_3712)
);

INVxp67_ASAP7_75t_SL g3713 ( 
.A(n_3638),
.Y(n_3713)
);

INVxp67_ASAP7_75t_L g3714 ( 
.A(n_3677),
.Y(n_3714)
);

AND2x2_ASAP7_75t_L g3715 ( 
.A(n_3601),
.B(n_3468),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3563),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_L g3717 ( 
.A(n_3629),
.B(n_3450),
.Y(n_3717)
);

AOI222xp33_ASAP7_75t_L g3718 ( 
.A1(n_3634),
.A2(n_3506),
.B1(n_3500),
.B2(n_3377),
.C1(n_3402),
.C2(n_3476),
.Y(n_3718)
);

INVx1_ASAP7_75t_SL g3719 ( 
.A(n_3573),
.Y(n_3719)
);

NAND3xp33_ASAP7_75t_L g3720 ( 
.A(n_3554),
.B(n_3568),
.C(n_3569),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_3590),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_3644),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_L g3723 ( 
.A(n_3633),
.B(n_3452),
.Y(n_3723)
);

INVx2_ASAP7_75t_L g3724 ( 
.A(n_3679),
.Y(n_3724)
);

INVx2_ASAP7_75t_L g3725 ( 
.A(n_3571),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3564),
.Y(n_3726)
);

AND2x2_ASAP7_75t_L g3727 ( 
.A(n_3639),
.B(n_3458),
.Y(n_3727)
);

AND2x2_ASAP7_75t_L g3728 ( 
.A(n_3636),
.B(n_3427),
.Y(n_3728)
);

OR2x6_ASAP7_75t_L g3729 ( 
.A(n_3645),
.B(n_3464),
.Y(n_3729)
);

OR2x2_ASAP7_75t_L g3730 ( 
.A(n_3598),
.B(n_3511),
.Y(n_3730)
);

INVx2_ASAP7_75t_L g3731 ( 
.A(n_3583),
.Y(n_3731)
);

AOI22xp33_ASAP7_75t_L g3732 ( 
.A1(n_3667),
.A2(n_3512),
.B1(n_3535),
.B2(n_3520),
.Y(n_3732)
);

OA21x2_ASAP7_75t_L g3733 ( 
.A1(n_3553),
.A2(n_3548),
.B(n_3545),
.Y(n_3733)
);

INVx2_ASAP7_75t_L g3734 ( 
.A(n_3584),
.Y(n_3734)
);

AND2x2_ASAP7_75t_L g3735 ( 
.A(n_3665),
.B(n_3429),
.Y(n_3735)
);

AND2x2_ASAP7_75t_L g3736 ( 
.A(n_3666),
.B(n_3430),
.Y(n_3736)
);

INVx1_ASAP7_75t_SL g3737 ( 
.A(n_3565),
.Y(n_3737)
);

INVx1_ASAP7_75t_SL g3738 ( 
.A(n_3570),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3578),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3643),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3671),
.Y(n_3741)
);

AND2x2_ASAP7_75t_L g3742 ( 
.A(n_3678),
.B(n_3431),
.Y(n_3742)
);

OR2x2_ASAP7_75t_L g3743 ( 
.A(n_3640),
.B(n_3425),
.Y(n_3743)
);

INVx2_ASAP7_75t_L g3744 ( 
.A(n_3596),
.Y(n_3744)
);

INVx2_ASAP7_75t_L g3745 ( 
.A(n_3680),
.Y(n_3745)
);

OR2x2_ASAP7_75t_L g3746 ( 
.A(n_3646),
.B(n_3369),
.Y(n_3746)
);

OAI21xp5_ASAP7_75t_L g3747 ( 
.A1(n_3617),
.A2(n_3486),
.B(n_3474),
.Y(n_3747)
);

AOI33xp33_ASAP7_75t_L g3748 ( 
.A1(n_3588),
.A2(n_3493),
.A3(n_3482),
.B1(n_3456),
.B2(n_3412),
.B3(n_185),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3681),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_3626),
.Y(n_3750)
);

INVx1_ASAP7_75t_L g3751 ( 
.A(n_3589),
.Y(n_3751)
);

NAND2xp5_ASAP7_75t_L g3752 ( 
.A(n_3658),
.B(n_3412),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3654),
.Y(n_3753)
);

OR2x6_ASAP7_75t_L g3754 ( 
.A(n_3659),
.B(n_182),
.Y(n_3754)
);

HB1xp67_ASAP7_75t_L g3755 ( 
.A(n_3561),
.Y(n_3755)
);

AND2x2_ASAP7_75t_L g3756 ( 
.A(n_3685),
.B(n_183),
.Y(n_3756)
);

OR2x2_ASAP7_75t_L g3757 ( 
.A(n_3566),
.B(n_3591),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_L g3758 ( 
.A(n_3630),
.B(n_3607),
.Y(n_3758)
);

NAND2xp5_ASAP7_75t_L g3759 ( 
.A(n_3660),
.B(n_183),
.Y(n_3759)
);

OAI22xp5_ASAP7_75t_L g3760 ( 
.A1(n_3587),
.A2(n_1709),
.B1(n_1717),
.B2(n_1683),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3661),
.Y(n_3761)
);

NAND2xp5_ASAP7_75t_L g3762 ( 
.A(n_3657),
.B(n_3641),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3597),
.Y(n_3763)
);

OR2x6_ASAP7_75t_L g3764 ( 
.A(n_3567),
.B(n_185),
.Y(n_3764)
);

AND2x2_ASAP7_75t_L g3765 ( 
.A(n_3647),
.B(n_186),
.Y(n_3765)
);

HB1xp67_ASAP7_75t_L g3766 ( 
.A(n_3586),
.Y(n_3766)
);

AND2x2_ASAP7_75t_L g3767 ( 
.A(n_3623),
.B(n_186),
.Y(n_3767)
);

BUFx2_ASAP7_75t_L g3768 ( 
.A(n_3609),
.Y(n_3768)
);

AOI22xp33_ASAP7_75t_L g3769 ( 
.A1(n_3635),
.A2(n_1408),
.B1(n_1410),
.B2(n_1404),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_3600),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_3604),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3614),
.Y(n_3772)
);

BUFx2_ASAP7_75t_L g3773 ( 
.A(n_3603),
.Y(n_3773)
);

AND2x2_ASAP7_75t_L g3774 ( 
.A(n_3624),
.B(n_188),
.Y(n_3774)
);

OAI33xp33_ASAP7_75t_L g3775 ( 
.A1(n_3618),
.A2(n_1429),
.A3(n_1416),
.B1(n_1441),
.B2(n_1420),
.B3(n_1412),
.Y(n_3775)
);

BUFx3_ASAP7_75t_L g3776 ( 
.A(n_3692),
.Y(n_3776)
);

AND2x2_ASAP7_75t_L g3777 ( 
.A(n_3719),
.B(n_3572),
.Y(n_3777)
);

OR2x2_ASAP7_75t_L g3778 ( 
.A(n_3714),
.B(n_3592),
.Y(n_3778)
);

AND2x2_ASAP7_75t_L g3779 ( 
.A(n_3699),
.B(n_3648),
.Y(n_3779)
);

INVx2_ASAP7_75t_L g3780 ( 
.A(n_3702),
.Y(n_3780)
);

AO21x2_ASAP7_75t_L g3781 ( 
.A1(n_3752),
.A2(n_3625),
.B(n_3608),
.Y(n_3781)
);

AND2x2_ASAP7_75t_L g3782 ( 
.A(n_3695),
.B(n_3653),
.Y(n_3782)
);

INVx2_ASAP7_75t_L g3783 ( 
.A(n_3710),
.Y(n_3783)
);

NAND2xp5_ASAP7_75t_L g3784 ( 
.A(n_3713),
.B(n_3593),
.Y(n_3784)
);

INVx1_ASAP7_75t_L g3785 ( 
.A(n_3701),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_3688),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3689),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3756),
.Y(n_3788)
);

OR2x2_ASAP7_75t_L g3789 ( 
.A(n_3737),
.B(n_3631),
.Y(n_3789)
);

INVx2_ASAP7_75t_L g3790 ( 
.A(n_3700),
.Y(n_3790)
);

AND2x4_ASAP7_75t_L g3791 ( 
.A(n_3697),
.B(n_3683),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_3755),
.B(n_3627),
.Y(n_3792)
);

INVx2_ASAP7_75t_L g3793 ( 
.A(n_3729),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_3727),
.Y(n_3794)
);

INVx3_ASAP7_75t_L g3795 ( 
.A(n_3724),
.Y(n_3795)
);

INVx2_ASAP7_75t_L g3796 ( 
.A(n_3729),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_L g3797 ( 
.A(n_3748),
.B(n_3715),
.Y(n_3797)
);

OR2x2_ASAP7_75t_L g3798 ( 
.A(n_3762),
.B(n_3580),
.Y(n_3798)
);

INVx2_ASAP7_75t_L g3799 ( 
.A(n_3773),
.Y(n_3799)
);

INVx3_ASAP7_75t_L g3800 ( 
.A(n_3703),
.Y(n_3800)
);

INVx2_ASAP7_75t_L g3801 ( 
.A(n_3693),
.Y(n_3801)
);

NAND2xp5_ASAP7_75t_L g3802 ( 
.A(n_3709),
.B(n_3611),
.Y(n_3802)
);

OR2x6_ASAP7_75t_L g3803 ( 
.A(n_3764),
.B(n_3672),
.Y(n_3803)
);

HB1xp67_ASAP7_75t_L g3804 ( 
.A(n_3712),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3757),
.Y(n_3805)
);

NAND2xp5_ASAP7_75t_L g3806 ( 
.A(n_3707),
.B(n_3620),
.Y(n_3806)
);

INVxp67_ASAP7_75t_SL g3807 ( 
.A(n_3723),
.Y(n_3807)
);

AND2x2_ASAP7_75t_L g3808 ( 
.A(n_3728),
.B(n_3686),
.Y(n_3808)
);

INVx2_ASAP7_75t_L g3809 ( 
.A(n_3725),
.Y(n_3809)
);

OR2x2_ASAP7_75t_L g3810 ( 
.A(n_3738),
.B(n_3622),
.Y(n_3810)
);

AND2x2_ASAP7_75t_L g3811 ( 
.A(n_3735),
.B(n_3605),
.Y(n_3811)
);

OR2x2_ASAP7_75t_L g3812 ( 
.A(n_3717),
.B(n_3664),
.Y(n_3812)
);

AND2x2_ASAP7_75t_L g3813 ( 
.A(n_3736),
.B(n_3595),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_L g3814 ( 
.A(n_3768),
.B(n_3619),
.Y(n_3814)
);

INVx1_ASAP7_75t_L g3815 ( 
.A(n_3750),
.Y(n_3815)
);

AND2x2_ASAP7_75t_L g3816 ( 
.A(n_3742),
.B(n_3628),
.Y(n_3816)
);

AND2x4_ASAP7_75t_L g3817 ( 
.A(n_3705),
.B(n_3632),
.Y(n_3817)
);

AND2x2_ASAP7_75t_L g3818 ( 
.A(n_3745),
.B(n_3652),
.Y(n_3818)
);

BUFx2_ASAP7_75t_SL g3819 ( 
.A(n_3767),
.Y(n_3819)
);

OAI22xp5_ASAP7_75t_L g3820 ( 
.A1(n_3708),
.A2(n_3621),
.B1(n_3670),
.B2(n_3575),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_L g3821 ( 
.A(n_3698),
.B(n_3655),
.Y(n_3821)
);

NAND2x1p5_ASAP7_75t_L g3822 ( 
.A(n_3774),
.B(n_3676),
.Y(n_3822)
);

BUFx2_ASAP7_75t_L g3823 ( 
.A(n_3754),
.Y(n_3823)
);

INVx1_ASAP7_75t_L g3824 ( 
.A(n_3740),
.Y(n_3824)
);

NOR2xp33_ASAP7_75t_L g3825 ( 
.A(n_3731),
.B(n_3642),
.Y(n_3825)
);

OR2x2_ASAP7_75t_L g3826 ( 
.A(n_3690),
.B(n_3694),
.Y(n_3826)
);

OR2x2_ASAP7_75t_L g3827 ( 
.A(n_3704),
.B(n_3656),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3721),
.Y(n_3828)
);

NOR2xp67_ASAP7_75t_L g3829 ( 
.A(n_3751),
.B(n_3662),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_3786),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_L g3831 ( 
.A(n_3823),
.B(n_3734),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_L g3832 ( 
.A(n_3776),
.B(n_3744),
.Y(n_3832)
);

AOI22xp5_ASAP7_75t_SL g3833 ( 
.A1(n_3819),
.A2(n_3733),
.B1(n_3760),
.B2(n_3691),
.Y(n_3833)
);

OA22x2_ASAP7_75t_L g3834 ( 
.A1(n_3803),
.A2(n_3696),
.B1(n_3711),
.B2(n_3706),
.Y(n_3834)
);

AOI21xp33_ASAP7_75t_L g3835 ( 
.A1(n_3793),
.A2(n_3687),
.B(n_3720),
.Y(n_3835)
);

AOI21xp5_ASAP7_75t_L g3836 ( 
.A1(n_3820),
.A2(n_3747),
.B(n_3718),
.Y(n_3836)
);

AOI21xp33_ASAP7_75t_SL g3837 ( 
.A1(n_3826),
.A2(n_3749),
.B(n_3741),
.Y(n_3837)
);

INVxp67_ASAP7_75t_SL g3838 ( 
.A(n_3804),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3783),
.Y(n_3839)
);

OAI321xp33_ASAP7_75t_L g3840 ( 
.A1(n_3785),
.A2(n_3716),
.A3(n_3730),
.B1(n_3758),
.B2(n_3770),
.C(n_3763),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_3796),
.B(n_3753),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_SL g3842 ( 
.A(n_3791),
.B(n_3722),
.Y(n_3842)
);

INVx2_ASAP7_75t_L g3843 ( 
.A(n_3790),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3799),
.Y(n_3844)
);

O2A1O1Ixp33_ASAP7_75t_L g3845 ( 
.A1(n_3814),
.A2(n_3766),
.B(n_3754),
.C(n_3615),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3794),
.Y(n_3846)
);

OR2x2_ASAP7_75t_L g3847 ( 
.A(n_3792),
.B(n_3743),
.Y(n_3847)
);

INVx3_ASAP7_75t_L g3848 ( 
.A(n_3780),
.Y(n_3848)
);

OAI31xp33_ASAP7_75t_L g3849 ( 
.A1(n_3784),
.A2(n_3649),
.A3(n_3761),
.B(n_3577),
.Y(n_3849)
);

INVx1_ASAP7_75t_L g3850 ( 
.A(n_3829),
.Y(n_3850)
);

AOI221xp5_ASAP7_75t_L g3851 ( 
.A1(n_3787),
.A2(n_3732),
.B1(n_3650),
.B2(n_3739),
.C(n_3726),
.Y(n_3851)
);

OAI22xp5_ASAP7_75t_L g3852 ( 
.A1(n_3803),
.A2(n_3746),
.B1(n_3764),
.B2(n_3759),
.Y(n_3852)
);

OAI211xp5_ASAP7_75t_L g3853 ( 
.A1(n_3797),
.A2(n_3772),
.B(n_3771),
.C(n_3674),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3809),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_SL g3855 ( 
.A(n_3777),
.B(n_3795),
.Y(n_3855)
);

AOI22xp5_ASAP7_75t_L g3856 ( 
.A1(n_3800),
.A2(n_3775),
.B1(n_3675),
.B2(n_3684),
.Y(n_3856)
);

AOI222xp33_ASAP7_75t_L g3857 ( 
.A1(n_3821),
.A2(n_3682),
.B1(n_3765),
.B2(n_3769),
.C1(n_3668),
.C2(n_1480),
.Y(n_3857)
);

OAI221xp5_ASAP7_75t_L g3858 ( 
.A1(n_3807),
.A2(n_1464),
.B1(n_1484),
.B2(n_1462),
.C(n_1457),
.Y(n_3858)
);

AOI222xp33_ASAP7_75t_L g3859 ( 
.A1(n_3805),
.A2(n_3824),
.B1(n_3828),
.B2(n_3815),
.C1(n_3788),
.C2(n_3808),
.Y(n_3859)
);

AOI21xp33_ASAP7_75t_L g3860 ( 
.A1(n_3778),
.A2(n_189),
.B(n_190),
.Y(n_3860)
);

INVx1_ASAP7_75t_SL g3861 ( 
.A(n_3779),
.Y(n_3861)
);

NOR2xp33_ASAP7_75t_L g3862 ( 
.A(n_3802),
.B(n_189),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_L g3863 ( 
.A(n_3782),
.B(n_190),
.Y(n_3863)
);

INVxp67_ASAP7_75t_L g3864 ( 
.A(n_3811),
.Y(n_3864)
);

INVx1_ASAP7_75t_L g3865 ( 
.A(n_3816),
.Y(n_3865)
);

NOR2xp33_ASAP7_75t_L g3866 ( 
.A(n_3806),
.B(n_192),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3827),
.Y(n_3867)
);

NOR2x1_ASAP7_75t_L g3868 ( 
.A(n_3781),
.B(n_192),
.Y(n_3868)
);

INVx1_ASAP7_75t_SL g3869 ( 
.A(n_3789),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_L g3870 ( 
.A(n_3838),
.B(n_3801),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_3831),
.Y(n_3871)
);

INVx1_ASAP7_75t_L g3872 ( 
.A(n_3832),
.Y(n_3872)
);

AOI22xp33_ASAP7_75t_L g3873 ( 
.A1(n_3836),
.A2(n_3813),
.B1(n_3812),
.B2(n_3798),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_3865),
.Y(n_3874)
);

NAND2xp5_ASAP7_75t_L g3875 ( 
.A(n_3861),
.B(n_3818),
.Y(n_3875)
);

OR2x2_ASAP7_75t_L g3876 ( 
.A(n_3847),
.B(n_3822),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3841),
.Y(n_3877)
);

INVxp67_ASAP7_75t_L g3878 ( 
.A(n_3868),
.Y(n_3878)
);

AND2x2_ASAP7_75t_L g3879 ( 
.A(n_3848),
.B(n_3825),
.Y(n_3879)
);

INVx1_ASAP7_75t_L g3880 ( 
.A(n_3863),
.Y(n_3880)
);

NAND2xp5_ASAP7_75t_L g3881 ( 
.A(n_3848),
.B(n_3850),
.Y(n_3881)
);

HB1xp67_ASAP7_75t_L g3882 ( 
.A(n_3834),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_3864),
.B(n_3817),
.Y(n_3883)
);

OAI22xp33_ASAP7_75t_L g3884 ( 
.A1(n_3869),
.A2(n_3810),
.B1(n_1486),
.B2(n_1489),
.Y(n_3884)
);

NOR2xp33_ASAP7_75t_L g3885 ( 
.A(n_3855),
.B(n_193),
.Y(n_3885)
);

NAND2xp5_ASAP7_75t_L g3886 ( 
.A(n_3843),
.B(n_194),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3867),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3844),
.Y(n_3888)
);

AND2x2_ASAP7_75t_L g3889 ( 
.A(n_3839),
.B(n_194),
.Y(n_3889)
);

NAND2xp5_ASAP7_75t_L g3890 ( 
.A(n_3833),
.B(n_195),
.Y(n_3890)
);

AND2x2_ASAP7_75t_L g3891 ( 
.A(n_3842),
.B(n_197),
.Y(n_3891)
);

INVx1_ASAP7_75t_SL g3892 ( 
.A(n_3830),
.Y(n_3892)
);

INVx1_ASAP7_75t_L g3893 ( 
.A(n_3846),
.Y(n_3893)
);

INVx1_ASAP7_75t_L g3894 ( 
.A(n_3854),
.Y(n_3894)
);

INVxp67_ASAP7_75t_L g3895 ( 
.A(n_3862),
.Y(n_3895)
);

NAND2xp5_ASAP7_75t_L g3896 ( 
.A(n_3859),
.B(n_198),
.Y(n_3896)
);

OAI22xp5_ASAP7_75t_L g3897 ( 
.A1(n_3851),
.A2(n_1503),
.B1(n_1504),
.B2(n_1485),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_L g3898 ( 
.A(n_3837),
.B(n_198),
.Y(n_3898)
);

NAND2xp5_ASAP7_75t_L g3899 ( 
.A(n_3866),
.B(n_199),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_SL g3900 ( 
.A(n_3852),
.B(n_1514),
.Y(n_3900)
);

AND2x2_ASAP7_75t_L g3901 ( 
.A(n_3835),
.B(n_199),
.Y(n_3901)
);

OAI22xp5_ASAP7_75t_L g3902 ( 
.A1(n_3856),
.A2(n_1521),
.B1(n_1527),
.B2(n_1519),
.Y(n_3902)
);

AOI21xp5_ASAP7_75t_L g3903 ( 
.A1(n_3845),
.A2(n_3840),
.B(n_3849),
.Y(n_3903)
);

INVx1_ASAP7_75t_L g3904 ( 
.A(n_3853),
.Y(n_3904)
);

NAND2xp5_ASAP7_75t_SL g3905 ( 
.A(n_3860),
.B(n_3857),
.Y(n_3905)
);

INVx1_ASAP7_75t_L g3906 ( 
.A(n_3858),
.Y(n_3906)
);

AND2x2_ASAP7_75t_L g3907 ( 
.A(n_3861),
.B(n_200),
.Y(n_3907)
);

NAND2xp33_ASAP7_75t_R g3908 ( 
.A(n_3848),
.B(n_201),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3838),
.Y(n_3909)
);

AND2x2_ASAP7_75t_L g3910 ( 
.A(n_3861),
.B(n_202),
.Y(n_3910)
);

AND2x2_ASAP7_75t_L g3911 ( 
.A(n_3879),
.B(n_202),
.Y(n_3911)
);

NAND2xp5_ASAP7_75t_L g3912 ( 
.A(n_3878),
.B(n_203),
.Y(n_3912)
);

INVx2_ASAP7_75t_SL g3913 ( 
.A(n_3876),
.Y(n_3913)
);

AND2x2_ASAP7_75t_L g3914 ( 
.A(n_3891),
.B(n_203),
.Y(n_3914)
);

NAND2xp5_ASAP7_75t_L g3915 ( 
.A(n_3909),
.B(n_3907),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3875),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_L g3917 ( 
.A(n_3910),
.B(n_204),
.Y(n_3917)
);

INVxp67_ASAP7_75t_SL g3918 ( 
.A(n_3908),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3870),
.Y(n_3919)
);

BUFx3_ASAP7_75t_L g3920 ( 
.A(n_3881),
.Y(n_3920)
);

NAND2xp5_ASAP7_75t_L g3921 ( 
.A(n_3882),
.B(n_204),
.Y(n_3921)
);

AND2x2_ASAP7_75t_L g3922 ( 
.A(n_3901),
.B(n_206),
.Y(n_3922)
);

AND2x2_ASAP7_75t_L g3923 ( 
.A(n_3871),
.B(n_207),
.Y(n_3923)
);

OR2x2_ASAP7_75t_L g3924 ( 
.A(n_3896),
.B(n_207),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3883),
.Y(n_3925)
);

NOR2xp33_ASAP7_75t_L g3926 ( 
.A(n_3892),
.B(n_208),
.Y(n_3926)
);

NAND2xp5_ASAP7_75t_SL g3927 ( 
.A(n_3873),
.B(n_1775),
.Y(n_3927)
);

INVx2_ASAP7_75t_SL g3928 ( 
.A(n_3889),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3886),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3904),
.B(n_208),
.Y(n_3930)
);

AND2x2_ASAP7_75t_L g3931 ( 
.A(n_3872),
.B(n_211),
.Y(n_3931)
);

NAND2xp5_ASAP7_75t_L g3932 ( 
.A(n_3885),
.B(n_211),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_L g3933 ( 
.A(n_3887),
.B(n_212),
.Y(n_3933)
);

NOR2xp33_ASAP7_75t_L g3934 ( 
.A(n_3890),
.B(n_212),
.Y(n_3934)
);

INVx1_ASAP7_75t_SL g3935 ( 
.A(n_3898),
.Y(n_3935)
);

NAND2xp5_ASAP7_75t_L g3936 ( 
.A(n_3874),
.B(n_213),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3888),
.Y(n_3937)
);

OAI221xp5_ASAP7_75t_L g3938 ( 
.A1(n_3903),
.A2(n_1676),
.B1(n_1726),
.B2(n_1674),
.C(n_1670),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_L g3939 ( 
.A(n_3895),
.B(n_213),
.Y(n_3939)
);

AND2x2_ASAP7_75t_L g3940 ( 
.A(n_3877),
.B(n_214),
.Y(n_3940)
);

INVxp67_ASAP7_75t_SL g3941 ( 
.A(n_3899),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3893),
.Y(n_3942)
);

OR2x2_ASAP7_75t_L g3943 ( 
.A(n_3894),
.B(n_215),
.Y(n_3943)
);

NAND3xp33_ASAP7_75t_L g3944 ( 
.A(n_3902),
.B(n_1544),
.C(n_1540),
.Y(n_3944)
);

NAND2xp5_ASAP7_75t_L g3945 ( 
.A(n_3880),
.B(n_215),
.Y(n_3945)
);

NAND2xp5_ASAP7_75t_L g3946 ( 
.A(n_3906),
.B(n_216),
.Y(n_3946)
);

OR2x2_ASAP7_75t_L g3947 ( 
.A(n_3905),
.B(n_218),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_L g3948 ( 
.A(n_3884),
.B(n_218),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_SL g3949 ( 
.A(n_3897),
.B(n_1757),
.Y(n_3949)
);

HB1xp67_ASAP7_75t_L g3950 ( 
.A(n_3900),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3875),
.Y(n_3951)
);

INVxp67_ASAP7_75t_L g3952 ( 
.A(n_3908),
.Y(n_3952)
);

INVxp67_ASAP7_75t_L g3953 ( 
.A(n_3908),
.Y(n_3953)
);

INVxp67_ASAP7_75t_L g3954 ( 
.A(n_3908),
.Y(n_3954)
);

NAND2xp5_ASAP7_75t_L g3955 ( 
.A(n_3878),
.B(n_219),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3878),
.B(n_220),
.Y(n_3956)
);

INVxp67_ASAP7_75t_L g3957 ( 
.A(n_3908),
.Y(n_3957)
);

OR2x2_ASAP7_75t_L g3958 ( 
.A(n_3878),
.B(n_220),
.Y(n_3958)
);

OR2x2_ASAP7_75t_L g3959 ( 
.A(n_3878),
.B(n_221),
.Y(n_3959)
);

NAND2xp5_ASAP7_75t_L g3960 ( 
.A(n_3878),
.B(n_222),
.Y(n_3960)
);

AOI222xp33_ASAP7_75t_L g3961 ( 
.A1(n_3921),
.A2(n_1577),
.B1(n_1552),
.B2(n_1584),
.C1(n_1566),
.C2(n_1547),
.Y(n_3961)
);

NOR3xp33_ASAP7_75t_L g3962 ( 
.A(n_3918),
.B(n_1593),
.C(n_1588),
.Y(n_3962)
);

AO21x1_ASAP7_75t_L g3963 ( 
.A1(n_3926),
.A2(n_223),
.B(n_224),
.Y(n_3963)
);

NOR2xp33_ASAP7_75t_R g3964 ( 
.A(n_3913),
.B(n_3952),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3911),
.Y(n_3965)
);

AND2x2_ASAP7_75t_L g3966 ( 
.A(n_3953),
.B(n_223),
.Y(n_3966)
);

AOI221xp5_ASAP7_75t_L g3967 ( 
.A1(n_3930),
.A2(n_1604),
.B1(n_1606),
.B2(n_1596),
.C(n_1594),
.Y(n_3967)
);

NAND2xp5_ASAP7_75t_SL g3968 ( 
.A(n_3954),
.B(n_1614),
.Y(n_3968)
);

AOI211x1_ASAP7_75t_L g3969 ( 
.A1(n_3915),
.A2(n_228),
.B(n_225),
.C(n_226),
.Y(n_3969)
);

NOR2x1_ASAP7_75t_L g3970 ( 
.A(n_3920),
.B(n_225),
.Y(n_3970)
);

NAND2x1p5_ASAP7_75t_L g3971 ( 
.A(n_3928),
.B(n_226),
.Y(n_3971)
);

NOR2x1_ASAP7_75t_L g3972 ( 
.A(n_3958),
.B(n_228),
.Y(n_3972)
);

NAND2xp5_ASAP7_75t_L g3973 ( 
.A(n_3957),
.B(n_229),
.Y(n_3973)
);

OAI21xp5_ASAP7_75t_SL g3974 ( 
.A1(n_3916),
.A2(n_229),
.B(n_230),
.Y(n_3974)
);

XNOR2x1_ASAP7_75t_L g3975 ( 
.A(n_3947),
.B(n_230),
.Y(n_3975)
);

OAI211xp5_ASAP7_75t_L g3976 ( 
.A1(n_3951),
.A2(n_233),
.B(n_231),
.C(n_232),
.Y(n_3976)
);

NOR2xp33_ASAP7_75t_L g3977 ( 
.A(n_3917),
.B(n_231),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_SL g3978 ( 
.A(n_3959),
.B(n_3922),
.Y(n_3978)
);

AND2x2_ASAP7_75t_L g3979 ( 
.A(n_3914),
.B(n_232),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_L g3980 ( 
.A(n_3934),
.B(n_233),
.Y(n_3980)
);

NOR3x1_ASAP7_75t_L g3981 ( 
.A(n_3946),
.B(n_234),
.C(n_235),
.Y(n_3981)
);

NAND2xp5_ASAP7_75t_L g3982 ( 
.A(n_3923),
.B(n_235),
.Y(n_3982)
);

NAND4xp75_ASAP7_75t_L g3983 ( 
.A(n_3919),
.B(n_238),
.C(n_236),
.D(n_237),
.Y(n_3983)
);

NAND2xp5_ASAP7_75t_SL g3984 ( 
.A(n_3912),
.B(n_3955),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3960),
.Y(n_3985)
);

OR2x6_ASAP7_75t_L g3986 ( 
.A(n_3956),
.B(n_239),
.Y(n_3986)
);

NAND2xp5_ASAP7_75t_L g3987 ( 
.A(n_3935),
.B(n_237),
.Y(n_3987)
);

INVx1_ASAP7_75t_L g3988 ( 
.A(n_3943),
.Y(n_3988)
);

NOR2xp33_ASAP7_75t_L g3989 ( 
.A(n_3924),
.B(n_239),
.Y(n_3989)
);

NAND3xp33_ASAP7_75t_L g3990 ( 
.A(n_3925),
.B(n_1622),
.C(n_1618),
.Y(n_3990)
);

INVx1_ASAP7_75t_L g3991 ( 
.A(n_3931),
.Y(n_3991)
);

NOR3xp33_ASAP7_75t_L g3992 ( 
.A(n_3927),
.B(n_1640),
.C(n_1626),
.Y(n_3992)
);

NOR2xp33_ASAP7_75t_L g3993 ( 
.A(n_3932),
.B(n_240),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_SL g3994 ( 
.A(n_3940),
.B(n_1649),
.Y(n_3994)
);

INVxp67_ASAP7_75t_L g3995 ( 
.A(n_3936),
.Y(n_3995)
);

INVx1_ASAP7_75t_L g3996 ( 
.A(n_3933),
.Y(n_3996)
);

AOI211xp5_ASAP7_75t_L g3997 ( 
.A1(n_3937),
.A2(n_242),
.B(n_240),
.C(n_241),
.Y(n_3997)
);

AND2x2_ASAP7_75t_L g3998 ( 
.A(n_3941),
.B(n_242),
.Y(n_3998)
);

AOI21xp33_ASAP7_75t_L g3999 ( 
.A1(n_3929),
.A2(n_246),
.B(n_245),
.Y(n_3999)
);

AOI221xp5_ASAP7_75t_L g4000 ( 
.A1(n_3942),
.A2(n_1735),
.B1(n_1744),
.B2(n_1669),
.C(n_1668),
.Y(n_4000)
);

NOR3xp33_ASAP7_75t_L g4001 ( 
.A(n_3950),
.B(n_1753),
.C(n_1750),
.Y(n_4001)
);

AND3x4_ASAP7_75t_L g4002 ( 
.A(n_3939),
.B(n_3945),
.C(n_3948),
.Y(n_4002)
);

NAND5xp2_ASAP7_75t_L g4003 ( 
.A(n_3938),
.B(n_3949),
.C(n_3944),
.D(n_247),
.E(n_243),
.Y(n_4003)
);

AND2x2_ASAP7_75t_L g4004 ( 
.A(n_3918),
.B(n_243),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_L g4005 ( 
.A(n_3918),
.B(n_246),
.Y(n_4005)
);

INVx1_ASAP7_75t_L g4006 ( 
.A(n_3918),
.Y(n_4006)
);

AOI21xp33_ASAP7_75t_SL g4007 ( 
.A1(n_3952),
.A2(n_249),
.B(n_248),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_3918),
.Y(n_4008)
);

INVx1_ASAP7_75t_L g4009 ( 
.A(n_3918),
.Y(n_4009)
);

OAI22xp5_ASAP7_75t_L g4010 ( 
.A1(n_3952),
.A2(n_1756),
.B1(n_1773),
.B2(n_1754),
.Y(n_4010)
);

NAND3xp33_ASAP7_75t_L g4011 ( 
.A(n_3952),
.B(n_247),
.C(n_249),
.Y(n_4011)
);

INVx1_ASAP7_75t_L g4012 ( 
.A(n_3918),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_L g4013 ( 
.A(n_3918),
.B(n_250),
.Y(n_4013)
);

INVxp67_ASAP7_75t_SL g4014 ( 
.A(n_3952),
.Y(n_4014)
);

INVx1_ASAP7_75t_L g4015 ( 
.A(n_3918),
.Y(n_4015)
);

NOR3xp33_ASAP7_75t_L g4016 ( 
.A(n_3918),
.B(n_259),
.C(n_250),
.Y(n_4016)
);

OAI21xp5_ASAP7_75t_L g4017 ( 
.A1(n_3952),
.A2(n_251),
.B(n_252),
.Y(n_4017)
);

CKINVDCx20_ASAP7_75t_L g4018 ( 
.A(n_3918),
.Y(n_4018)
);

AND2x2_ASAP7_75t_L g4019 ( 
.A(n_3918),
.B(n_252),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_3918),
.Y(n_4020)
);

NAND2xp5_ASAP7_75t_L g4021 ( 
.A(n_3918),
.B(n_253),
.Y(n_4021)
);

INVxp67_ASAP7_75t_SL g4022 ( 
.A(n_3952),
.Y(n_4022)
);

NAND4xp25_ASAP7_75t_L g4023 ( 
.A(n_3915),
.B(n_255),
.C(n_253),
.D(n_254),
.Y(n_4023)
);

INVx1_ASAP7_75t_L g4024 ( 
.A(n_3918),
.Y(n_4024)
);

NAND2xp5_ASAP7_75t_SL g4025 ( 
.A(n_3952),
.B(n_254),
.Y(n_4025)
);

INVxp67_ASAP7_75t_SL g4026 ( 
.A(n_3952),
.Y(n_4026)
);

OR2x2_ASAP7_75t_L g4027 ( 
.A(n_3918),
.B(n_255),
.Y(n_4027)
);

NOR2xp33_ASAP7_75t_L g4028 ( 
.A(n_3952),
.B(n_256),
.Y(n_4028)
);

NOR2x1_ASAP7_75t_SL g4029 ( 
.A(n_3913),
.B(n_256),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_SL g4030 ( 
.A(n_3952),
.B(n_258),
.Y(n_4030)
);

AOI31xp33_ASAP7_75t_L g4031 ( 
.A1(n_3918),
.A2(n_261),
.A3(n_262),
.B(n_260),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_3918),
.Y(n_4032)
);

AOI21xp5_ASAP7_75t_L g4033 ( 
.A1(n_3918),
.A2(n_259),
.B(n_261),
.Y(n_4033)
);

AOI22xp5_ASAP7_75t_L g4034 ( 
.A1(n_3913),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.Y(n_4034)
);

NAND2xp5_ASAP7_75t_L g4035 ( 
.A(n_3918),
.B(n_265),
.Y(n_4035)
);

AND2x2_ASAP7_75t_L g4036 ( 
.A(n_3918),
.B(n_265),
.Y(n_4036)
);

INVxp67_ASAP7_75t_L g4037 ( 
.A(n_3918),
.Y(n_4037)
);

AOI211xp5_ASAP7_75t_L g4038 ( 
.A1(n_3952),
.A2(n_268),
.B(n_266),
.C(n_267),
.Y(n_4038)
);

NOR3xp33_ASAP7_75t_L g4039 ( 
.A(n_3918),
.B(n_276),
.C(n_267),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_SL g4040 ( 
.A(n_3952),
.B(n_269),
.Y(n_4040)
);

NOR3xp33_ASAP7_75t_L g4041 ( 
.A(n_3918),
.B(n_278),
.C(n_269),
.Y(n_4041)
);

NOR2xp67_ASAP7_75t_L g4042 ( 
.A(n_3952),
.B(n_270),
.Y(n_4042)
);

AOI211xp5_ASAP7_75t_L g4043 ( 
.A1(n_3952),
.A2(n_273),
.B(n_271),
.C(n_272),
.Y(n_4043)
);

AOI221x1_ASAP7_75t_L g4044 ( 
.A1(n_4016),
.A2(n_273),
.B1(n_271),
.B2(n_272),
.C(n_274),
.Y(n_4044)
);

NOR2xp33_ASAP7_75t_L g4045 ( 
.A(n_4037),
.B(n_274),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_4029),
.Y(n_4046)
);

OAI211xp5_ASAP7_75t_L g4047 ( 
.A1(n_3964),
.A2(n_286),
.B(n_294),
.C(n_275),
.Y(n_4047)
);

NOR3xp33_ASAP7_75t_L g4048 ( 
.A(n_4006),
.B(n_275),
.C(n_277),
.Y(n_4048)
);

INVx2_ASAP7_75t_L g4049 ( 
.A(n_3971),
.Y(n_4049)
);

AOI221xp5_ASAP7_75t_L g4050 ( 
.A1(n_4008),
.A2(n_280),
.B1(n_278),
.B2(n_279),
.C(n_281),
.Y(n_4050)
);

NAND4xp75_ASAP7_75t_L g4051 ( 
.A(n_3970),
.B(n_281),
.C(n_279),
.D(n_280),
.Y(n_4051)
);

INVx2_ASAP7_75t_L g4052 ( 
.A(n_4018),
.Y(n_4052)
);

NAND4xp25_ASAP7_75t_L g4053 ( 
.A(n_4009),
.B(n_287),
.C(n_282),
.D(n_285),
.Y(n_4053)
);

OAI211xp5_ASAP7_75t_L g4054 ( 
.A1(n_3969),
.A2(n_4014),
.B(n_4026),
.C(n_4022),
.Y(n_4054)
);

INVxp67_ASAP7_75t_L g4055 ( 
.A(n_3972),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_L g4056 ( 
.A(n_4042),
.B(n_285),
.Y(n_4056)
);

AOI221xp5_ASAP7_75t_L g4057 ( 
.A1(n_4012),
.A2(n_289),
.B1(n_287),
.B2(n_288),
.C(n_290),
.Y(n_4057)
);

OAI321xp33_ASAP7_75t_L g4058 ( 
.A1(n_4015),
.A2(n_290),
.A3(n_292),
.B1(n_288),
.B2(n_289),
.C(n_291),
.Y(n_4058)
);

INVx1_ASAP7_75t_L g4059 ( 
.A(n_4004),
.Y(n_4059)
);

AOI221xp5_ASAP7_75t_L g4060 ( 
.A1(n_4020),
.A2(n_295),
.B1(n_292),
.B2(n_293),
.C(n_296),
.Y(n_4060)
);

AOI21xp5_ASAP7_75t_L g4061 ( 
.A1(n_3978),
.A2(n_293),
.B(n_295),
.Y(n_4061)
);

AOI31xp33_ASAP7_75t_L g4062 ( 
.A1(n_3963),
.A2(n_300),
.A3(n_297),
.B(n_298),
.Y(n_4062)
);

OAI21xp33_ASAP7_75t_L g4063 ( 
.A1(n_4024),
.A2(n_298),
.B(n_301),
.Y(n_4063)
);

NOR2xp33_ASAP7_75t_L g4064 ( 
.A(n_4032),
.B(n_301),
.Y(n_4064)
);

O2A1O1Ixp33_ASAP7_75t_L g4065 ( 
.A1(n_4031),
.A2(n_304),
.B(n_302),
.C(n_303),
.Y(n_4065)
);

AND2x2_ASAP7_75t_SL g4066 ( 
.A(n_3981),
.B(n_4019),
.Y(n_4066)
);

AOI21x1_ASAP7_75t_L g4067 ( 
.A1(n_4033),
.A2(n_311),
.B(n_303),
.Y(n_4067)
);

AOI221xp5_ASAP7_75t_L g4068 ( 
.A1(n_4028),
.A2(n_3965),
.B1(n_4036),
.B2(n_4041),
.C(n_4039),
.Y(n_4068)
);

AOI221xp5_ASAP7_75t_L g4069 ( 
.A1(n_4005),
.A2(n_306),
.B1(n_304),
.B2(n_305),
.C(n_307),
.Y(n_4069)
);

XNOR2x1_ASAP7_75t_L g4070 ( 
.A(n_3975),
.B(n_305),
.Y(n_4070)
);

NOR4xp25_ASAP7_75t_L g4071 ( 
.A(n_3984),
.B(n_3991),
.C(n_3988),
.D(n_4013),
.Y(n_4071)
);

NOR5xp2_ASAP7_75t_L g4072 ( 
.A(n_4011),
.B(n_309),
.C(n_307),
.D(n_308),
.E(n_310),
.Y(n_4072)
);

AOI21xp5_ASAP7_75t_L g4073 ( 
.A1(n_4025),
.A2(n_309),
.B(n_311),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_4027),
.Y(n_4074)
);

AOI221xp5_ASAP7_75t_L g4075 ( 
.A1(n_4021),
.A2(n_315),
.B1(n_312),
.B2(n_314),
.C(n_316),
.Y(n_4075)
);

AOI21xp33_ASAP7_75t_L g4076 ( 
.A1(n_4035),
.A2(n_312),
.B(n_315),
.Y(n_4076)
);

INVx1_ASAP7_75t_L g4077 ( 
.A(n_3966),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_3979),
.Y(n_4078)
);

OAI21xp5_ASAP7_75t_SL g4079 ( 
.A1(n_3973),
.A2(n_316),
.B(n_317),
.Y(n_4079)
);

OAI321xp33_ASAP7_75t_L g4080 ( 
.A1(n_3995),
.A2(n_319),
.A3(n_322),
.B1(n_317),
.B2(n_318),
.C(n_321),
.Y(n_4080)
);

AOI22xp5_ASAP7_75t_L g4081 ( 
.A1(n_4002),
.A2(n_321),
.B1(n_318),
.B2(n_319),
.Y(n_4081)
);

AOI222xp33_ASAP7_75t_L g4082 ( 
.A1(n_3985),
.A2(n_324),
.B1(n_326),
.B2(n_322),
.C1(n_323),
.C2(n_325),
.Y(n_4082)
);

AOI221xp5_ASAP7_75t_L g4083 ( 
.A1(n_4007),
.A2(n_327),
.B1(n_323),
.B2(n_325),
.C(n_328),
.Y(n_4083)
);

NAND2xp5_ASAP7_75t_L g4084 ( 
.A(n_3998),
.B(n_329),
.Y(n_4084)
);

AOI221xp5_ASAP7_75t_L g4085 ( 
.A1(n_4003),
.A2(n_333),
.B1(n_330),
.B2(n_332),
.C(n_334),
.Y(n_4085)
);

AOI222xp33_ASAP7_75t_L g4086 ( 
.A1(n_3996),
.A2(n_335),
.B1(n_337),
.B2(n_332),
.C1(n_334),
.C2(n_336),
.Y(n_4086)
);

AOI221xp5_ASAP7_75t_L g4087 ( 
.A1(n_3962),
.A2(n_338),
.B1(n_336),
.B2(n_337),
.C(n_339),
.Y(n_4087)
);

AOI321xp33_ASAP7_75t_L g4088 ( 
.A1(n_4030),
.A2(n_341),
.A3(n_345),
.B1(n_338),
.B2(n_340),
.C(n_344),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_3983),
.Y(n_4089)
);

NAND3x1_ASAP7_75t_L g4090 ( 
.A(n_4017),
.B(n_341),
.C(n_344),
.Y(n_4090)
);

AOI211xp5_ASAP7_75t_L g4091 ( 
.A1(n_4040),
.A2(n_347),
.B(n_345),
.C(n_346),
.Y(n_4091)
);

NAND3xp33_ASAP7_75t_L g4092 ( 
.A(n_4038),
.B(n_347),
.C(n_349),
.Y(n_4092)
);

AOI32xp33_ASAP7_75t_L g4093 ( 
.A1(n_3989),
.A2(n_3977),
.A3(n_3987),
.B1(n_4043),
.B2(n_3993),
.Y(n_4093)
);

AOI32xp33_ASAP7_75t_L g4094 ( 
.A1(n_4001),
.A2(n_3992),
.A3(n_3997),
.B1(n_3980),
.B2(n_3982),
.Y(n_4094)
);

NAND2xp5_ASAP7_75t_L g4095 ( 
.A(n_4034),
.B(n_350),
.Y(n_4095)
);

OAI221xp5_ASAP7_75t_L g4096 ( 
.A1(n_3974),
.A2(n_353),
.B1(n_351),
.B2(n_352),
.C(n_354),
.Y(n_4096)
);

AOI22xp5_ASAP7_75t_L g4097 ( 
.A1(n_4023),
.A2(n_353),
.B1(n_351),
.B2(n_352),
.Y(n_4097)
);

AOI221xp5_ASAP7_75t_L g4098 ( 
.A1(n_3999),
.A2(n_358),
.B1(n_355),
.B2(n_357),
.C(n_359),
.Y(n_4098)
);

NOR2xp33_ASAP7_75t_R g4099 ( 
.A(n_3976),
.B(n_3986),
.Y(n_4099)
);

AOI211xp5_ASAP7_75t_L g4100 ( 
.A1(n_3994),
.A2(n_358),
.B(n_355),
.C(n_357),
.Y(n_4100)
);

AOI221xp5_ASAP7_75t_L g4101 ( 
.A1(n_3968),
.A2(n_361),
.B1(n_359),
.B2(n_360),
.C(n_362),
.Y(n_4101)
);

AOI33xp33_ASAP7_75t_L g4102 ( 
.A1(n_3967),
.A2(n_364),
.A3(n_366),
.B1(n_360),
.B2(n_363),
.B3(n_365),
.Y(n_4102)
);

OAI221xp5_ASAP7_75t_L g4103 ( 
.A1(n_3986),
.A2(n_365),
.B1(n_363),
.B2(n_364),
.C(n_366),
.Y(n_4103)
);

NAND2xp33_ASAP7_75t_R g4104 ( 
.A(n_3961),
.B(n_367),
.Y(n_4104)
);

NOR2xp33_ASAP7_75t_L g4105 ( 
.A(n_3990),
.B(n_367),
.Y(n_4105)
);

AOI21xp5_ASAP7_75t_L g4106 ( 
.A1(n_4010),
.A2(n_368),
.B(n_370),
.Y(n_4106)
);

AOI221xp5_ASAP7_75t_L g4107 ( 
.A1(n_4000),
.A2(n_372),
.B1(n_370),
.B2(n_371),
.C(n_373),
.Y(n_4107)
);

AOI22xp5_ASAP7_75t_L g4108 ( 
.A1(n_4014),
.A2(n_374),
.B1(n_372),
.B2(n_373),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_L g4109 ( 
.A(n_4042),
.B(n_374),
.Y(n_4109)
);

AOI22xp5_ASAP7_75t_L g4110 ( 
.A1(n_4014),
.A2(n_377),
.B1(n_375),
.B2(n_376),
.Y(n_4110)
);

XNOR2xp5_ASAP7_75t_L g4111 ( 
.A(n_3975),
.B(n_375),
.Y(n_4111)
);

AOI31xp33_ASAP7_75t_L g4112 ( 
.A1(n_3963),
.A2(n_378),
.A3(n_376),
.B(n_377),
.Y(n_4112)
);

AOI22xp33_ASAP7_75t_L g4113 ( 
.A1(n_4018),
.A2(n_381),
.B1(n_378),
.B2(n_379),
.Y(n_4113)
);

AOI321xp33_ASAP7_75t_L g4114 ( 
.A1(n_4014),
.A2(n_382),
.A3(n_384),
.B1(n_379),
.B2(n_381),
.C(n_383),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_L g4115 ( 
.A(n_4042),
.B(n_382),
.Y(n_4115)
);

NAND2xp33_ASAP7_75t_R g4116 ( 
.A(n_3964),
.B(n_383),
.Y(n_4116)
);

AOI221xp5_ASAP7_75t_L g4117 ( 
.A1(n_4037),
.A2(n_387),
.B1(n_385),
.B2(n_386),
.C(n_388),
.Y(n_4117)
);

AOI221x1_ASAP7_75t_L g4118 ( 
.A1(n_4016),
.A2(n_387),
.B1(n_385),
.B2(n_386),
.C(n_389),
.Y(n_4118)
);

INVx2_ASAP7_75t_L g4119 ( 
.A(n_4029),
.Y(n_4119)
);

OAI21xp5_ASAP7_75t_SL g4120 ( 
.A1(n_4037),
.A2(n_389),
.B(n_391),
.Y(n_4120)
);

AOI22xp5_ASAP7_75t_L g4121 ( 
.A1(n_4014),
.A2(n_395),
.B1(n_393),
.B2(n_394),
.Y(n_4121)
);

NOR3xp33_ASAP7_75t_SL g4122 ( 
.A(n_3978),
.B(n_395),
.C(n_396),
.Y(n_4122)
);

AOI311xp33_ASAP7_75t_L g4123 ( 
.A1(n_4006),
.A2(n_398),
.A3(n_396),
.B(n_397),
.C(n_399),
.Y(n_4123)
);

OAI221xp5_ASAP7_75t_SL g4124 ( 
.A1(n_4037),
.A2(n_400),
.B1(n_397),
.B2(n_398),
.C(n_401),
.Y(n_4124)
);

AOI21xp33_ASAP7_75t_L g4125 ( 
.A1(n_4037),
.A2(n_400),
.B(n_402),
.Y(n_4125)
);

INVxp67_ASAP7_75t_L g4126 ( 
.A(n_4029),
.Y(n_4126)
);

NOR3xp33_ASAP7_75t_L g4127 ( 
.A(n_4054),
.B(n_4126),
.C(n_4052),
.Y(n_4127)
);

AOI221xp5_ASAP7_75t_L g4128 ( 
.A1(n_4062),
.A2(n_405),
.B1(n_402),
.B2(n_404),
.C(n_406),
.Y(n_4128)
);

OAI211xp5_ASAP7_75t_L g4129 ( 
.A1(n_4055),
.A2(n_406),
.B(n_404),
.C(n_405),
.Y(n_4129)
);

AND2x2_ASAP7_75t_L g4130 ( 
.A(n_4066),
.B(n_407),
.Y(n_4130)
);

OAI21xp33_ASAP7_75t_L g4131 ( 
.A1(n_4089),
.A2(n_408),
.B(n_409),
.Y(n_4131)
);

AOI222xp33_ASAP7_75t_L g4132 ( 
.A1(n_4046),
.A2(n_411),
.B1(n_414),
.B2(n_408),
.C1(n_410),
.C2(n_413),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_4119),
.Y(n_4133)
);

OAI221xp5_ASAP7_75t_L g4134 ( 
.A1(n_4068),
.A2(n_413),
.B1(n_410),
.B2(n_411),
.C(n_415),
.Y(n_4134)
);

OAI211xp5_ASAP7_75t_SL g4135 ( 
.A1(n_4093),
.A2(n_417),
.B(n_415),
.C(n_416),
.Y(n_4135)
);

AOI21xp5_ASAP7_75t_L g4136 ( 
.A1(n_4056),
.A2(n_416),
.B(n_418),
.Y(n_4136)
);

AOI21xp5_ASAP7_75t_L g4137 ( 
.A1(n_4109),
.A2(n_418),
.B(n_419),
.Y(n_4137)
);

AOI221xp5_ASAP7_75t_L g4138 ( 
.A1(n_4112),
.A2(n_422),
.B1(n_420),
.B2(n_421),
.C(n_423),
.Y(n_4138)
);

AOI222xp33_ASAP7_75t_L g4139 ( 
.A1(n_4059),
.A2(n_426),
.B1(n_428),
.B2(n_420),
.C1(n_425),
.C2(n_427),
.Y(n_4139)
);

INVx1_ASAP7_75t_L g4140 ( 
.A(n_4115),
.Y(n_4140)
);

AOI211xp5_ASAP7_75t_L g4141 ( 
.A1(n_4071),
.A2(n_431),
.B(n_429),
.C(n_430),
.Y(n_4141)
);

AOI22xp33_ASAP7_75t_SL g4142 ( 
.A1(n_4099),
.A2(n_4049),
.B1(n_4074),
.B2(n_4078),
.Y(n_4142)
);

NAND4xp25_ASAP7_75t_L g4143 ( 
.A(n_4085),
.B(n_431),
.C(n_429),
.D(n_430),
.Y(n_4143)
);

NOR2xp33_ASAP7_75t_SL g4144 ( 
.A(n_4051),
.B(n_433),
.Y(n_4144)
);

BUFx2_ASAP7_75t_L g4145 ( 
.A(n_4090),
.Y(n_4145)
);

OR2x2_ASAP7_75t_L g4146 ( 
.A(n_4084),
.B(n_4077),
.Y(n_4146)
);

AOI21xp5_ASAP7_75t_L g4147 ( 
.A1(n_4065),
.A2(n_433),
.B(n_434),
.Y(n_4147)
);

OAI221xp5_ASAP7_75t_L g4148 ( 
.A1(n_4116),
.A2(n_436),
.B1(n_434),
.B2(n_435),
.C(n_437),
.Y(n_4148)
);

O2A1O1Ixp33_ASAP7_75t_L g4149 ( 
.A1(n_4058),
.A2(n_438),
.B(n_435),
.C(n_437),
.Y(n_4149)
);

OAI21xp33_ASAP7_75t_L g4150 ( 
.A1(n_4070),
.A2(n_438),
.B(n_440),
.Y(n_4150)
);

AOI221xp5_ASAP7_75t_SL g4151 ( 
.A1(n_4061),
.A2(n_442),
.B1(n_440),
.B2(n_441),
.C(n_443),
.Y(n_4151)
);

INVx1_ASAP7_75t_L g4152 ( 
.A(n_4111),
.Y(n_4152)
);

AOI211xp5_ASAP7_75t_L g4153 ( 
.A1(n_4092),
.A2(n_445),
.B(n_442),
.C(n_444),
.Y(n_4153)
);

NAND5xp2_ASAP7_75t_SL g4154 ( 
.A(n_4088),
.B(n_4047),
.C(n_4114),
.D(n_4097),
.E(n_4096),
.Y(n_4154)
);

AOI211xp5_ASAP7_75t_L g4155 ( 
.A1(n_4045),
.A2(n_448),
.B(n_445),
.C(n_447),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_L g4156 ( 
.A(n_4113),
.B(n_447),
.Y(n_4156)
);

NAND3xp33_ASAP7_75t_L g4157 ( 
.A(n_4122),
.B(n_4118),
.C(n_4044),
.Y(n_4157)
);

AOI22xp5_ASAP7_75t_L g4158 ( 
.A1(n_4064),
.A2(n_450),
.B1(n_448),
.B2(n_449),
.Y(n_4158)
);

OAI211xp5_ASAP7_75t_L g4159 ( 
.A1(n_4094),
.A2(n_454),
.B(n_451),
.C(n_453),
.Y(n_4159)
);

AOI221xp5_ASAP7_75t_L g4160 ( 
.A1(n_4080),
.A2(n_455),
.B1(n_451),
.B2(n_454),
.C(n_456),
.Y(n_4160)
);

AOI211xp5_ASAP7_75t_L g4161 ( 
.A1(n_4120),
.A2(n_459),
.B(n_456),
.C(n_457),
.Y(n_4161)
);

OAI221xp5_ASAP7_75t_SL g4162 ( 
.A1(n_4079),
.A2(n_462),
.B1(n_460),
.B2(n_461),
.C(n_463),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_4067),
.Y(n_4163)
);

NOR3xp33_ASAP7_75t_SL g4164 ( 
.A(n_4104),
.B(n_460),
.C(n_461),
.Y(n_4164)
);

AOI211xp5_ASAP7_75t_L g4165 ( 
.A1(n_4124),
.A2(n_4076),
.B(n_4125),
.C(n_4073),
.Y(n_4165)
);

OAI21xp5_ASAP7_75t_L g4166 ( 
.A1(n_4106),
.A2(n_465),
.B(n_464),
.Y(n_4166)
);

AOI222xp33_ASAP7_75t_L g4167 ( 
.A1(n_4098),
.A2(n_465),
.B1(n_467),
.B2(n_462),
.C1(n_464),
.C2(n_466),
.Y(n_4167)
);

OAI221xp5_ASAP7_75t_L g4168 ( 
.A1(n_4083),
.A2(n_468),
.B1(n_466),
.B2(n_467),
.C(n_469),
.Y(n_4168)
);

AOI211xp5_ASAP7_75t_L g4169 ( 
.A1(n_4063),
.A2(n_470),
.B(n_468),
.C(n_469),
.Y(n_4169)
);

CKINVDCx6p67_ASAP7_75t_R g4170 ( 
.A(n_4095),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_4081),
.Y(n_4171)
);

OAI211xp5_ASAP7_75t_SL g4172 ( 
.A1(n_4091),
.A2(n_474),
.B(n_472),
.C(n_473),
.Y(n_4172)
);

AOI211xp5_ASAP7_75t_L g4173 ( 
.A1(n_4053),
.A2(n_475),
.B(n_473),
.C(n_474),
.Y(n_4173)
);

INVx2_ASAP7_75t_L g4174 ( 
.A(n_4103),
.Y(n_4174)
);

CKINVDCx16_ASAP7_75t_R g4175 ( 
.A(n_4108),
.Y(n_4175)
);

AOI221xp5_ASAP7_75t_L g4176 ( 
.A1(n_4048),
.A2(n_477),
.B1(n_475),
.B2(n_476),
.C(n_478),
.Y(n_4176)
);

OAI222xp33_ASAP7_75t_L g4177 ( 
.A1(n_4110),
.A2(n_481),
.B1(n_483),
.B2(n_476),
.C1(n_477),
.C2(n_482),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_4102),
.Y(n_4178)
);

OAI21xp5_ASAP7_75t_L g4179 ( 
.A1(n_4105),
.A2(n_484),
.B(n_483),
.Y(n_4179)
);

AOI22x1_ASAP7_75t_L g4180 ( 
.A1(n_4086),
.A2(n_485),
.B1(n_481),
.B2(n_484),
.Y(n_4180)
);

OAI211xp5_ASAP7_75t_L g4181 ( 
.A1(n_4123),
.A2(n_488),
.B(n_486),
.C(n_487),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_4121),
.Y(n_4182)
);

HB1xp67_ASAP7_75t_L g4183 ( 
.A(n_4100),
.Y(n_4183)
);

NAND2xp5_ASAP7_75t_L g4184 ( 
.A(n_4082),
.B(n_486),
.Y(n_4184)
);

AO22x2_ASAP7_75t_L g4185 ( 
.A1(n_4072),
.A2(n_490),
.B1(n_487),
.B2(n_489),
.Y(n_4185)
);

AOI221x1_ASAP7_75t_L g4186 ( 
.A1(n_4107),
.A2(n_492),
.B1(n_490),
.B2(n_491),
.C(n_493),
.Y(n_4186)
);

OAI211xp5_ASAP7_75t_SL g4187 ( 
.A1(n_4087),
.A2(n_496),
.B(n_492),
.C(n_494),
.Y(n_4187)
);

NAND2xp5_ASAP7_75t_L g4188 ( 
.A(n_4050),
.B(n_494),
.Y(n_4188)
);

NAND4xp25_ASAP7_75t_L g4189 ( 
.A(n_4069),
.B(n_499),
.C(n_496),
.D(n_498),
.Y(n_4189)
);

A2O1A1Ixp33_ASAP7_75t_SL g4190 ( 
.A1(n_4057),
.A2(n_502),
.B(n_500),
.C(n_501),
.Y(n_4190)
);

AOI211xp5_ASAP7_75t_SL g4191 ( 
.A1(n_4101),
.A2(n_505),
.B(n_500),
.C(n_504),
.Y(n_4191)
);

OAI211xp5_ASAP7_75t_L g4192 ( 
.A1(n_4117),
.A2(n_506),
.B(n_504),
.C(n_505),
.Y(n_4192)
);

HB1xp67_ASAP7_75t_L g4193 ( 
.A(n_4060),
.Y(n_4193)
);

OAI22xp5_ASAP7_75t_L g4194 ( 
.A1(n_4075),
.A2(n_508),
.B1(n_506),
.B2(n_507),
.Y(n_4194)
);

NOR3xp33_ASAP7_75t_L g4195 ( 
.A(n_4054),
.B(n_509),
.C(n_508),
.Y(n_4195)
);

INVxp67_ASAP7_75t_SL g4196 ( 
.A(n_4072),
.Y(n_4196)
);

AOI22xp5_ASAP7_75t_L g4197 ( 
.A1(n_4052),
.A2(n_510),
.B1(n_507),
.B2(n_509),
.Y(n_4197)
);

AOI222xp33_ASAP7_75t_L g4198 ( 
.A1(n_4126),
.A2(n_512),
.B1(n_514),
.B2(n_510),
.C1(n_511),
.C2(n_513),
.Y(n_4198)
);

AOI211x1_ASAP7_75t_SL g4199 ( 
.A1(n_4052),
.A2(n_515),
.B(n_511),
.C(n_513),
.Y(n_4199)
);

AOI211xp5_ASAP7_75t_L g4200 ( 
.A1(n_4054),
.A2(n_518),
.B(n_515),
.C(n_517),
.Y(n_4200)
);

AOI221xp5_ASAP7_75t_L g4201 ( 
.A1(n_4062),
.A2(n_521),
.B1(n_519),
.B2(n_520),
.C(n_522),
.Y(n_4201)
);

AND2x2_ASAP7_75t_L g4202 ( 
.A(n_4066),
.B(n_519),
.Y(n_4202)
);

O2A1O1Ixp33_ASAP7_75t_L g4203 ( 
.A1(n_4062),
.A2(n_524),
.B(n_520),
.C(n_521),
.Y(n_4203)
);

INVx2_ASAP7_75t_L g4204 ( 
.A(n_4119),
.Y(n_4204)
);

AO22x1_ASAP7_75t_SL g4205 ( 
.A1(n_4046),
.A2(n_526),
.B1(n_524),
.B2(n_525),
.Y(n_4205)
);

AOI221xp5_ASAP7_75t_L g4206 ( 
.A1(n_4062),
.A2(n_527),
.B1(n_525),
.B2(n_526),
.C(n_528),
.Y(n_4206)
);

NAND3xp33_ASAP7_75t_L g4207 ( 
.A(n_4122),
.B(n_527),
.C(n_528),
.Y(n_4207)
);

AOI221xp5_ASAP7_75t_L g4208 ( 
.A1(n_4062),
.A2(n_533),
.B1(n_530),
.B2(n_532),
.C(n_534),
.Y(n_4208)
);

OAI211xp5_ASAP7_75t_L g4209 ( 
.A1(n_4126),
.A2(n_535),
.B(n_532),
.C(n_534),
.Y(n_4209)
);

NOR4xp25_ASAP7_75t_L g4210 ( 
.A(n_4054),
.B(n_537),
.C(n_535),
.D(n_536),
.Y(n_4210)
);

NAND4xp25_ASAP7_75t_L g4211 ( 
.A(n_4068),
.B(n_540),
.C(n_538),
.D(n_539),
.Y(n_4211)
);

AND2x2_ASAP7_75t_L g4212 ( 
.A(n_4130),
.B(n_4202),
.Y(n_4212)
);

AOI22xp5_ASAP7_75t_L g4213 ( 
.A1(n_4127),
.A2(n_540),
.B1(n_538),
.B2(n_539),
.Y(n_4213)
);

INVx1_ASAP7_75t_L g4214 ( 
.A(n_4205),
.Y(n_4214)
);

OAI22xp5_ASAP7_75t_L g4215 ( 
.A1(n_4142),
.A2(n_543),
.B1(n_541),
.B2(n_542),
.Y(n_4215)
);

OAI32xp33_ASAP7_75t_L g4216 ( 
.A1(n_4199),
.A2(n_544),
.A3(n_541),
.B1(n_542),
.B2(n_546),
.Y(n_4216)
);

NOR2x1p5_ASAP7_75t_L g4217 ( 
.A(n_4196),
.B(n_547),
.Y(n_4217)
);

OAI22xp33_ASAP7_75t_L g4218 ( 
.A1(n_4144),
.A2(n_549),
.B1(n_547),
.B2(n_548),
.Y(n_4218)
);

INVxp67_ASAP7_75t_SL g4219 ( 
.A(n_4157),
.Y(n_4219)
);

AND2x2_ASAP7_75t_L g4220 ( 
.A(n_4204),
.B(n_550),
.Y(n_4220)
);

AND2x2_ASAP7_75t_L g4221 ( 
.A(n_4164),
.B(n_4133),
.Y(n_4221)
);

OAI22xp5_ASAP7_75t_L g4222 ( 
.A1(n_4207),
.A2(n_553),
.B1(n_550),
.B2(n_552),
.Y(n_4222)
);

AND2x2_ASAP7_75t_L g4223 ( 
.A(n_4145),
.B(n_552),
.Y(n_4223)
);

NAND2xp5_ASAP7_75t_L g4224 ( 
.A(n_4210),
.B(n_553),
.Y(n_4224)
);

NAND3x1_ASAP7_75t_SL g4225 ( 
.A(n_4128),
.B(n_554),
.C(n_555),
.Y(n_4225)
);

INVxp67_ASAP7_75t_L g4226 ( 
.A(n_4185),
.Y(n_4226)
);

OR2x2_ASAP7_75t_L g4227 ( 
.A(n_4211),
.B(n_4143),
.Y(n_4227)
);

INVxp67_ASAP7_75t_L g4228 ( 
.A(n_4185),
.Y(n_4228)
);

HB1xp67_ASAP7_75t_L g4229 ( 
.A(n_4163),
.Y(n_4229)
);

NAND3xp33_ASAP7_75t_SL g4230 ( 
.A(n_4141),
.B(n_554),
.C(n_555),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_4203),
.Y(n_4231)
);

AOI22xp33_ASAP7_75t_L g4232 ( 
.A1(n_4195),
.A2(n_558),
.B1(n_556),
.B2(n_557),
.Y(n_4232)
);

OAI322xp33_ASAP7_75t_L g4233 ( 
.A1(n_4178),
.A2(n_566),
.A3(n_565),
.B1(n_562),
.B2(n_559),
.C1(n_561),
.C2(n_564),
.Y(n_4233)
);

AND2x4_ASAP7_75t_L g4234 ( 
.A(n_4152),
.B(n_559),
.Y(n_4234)
);

NOR3xp33_ASAP7_75t_L g4235 ( 
.A(n_4175),
.B(n_561),
.C(n_562),
.Y(n_4235)
);

NOR2xp33_ASAP7_75t_L g4236 ( 
.A(n_4148),
.B(n_4162),
.Y(n_4236)
);

NAND2xp5_ASAP7_75t_SL g4237 ( 
.A(n_4138),
.B(n_564),
.Y(n_4237)
);

NAND2x1p5_ASAP7_75t_L g4238 ( 
.A(n_4146),
.B(n_567),
.Y(n_4238)
);

OAI221xp5_ASAP7_75t_L g4239 ( 
.A1(n_4200),
.A2(n_568),
.B1(n_565),
.B2(n_567),
.C(n_569),
.Y(n_4239)
);

A2O1A1Ixp33_ASAP7_75t_SL g4240 ( 
.A1(n_4140),
.A2(n_570),
.B(n_568),
.C(n_569),
.Y(n_4240)
);

NAND2xp5_ASAP7_75t_SL g4241 ( 
.A(n_4201),
.B(n_570),
.Y(n_4241)
);

NOR3xp33_ASAP7_75t_L g4242 ( 
.A(n_4150),
.B(n_571),
.C(n_572),
.Y(n_4242)
);

NOR3xp33_ASAP7_75t_L g4243 ( 
.A(n_4134),
.B(n_573),
.C(n_574),
.Y(n_4243)
);

NOR2xp33_ASAP7_75t_SL g4244 ( 
.A(n_4177),
.B(n_575),
.Y(n_4244)
);

AND2x4_ASAP7_75t_L g4245 ( 
.A(n_4171),
.B(n_573),
.Y(n_4245)
);

AOI22xp5_ASAP7_75t_L g4246 ( 
.A1(n_4181),
.A2(n_578),
.B1(n_576),
.B2(n_577),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_4180),
.Y(n_4247)
);

O2A1O1Ixp33_ASAP7_75t_L g4248 ( 
.A1(n_4190),
.A2(n_580),
.B(n_577),
.C(n_578),
.Y(n_4248)
);

AOI21xp5_ASAP7_75t_L g4249 ( 
.A1(n_4136),
.A2(n_580),
.B(n_581),
.Y(n_4249)
);

HB1xp67_ASAP7_75t_L g4250 ( 
.A(n_4166),
.Y(n_4250)
);

AOI221xp5_ASAP7_75t_L g4251 ( 
.A1(n_4154),
.A2(n_583),
.B1(n_581),
.B2(n_582),
.C(n_584),
.Y(n_4251)
);

OAI221xp5_ASAP7_75t_L g4252 ( 
.A1(n_4160),
.A2(n_587),
.B1(n_582),
.B2(n_586),
.C(n_588),
.Y(n_4252)
);

NAND2xp5_ASAP7_75t_L g4253 ( 
.A(n_4198),
.B(n_588),
.Y(n_4253)
);

NAND2x1p5_ASAP7_75t_L g4254 ( 
.A(n_4182),
.B(n_591),
.Y(n_4254)
);

AOI222xp33_ASAP7_75t_L g4255 ( 
.A1(n_4193),
.A2(n_4183),
.B1(n_4174),
.B2(n_4184),
.C1(n_4208),
.C2(n_4206),
.Y(n_4255)
);

AND2x4_ASAP7_75t_L g4256 ( 
.A(n_4179),
.B(n_590),
.Y(n_4256)
);

NOR3xp33_ASAP7_75t_L g4257 ( 
.A(n_4188),
.B(n_591),
.C(n_593),
.Y(n_4257)
);

OAI21xp33_ASAP7_75t_L g4258 ( 
.A1(n_4189),
.A2(n_593),
.B(n_594),
.Y(n_4258)
);

OAI221xp5_ASAP7_75t_L g4259 ( 
.A1(n_4151),
.A2(n_596),
.B1(n_594),
.B2(n_595),
.C(n_597),
.Y(n_4259)
);

OAI22xp33_ASAP7_75t_L g4260 ( 
.A1(n_4191),
.A2(n_598),
.B1(n_596),
.B2(n_597),
.Y(n_4260)
);

NAND3xp33_ASAP7_75t_L g4261 ( 
.A(n_4153),
.B(n_598),
.C(n_599),
.Y(n_4261)
);

NAND2xp5_ASAP7_75t_SL g4262 ( 
.A(n_4132),
.B(n_4161),
.Y(n_4262)
);

AND2x2_ASAP7_75t_L g4263 ( 
.A(n_4170),
.B(n_600),
.Y(n_4263)
);

INVx1_ASAP7_75t_SL g4264 ( 
.A(n_4156),
.Y(n_4264)
);

NOR3xp33_ASAP7_75t_L g4265 ( 
.A(n_4168),
.B(n_600),
.C(n_602),
.Y(n_4265)
);

NAND2xp5_ASAP7_75t_L g4266 ( 
.A(n_4147),
.B(n_604),
.Y(n_4266)
);

O2A1O1Ixp33_ASAP7_75t_L g4267 ( 
.A1(n_4135),
.A2(n_606),
.B(n_604),
.C(n_605),
.Y(n_4267)
);

NOR2x1_ASAP7_75t_L g4268 ( 
.A(n_4209),
.B(n_605),
.Y(n_4268)
);

NOR2x1p5_ASAP7_75t_L g4269 ( 
.A(n_4172),
.B(n_606),
.Y(n_4269)
);

NAND3xp33_ASAP7_75t_L g4270 ( 
.A(n_4173),
.B(n_607),
.C(n_608),
.Y(n_4270)
);

XNOR2x1_ASAP7_75t_L g4271 ( 
.A(n_4194),
.B(n_609),
.Y(n_4271)
);

AOI221x1_ASAP7_75t_L g4272 ( 
.A1(n_4137),
.A2(n_612),
.B1(n_609),
.B2(n_611),
.C(n_613),
.Y(n_4272)
);

A2O1A1Ixp33_ASAP7_75t_L g4273 ( 
.A1(n_4149),
.A2(n_4131),
.B(n_4176),
.C(n_4159),
.Y(n_4273)
);

NOR2xp67_ASAP7_75t_L g4274 ( 
.A(n_4129),
.B(n_611),
.Y(n_4274)
);

NOR3xp33_ASAP7_75t_L g4275 ( 
.A(n_4192),
.B(n_612),
.C(n_613),
.Y(n_4275)
);

NAND2xp5_ASAP7_75t_SL g4276 ( 
.A(n_4139),
.B(n_615),
.Y(n_4276)
);

NAND3xp33_ASAP7_75t_SL g4277 ( 
.A(n_4165),
.B(n_615),
.C(n_616),
.Y(n_4277)
);

NOR2x1_ASAP7_75t_L g4278 ( 
.A(n_4187),
.B(n_617),
.Y(n_4278)
);

AND2x4_ASAP7_75t_L g4279 ( 
.A(n_4186),
.B(n_618),
.Y(n_4279)
);

AOI22xp5_ASAP7_75t_L g4280 ( 
.A1(n_4167),
.A2(n_620),
.B1(n_618),
.B2(n_619),
.Y(n_4280)
);

CKINVDCx16_ASAP7_75t_R g4281 ( 
.A(n_4197),
.Y(n_4281)
);

OAI22xp5_ASAP7_75t_L g4282 ( 
.A1(n_4169),
.A2(n_622),
.B1(n_619),
.B2(n_621),
.Y(n_4282)
);

AOI22xp5_ASAP7_75t_L g4283 ( 
.A1(n_4155),
.A2(n_625),
.B1(n_621),
.B2(n_624),
.Y(n_4283)
);

NOR3x1_ASAP7_75t_L g4284 ( 
.A(n_4158),
.B(n_624),
.C(n_625),
.Y(n_4284)
);

XOR2xp5_ASAP7_75t_L g4285 ( 
.A(n_4154),
.B(n_626),
.Y(n_4285)
);

AOI21xp5_ASAP7_75t_L g4286 ( 
.A1(n_4163),
.A2(n_626),
.B(n_627),
.Y(n_4286)
);

AND3x2_ASAP7_75t_L g4287 ( 
.A(n_4141),
.B(n_627),
.C(n_628),
.Y(n_4287)
);

INVx2_ASAP7_75t_L g4288 ( 
.A(n_4217),
.Y(n_4288)
);

OAI221xp5_ASAP7_75t_L g4289 ( 
.A1(n_4226),
.A2(n_644),
.B1(n_655),
.B2(n_636),
.C(n_628),
.Y(n_4289)
);

OR2x2_ASAP7_75t_L g4290 ( 
.A(n_4214),
.B(n_629),
.Y(n_4290)
);

OAI21xp5_ASAP7_75t_SL g4291 ( 
.A1(n_4246),
.A2(n_630),
.B(n_631),
.Y(n_4291)
);

NAND2xp5_ASAP7_75t_L g4292 ( 
.A(n_4287),
.B(n_631),
.Y(n_4292)
);

NAND3xp33_ASAP7_75t_L g4293 ( 
.A(n_4251),
.B(n_632),
.C(n_633),
.Y(n_4293)
);

OAI22xp5_ASAP7_75t_L g4294 ( 
.A1(n_4228),
.A2(n_634),
.B1(n_632),
.B2(n_633),
.Y(n_4294)
);

NOR2xp67_ASAP7_75t_L g4295 ( 
.A(n_4279),
.B(n_4277),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_4223),
.Y(n_4296)
);

NAND2xp5_ASAP7_75t_L g4297 ( 
.A(n_4245),
.B(n_4220),
.Y(n_4297)
);

NOR3xp33_ASAP7_75t_L g4298 ( 
.A(n_4219),
.B(n_4281),
.C(n_4231),
.Y(n_4298)
);

AND2x4_ASAP7_75t_L g4299 ( 
.A(n_4212),
.B(n_634),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_4285),
.Y(n_4300)
);

OR5x1_ASAP7_75t_L g4301 ( 
.A(n_4230),
.B(n_637),
.C(n_635),
.D(n_636),
.E(n_638),
.Y(n_4301)
);

NOR3x2_ASAP7_75t_L g4302 ( 
.A(n_4227),
.B(n_635),
.C(n_637),
.Y(n_4302)
);

NAND2x1p5_ASAP7_75t_L g4303 ( 
.A(n_4263),
.B(n_638),
.Y(n_4303)
);

NOR2x1_ASAP7_75t_L g4304 ( 
.A(n_4233),
.B(n_4224),
.Y(n_4304)
);

NAND2xp5_ASAP7_75t_L g4305 ( 
.A(n_4234),
.B(n_639),
.Y(n_4305)
);

AND3x4_ASAP7_75t_L g4306 ( 
.A(n_4278),
.B(n_639),
.C(n_640),
.Y(n_4306)
);

OAI22x1_ASAP7_75t_L g4307 ( 
.A1(n_4213),
.A2(n_642),
.B1(n_640),
.B2(n_641),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_4238),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_4254),
.Y(n_4309)
);

AND3x4_ASAP7_75t_L g4310 ( 
.A(n_4275),
.B(n_643),
.C(n_645),
.Y(n_4310)
);

CKINVDCx20_ASAP7_75t_R g4311 ( 
.A(n_4250),
.Y(n_4311)
);

AOI221xp5_ASAP7_75t_L g4312 ( 
.A1(n_4216),
.A2(n_648),
.B1(n_643),
.B2(n_645),
.C(n_649),
.Y(n_4312)
);

NAND4xp25_ASAP7_75t_L g4313 ( 
.A(n_4255),
.B(n_652),
.C(n_649),
.D(n_651),
.Y(n_4313)
);

NOR3xp33_ASAP7_75t_L g4314 ( 
.A(n_4215),
.B(n_651),
.C(n_653),
.Y(n_4314)
);

XNOR2xp5_ASAP7_75t_L g4315 ( 
.A(n_4225),
.B(n_653),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_4234),
.Y(n_4316)
);

OAI211xp5_ASAP7_75t_L g4317 ( 
.A1(n_4280),
.A2(n_4258),
.B(n_4232),
.C(n_4248),
.Y(n_4317)
);

O2A1O1Ixp33_ASAP7_75t_L g4318 ( 
.A1(n_4240),
.A2(n_657),
.B(n_654),
.C(n_656),
.Y(n_4318)
);

AOI221xp5_ASAP7_75t_L g4319 ( 
.A1(n_4260),
.A2(n_659),
.B1(n_654),
.B2(n_656),
.C(n_660),
.Y(n_4319)
);

HB1xp67_ASAP7_75t_L g4320 ( 
.A(n_4274),
.Y(n_4320)
);

NOR2x1_ASAP7_75t_L g4321 ( 
.A(n_4218),
.B(n_659),
.Y(n_4321)
);

INVx2_ASAP7_75t_L g4322 ( 
.A(n_4284),
.Y(n_4322)
);

AND2x2_ASAP7_75t_L g4323 ( 
.A(n_4221),
.B(n_660),
.Y(n_4323)
);

AND2x2_ASAP7_75t_L g4324 ( 
.A(n_4269),
.B(n_661),
.Y(n_4324)
);

NOR3xp33_ASAP7_75t_L g4325 ( 
.A(n_4252),
.B(n_661),
.C(n_662),
.Y(n_4325)
);

NOR2xp33_ASAP7_75t_L g4326 ( 
.A(n_4259),
.B(n_662),
.Y(n_4326)
);

AND2x4_ASAP7_75t_L g4327 ( 
.A(n_4247),
.B(n_663),
.Y(n_4327)
);

NOR2xp33_ASAP7_75t_L g4328 ( 
.A(n_4244),
.B(n_4239),
.Y(n_4328)
);

NAND5xp2_ASAP7_75t_L g4329 ( 
.A(n_4236),
.B(n_665),
.C(n_663),
.D(n_664),
.E(n_670),
.Y(n_4329)
);

AOI211xp5_ASAP7_75t_L g4330 ( 
.A1(n_4222),
.A2(n_671),
.B(n_665),
.C(n_670),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_4229),
.Y(n_4331)
);

NOR3xp33_ASAP7_75t_L g4332 ( 
.A(n_4253),
.B(n_671),
.C(n_672),
.Y(n_4332)
);

AND2x4_ASAP7_75t_L g4333 ( 
.A(n_4268),
.B(n_672),
.Y(n_4333)
);

OAI21xp33_ASAP7_75t_L g4334 ( 
.A1(n_4273),
.A2(n_673),
.B(n_675),
.Y(n_4334)
);

A2O1A1Ixp33_ASAP7_75t_L g4335 ( 
.A1(n_4267),
.A2(n_4286),
.B(n_4249),
.C(n_4235),
.Y(n_4335)
);

INVx1_ASAP7_75t_L g4336 ( 
.A(n_4266),
.Y(n_4336)
);

HB1xp67_ASAP7_75t_L g4337 ( 
.A(n_4272),
.Y(n_4337)
);

BUFx4f_ASAP7_75t_L g4338 ( 
.A(n_4256),
.Y(n_4338)
);

NOR3x1_ASAP7_75t_SL g4339 ( 
.A(n_4264),
.B(n_4271),
.C(n_4257),
.Y(n_4339)
);

NOR3xp33_ASAP7_75t_L g4340 ( 
.A(n_4237),
.B(n_673),
.C(n_675),
.Y(n_4340)
);

NOR2x1_ASAP7_75t_L g4341 ( 
.A(n_4270),
.B(n_676),
.Y(n_4341)
);

AOI221xp5_ASAP7_75t_L g4342 ( 
.A1(n_4243),
.A2(n_682),
.B1(n_677),
.B2(n_678),
.C(n_683),
.Y(n_4342)
);

NOR2x1_ASAP7_75t_L g4343 ( 
.A(n_4313),
.B(n_4261),
.Y(n_4343)
);

CKINVDCx5p33_ASAP7_75t_R g4344 ( 
.A(n_4311),
.Y(n_4344)
);

CKINVDCx5p33_ASAP7_75t_R g4345 ( 
.A(n_4338),
.Y(n_4345)
);

INVxp67_ASAP7_75t_L g4346 ( 
.A(n_4329),
.Y(n_4346)
);

INVx2_ASAP7_75t_L g4347 ( 
.A(n_4303),
.Y(n_4347)
);

AOI211xp5_ASAP7_75t_L g4348 ( 
.A1(n_4318),
.A2(n_4282),
.B(n_4242),
.C(n_4276),
.Y(n_4348)
);

HB1xp67_ASAP7_75t_L g4349 ( 
.A(n_4337),
.Y(n_4349)
);

INVx1_ASAP7_75t_L g4350 ( 
.A(n_4290),
.Y(n_4350)
);

BUFx6f_ASAP7_75t_L g4351 ( 
.A(n_4327),
.Y(n_4351)
);

CKINVDCx20_ASAP7_75t_R g4352 ( 
.A(n_4300),
.Y(n_4352)
);

CKINVDCx20_ASAP7_75t_R g4353 ( 
.A(n_4320),
.Y(n_4353)
);

INVx1_ASAP7_75t_SL g4354 ( 
.A(n_4302),
.Y(n_4354)
);

CKINVDCx11_ASAP7_75t_R g4355 ( 
.A(n_4288),
.Y(n_4355)
);

BUFx2_ASAP7_75t_L g4356 ( 
.A(n_4333),
.Y(n_4356)
);

BUFx6f_ASAP7_75t_L g4357 ( 
.A(n_4331),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_4315),
.Y(n_4358)
);

XNOR2xp5_ASAP7_75t_L g4359 ( 
.A(n_4306),
.B(n_4283),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_4299),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_4305),
.Y(n_4361)
);

NOR2xp33_ASAP7_75t_L g4362 ( 
.A(n_4334),
.B(n_4262),
.Y(n_4362)
);

CKINVDCx5p33_ASAP7_75t_R g4363 ( 
.A(n_4296),
.Y(n_4363)
);

CKINVDCx5p33_ASAP7_75t_R g4364 ( 
.A(n_4323),
.Y(n_4364)
);

CKINVDCx6p67_ASAP7_75t_R g4365 ( 
.A(n_4333),
.Y(n_4365)
);

INVx1_ASAP7_75t_L g4366 ( 
.A(n_4324),
.Y(n_4366)
);

CKINVDCx5p33_ASAP7_75t_R g4367 ( 
.A(n_4322),
.Y(n_4367)
);

CKINVDCx5p33_ASAP7_75t_R g4368 ( 
.A(n_4316),
.Y(n_4368)
);

OAI22xp33_ASAP7_75t_L g4369 ( 
.A1(n_4292),
.A2(n_4241),
.B1(n_4256),
.B2(n_4265),
.Y(n_4369)
);

OR2x2_ASAP7_75t_L g4370 ( 
.A(n_4308),
.B(n_677),
.Y(n_4370)
);

NOR2x1_ASAP7_75t_L g4371 ( 
.A(n_4295),
.B(n_678),
.Y(n_4371)
);

CKINVDCx5p33_ASAP7_75t_R g4372 ( 
.A(n_4309),
.Y(n_4372)
);

INVx2_ASAP7_75t_SL g4373 ( 
.A(n_4321),
.Y(n_4373)
);

OA21x2_ASAP7_75t_L g4374 ( 
.A1(n_4297),
.A2(n_682),
.B(n_683),
.Y(n_4374)
);

NAND2xp5_ASAP7_75t_L g4375 ( 
.A(n_4312),
.B(n_684),
.Y(n_4375)
);

INVx2_ASAP7_75t_L g4376 ( 
.A(n_4307),
.Y(n_4376)
);

AOI22xp33_ASAP7_75t_L g4377 ( 
.A1(n_4357),
.A2(n_4298),
.B1(n_4325),
.B2(n_4332),
.Y(n_4377)
);

OAI22xp5_ASAP7_75t_SL g4378 ( 
.A1(n_4352),
.A2(n_4301),
.B1(n_4310),
.B2(n_4326),
.Y(n_4378)
);

AOI21xp5_ASAP7_75t_L g4379 ( 
.A1(n_4356),
.A2(n_4335),
.B(n_4291),
.Y(n_4379)
);

AOI22xp5_ASAP7_75t_L g4380 ( 
.A1(n_4344),
.A2(n_4328),
.B1(n_4340),
.B2(n_4314),
.Y(n_4380)
);

AOI22xp5_ASAP7_75t_L g4381 ( 
.A1(n_4353),
.A2(n_4304),
.B1(n_4317),
.B2(n_4293),
.Y(n_4381)
);

NOR3xp33_ASAP7_75t_L g4382 ( 
.A(n_4355),
.B(n_4336),
.C(n_4342),
.Y(n_4382)
);

AOI21xp5_ASAP7_75t_L g4383 ( 
.A1(n_4349),
.A2(n_4341),
.B(n_4319),
.Y(n_4383)
);

AOI211xp5_ASAP7_75t_SL g4384 ( 
.A1(n_4369),
.A2(n_4289),
.B(n_4294),
.C(n_4330),
.Y(n_4384)
);

INVx1_ASAP7_75t_L g4385 ( 
.A(n_4371),
.Y(n_4385)
);

INVx1_ASAP7_75t_L g4386 ( 
.A(n_4365),
.Y(n_4386)
);

NOR2xp33_ASAP7_75t_L g4387 ( 
.A(n_4346),
.B(n_4339),
.Y(n_4387)
);

OA21x2_ASAP7_75t_L g4388 ( 
.A1(n_4376),
.A2(n_684),
.B(n_685),
.Y(n_4388)
);

INVx2_ASAP7_75t_L g4389 ( 
.A(n_4374),
.Y(n_4389)
);

NAND3xp33_ASAP7_75t_L g4390 ( 
.A(n_4348),
.B(n_686),
.C(n_687),
.Y(n_4390)
);

OAI21xp5_ASAP7_75t_L g4391 ( 
.A1(n_4343),
.A2(n_686),
.B(n_688),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_4370),
.Y(n_4392)
);

OAI21xp5_ASAP7_75t_L g4393 ( 
.A1(n_4362),
.A2(n_689),
.B(n_690),
.Y(n_4393)
);

BUFx2_ASAP7_75t_L g4394 ( 
.A(n_4388),
.Y(n_4394)
);

HB1xp67_ASAP7_75t_L g4395 ( 
.A(n_4389),
.Y(n_4395)
);

INVx1_ASAP7_75t_L g4396 ( 
.A(n_4390),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4385),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4378),
.Y(n_4398)
);

NOR2x1_ASAP7_75t_L g4399 ( 
.A(n_4391),
.B(n_4374),
.Y(n_4399)
);

INVx1_ASAP7_75t_L g4400 ( 
.A(n_4386),
.Y(n_4400)
);

AOI22xp33_ASAP7_75t_L g4401 ( 
.A1(n_4387),
.A2(n_4357),
.B1(n_4351),
.B2(n_4373),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_4392),
.Y(n_4402)
);

NOR2x1p5_ASAP7_75t_L g4403 ( 
.A(n_4384),
.B(n_4360),
.Y(n_4403)
);

NOR4xp25_ASAP7_75t_L g4404 ( 
.A(n_4377),
.B(n_4354),
.C(n_4358),
.D(n_4366),
.Y(n_4404)
);

INVx1_ASAP7_75t_L g4405 ( 
.A(n_4394),
.Y(n_4405)
);

INVx1_ASAP7_75t_L g4406 ( 
.A(n_4395),
.Y(n_4406)
);

INVx1_ASAP7_75t_L g4407 ( 
.A(n_4399),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_4400),
.Y(n_4408)
);

INVx2_ASAP7_75t_SL g4409 ( 
.A(n_4403),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4402),
.Y(n_4410)
);

INVx1_ASAP7_75t_L g4411 ( 
.A(n_4397),
.Y(n_4411)
);

NAND4xp25_ASAP7_75t_SL g4412 ( 
.A(n_4406),
.B(n_4401),
.C(n_4381),
.D(n_4383),
.Y(n_4412)
);

OAI22xp5_ASAP7_75t_SL g4413 ( 
.A1(n_4409),
.A2(n_4364),
.B1(n_4345),
.B2(n_4368),
.Y(n_4413)
);

OR2x2_ASAP7_75t_L g4414 ( 
.A(n_4405),
.B(n_4375),
.Y(n_4414)
);

OAI322xp33_ASAP7_75t_L g4415 ( 
.A1(n_4407),
.A2(n_4398),
.A3(n_4380),
.B1(n_4379),
.B2(n_4350),
.C1(n_4396),
.C2(n_4347),
.Y(n_4415)
);

HB1xp67_ASAP7_75t_L g4416 ( 
.A(n_4408),
.Y(n_4416)
);

INVx1_ASAP7_75t_L g4417 ( 
.A(n_4416),
.Y(n_4417)
);

OAI21xp5_ASAP7_75t_L g4418 ( 
.A1(n_4412),
.A2(n_4404),
.B(n_4411),
.Y(n_4418)
);

AOI32xp33_ASAP7_75t_L g4419 ( 
.A1(n_4417),
.A2(n_4410),
.A3(n_4382),
.B1(n_4367),
.B2(n_4361),
.Y(n_4419)
);

AOI22xp33_ASAP7_75t_L g4420 ( 
.A1(n_4419),
.A2(n_4351),
.B1(n_4413),
.B2(n_4372),
.Y(n_4420)
);

OA22x2_ASAP7_75t_L g4421 ( 
.A1(n_4420),
.A2(n_4418),
.B1(n_4363),
.B2(n_4359),
.Y(n_4421)
);

AO21x2_ASAP7_75t_L g4422 ( 
.A1(n_4421),
.A2(n_4414),
.B(n_4415),
.Y(n_4422)
);

AOI22xp5_ASAP7_75t_L g4423 ( 
.A1(n_4422),
.A2(n_4393),
.B1(n_694),
.B2(n_691),
.Y(n_4423)
);

AOI211xp5_ASAP7_75t_L g4424 ( 
.A1(n_4423),
.A2(n_694),
.B(n_691),
.C(n_693),
.Y(n_4424)
);


endmodule