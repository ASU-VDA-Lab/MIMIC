module real_aes_6528_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g476 ( .A1(n_0), .A2(n_180), .B(n_477), .C(n_480), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_1), .B(n_471), .Y(n_482) );
INVx1_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
INVx1_ASAP7_75t_L g229 ( .A(n_3), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_4), .B(n_168), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_5), .A2(n_455), .B(n_525), .Y(n_524) );
OAI22xp5_ASAP7_75t_SL g751 ( .A1(n_6), .A2(n_9), .B1(n_438), .B2(n_752), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_6), .Y(n_752) );
AO21x2_ASAP7_75t_L g533 ( .A1(n_7), .A2(n_185), .B(n_534), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g179 ( .A1(n_8), .A2(n_38), .B1(n_141), .B2(n_153), .Y(n_179) );
AOI22xp5_ASAP7_75t_L g124 ( .A1(n_9), .A2(n_125), .B1(n_126), .B2(n_438), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_9), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_10), .B(n_185), .Y(n_218) );
AND2x6_ASAP7_75t_L g156 ( .A(n_11), .B(n_157), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_12), .A2(n_156), .B(n_458), .C(n_547), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_13), .B(n_39), .Y(n_111) );
INVx1_ASAP7_75t_L g137 ( .A(n_14), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_15), .B(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g223 ( .A(n_16), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_17), .B(n_168), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_18), .B(n_183), .Y(n_201) );
AO32x2_ASAP7_75t_L g177 ( .A1(n_19), .A2(n_178), .A3(n_182), .B1(n_184), .B2(n_185), .Y(n_177) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_20), .A2(n_101), .B1(n_112), .B2(n_755), .Y(n_100) );
AOI222xp33_ASAP7_75t_SL g121 ( .A1(n_21), .A2(n_92), .B1(n_122), .B2(n_737), .C1(n_738), .C2(n_740), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_21), .Y(n_737) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_22), .B(n_141), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_23), .B(n_183), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_24), .A2(n_54), .B1(n_141), .B2(n_153), .Y(n_181) );
AOI22xp33_ASAP7_75t_SL g194 ( .A1(n_25), .A2(n_79), .B1(n_141), .B2(n_145), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_26), .B(n_141), .Y(n_171) );
A2O1A1Ixp33_ASAP7_75t_L g457 ( .A1(n_27), .A2(n_184), .B(n_458), .C(n_460), .Y(n_457) );
A2O1A1Ixp33_ASAP7_75t_L g536 ( .A1(n_28), .A2(n_184), .B(n_458), .C(n_537), .Y(n_536) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_29), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_30), .B(n_133), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_31), .A2(n_455), .B(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_32), .B(n_133), .Y(n_175) );
INVx2_ASAP7_75t_L g143 ( .A(n_33), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_34), .A2(n_489), .B(n_490), .C(n_494), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_35), .B(n_141), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_36), .B(n_133), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_37), .B(n_148), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_40), .B(n_454), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_41), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_42), .B(n_168), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_43), .B(n_455), .Y(n_535) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_44), .A2(n_489), .B(n_494), .C(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_45), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_46), .B(n_141), .Y(n_211) );
INVx1_ASAP7_75t_L g478 ( .A(n_47), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g192 ( .A1(n_48), .A2(n_88), .B1(n_153), .B2(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g517 ( .A(n_49), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_50), .B(n_141), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_51), .B(n_141), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_52), .B(n_455), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_53), .B(n_216), .Y(n_215) );
AOI22xp33_ASAP7_75t_SL g205 ( .A1(n_55), .A2(n_59), .B1(n_141), .B2(n_145), .Y(n_205) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_56), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_57), .B(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_58), .B(n_141), .Y(n_242) );
INVx1_ASAP7_75t_L g157 ( .A(n_60), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_61), .B(n_455), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_62), .B(n_471), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_63), .A2(n_216), .B(n_226), .C(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_64), .B(n_141), .Y(n_230) );
INVx1_ASAP7_75t_L g136 ( .A(n_65), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_66), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_67), .B(n_168), .Y(n_492) );
AO32x2_ASAP7_75t_L g190 ( .A1(n_68), .A2(n_184), .A3(n_185), .B1(n_191), .B2(n_195), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_69), .B(n_169), .Y(n_548) );
INVx1_ASAP7_75t_L g241 ( .A(n_70), .Y(n_241) );
INVx1_ASAP7_75t_L g166 ( .A(n_71), .Y(n_166) );
CKINVDCx16_ASAP7_75t_R g474 ( .A(n_72), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_73), .B(n_462), .Y(n_461) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_74), .A2(n_458), .B(n_494), .C(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_75), .B(n_145), .Y(n_167) );
CKINVDCx16_ASAP7_75t_R g526 ( .A(n_76), .Y(n_526) );
INVx1_ASAP7_75t_L g105 ( .A(n_77), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_78), .B(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_80), .B(n_153), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_81), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_82), .B(n_145), .Y(n_172) );
INVx2_ASAP7_75t_L g134 ( .A(n_83), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_84), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_85), .B(n_155), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_86), .B(n_145), .Y(n_212) );
OR2x2_ASAP7_75t_L g107 ( .A(n_87), .B(n_108), .Y(n_107) );
OR2x2_ASAP7_75t_L g441 ( .A(n_87), .B(n_109), .Y(n_441) );
INVx2_ASAP7_75t_L g736 ( .A(n_87), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_89), .A2(n_99), .B1(n_145), .B2(n_146), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_90), .B(n_455), .Y(n_487) );
INVx1_ASAP7_75t_L g491 ( .A(n_91), .Y(n_491) );
INVxp67_ASAP7_75t_L g529 ( .A(n_93), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_94), .B(n_145), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_95), .B(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g504 ( .A(n_96), .Y(n_504) );
INVx1_ASAP7_75t_L g544 ( .A(n_97), .Y(n_544) );
AND2x2_ASAP7_75t_L g519 ( .A(n_98), .B(n_133), .Y(n_519) );
INVx1_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g756 ( .A(n_102), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_103), .B(n_106), .Y(n_102) );
INVx1_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_107), .Y(n_119) );
INVx1_ASAP7_75t_SL g754 ( .A(n_107), .Y(n_754) );
NOR2x2_ASAP7_75t_L g742 ( .A(n_108), .B(n_736), .Y(n_742) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g735 ( .A(n_109), .B(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
AOI22x1_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_121), .B1(n_743), .B2(n_744), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_118), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_SL g743 ( .A(n_116), .Y(n_743) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g744 ( .A1(n_118), .A2(n_745), .B(n_753), .Y(n_744) );
NOR2xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_120), .Y(n_118) );
OAI22x1_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_439), .B1(n_442), .B2(n_733), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI22xp5_ASAP7_75t_SL g738 ( .A1(n_124), .A2(n_443), .B1(n_733), .B2(n_739), .Y(n_738) );
OAI22xp5_ASAP7_75t_SL g749 ( .A1(n_125), .A2(n_126), .B1(n_750), .B2(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_360), .Y(n_126) );
NAND5xp2_ASAP7_75t_L g127 ( .A(n_128), .B(n_279), .C(n_294), .D(n_320), .E(n_342), .Y(n_127) );
NOR2xp33_ASAP7_75t_SL g128 ( .A(n_129), .B(n_259), .Y(n_128) );
OAI221xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_196), .B1(n_232), .B2(n_248), .C(n_249), .Y(n_129) );
NOR2xp33_ASAP7_75t_SL g130 ( .A(n_131), .B(n_186), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_131), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_SL g436 ( .A(n_131), .Y(n_436) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_159), .Y(n_131) );
INVx1_ASAP7_75t_L g276 ( .A(n_132), .Y(n_276) );
AND2x2_ASAP7_75t_L g278 ( .A(n_132), .B(n_177), .Y(n_278) );
AND2x2_ASAP7_75t_L g288 ( .A(n_132), .B(n_176), .Y(n_288) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_132), .Y(n_306) );
INVx1_ASAP7_75t_L g316 ( .A(n_132), .Y(n_316) );
OR2x2_ASAP7_75t_L g354 ( .A(n_132), .B(n_253), .Y(n_354) );
INVx2_ASAP7_75t_L g404 ( .A(n_132), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_132), .B(n_252), .Y(n_421) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_138), .B(n_158), .Y(n_132) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_133), .A2(n_163), .B(n_175), .Y(n_162) );
INVx2_ASAP7_75t_L g195 ( .A(n_133), .Y(n_195) );
INVx1_ASAP7_75t_L g468 ( .A(n_133), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_133), .A2(n_487), .B(n_488), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_133), .A2(n_514), .B(n_515), .Y(n_513) );
AND2x2_ASAP7_75t_SL g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AND2x2_ASAP7_75t_L g183 ( .A(n_134), .B(n_135), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
OAI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_150), .B(n_156), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_144), .B(n_147), .Y(n_139) );
INVx3_ASAP7_75t_L g165 ( .A(n_141), .Y(n_165) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_141), .Y(n_506) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g153 ( .A(n_142), .Y(n_153) );
BUFx3_ASAP7_75t_L g193 ( .A(n_142), .Y(n_193) );
AND2x6_ASAP7_75t_L g458 ( .A(n_142), .B(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g146 ( .A(n_143), .Y(n_146) );
INVx1_ASAP7_75t_L g217 ( .A(n_143), .Y(n_217) );
INVx2_ASAP7_75t_L g224 ( .A(n_145), .Y(n_224) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_149), .Y(n_155) );
INVx3_ASAP7_75t_L g169 ( .A(n_149), .Y(n_169) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_149), .Y(n_174) );
AND2x2_ASAP7_75t_L g456 ( .A(n_149), .B(n_217), .Y(n_456) );
INVx1_ASAP7_75t_L g459 ( .A(n_149), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_154), .Y(n_150) );
O2A1O1Ixp5_ASAP7_75t_L g240 ( .A1(n_154), .A2(n_228), .B(n_241), .C(n_242), .Y(n_240) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
OAI22xp5_ASAP7_75t_L g178 ( .A1(n_155), .A2(n_179), .B1(n_180), .B2(n_181), .Y(n_178) );
OAI22xp5_ASAP7_75t_SL g191 ( .A1(n_155), .A2(n_169), .B1(n_192), .B2(n_194), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g203 ( .A1(n_155), .A2(n_180), .B1(n_204), .B2(n_205), .Y(n_203) );
INVx4_ASAP7_75t_L g479 ( .A(n_155), .Y(n_479) );
OAI21xp5_ASAP7_75t_L g163 ( .A1(n_156), .A2(n_164), .B(n_170), .Y(n_163) );
BUFx3_ASAP7_75t_L g184 ( .A(n_156), .Y(n_184) );
OAI21xp5_ASAP7_75t_L g209 ( .A1(n_156), .A2(n_210), .B(n_213), .Y(n_209) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_156), .A2(n_222), .B(n_227), .Y(n_221) );
AND2x4_ASAP7_75t_L g455 ( .A(n_156), .B(n_456), .Y(n_455) );
INVx4_ASAP7_75t_SL g481 ( .A(n_156), .Y(n_481) );
NAND2x1p5_ASAP7_75t_L g545 ( .A(n_156), .B(n_456), .Y(n_545) );
NOR2xp67_ASAP7_75t_L g159 ( .A(n_160), .B(n_176), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_161), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_161), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_SL g336 ( .A(n_161), .B(n_276), .Y(n_336) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_162), .Y(n_188) );
INVx2_ASAP7_75t_L g253 ( .A(n_162), .Y(n_253) );
OR2x2_ASAP7_75t_L g315 ( .A(n_162), .B(n_316), .Y(n_315) );
O2A1O1Ixp5_ASAP7_75t_SL g164 ( .A1(n_165), .A2(n_166), .B(n_167), .C(n_168), .Y(n_164) );
INVx2_ASAP7_75t_L g180 ( .A(n_168), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_168), .A2(n_211), .B(n_212), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_168), .A2(n_238), .B(n_239), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_168), .B(n_529), .Y(n_528) );
INVx5_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_173), .Y(n_170) );
INVx1_ASAP7_75t_L g226 ( .A(n_173), .Y(n_226) );
INVx4_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g462 ( .A(n_174), .Y(n_462) );
AND2x2_ASAP7_75t_L g254 ( .A(n_176), .B(n_190), .Y(n_254) );
AND2x2_ASAP7_75t_L g271 ( .A(n_176), .B(n_251), .Y(n_271) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g189 ( .A(n_177), .B(n_190), .Y(n_189) );
BUFx2_ASAP7_75t_L g274 ( .A(n_177), .Y(n_274) );
AND2x2_ASAP7_75t_L g403 ( .A(n_177), .B(n_404), .Y(n_403) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_180), .A2(n_214), .B(n_215), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_L g227 ( .A1(n_180), .A2(n_228), .B(n_229), .C(n_230), .Y(n_227) );
INVx2_ASAP7_75t_L g220 ( .A(n_182), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_182), .B(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_183), .Y(n_185) );
NAND3xp33_ASAP7_75t_L g202 ( .A(n_184), .B(n_203), .C(n_206), .Y(n_202) );
OAI21xp5_ASAP7_75t_L g236 ( .A1(n_184), .A2(n_237), .B(n_240), .Y(n_236) );
INVx4_ASAP7_75t_L g206 ( .A(n_185), .Y(n_206) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_185), .A2(n_209), .B(n_218), .Y(n_208) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_185), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_185), .A2(n_535), .B(n_536), .Y(n_534) );
INVx1_ASAP7_75t_L g248 ( .A(n_186), .Y(n_248) );
AND2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_189), .Y(n_186) );
AND2x2_ASAP7_75t_L g366 ( .A(n_187), .B(n_254), .Y(n_366) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g367 ( .A(n_188), .B(n_278), .Y(n_367) );
O2A1O1Ixp33_ASAP7_75t_L g334 ( .A1(n_189), .A2(n_335), .B(n_337), .C(n_339), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_189), .B(n_335), .Y(n_344) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_189), .A2(n_265), .B1(n_408), .B2(n_409), .C(n_411), .Y(n_407) );
INVx1_ASAP7_75t_L g251 ( .A(n_190), .Y(n_251) );
INVx1_ASAP7_75t_L g287 ( .A(n_190), .Y(n_287) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_190), .Y(n_296) );
INVx2_ASAP7_75t_L g480 ( .A(n_193), .Y(n_480) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_193), .Y(n_493) );
INVx1_ASAP7_75t_L g465 ( .A(n_195), .Y(n_465) );
INVx1_ASAP7_75t_SL g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_207), .Y(n_197) );
AND2x2_ASAP7_75t_L g313 ( .A(n_198), .B(n_258), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_198), .B(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_199), .B(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g405 ( .A(n_199), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g437 ( .A(n_199), .Y(n_437) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx3_ASAP7_75t_L g267 ( .A(n_200), .Y(n_267) );
AND2x2_ASAP7_75t_L g293 ( .A(n_200), .B(n_247), .Y(n_293) );
NOR2x1_ASAP7_75t_L g302 ( .A(n_200), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g309 ( .A(n_200), .B(n_310), .Y(n_309) );
AND2x4_ASAP7_75t_L g200 ( .A(n_201), .B(n_202), .Y(n_200) );
INVx1_ASAP7_75t_L g245 ( .A(n_201), .Y(n_245) );
AO21x1_ASAP7_75t_L g244 ( .A1(n_203), .A2(n_206), .B(n_245), .Y(n_244) );
INVx3_ASAP7_75t_L g471 ( .A(n_206), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_206), .B(n_496), .Y(n_495) );
AO21x2_ASAP7_75t_L g500 ( .A1(n_206), .A2(n_501), .B(n_508), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_206), .B(n_509), .Y(n_508) );
AO21x2_ASAP7_75t_L g542 ( .A1(n_206), .A2(n_543), .B(n_550), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_207), .B(n_349), .Y(n_384) );
INVx1_ASAP7_75t_SL g388 ( .A(n_207), .Y(n_388) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_219), .Y(n_207) );
INVx3_ASAP7_75t_L g247 ( .A(n_208), .Y(n_247) );
AND2x2_ASAP7_75t_L g258 ( .A(n_208), .B(n_235), .Y(n_258) );
AND2x2_ASAP7_75t_L g280 ( .A(n_208), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g325 ( .A(n_208), .B(n_319), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_208), .B(n_257), .Y(n_406) );
INVx2_ASAP7_75t_L g228 ( .A(n_216), .Y(n_228) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g246 ( .A(n_219), .B(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g257 ( .A(n_219), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_219), .B(n_235), .Y(n_282) );
AND2x2_ASAP7_75t_L g318 ( .A(n_219), .B(n_319), .Y(n_318) );
OA21x2_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_231), .Y(n_219) );
OA21x2_ASAP7_75t_L g235 ( .A1(n_220), .A2(n_236), .B(n_243), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_225), .C(n_226), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_224), .A2(n_538), .B(n_539), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_224), .A2(n_548), .B(n_549), .Y(n_547) );
O2A1O1Ixp33_ASAP7_75t_L g503 ( .A1(n_226), .A2(n_504), .B(n_505), .C(n_506), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_228), .A2(n_461), .B(n_463), .Y(n_460) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_246), .Y(n_233) );
INVx1_ASAP7_75t_L g298 ( .A(n_234), .Y(n_298) );
AND2x2_ASAP7_75t_L g340 ( .A(n_234), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_SL g346 ( .A(n_234), .B(n_261), .Y(n_346) );
AOI21xp5_ASAP7_75t_SL g420 ( .A1(n_234), .A2(n_252), .B(n_275), .Y(n_420) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_244), .Y(n_234) );
OR2x2_ASAP7_75t_L g263 ( .A(n_235), .B(n_244), .Y(n_263) );
AND2x2_ASAP7_75t_L g310 ( .A(n_235), .B(n_247), .Y(n_310) );
INVx2_ASAP7_75t_L g319 ( .A(n_235), .Y(n_319) );
INVx1_ASAP7_75t_L g425 ( .A(n_235), .Y(n_425) );
AND2x2_ASAP7_75t_L g349 ( .A(n_244), .B(n_319), .Y(n_349) );
INVx1_ASAP7_75t_L g374 ( .A(n_244), .Y(n_374) );
AND2x2_ASAP7_75t_L g283 ( .A(n_246), .B(n_267), .Y(n_283) );
AND2x2_ASAP7_75t_L g295 ( .A(n_246), .B(n_296), .Y(n_295) );
INVx2_ASAP7_75t_SL g413 ( .A(n_246), .Y(n_413) );
INVx2_ASAP7_75t_L g303 ( .A(n_247), .Y(n_303) );
AND2x2_ASAP7_75t_L g341 ( .A(n_247), .B(n_257), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_247), .B(n_425), .Y(n_424) );
OAI21xp33_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_254), .B(n_255), .Y(n_249) );
AND2x2_ASAP7_75t_L g356 ( .A(n_250), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g410 ( .A(n_250), .Y(n_410) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
INVx1_ASAP7_75t_L g330 ( .A(n_251), .Y(n_330) );
BUFx2_ASAP7_75t_L g429 ( .A(n_251), .Y(n_429) );
BUFx2_ASAP7_75t_L g300 ( .A(n_252), .Y(n_300) );
AND2x2_ASAP7_75t_L g402 ( .A(n_252), .B(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g385 ( .A(n_253), .Y(n_385) );
AND2x4_ASAP7_75t_L g312 ( .A(n_254), .B(n_275), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g348 ( .A(n_254), .B(n_336), .Y(n_348) );
AOI32xp33_ASAP7_75t_L g272 ( .A1(n_255), .A2(n_273), .A3(n_275), .B1(n_277), .B2(n_278), .Y(n_272) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_258), .Y(n_255) );
INVx3_ASAP7_75t_L g261 ( .A(n_256), .Y(n_261) );
OR2x2_ASAP7_75t_L g397 ( .A(n_256), .B(n_353), .Y(n_397) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g266 ( .A(n_257), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g373 ( .A(n_257), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g265 ( .A(n_258), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g277 ( .A(n_258), .B(n_267), .Y(n_277) );
INVx1_ASAP7_75t_L g398 ( .A(n_258), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_258), .B(n_373), .Y(n_431) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_264), .B(n_268), .C(n_272), .Y(n_259) );
OAI322xp33_ASAP7_75t_L g368 ( .A1(n_260), .A2(n_305), .A3(n_369), .B1(n_371), .B2(n_375), .C1(n_376), .C2(n_380), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVxp67_ASAP7_75t_L g333 ( .A(n_261), .Y(n_333) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g387 ( .A(n_263), .B(n_388), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_263), .B(n_303), .Y(n_434) );
INVxp67_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g326 ( .A(n_266), .Y(n_326) );
OR2x2_ASAP7_75t_L g412 ( .A(n_267), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_270), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g321 ( .A(n_271), .B(n_300), .Y(n_321) );
AND2x2_ASAP7_75t_L g392 ( .A(n_271), .B(n_305), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_271), .B(n_379), .Y(n_414) );
AOI221xp5_ASAP7_75t_L g279 ( .A1(n_273), .A2(n_280), .B1(n_283), .B2(n_284), .C(n_289), .Y(n_279) );
OR2x2_ASAP7_75t_L g290 ( .A(n_273), .B(n_286), .Y(n_290) );
AND2x2_ASAP7_75t_L g378 ( .A(n_273), .B(n_379), .Y(n_378) );
AOI32xp33_ASAP7_75t_L g417 ( .A1(n_273), .A2(n_303), .A3(n_418), .B1(n_419), .B2(n_422), .Y(n_417) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND3xp33_ASAP7_75t_L g351 ( .A(n_274), .B(n_310), .C(n_333), .Y(n_351) );
AND2x2_ASAP7_75t_L g377 ( .A(n_274), .B(n_370), .Y(n_377) );
INVxp67_ASAP7_75t_L g357 ( .A(n_275), .Y(n_357) );
BUFx3_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g386 ( .A(n_278), .B(n_330), .Y(n_386) );
INVx2_ASAP7_75t_L g396 ( .A(n_278), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_278), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g365 ( .A(n_281), .Y(n_365) );
OR2x2_ASAP7_75t_L g291 ( .A(n_282), .B(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_284), .B(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_288), .Y(n_284) );
INVx1_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_287), .Y(n_370) );
AND2x2_ASAP7_75t_L g329 ( .A(n_288), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g375 ( .A(n_288), .Y(n_375) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_288), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
AOI21xp33_ASAP7_75t_SL g314 ( .A1(n_290), .A2(n_315), .B(n_317), .Y(n_314) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g408 ( .A(n_293), .B(n_318), .Y(n_408) );
AOI211xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_297), .B(n_307), .C(n_314), .Y(n_294) );
AND2x2_ASAP7_75t_L g338 ( .A(n_296), .B(n_306), .Y(n_338) );
INVx2_ASAP7_75t_L g353 ( .A(n_296), .Y(n_353) );
OR2x2_ASAP7_75t_L g391 ( .A(n_296), .B(n_354), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_296), .B(n_434), .Y(n_433) );
AOI211xp5_ASAP7_75t_SL g297 ( .A1(n_298), .A2(n_299), .B(n_301), .C(n_304), .Y(n_297) );
INVxp67_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_300), .B(n_338), .Y(n_337) );
OAI211xp5_ASAP7_75t_L g419 ( .A1(n_301), .A2(n_396), .B(n_420), .C(n_421), .Y(n_419) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2x1p5_ASAP7_75t_L g317 ( .A(n_302), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g359 ( .A(n_303), .B(n_349), .Y(n_359) );
INVx1_ASAP7_75t_L g364 ( .A(n_303), .Y(n_364) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_308), .B(n_311), .Y(n_307) );
INVxp33_ASAP7_75t_L g415 ( .A(n_309), .Y(n_415) );
AND2x2_ASAP7_75t_L g394 ( .A(n_310), .B(n_373), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_315), .A2(n_377), .B(n_378), .Y(n_376) );
OAI322xp33_ASAP7_75t_L g395 ( .A1(n_317), .A2(n_396), .A3(n_397), .B1(n_398), .B2(n_399), .C1(n_401), .C2(n_405), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_322), .B1(n_327), .B2(n_331), .C(n_334), .Y(n_320) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g372 ( .A(n_325), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g416 ( .A(n_329), .Y(n_416) );
INVxp67_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_332), .B(n_352), .Y(n_418) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g381 ( .A(n_341), .B(n_349), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_345), .B1(n_347), .B2(n_349), .C(n_350), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g361 ( .A1(n_345), .A2(n_362), .B1(n_366), .B2(n_367), .C(n_368), .Y(n_361) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVxp67_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_349), .B(n_364), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_352), .B1(n_355), .B2(n_358), .Y(n_350) );
OR2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx2_ASAP7_75t_SL g379 ( .A(n_354), .Y(n_379) );
INVxp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND5xp2_ASAP7_75t_L g360 ( .A(n_361), .B(n_382), .C(n_407), .D(n_417), .E(n_427), .Y(n_360) );
NAND2xp5_ASAP7_75t_SL g362 ( .A(n_363), .B(n_365), .Y(n_362) );
NOR4xp25_ASAP7_75t_L g435 ( .A(n_364), .B(n_370), .C(n_436), .D(n_437), .Y(n_435) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_367), .A2(n_428), .B1(n_430), .B2(n_432), .C(n_435), .Y(n_427) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g426 ( .A(n_373), .Y(n_426) );
OAI322xp33_ASAP7_75t_L g383 ( .A1(n_377), .A2(n_384), .A3(n_385), .B1(n_386), .B2(n_387), .C1(n_389), .C2(n_393), .Y(n_383) );
INVx1_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_383), .B(n_395), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g428 ( .A(n_403), .B(n_429), .Y(n_428) );
OAI22xp33_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_414), .B1(n_415), .B2(n_416), .Y(n_411) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_426), .Y(n_423) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVxp67_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g739 ( .A(n_440), .Y(n_739) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_SL g443 ( .A(n_444), .B(n_688), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_445), .B(n_623), .Y(n_444) );
NAND4xp25_ASAP7_75t_SL g445 ( .A(n_446), .B(n_568), .C(n_592), .D(n_615), .Y(n_445) );
AOI221xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_510), .B1(n_540), .B2(n_552), .C(n_555), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_483), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_449), .A2(n_469), .B1(n_511), .B2(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_449), .B(n_484), .Y(n_626) );
AND2x2_ASAP7_75t_L g645 ( .A(n_449), .B(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_449), .B(n_629), .Y(n_715) );
AND2x4_ASAP7_75t_L g449 ( .A(n_450), .B(n_469), .Y(n_449) );
AND2x2_ASAP7_75t_L g583 ( .A(n_450), .B(n_484), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_450), .B(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g606 ( .A(n_450), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g611 ( .A(n_450), .B(n_470), .Y(n_611) );
INVx2_ASAP7_75t_L g643 ( .A(n_450), .Y(n_643) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_450), .Y(n_687) );
AND2x2_ASAP7_75t_L g704 ( .A(n_450), .B(n_581), .Y(n_704) );
INVx5_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g622 ( .A(n_451), .B(n_581), .Y(n_622) );
AND2x4_ASAP7_75t_L g636 ( .A(n_451), .B(n_469), .Y(n_636) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_451), .Y(n_640) );
AND2x2_ASAP7_75t_L g660 ( .A(n_451), .B(n_575), .Y(n_660) );
AND2x2_ASAP7_75t_L g710 ( .A(n_451), .B(n_485), .Y(n_710) );
AND2x2_ASAP7_75t_L g720 ( .A(n_451), .B(n_470), .Y(n_720) );
OR2x6_ASAP7_75t_L g451 ( .A(n_452), .B(n_466), .Y(n_451) );
AOI21xp5_ASAP7_75t_SL g452 ( .A1(n_453), .A2(n_457), .B(n_465), .Y(n_452) );
BUFx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx5_ASAP7_75t_L g475 ( .A(n_458), .Y(n_475) );
INVx2_ASAP7_75t_L g464 ( .A(n_462), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_464), .A2(n_491), .B(n_492), .C(n_493), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_L g516 ( .A1(n_464), .A2(n_493), .B(n_517), .C(n_518), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
AND2x2_ASAP7_75t_L g576 ( .A(n_469), .B(n_484), .Y(n_576) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_469), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_469), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g666 ( .A(n_469), .Y(n_666) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g554 ( .A(n_470), .B(n_499), .Y(n_554) );
AND2x2_ASAP7_75t_L g581 ( .A(n_470), .B(n_500), .Y(n_581) );
OA21x2_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B(n_482), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_SL g473 ( .A1(n_474), .A2(n_475), .B(n_476), .C(n_481), .Y(n_473) );
INVx2_ASAP7_75t_L g489 ( .A(n_475), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_L g525 ( .A1(n_475), .A2(n_481), .B(n_526), .C(n_527), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
INVx1_ASAP7_75t_L g494 ( .A(n_481), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_483), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_497), .Y(n_483) );
OR2x2_ASAP7_75t_L g607 ( .A(n_484), .B(n_498), .Y(n_607) );
AND2x2_ASAP7_75t_L g644 ( .A(n_484), .B(n_554), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_484), .B(n_575), .Y(n_655) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_484), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_484), .B(n_611), .Y(n_728) );
INVx5_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx2_ASAP7_75t_L g553 ( .A(n_485), .Y(n_553) );
AND2x2_ASAP7_75t_L g562 ( .A(n_485), .B(n_498), .Y(n_562) );
AND2x2_ASAP7_75t_L g678 ( .A(n_485), .B(n_573), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_485), .B(n_611), .Y(n_700) );
OR2x6_ASAP7_75t_L g485 ( .A(n_486), .B(n_495), .Y(n_485) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_498), .Y(n_646) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_499), .Y(n_598) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx2_ASAP7_75t_L g575 ( .A(n_500), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_507), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_511), .B(n_520), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_511), .B(n_588), .Y(n_707) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_512), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g559 ( .A(n_512), .B(n_560), .Y(n_559) );
INVx5_ASAP7_75t_SL g567 ( .A(n_512), .Y(n_567) );
OR2x2_ASAP7_75t_L g590 ( .A(n_512), .B(n_560), .Y(n_590) );
OR2x2_ASAP7_75t_L g600 ( .A(n_512), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g663 ( .A(n_512), .B(n_522), .Y(n_663) );
AND2x2_ASAP7_75t_SL g701 ( .A(n_512), .B(n_521), .Y(n_701) );
NOR4xp25_ASAP7_75t_L g722 ( .A(n_512), .B(n_643), .C(n_723), .D(n_724), .Y(n_722) );
AND2x2_ASAP7_75t_L g732 ( .A(n_512), .B(n_564), .Y(n_732) );
OR2x6_ASAP7_75t_L g512 ( .A(n_513), .B(n_519), .Y(n_512) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g557 ( .A(n_521), .B(n_553), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_521), .B(n_559), .Y(n_726) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_531), .Y(n_521) );
OR2x2_ASAP7_75t_L g566 ( .A(n_522), .B(n_567), .Y(n_566) );
INVx3_ASAP7_75t_L g573 ( .A(n_522), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_522), .B(n_542), .Y(n_585) );
INVxp67_ASAP7_75t_L g588 ( .A(n_522), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_522), .B(n_560), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_522), .B(n_532), .Y(n_654) );
AND2x2_ASAP7_75t_L g669 ( .A(n_522), .B(n_564), .Y(n_669) );
OR2x2_ASAP7_75t_L g698 ( .A(n_522), .B(n_532), .Y(n_698) );
OA21x2_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_524), .B(n_530), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_531), .B(n_603), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_531), .B(n_567), .Y(n_706) );
OR2x2_ASAP7_75t_L g727 ( .A(n_531), .B(n_604), .Y(n_727) );
INVx1_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
OR2x2_ASAP7_75t_L g541 ( .A(n_532), .B(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g564 ( .A(n_532), .B(n_560), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_532), .B(n_542), .Y(n_579) );
AND2x2_ASAP7_75t_L g649 ( .A(n_532), .B(n_573), .Y(n_649) );
AND2x2_ASAP7_75t_L g683 ( .A(n_532), .B(n_567), .Y(n_683) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_533), .B(n_567), .Y(n_586) );
AND2x2_ASAP7_75t_L g614 ( .A(n_533), .B(n_542), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_540), .B(n_622), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_541), .A2(n_629), .B1(n_665), .B2(n_682), .C(n_684), .Y(n_681) );
INVx5_ASAP7_75t_SL g560 ( .A(n_542), .Y(n_560) );
OAI21xp5_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_545), .B(n_546), .Y(n_543) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
OAI33xp33_ASAP7_75t_L g580 ( .A1(n_553), .A2(n_581), .A3(n_582), .B1(n_584), .B2(n_587), .B3(n_591), .Y(n_580) );
OR2x2_ASAP7_75t_L g596 ( .A(n_553), .B(n_597), .Y(n_596) );
AOI322xp5_ASAP7_75t_L g705 ( .A1(n_553), .A2(n_622), .A3(n_629), .B1(n_706), .B2(n_707), .C1(n_708), .C2(n_711), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_553), .B(n_581), .Y(n_723) );
A2O1A1Ixp33_ASAP7_75t_SL g729 ( .A1(n_553), .A2(n_581), .B(n_730), .C(n_732), .Y(n_729) );
AOI221xp5_ASAP7_75t_L g568 ( .A1(n_554), .A2(n_569), .B1(n_574), .B2(n_577), .C(n_580), .Y(n_568) );
INVx1_ASAP7_75t_L g661 ( .A(n_554), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_554), .B(n_710), .Y(n_709) );
OAI22xp33_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_558), .B1(n_561), .B2(n_563), .Y(n_555) );
INVx1_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g638 ( .A(n_559), .B(n_573), .Y(n_638) );
AND2x2_ASAP7_75t_L g696 ( .A(n_559), .B(n_697), .Y(n_696) );
OR2x2_ASAP7_75t_L g604 ( .A(n_560), .B(n_567), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_560), .B(n_573), .Y(n_632) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_562), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_562), .B(n_640), .Y(n_694) );
OAI321xp33_ASAP7_75t_L g713 ( .A1(n_562), .A2(n_635), .A3(n_714), .B1(n_715), .B2(n_716), .C(n_717), .Y(n_713) );
INVx1_ASAP7_75t_L g680 ( .A(n_563), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_564), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g619 ( .A(n_564), .B(n_567), .Y(n_619) );
AOI321xp33_ASAP7_75t_L g677 ( .A1(n_564), .A2(n_581), .A3(n_678), .B1(n_679), .B2(n_680), .C(n_681), .Y(n_677) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g594 ( .A(n_566), .B(n_579), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_567), .B(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_567), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_567), .B(n_653), .Y(n_690) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x4_ASAP7_75t_L g613 ( .A(n_571), .B(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OR2x2_ASAP7_75t_L g578 ( .A(n_572), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g686 ( .A(n_573), .Y(n_686) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_576), .B(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g609 ( .A(n_581), .Y(n_609) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_583), .B(n_618), .Y(n_667) );
OR2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
OR2x2_ASAP7_75t_L g631 ( .A(n_586), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_SL g676 ( .A(n_586), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_587), .A2(n_634), .B1(n_637), .B2(n_639), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g731 ( .A(n_590), .B(n_654), .Y(n_731) );
AOI221xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_595), .B1(n_599), .B2(n_605), .C(n_608), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
BUFx2_ASAP7_75t_L g629 ( .A(n_598), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_602), .Y(n_599) );
INVx1_ASAP7_75t_SL g675 ( .A(n_601), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_603), .B(n_653), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_603), .A2(n_671), .B(n_673), .Y(n_670) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g716 ( .A(n_604), .B(n_698), .Y(n_716) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx2_ASAP7_75t_SL g618 ( .A(n_607), .Y(n_618) );
AOI21xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B(n_612), .Y(n_608) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g662 ( .A(n_614), .B(n_663), .Y(n_662) );
INVxp67_ASAP7_75t_L g724 ( .A(n_614), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_619), .B(n_620), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_618), .B(n_636), .Y(n_672) );
INVxp67_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g693 ( .A(n_622), .Y(n_693) );
NAND5xp2_ASAP7_75t_L g623 ( .A(n_624), .B(n_641), .C(n_650), .D(n_670), .E(n_677), .Y(n_623) );
O2A1O1Ixp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_627), .B(n_630), .C(n_633), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g665 ( .A(n_629), .Y(n_665) );
CKINVDCx16_ASAP7_75t_R g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_637), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g679 ( .A(n_639), .Y(n_679) );
OAI21xp5_ASAP7_75t_SL g641 ( .A1(n_642), .A2(n_645), .B(n_647), .Y(n_641) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_642), .A2(n_696), .B1(n_699), .B2(n_701), .C(n_702), .Y(n_695) );
AND2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
AOI321xp33_ASAP7_75t_L g650 ( .A1(n_643), .A2(n_651), .A3(n_655), .B1(n_656), .B2(n_662), .C(n_664), .Y(n_650) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g721 ( .A(n_655), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_657), .B(n_661), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g673 ( .A(n_658), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
NOR2xp67_ASAP7_75t_SL g685 ( .A(n_659), .B(n_666), .Y(n_685) );
AOI321xp33_ASAP7_75t_SL g717 ( .A1(n_662), .A2(n_718), .A3(n_719), .B1(n_720), .B2(n_721), .C(n_722), .Y(n_717) );
O2A1O1Ixp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_666), .B(n_667), .C(n_668), .Y(n_664) );
INVx1_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_675), .B(n_683), .Y(n_712) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND3xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .C(n_687), .Y(n_684) );
NOR3xp33_ASAP7_75t_L g688 ( .A(n_689), .B(n_713), .C(n_725), .Y(n_688) );
OAI211xp5_ASAP7_75t_SL g689 ( .A1(n_690), .A2(n_691), .B(n_695), .C(n_705), .Y(n_689) );
INVxp67_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_693), .B(n_694), .Y(n_692) );
OAI221xp5_ASAP7_75t_L g725 ( .A1(n_694), .A2(n_726), .B1(n_727), .B2(n_728), .C(n_729), .Y(n_725) );
INVx1_ASAP7_75t_L g714 ( .A(n_696), .Y(n_714) );
INVx1_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g718 ( .A(n_716), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
CKINVDCx14_ASAP7_75t_R g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
endmodule