module fake_netlist_1_5257_n_806 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_113, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_111, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_112, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_806);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_113;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_112;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_806;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_637;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_659;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_476;
wire n_227;
wire n_384;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_228;
wire n_786;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_769;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_482;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_699;
wire n_519;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_276;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
NOR2xp67_ASAP7_75t_L g114 ( .A(n_11), .B(n_95), .Y(n_114) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_35), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_88), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_71), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_31), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_94), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_65), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_5), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_90), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_112), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_9), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_55), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_45), .Y(n_126) );
INVx1_ASAP7_75t_SL g127 ( .A(n_41), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_78), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_33), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_11), .Y(n_130) );
INVxp67_ASAP7_75t_SL g131 ( .A(n_17), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_97), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_69), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_68), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_17), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_109), .Y(n_136) );
NOR2xp67_ASAP7_75t_L g137 ( .A(n_18), .B(n_62), .Y(n_137) );
CKINVDCx14_ASAP7_75t_R g138 ( .A(n_60), .Y(n_138) );
BUFx3_ASAP7_75t_L g139 ( .A(n_73), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_58), .Y(n_140) );
BUFx10_ASAP7_75t_L g141 ( .A(n_108), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_106), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_84), .Y(n_143) );
CKINVDCx16_ASAP7_75t_R g144 ( .A(n_83), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_43), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_15), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_76), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_6), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_50), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_85), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g151 ( .A(n_113), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g152 ( .A(n_82), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_61), .Y(n_153) );
INVx1_ASAP7_75t_SL g154 ( .A(n_92), .Y(n_154) );
INVxp67_ASAP7_75t_L g155 ( .A(n_27), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_72), .Y(n_156) );
CKINVDCx16_ASAP7_75t_R g157 ( .A(n_99), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_28), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_80), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_37), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_115), .Y(n_161) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_129), .A2(n_0), .B(n_1), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_115), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_121), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_141), .Y(n_165) );
BUFx12f_ASAP7_75t_L g166 ( .A(n_141), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_115), .Y(n_167) );
HB1xp67_ASAP7_75t_L g168 ( .A(n_124), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_124), .Y(n_169) );
AND2x2_ASAP7_75t_L g170 ( .A(n_144), .B(n_0), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_121), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_115), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_119), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_122), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_115), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_141), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_123), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_139), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_129), .B(n_1), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_125), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_139), .Y(n_181) );
CKINVDCx16_ASAP7_75t_R g182 ( .A(n_166), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_178), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_162), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_162), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_165), .B(n_157), .Y(n_186) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_179), .A2(n_148), .B1(n_135), .B2(n_130), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_162), .Y(n_188) );
OAI22xp5_ASAP7_75t_L g189 ( .A1(n_168), .A2(n_146), .B1(n_156), .B2(n_128), .Y(n_189) );
OAI22xp5_ASAP7_75t_L g190 ( .A1(n_168), .A2(n_146), .B1(n_151), .B2(n_152), .Y(n_190) );
NAND3xp33_ASAP7_75t_L g191 ( .A(n_173), .B(n_160), .C(n_116), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_165), .B(n_116), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_165), .B(n_117), .Y(n_193) );
OR2x6_ASAP7_75t_L g194 ( .A(n_166), .B(n_114), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_166), .A2(n_131), .B1(n_117), .B2(n_136), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_178), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_178), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_165), .B(n_155), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_165), .B(n_118), .Y(n_199) );
OR2x6_ASAP7_75t_L g200 ( .A(n_170), .B(n_137), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_178), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_176), .B(n_118), .Y(n_202) );
INVx1_ASAP7_75t_SL g203 ( .A(n_169), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_179), .Y(n_204) );
INVx3_ASAP7_75t_L g205 ( .A(n_179), .Y(n_205) );
AO22x2_ASAP7_75t_L g206 ( .A1(n_179), .A2(n_149), .B1(n_133), .B2(n_134), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g207 ( .A1(n_170), .A2(n_169), .B1(n_179), .B2(n_176), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_178), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_162), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_170), .Y(n_210) );
NAND2xp33_ASAP7_75t_L g211 ( .A(n_173), .B(n_120), .Y(n_211) );
CKINVDCx6p67_ASAP7_75t_R g212 ( .A(n_174), .Y(n_212) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_161), .Y(n_213) );
AO22x1_ASAP7_75t_L g214 ( .A1(n_176), .A2(n_159), .B1(n_158), .B2(n_153), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_205), .A2(n_174), .B(n_180), .C(n_177), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_186), .B(n_176), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_202), .B(n_176), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_206), .A2(n_180), .B1(n_177), .B2(n_162), .Y(n_218) );
BUFx3_ASAP7_75t_L g219 ( .A(n_212), .Y(n_219) );
AOI22x1_ASAP7_75t_L g220 ( .A1(n_184), .A2(n_181), .B1(n_178), .B2(n_175), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_195), .B(n_120), .Y(n_221) );
AOI22xp33_ASAP7_75t_L g222 ( .A1(n_206), .A2(n_162), .B1(n_138), .B2(n_181), .Y(n_222) );
INVxp67_ASAP7_75t_L g223 ( .A(n_189), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_205), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_192), .B(n_136), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_198), .B(n_142), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_212), .B(n_142), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_205), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_187), .B(n_191), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g230 ( .A1(n_206), .A2(n_160), .B1(n_143), .B2(n_145), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_211), .B(n_143), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_207), .B(n_145), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_206), .B(n_164), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_204), .B(n_126), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_184), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_182), .Y(n_236) );
OAI21xp5_ASAP7_75t_L g237 ( .A1(n_185), .A2(n_150), .B(n_147), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_211), .B(n_164), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_193), .B(n_171), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_210), .B(n_171), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_199), .B(n_127), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_209), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_214), .B(n_132), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_214), .B(n_154), .Y(n_244) );
BUFx8_ASAP7_75t_L g245 ( .A(n_185), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_209), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_188), .Y(n_247) );
AND2x6_ASAP7_75t_SL g248 ( .A(n_194), .B(n_2), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_188), .A2(n_181), .B1(n_178), .B2(n_140), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_209), .A2(n_181), .B1(n_178), .B2(n_140), .Y(n_250) );
INVx2_ASAP7_75t_SL g251 ( .A(n_194), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_210), .B(n_181), .Y(n_252) );
BUFx6f_ASAP7_75t_SL g253 ( .A(n_194), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_190), .B(n_181), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_203), .B(n_181), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_183), .B(n_181), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_200), .B(n_167), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_200), .B(n_2), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_194), .B(n_24), .Y(n_259) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_219), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_240), .B(n_200), .Y(n_261) );
AOI21x1_ASAP7_75t_L g262 ( .A1(n_235), .A2(n_183), .B(n_208), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_232), .B(n_200), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_224), .Y(n_264) );
AOI21xp33_ASAP7_75t_L g265 ( .A1(n_223), .A2(n_196), .B(n_197), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_240), .B(n_3), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_235), .A2(n_208), .B(n_201), .Y(n_267) );
INVx3_ASAP7_75t_L g268 ( .A(n_245), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_221), .B(n_3), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_247), .A2(n_201), .B(n_197), .Y(n_270) );
NOR2x1_ASAP7_75t_L g271 ( .A(n_219), .B(n_196), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_247), .A2(n_175), .B(n_167), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_258), .B(n_4), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_229), .B(n_4), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_224), .Y(n_275) );
AND2x4_ASAP7_75t_L g276 ( .A(n_219), .B(n_5), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_233), .B(n_6), .Y(n_277) );
AO22x1_ASAP7_75t_L g278 ( .A1(n_245), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_233), .A2(n_258), .B1(n_245), .B2(n_254), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_227), .B(n_7), .Y(n_280) );
AOI21x1_ASAP7_75t_L g281 ( .A1(n_256), .A2(n_175), .B(n_167), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_242), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_245), .B(n_161), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_251), .B(n_8), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_228), .Y(n_285) );
O2A1O1Ixp33_ASAP7_75t_SL g286 ( .A1(n_218), .A2(n_167), .B(n_175), .C(n_49), .Y(n_286) );
INVx4_ASAP7_75t_L g287 ( .A(n_253), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_216), .B(n_10), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_242), .Y(n_289) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_230), .A2(n_161), .B1(n_163), .B2(n_172), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_242), .A2(n_213), .B(n_172), .Y(n_291) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_236), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g293 ( .A1(n_230), .A2(n_172), .B1(n_163), .B2(n_161), .Y(n_293) );
AOI22xp5_ASAP7_75t_L g294 ( .A1(n_251), .A2(n_172), .B1(n_163), .B2(n_161), .Y(n_294) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_253), .A2(n_172), .B1(n_163), .B2(n_161), .C(n_213), .Y(n_295) );
AND2x6_ASAP7_75t_L g296 ( .A(n_218), .B(n_161), .Y(n_296) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_246), .Y(n_297) );
AND2x2_ASAP7_75t_SL g298 ( .A(n_222), .B(n_259), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_266), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_267), .A2(n_217), .B(n_246), .Y(n_300) );
AOI21x1_ASAP7_75t_SL g301 ( .A1(n_288), .A2(n_252), .B(n_257), .Y(n_301) );
INVx5_ASAP7_75t_L g302 ( .A(n_268), .Y(n_302) );
NOR2xp67_ASAP7_75t_SL g303 ( .A(n_268), .B(n_236), .Y(n_303) );
AOI21xp33_ASAP7_75t_L g304 ( .A1(n_263), .A2(n_225), .B(n_231), .Y(n_304) );
AOI21x1_ASAP7_75t_L g305 ( .A1(n_262), .A2(n_237), .B(n_238), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g306 ( .A1(n_298), .A2(n_237), .B1(n_215), .B2(n_244), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_270), .A2(n_228), .B(n_234), .Y(n_307) );
AOI21xp5_ASAP7_75t_SL g308 ( .A1(n_276), .A2(n_253), .B(n_255), .Y(n_308) );
NOR2xp33_ASAP7_75t_R g309 ( .A(n_268), .B(n_248), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_261), .B(n_239), .Y(n_310) );
O2A1O1Ixp5_ASAP7_75t_SL g311 ( .A1(n_290), .A2(n_243), .B(n_226), .C(n_172), .Y(n_311) );
AO31x2_ASAP7_75t_L g312 ( .A1(n_274), .A2(n_241), .A3(n_220), .B(n_249), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_276), .B(n_250), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_282), .A2(n_220), .B(n_213), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_276), .B(n_248), .Y(n_315) );
OAI22xp5_ASAP7_75t_L g316 ( .A1(n_298), .A2(n_172), .B1(n_163), .B2(n_161), .Y(n_316) );
OAI21x1_ASAP7_75t_L g317 ( .A1(n_291), .A2(n_172), .B(n_163), .Y(n_317) );
A2O1A1Ixp33_ASAP7_75t_L g318 ( .A1(n_274), .A2(n_269), .B(n_284), .C(n_293), .Y(n_318) );
OAI21x1_ASAP7_75t_L g319 ( .A1(n_281), .A2(n_163), .B(n_213), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_263), .B(n_10), .Y(n_320) );
AOI221xp5_ASAP7_75t_SL g321 ( .A1(n_269), .A2(n_163), .B1(n_213), .B2(n_14), .C(n_15), .Y(n_321) );
AO31x2_ASAP7_75t_L g322 ( .A1(n_282), .A2(n_12), .A3(n_13), .B(n_14), .Y(n_322) );
INVx5_ASAP7_75t_L g323 ( .A(n_287), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_273), .B(n_12), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_284), .B(n_13), .Y(n_325) );
BUFx10_ASAP7_75t_L g326 ( .A(n_292), .Y(n_326) );
OAI21x1_ASAP7_75t_L g327 ( .A1(n_301), .A2(n_283), .B(n_289), .Y(n_327) );
OAI21x1_ASAP7_75t_L g328 ( .A1(n_319), .A2(n_283), .B(n_289), .Y(n_328) );
OA21x2_ASAP7_75t_L g329 ( .A1(n_321), .A2(n_265), .B(n_272), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_322), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_323), .B(n_264), .Y(n_331) );
BUFx3_ASAP7_75t_L g332 ( .A(n_323), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_322), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_300), .A2(n_286), .B(n_280), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_318), .A2(n_286), .B(n_275), .Y(n_335) );
CKINVDCx11_ASAP7_75t_R g336 ( .A(n_326), .Y(n_336) );
O2A1O1Ixp33_ASAP7_75t_L g337 ( .A1(n_304), .A2(n_277), .B(n_260), .C(n_285), .Y(n_337) );
OAI21x1_ASAP7_75t_L g338 ( .A1(n_314), .A2(n_271), .B(n_294), .Y(n_338) );
AO31x2_ASAP7_75t_L g339 ( .A1(n_316), .A2(n_296), .A3(n_287), .B(n_278), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_310), .B(n_279), .Y(n_340) );
BUFx6f_ASAP7_75t_L g341 ( .A(n_323), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_299), .B(n_296), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_320), .B(n_287), .Y(n_343) );
BUFx8_ASAP7_75t_L g344 ( .A(n_303), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_322), .Y(n_345) );
OAI21x1_ASAP7_75t_L g346 ( .A1(n_311), .A2(n_295), .B(n_296), .Y(n_346) );
OR2x6_ASAP7_75t_L g347 ( .A(n_308), .B(n_297), .Y(n_347) );
NOR2xp67_ASAP7_75t_SL g348 ( .A(n_302), .B(n_296), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_302), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_307), .Y(n_350) );
BUFx2_ASAP7_75t_L g351 ( .A(n_339), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_342), .B(n_321), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_340), .B(n_315), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_339), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_330), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_330), .Y(n_356) );
INVxp67_ASAP7_75t_SL g357 ( .A(n_348), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_350), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_333), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_350), .Y(n_360) );
CKINVDCx11_ASAP7_75t_R g361 ( .A(n_336), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_347), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_333), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_339), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_345), .Y(n_365) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_339), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_345), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_342), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_327), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_327), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_334), .A2(n_316), .B(n_317), .Y(n_371) );
NAND2xp5_ASAP7_75t_SL g372 ( .A(n_341), .B(n_302), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_328), .Y(n_373) );
AO21x2_ASAP7_75t_L g374 ( .A1(n_335), .A2(n_306), .B(n_305), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_339), .B(n_306), .Y(n_375) );
INVx3_ASAP7_75t_L g376 ( .A(n_341), .Y(n_376) );
INVxp33_ASAP7_75t_L g377 ( .A(n_341), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_328), .Y(n_378) );
AND2x4_ASAP7_75t_L g379 ( .A(n_347), .B(n_296), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_343), .B(n_324), .Y(n_380) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_347), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_375), .B(n_329), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_368), .B(n_332), .Y(n_383) );
NOR2x1_ASAP7_75t_SL g384 ( .A(n_372), .B(n_347), .Y(n_384) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_365), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_375), .B(n_329), .Y(n_386) );
INVx2_ASAP7_75t_SL g387 ( .A(n_362), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_368), .B(n_332), .Y(n_388) );
INVx3_ASAP7_75t_L g389 ( .A(n_362), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_355), .Y(n_390) );
OA21x2_ASAP7_75t_L g391 ( .A1(n_371), .A2(n_346), .B(n_338), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_358), .Y(n_392) );
BUFx2_ASAP7_75t_L g393 ( .A(n_357), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_355), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_375), .B(n_329), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_356), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_358), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_356), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_358), .Y(n_399) );
BUFx2_ASAP7_75t_L g400 ( .A(n_357), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_359), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_359), .B(n_349), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_352), .B(n_337), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_360), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_363), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_365), .B(n_329), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_365), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_360), .B(n_347), .Y(n_408) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_360), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_353), .B(n_326), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_363), .B(n_343), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_376), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_352), .B(n_348), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_367), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_381), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_352), .B(n_346), .Y(n_416) );
BUFx2_ASAP7_75t_L g417 ( .A(n_381), .Y(n_417) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_367), .Y(n_418) );
INVx2_ASAP7_75t_SL g419 ( .A(n_362), .Y(n_419) );
AO31x2_ASAP7_75t_L g420 ( .A1(n_351), .A2(n_325), .A3(n_296), .B(n_312), .Y(n_420) );
AO21x2_ASAP7_75t_L g421 ( .A1(n_371), .A2(n_338), .B(n_313), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_354), .Y(n_422) );
AOI222xp33_ASAP7_75t_L g423 ( .A1(n_353), .A2(n_344), .B1(n_309), .B2(n_331), .C1(n_341), .C2(n_21), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_354), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_351), .B(n_341), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_380), .B(n_331), .Y(n_426) );
AND2x4_ASAP7_75t_SL g427 ( .A(n_376), .B(n_331), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_378), .Y(n_428) );
AND2x4_ASAP7_75t_L g429 ( .A(n_362), .B(n_331), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_364), .B(n_366), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_364), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_385), .B(n_366), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_428), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_416), .B(n_362), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_414), .Y(n_435) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_391), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_416), .B(n_362), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_414), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_416), .B(n_362), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_402), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_411), .B(n_380), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_414), .Y(n_442) );
INVx2_ASAP7_75t_SL g443 ( .A(n_427), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_390), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_382), .B(n_373), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_428), .Y(n_446) );
BUFx3_ASAP7_75t_L g447 ( .A(n_427), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_382), .B(n_373), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_428), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_382), .B(n_374), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_386), .B(n_374), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_386), .B(n_374), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_402), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_392), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_390), .Y(n_455) );
BUFx2_ASAP7_75t_L g456 ( .A(n_393), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_392), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_386), .B(n_374), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_385), .B(n_380), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_394), .Y(n_460) );
AND2x4_ASAP7_75t_L g461 ( .A(n_389), .B(n_379), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_394), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_410), .B(n_361), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_392), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_396), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_396), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_407), .B(n_369), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_395), .B(n_369), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_395), .B(n_370), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_398), .Y(n_470) );
BUFx2_ASAP7_75t_SL g471 ( .A(n_429), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_397), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_395), .B(n_370), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_411), .B(n_376), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_407), .B(n_376), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_398), .Y(n_476) );
OR2x6_ASAP7_75t_SL g477 ( .A(n_426), .B(n_344), .Y(n_477) );
BUFx2_ASAP7_75t_L g478 ( .A(n_393), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_418), .B(n_376), .Y(n_479) );
INVx2_ASAP7_75t_SL g480 ( .A(n_427), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_397), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_413), .B(n_379), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_413), .B(n_379), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_389), .B(n_379), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_413), .B(n_379), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_401), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_401), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_405), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_426), .B(n_377), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_403), .B(n_377), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_397), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_423), .B(n_344), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_403), .B(n_344), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_408), .B(n_378), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_405), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_408), .B(n_378), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_418), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_408), .B(n_371), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_409), .B(n_372), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_409), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_399), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_423), .B(n_297), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_430), .B(n_16), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_383), .B(n_16), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_399), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_399), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_440), .B(n_430), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_433), .Y(n_508) );
INVxp67_ASAP7_75t_L g509 ( .A(n_453), .Y(n_509) );
INVx3_ASAP7_75t_L g510 ( .A(n_447), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_444), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_482), .B(n_425), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_444), .Y(n_513) );
BUFx2_ASAP7_75t_L g514 ( .A(n_477), .Y(n_514) );
NAND2xp33_ASAP7_75t_L g515 ( .A(n_492), .B(n_415), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_434), .B(n_430), .Y(n_516) );
INVxp67_ASAP7_75t_L g517 ( .A(n_477), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_434), .B(n_406), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_455), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_455), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_437), .B(n_439), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_460), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_460), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_503), .B(n_422), .Y(n_524) );
AND3x2_ASAP7_75t_L g525 ( .A(n_456), .B(n_400), .C(n_417), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_462), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_462), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_465), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_482), .B(n_425), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_437), .B(n_406), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_439), .B(n_406), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_465), .Y(n_532) );
INVx2_ASAP7_75t_SL g533 ( .A(n_447), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_433), .Y(n_534) );
CKINVDCx16_ASAP7_75t_R g535 ( .A(n_447), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_450), .B(n_425), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_503), .B(n_422), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_466), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_490), .B(n_424), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_433), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_450), .B(n_389), .Y(n_541) );
INVxp67_ASAP7_75t_SL g542 ( .A(n_456), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_441), .B(n_424), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_466), .Y(n_544) );
AND2x4_ASAP7_75t_L g545 ( .A(n_461), .B(n_389), .Y(n_545) );
AND2x4_ASAP7_75t_L g546 ( .A(n_461), .B(n_387), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_459), .B(n_417), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_470), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_459), .B(n_415), .Y(n_549) );
BUFx2_ASAP7_75t_L g550 ( .A(n_478), .Y(n_550) );
INVx3_ASAP7_75t_R g551 ( .A(n_478), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_432), .B(n_431), .Y(n_552) );
AND3x2_ASAP7_75t_L g553 ( .A(n_463), .B(n_400), .C(n_412), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_432), .B(n_431), .Y(n_554) );
NAND2x1p5_ASAP7_75t_L g555 ( .A(n_443), .B(n_429), .Y(n_555) );
INVxp67_ASAP7_75t_L g556 ( .A(n_493), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_470), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_483), .B(n_429), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_483), .B(n_429), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_446), .Y(n_560) );
INVx3_ASAP7_75t_L g561 ( .A(n_436), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_451), .B(n_387), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_476), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_451), .B(n_387), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_504), .B(n_383), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_452), .B(n_419), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_446), .Y(n_567) );
AND3x2_ASAP7_75t_L g568 ( .A(n_499), .B(n_404), .C(n_384), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_452), .B(n_419), .Y(n_569) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_502), .A2(n_388), .B1(n_419), .B2(n_404), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_445), .B(n_388), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_476), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_474), .B(n_404), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_486), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_486), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_446), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_458), .B(n_421), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_445), .B(n_384), .Y(n_578) );
INVxp67_ASAP7_75t_SL g579 ( .A(n_475), .Y(n_579) );
BUFx2_ASAP7_75t_SL g580 ( .A(n_443), .Y(n_580) );
NAND3xp33_ASAP7_75t_L g581 ( .A(n_497), .B(n_391), .C(n_297), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_449), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_487), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_458), .B(n_421), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_448), .B(n_421), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_498), .B(n_421), .Y(n_586) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_500), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_498), .B(n_391), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_487), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_488), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_479), .B(n_391), .Y(n_591) );
AND2x4_ASAP7_75t_L g592 ( .A(n_461), .B(n_420), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_449), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_485), .B(n_391), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_448), .B(n_420), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_449), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_587), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_521), .B(n_485), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_509), .B(n_497), .Y(n_599) );
INVxp67_ASAP7_75t_L g600 ( .A(n_514), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_550), .Y(n_601) );
AND2x4_ASAP7_75t_L g602 ( .A(n_510), .B(n_461), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_521), .B(n_484), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_587), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_507), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_571), .B(n_468), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_511), .Y(n_607) );
A2O1A1Ixp33_ASAP7_75t_L g608 ( .A1(n_517), .A2(n_480), .B(n_471), .C(n_499), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_536), .B(n_484), .Y(n_609) );
AND2x4_ASAP7_75t_L g610 ( .A(n_510), .B(n_484), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_513), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_595), .B(n_500), .Y(n_612) );
INVx2_ASAP7_75t_SL g613 ( .A(n_535), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_519), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_520), .Y(n_615) );
BUFx2_ASAP7_75t_L g616 ( .A(n_542), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_536), .B(n_484), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_549), .B(n_468), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_516), .B(n_469), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_595), .B(n_469), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_522), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_577), .B(n_473), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_570), .A2(n_480), .B1(n_479), .B2(n_471), .Y(n_623) );
AND2x4_ASAP7_75t_L g624 ( .A(n_510), .B(n_473), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_579), .B(n_475), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_508), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_523), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_577), .B(n_584), .Y(n_628) );
NOR2xp33_ASAP7_75t_SL g629 ( .A(n_580), .B(n_501), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_547), .B(n_494), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_508), .Y(n_631) );
INVx1_ASAP7_75t_SL g632 ( .A(n_533), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_573), .B(n_494), .Y(n_633) );
OR2x2_ASAP7_75t_L g634 ( .A(n_516), .B(n_496), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_526), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_534), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_534), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_584), .B(n_488), .Y(n_638) );
AND2x2_ASAP7_75t_SL g639 ( .A(n_515), .B(n_435), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_588), .B(n_495), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_588), .B(n_495), .Y(n_641) );
AND2x4_ASAP7_75t_L g642 ( .A(n_533), .B(n_496), .Y(n_642) );
NOR2x1_ASAP7_75t_L g643 ( .A(n_515), .B(n_435), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_512), .B(n_438), .Y(n_644) );
AND2x4_ASAP7_75t_L g645 ( .A(n_545), .B(n_438), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_529), .B(n_442), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_527), .Y(n_647) );
INVx2_ASAP7_75t_SL g648 ( .A(n_555), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_558), .B(n_442), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_528), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_532), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_540), .Y(n_652) );
INVx5_ASAP7_75t_L g653 ( .A(n_561), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_559), .B(n_489), .Y(n_654) );
OAI31xp33_ASAP7_75t_L g655 ( .A1(n_565), .A2(n_506), .A3(n_505), .B(n_501), .Y(n_655) );
NAND2x1_ASAP7_75t_L g656 ( .A(n_551), .B(n_505), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_552), .B(n_467), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_586), .B(n_506), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_538), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_562), .B(n_454), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_562), .B(n_454), .Y(n_661) );
NOR5xp2_ASAP7_75t_L g662 ( .A(n_556), .B(n_436), .C(n_420), .D(n_20), .E(n_21), .Y(n_662) );
OR2x6_ASAP7_75t_L g663 ( .A(n_555), .B(n_467), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_540), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_586), .B(n_491), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_544), .B(n_491), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_548), .B(n_491), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_560), .Y(n_668) );
NAND2xp33_ASAP7_75t_SL g669 ( .A(n_578), .B(n_481), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_557), .B(n_481), .Y(n_670) );
NOR2x1p5_ASAP7_75t_L g671 ( .A(n_592), .B(n_436), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_564), .B(n_481), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_565), .B(n_18), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_560), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_592), .B(n_472), .Y(n_675) );
AND2x4_ASAP7_75t_L g676 ( .A(n_545), .B(n_472), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_563), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_564), .B(n_472), .Y(n_678) );
OAI322xp33_ASAP7_75t_L g679 ( .A1(n_600), .A2(n_537), .A3(n_524), .B1(n_543), .B2(n_539), .C1(n_585), .C2(n_591), .Y(n_679) );
BUFx2_ASAP7_75t_L g680 ( .A(n_656), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_640), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_640), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_641), .Y(n_683) );
INVx2_ASAP7_75t_SL g684 ( .A(n_613), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_616), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_641), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_626), .Y(n_687) );
OA21x2_ASAP7_75t_L g688 ( .A1(n_608), .A2(n_581), .B(n_592), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_639), .A2(n_594), .B1(n_541), .B2(n_569), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_603), .B(n_566), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_599), .Y(n_691) );
OAI21xp33_ASAP7_75t_SL g692 ( .A1(n_671), .A2(n_566), .B(n_569), .Y(n_692) );
OR2x2_ASAP7_75t_L g693 ( .A(n_628), .B(n_518), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_673), .A2(n_541), .B1(n_545), .B2(n_546), .Y(n_694) );
OR2x2_ASAP7_75t_L g695 ( .A(n_628), .B(n_518), .Y(n_695) );
OAI22xp33_ASAP7_75t_L g696 ( .A1(n_629), .A2(n_554), .B1(n_553), .B2(n_568), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_597), .Y(n_697) );
AOI222xp33_ASAP7_75t_L g698 ( .A1(n_623), .A2(n_583), .B1(n_575), .B2(n_590), .C1(n_589), .C2(n_574), .Y(n_698) );
INVx1_ASAP7_75t_SL g699 ( .A(n_632), .Y(n_699) );
INVx1_ASAP7_75t_SL g700 ( .A(n_632), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_604), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_655), .B(n_530), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_629), .A2(n_546), .B1(n_553), .B2(n_530), .Y(n_703) );
INVx3_ASAP7_75t_L g704 ( .A(n_663), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_655), .B(n_531), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_657), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_623), .A2(n_546), .B1(n_531), .B2(n_572), .Y(n_707) );
OR2x2_ASAP7_75t_L g708 ( .A(n_612), .B(n_567), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_607), .Y(n_709) );
NOR2xp67_ASAP7_75t_L g710 ( .A(n_653), .B(n_561), .Y(n_710) );
NOR3xp33_ASAP7_75t_SL g711 ( .A(n_669), .B(n_525), .C(n_568), .Y(n_711) );
A2O1A1Ixp33_ASAP7_75t_L g712 ( .A1(n_643), .A2(n_561), .B(n_525), .C(n_582), .Y(n_712) );
AOI22xp33_ASAP7_75t_SL g713 ( .A1(n_624), .A2(n_436), .B1(n_593), .B2(n_582), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_631), .Y(n_714) );
BUFx2_ASAP7_75t_L g715 ( .A(n_663), .Y(n_715) );
BUFx2_ASAP7_75t_L g716 ( .A(n_663), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_638), .B(n_596), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_611), .Y(n_718) );
AOI21xp5_ASAP7_75t_L g719 ( .A1(n_675), .A2(n_596), .B(n_593), .Y(n_719) );
NOR2xp67_ASAP7_75t_L g720 ( .A(n_653), .B(n_576), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_638), .B(n_576), .Y(n_721) );
OAI22xp33_ASAP7_75t_L g722 ( .A1(n_648), .A2(n_567), .B1(n_464), .B2(n_457), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_614), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_615), .Y(n_724) );
OAI222xp33_ASAP7_75t_L g725 ( .A1(n_620), .A2(n_464), .B1(n_457), .B2(n_454), .C1(n_420), .C2(n_436), .Y(n_725) );
NOR2xp33_ASAP7_75t_SL g726 ( .A(n_653), .B(n_464), .Y(n_726) );
AND2x2_ASAP7_75t_L g727 ( .A(n_609), .B(n_457), .Y(n_727) );
OA21x2_ASAP7_75t_L g728 ( .A1(n_665), .A2(n_436), .B(n_420), .Y(n_728) );
OAI32xp33_ASAP7_75t_L g729 ( .A1(n_620), .A2(n_420), .A3(n_20), .B1(n_22), .B2(n_23), .Y(n_729) );
INVxp67_ASAP7_75t_L g730 ( .A(n_601), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_605), .B(n_19), .Y(n_731) );
NAND3xp33_ASAP7_75t_L g732 ( .A(n_662), .B(n_19), .C(n_22), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_715), .A2(n_624), .B1(n_642), .B2(n_618), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g734 ( .A1(n_707), .A2(n_642), .B1(n_612), .B2(n_645), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_681), .Y(n_735) );
AOI322xp5_ASAP7_75t_L g736 ( .A1(n_692), .A2(n_622), .A3(n_619), .B1(n_598), .B2(n_646), .C1(n_644), .C2(n_617), .Y(n_736) );
OAI32xp33_ASAP7_75t_L g737 ( .A1(n_704), .A2(n_625), .A3(n_634), .B1(n_606), .B2(n_622), .Y(n_737) );
NAND3xp33_ASAP7_75t_L g738 ( .A(n_698), .B(n_621), .C(n_677), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_702), .A2(n_645), .B1(n_602), .B2(n_610), .Y(n_739) );
AOI222xp33_ASAP7_75t_L g740 ( .A1(n_705), .A2(n_658), .B1(n_665), .B2(n_627), .C1(n_635), .C2(n_647), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_708), .Y(n_741) );
OAI22xp33_ASAP7_75t_SL g742 ( .A1(n_680), .A2(n_610), .B1(n_602), .B2(n_630), .Y(n_742) );
AOI221xp5_ASAP7_75t_L g743 ( .A1(n_679), .A2(n_658), .B1(n_650), .B2(n_651), .C(n_659), .Y(n_743) );
AOI221xp5_ASAP7_75t_L g744 ( .A1(n_679), .A2(n_649), .B1(n_654), .B2(n_678), .C(n_672), .Y(n_744) );
INVxp33_ASAP7_75t_L g745 ( .A(n_716), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_682), .Y(n_746) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_684), .B(n_633), .Y(n_747) );
NAND3xp33_ASAP7_75t_L g748 ( .A(n_698), .B(n_667), .C(n_666), .Y(n_748) );
NAND4xp25_ASAP7_75t_L g749 ( .A(n_731), .B(n_703), .C(n_732), .D(n_694), .Y(n_749) );
OAI321xp33_ASAP7_75t_L g750 ( .A1(n_696), .A2(n_670), .A3(n_666), .B1(n_667), .B2(n_661), .C(n_660), .Y(n_750) );
NAND3xp33_ASAP7_75t_L g751 ( .A(n_732), .B(n_670), .C(n_674), .Y(n_751) );
AOI21xp5_ASAP7_75t_L g752 ( .A1(n_712), .A2(n_676), .B(n_668), .Y(n_752) );
AOI21xp33_ASAP7_75t_SL g753 ( .A1(n_688), .A2(n_676), .B(n_23), .Y(n_753) );
OAI221xp5_ASAP7_75t_L g754 ( .A1(n_689), .A2(n_664), .B1(n_652), .B2(n_637), .C(n_636), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_683), .B(n_420), .Y(n_755) );
OAI32xp33_ASAP7_75t_L g756 ( .A1(n_704), .A2(n_25), .A3(n_26), .B1(n_29), .B2(n_30), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_686), .Y(n_757) );
OAI21xp5_ASAP7_75t_L g758 ( .A1(n_699), .A2(n_312), .B(n_34), .Y(n_758) );
OAI22xp33_ASAP7_75t_L g759 ( .A1(n_688), .A2(n_297), .B1(n_312), .B2(n_38), .Y(n_759) );
NAND2x1_ASAP7_75t_L g760 ( .A(n_711), .B(n_32), .Y(n_760) );
OAI221xp5_ASAP7_75t_L g761 ( .A1(n_713), .A2(n_36), .B1(n_39), .B2(n_40), .C(n_42), .Y(n_761) );
OAI222xp33_ASAP7_75t_L g762 ( .A1(n_699), .A2(n_44), .B1(n_46), .B2(n_47), .C1(n_48), .C2(n_51), .Y(n_762) );
AOI221xp5_ASAP7_75t_L g763 ( .A1(n_743), .A2(n_725), .B1(n_691), .B2(n_729), .C(n_706), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_740), .B(n_709), .Y(n_764) );
NOR4xp75_ASAP7_75t_L g765 ( .A(n_760), .B(n_717), .C(n_721), .D(n_690), .Y(n_765) );
NOR3xp33_ASAP7_75t_L g766 ( .A(n_753), .B(n_700), .C(n_685), .Y(n_766) );
XOR2xp5_ASAP7_75t_L g767 ( .A(n_749), .B(n_700), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_745), .A2(n_728), .B1(n_730), .B2(n_697), .Y(n_768) );
AOI221xp5_ASAP7_75t_SL g769 ( .A1(n_737), .A2(n_722), .B1(n_718), .B2(n_724), .C(n_723), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_739), .A2(n_693), .B1(n_695), .B2(n_720), .Y(n_770) );
NAND2xp5_ASAP7_75t_SL g771 ( .A(n_742), .B(n_726), .Y(n_771) );
NAND4xp25_ASAP7_75t_L g772 ( .A(n_751), .B(n_726), .C(n_710), .D(n_719), .Y(n_772) );
NOR2x1p5_ASAP7_75t_SL g773 ( .A(n_750), .B(n_714), .Y(n_773) );
A2O1A1Ixp33_ASAP7_75t_L g774 ( .A1(n_736), .A2(n_701), .B(n_727), .C(n_687), .Y(n_774) );
NOR4xp25_ASAP7_75t_L g775 ( .A(n_750), .B(n_728), .C(n_53), .D(n_54), .Y(n_775) );
AOI211xp5_ASAP7_75t_L g776 ( .A1(n_759), .A2(n_52), .B(n_56), .C(n_57), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_748), .B(n_59), .Y(n_777) );
O2A1O1Ixp33_ASAP7_75t_L g778 ( .A1(n_754), .A2(n_63), .B(n_64), .C(n_66), .Y(n_778) );
OAI211xp5_ASAP7_75t_L g779 ( .A1(n_767), .A2(n_734), .B(n_761), .C(n_752), .Y(n_779) );
OAI22xp33_ASAP7_75t_L g780 ( .A1(n_772), .A2(n_733), .B1(n_738), .B2(n_744), .Y(n_780) );
NOR3xp33_ASAP7_75t_SL g781 ( .A(n_771), .B(n_762), .C(n_756), .Y(n_781) );
NOR3xp33_ASAP7_75t_L g782 ( .A(n_777), .B(n_758), .C(n_755), .Y(n_782) );
AOI221xp5_ASAP7_75t_L g783 ( .A1(n_764), .A2(n_757), .B1(n_746), .B2(n_735), .C(n_747), .Y(n_783) );
NOR2x1_ASAP7_75t_SL g784 ( .A(n_770), .B(n_741), .Y(n_784) );
AOI221xp5_ASAP7_75t_L g785 ( .A1(n_769), .A2(n_67), .B1(n_70), .B2(n_74), .C(n_75), .Y(n_785) );
NAND3xp33_ASAP7_75t_L g786 ( .A(n_766), .B(n_77), .C(n_79), .Y(n_786) );
NAND3xp33_ASAP7_75t_L g787 ( .A(n_785), .B(n_766), .C(n_763), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_783), .B(n_774), .Y(n_788) );
NAND3xp33_ASAP7_75t_L g789 ( .A(n_781), .B(n_768), .C(n_775), .Y(n_789) );
NAND4xp25_ASAP7_75t_L g790 ( .A(n_779), .B(n_778), .C(n_776), .D(n_773), .Y(n_790) );
NAND3xp33_ASAP7_75t_L g791 ( .A(n_780), .B(n_765), .C(n_86), .Y(n_791) );
NAND3xp33_ASAP7_75t_L g792 ( .A(n_787), .B(n_786), .C(n_782), .Y(n_792) );
NAND4xp25_ASAP7_75t_L g793 ( .A(n_790), .B(n_784), .C(n_87), .D(n_89), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_789), .Y(n_794) );
AOI21xp5_ASAP7_75t_L g795 ( .A1(n_793), .A2(n_788), .B(n_791), .Y(n_795) );
OAI21xp5_ASAP7_75t_L g796 ( .A1(n_792), .A2(n_81), .B(n_91), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_796), .Y(n_797) );
INVx2_ASAP7_75t_L g798 ( .A(n_795), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_798), .Y(n_799) );
OAI21xp5_ASAP7_75t_SL g800 ( .A1(n_797), .A2(n_794), .B(n_96), .Y(n_800) );
OAI21xp5_ASAP7_75t_L g801 ( .A1(n_800), .A2(n_93), .B(n_98), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_799), .Y(n_802) );
INVxp67_ASAP7_75t_L g803 ( .A(n_802), .Y(n_803) );
OAI222xp33_ASAP7_75t_L g804 ( .A1(n_803), .A2(n_801), .B1(n_101), .B2(n_102), .C1(n_103), .C2(n_104), .Y(n_804) );
AO22x1_ASAP7_75t_L g805 ( .A1(n_804), .A2(n_100), .B1(n_105), .B2(n_107), .Y(n_805) );
AOI21xp5_ASAP7_75t_L g806 ( .A1(n_805), .A2(n_110), .B(n_111), .Y(n_806) );
endmodule