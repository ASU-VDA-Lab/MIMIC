module fake_jpeg_14631_n_326 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_38),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_18),
.Y(n_44)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_41),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_7),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_42),
.B(n_34),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_18),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_44),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_45),
.B(n_28),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_47),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_19),
.B1(n_15),
.B2(n_22),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_49),
.A2(n_22),
.B1(n_20),
.B2(n_28),
.Y(n_83)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_33),
.Y(n_56)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_62),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_19),
.B1(n_20),
.B2(n_15),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_63),
.A2(n_73),
.B1(n_51),
.B2(n_27),
.Y(n_94)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_67),
.Y(n_112)
);

OAI32xp33_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_43),
.A3(n_44),
.B1(n_42),
.B2(n_48),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_66),
.A2(n_58),
.B(n_21),
.C(n_41),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_33),
.Y(n_67)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_49),
.A2(n_36),
.B1(n_40),
.B2(n_35),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_72),
.A2(n_79),
.B1(n_57),
.B2(n_55),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_47),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

AND2x4_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_58),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_84),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_39),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_39),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_40),
.B1(n_35),
.B2(n_37),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_82),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g101 ( 
.A1(n_83),
.A2(n_56),
.B1(n_46),
.B2(n_59),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_85),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_52),
.B(n_27),
.Y(n_86)
);

NAND3xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_25),
.C(n_29),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_98),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_52),
.B(n_38),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_106),
.Y(n_132)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_93),
.A2(n_96),
.B1(n_103),
.B2(n_76),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_75),
.A2(n_46),
.B1(n_37),
.B2(n_35),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_75),
.A2(n_56),
.B1(n_51),
.B2(n_65),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_97),
.A2(n_101),
.B1(n_76),
.B2(n_85),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_66),
.Y(n_102)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_75),
.A2(n_38),
.B1(n_46),
.B2(n_56),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_39),
.Y(n_107)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

AO22x1_ASAP7_75t_L g109 ( 
.A1(n_72),
.A2(n_59),
.B1(n_58),
.B2(n_47),
.Y(n_109)
);

AND2x4_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_79),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_60),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_105),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_L g114 ( 
.A1(n_80),
.A2(n_54),
.B1(n_58),
.B2(n_47),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_114),
.A2(n_73),
.B1(n_69),
.B2(n_64),
.Y(n_129)
);

INVx4_ASAP7_75t_SL g115 ( 
.A(n_87),
.Y(n_115)
);

INVxp67_ASAP7_75t_SL g143 ( 
.A(n_115),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_102),
.A2(n_106),
.B1(n_107),
.B2(n_90),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_117),
.A2(n_119),
.B1(n_91),
.B2(n_104),
.Y(n_156)
);

OAI21x1_ASAP7_75t_SL g140 ( 
.A1(n_118),
.A2(n_109),
.B(n_130),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_106),
.A2(n_78),
.B1(n_60),
.B2(n_64),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_113),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_120),
.B(n_123),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_109),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_127),
.B(n_135),
.Y(n_149)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_129),
.A2(n_130),
.B1(n_138),
.B2(n_100),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_93),
.A2(n_70),
.B1(n_69),
.B2(n_61),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_92),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_92),
.A2(n_81),
.B1(n_77),
.B2(n_31),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_136),
.A2(n_81),
.B(n_110),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_89),
.A2(n_54),
.B1(n_68),
.B2(n_62),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_140),
.A2(n_162),
.B(n_168),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_99),
.Y(n_141)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_99),
.C(n_111),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_142),
.B(n_151),
.C(n_158),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_132),
.B(n_99),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_167),
.Y(n_182)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_145),
.B(n_146),
.Y(n_190)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_147),
.A2(n_121),
.B1(n_13),
.B2(n_2),
.Y(n_183)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_105),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_153),
.A2(n_155),
.B1(n_160),
.B2(n_161),
.Y(n_170)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_154),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_91),
.B1(n_104),
.B2(n_100),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_156),
.B(n_17),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_113),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_165),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_41),
.C(n_81),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_138),
.B(n_108),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_159),
.B(n_26),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_118),
.A2(n_95),
.B1(n_87),
.B2(n_88),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_118),
.A2(n_88),
.B1(n_62),
.B2(n_2),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_13),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_164),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_25),
.Y(n_165)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_116),
.B(n_21),
.Y(n_167)
);

AND2x4_ASAP7_75t_SL g169 ( 
.A(n_149),
.B(n_137),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_169),
.A2(n_175),
.B(n_151),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_124),
.B1(n_122),
.B2(n_116),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_174),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_157),
.A2(n_137),
.B(n_120),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_176),
.Y(n_221)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_165),
.A2(n_129),
.B1(n_115),
.B2(n_85),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_179),
.A2(n_191),
.B1(n_158),
.B2(n_142),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_163),
.A2(n_115),
.B1(n_16),
.B2(n_17),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_194),
.B1(n_12),
.B2(n_14),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_183),
.A2(n_187),
.B1(n_188),
.B2(n_195),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_139),
.B(n_121),
.Y(n_184)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_184),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_29),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_193),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_147),
.A2(n_71),
.B1(n_110),
.B2(n_3),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_147),
.A2(n_71),
.B1(n_110),
.B2(n_3),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_163),
.A2(n_30),
.B1(n_31),
.B2(n_16),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_141),
.B(n_162),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_17),
.B1(n_30),
.B2(n_21),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_162),
.A2(n_10),
.B1(n_14),
.B2(n_3),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_144),
.B(n_29),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_29),
.C(n_25),
.Y(n_217)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_198),
.B(n_199),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_200),
.B(n_8),
.Y(n_227)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_143),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_201),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_172),
.A2(n_155),
.B1(n_160),
.B2(n_168),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_203),
.A2(n_212),
.B1(n_200),
.B2(n_188),
.Y(n_231)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_205),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_156),
.Y(n_208)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_208),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_210),
.B(n_227),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_171),
.A2(n_167),
.B(n_1),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_211),
.A2(n_216),
.B(n_187),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_172),
.A2(n_175),
.B1(n_173),
.B2(n_170),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_213),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_29),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_191),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_171),
.A2(n_0),
.B(n_1),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_220),
.C(n_222),
.Y(n_247)
);

OAI21xp33_ASAP7_75t_L g218 ( 
.A1(n_169),
.A2(n_9),
.B(n_3),
.Y(n_218)
);

NOR3xp33_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_228),
.C(n_195),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_173),
.A2(n_178),
.B1(n_179),
.B2(n_201),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_224),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_182),
.B(n_25),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_26),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_178),
.B(n_26),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_198),
.Y(n_234)
);

BUFx5_ASAP7_75t_L g226 ( 
.A(n_192),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_226),
.Y(n_236)
);

AOI21xp33_ASAP7_75t_L g228 ( 
.A1(n_193),
.A2(n_8),
.B(n_4),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_231),
.A2(n_233),
.B1(n_235),
.B2(n_241),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_203),
.A2(n_185),
.B1(n_192),
.B2(n_181),
.Y(n_233)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_209),
.A2(n_185),
.B1(n_181),
.B2(n_176),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_196),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_240),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_190),
.Y(n_238)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_238),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_197),
.Y(n_239)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_186),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_189),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_249),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_183),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_247),
.C(n_217),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_216),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_256),
.C(n_263),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_245),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_222),
.Y(n_253)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_233),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_232),
.A2(n_223),
.B(n_208),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_257),
.A2(n_261),
.B1(n_248),
.B2(n_221),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_230),
.A2(n_219),
.B1(n_210),
.B2(n_206),
.Y(n_258)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_258),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_225),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_260),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_231),
.A2(n_213),
.B(n_206),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_205),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_214),
.Y(n_264)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

AOI22x1_ASAP7_75t_L g265 ( 
.A1(n_248),
.A2(n_246),
.B1(n_202),
.B2(n_249),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_265),
.A2(n_243),
.B1(n_226),
.B2(n_242),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_211),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_4),
.C(n_5),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_265),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_281),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_273),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_266),
.A2(n_229),
.B1(n_247),
.B2(n_204),
.Y(n_275)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_265),
.A2(n_221),
.B1(n_214),
.B2(n_202),
.Y(n_276)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_277),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_259),
.A2(n_243),
.B1(n_242),
.B2(n_227),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_261),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_255),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_250),
.C(n_263),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_283),
.B(n_289),
.Y(n_302)
);

NOR2xp67_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_262),
.Y(n_286)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_286),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_293),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_251),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_269),
.A2(n_257),
.B1(n_256),
.B2(n_252),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_291),
.A2(n_273),
.B1(n_278),
.B2(n_270),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_258),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_254),
.C(n_267),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_284),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_254),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_305),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_295),
.A2(n_269),
.B1(n_274),
.B2(n_277),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_299),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_300),
.B(n_303),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_285),
.A2(n_279),
.B(n_281),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_301),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_290),
.A2(n_280),
.B1(n_7),
.B2(n_8),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_288),
.B1(n_284),
.B2(n_283),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_6),
.Y(n_309)
);

AOI31xp33_ASAP7_75t_L g306 ( 
.A1(n_297),
.A2(n_288),
.A3(n_291),
.B(n_287),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_306),
.B(n_309),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_6),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_308),
.B(n_312),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_310),
.A2(n_301),
.B1(n_296),
.B2(n_12),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_302),
.B(n_7),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_305),
.C(n_298),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_316),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_311),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_318),
.A2(n_307),
.B(n_313),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_319),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_314),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_308),
.B(n_310),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_10),
.B(n_11),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_13),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_325),
.A2(n_10),
.B1(n_11),
.B2(n_307),
.Y(n_326)
);


endmodule