module fake_jpeg_12234_n_562 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_562);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_562;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_17),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx11_ASAP7_75t_L g169 ( 
.A(n_58),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_59),
.Y(n_201)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_61),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_62),
.Y(n_205)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_63),
.Y(n_174)
);

INVxp67_ASAP7_75t_SL g64 ( 
.A(n_24),
.Y(n_64)
);

CKINVDCx6p67_ASAP7_75t_R g159 ( 
.A(n_64),
.Y(n_159)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_66),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_19),
.B(n_18),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_67),
.B(n_73),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_68),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_19),
.B(n_16),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_69),
.B(n_13),
.Y(n_145)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_70),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_20),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_75),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_20),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_76),
.B(n_99),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_78),
.Y(n_197)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_79),
.Y(n_160)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_82),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_83),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_40),
.B(n_0),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_84),
.B(n_95),
.C(n_103),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_85),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_86),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_87),
.Y(n_210)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_88),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_89),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_90),
.Y(n_143)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_91),
.Y(n_208)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_21),
.B(n_15),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_93),
.B(n_98),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_94),
.Y(n_148)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_40),
.B(n_0),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_96),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_21),
.B(n_14),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_41),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_100),
.B(n_101),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_41),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_40),
.B(n_0),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_32),
.B(n_14),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_105),
.B(n_108),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_106),
.B(n_110),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_107),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_51),
.B(n_40),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_109),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_51),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_40),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_111),
.B(n_46),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_38),
.B(n_13),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_112),
.B(n_3),
.Y(n_200)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_25),
.Y(n_113)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_113),
.Y(n_188)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_52),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_42),
.Y(n_134)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_117),
.Y(n_180)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_24),
.Y(n_118)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_118),
.Y(n_182)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_29),
.Y(n_119)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_119),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_29),
.Y(n_120)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_120),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_29),
.Y(n_121)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_121),
.Y(n_194)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_25),
.Y(n_122)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_122),
.Y(n_196)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_34),
.Y(n_123)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_123),
.Y(n_199)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_34),
.Y(n_124)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_124),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_34),
.Y(n_125)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_125),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_58),
.B(n_38),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_126),
.B(n_136),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_59),
.A2(n_46),
.B1(n_42),
.B2(n_38),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_129),
.A2(n_141),
.B1(n_156),
.B2(n_168),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_92),
.A2(n_57),
.B1(n_56),
.B2(n_53),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_131),
.A2(n_133),
.B1(n_167),
.B2(n_187),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_87),
.A2(n_57),
.B1(n_56),
.B2(n_53),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_134),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_70),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_135),
.B(n_149),
.Y(n_236)
);

NOR2x1_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_50),
.Y(n_136)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_84),
.B(n_42),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_139),
.B(n_185),
.C(n_207),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_94),
.A2(n_46),
.B1(n_43),
.B2(n_49),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_145),
.B(n_4),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_115),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_97),
.A2(n_26),
.B1(n_49),
.B2(n_44),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_60),
.B(n_30),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_157),
.B(n_163),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_118),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_161),
.B(n_166),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_95),
.B(n_30),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_164),
.B(n_173),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_103),
.B(n_54),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_64),
.A2(n_50),
.B1(n_54),
.B2(n_44),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_104),
.A2(n_43),
.B1(n_39),
.B2(n_28),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_89),
.B(n_39),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_109),
.A2(n_28),
.B1(n_26),
.B2(n_12),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_181),
.A2(n_203),
.B1(n_209),
.B2(n_140),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_116),
.B(n_1),
.C(n_2),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_65),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_63),
.B(n_1),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_192),
.B(n_200),
.Y(n_249)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_124),
.Y(n_195)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_107),
.Y(n_202)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_62),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_203)
);

NAND2x1_ASAP7_75t_L g207 ( 
.A(n_119),
.B(n_123),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_66),
.A2(n_11),
.B1(n_5),
.B2(n_7),
.Y(n_209)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_169),
.Y(n_212)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_212),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_4),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_214),
.B(n_228),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_215),
.B(n_248),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_157),
.A2(n_72),
.B1(n_82),
.B2(n_77),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_217),
.A2(n_272),
.B1(n_275),
.B2(n_282),
.Y(n_326)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_144),
.Y(n_218)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_218),
.Y(n_286)
);

AOI22x1_ASAP7_75t_L g219 ( 
.A1(n_129),
.A2(n_68),
.B1(n_71),
.B2(n_125),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_219),
.A2(n_220),
.B(n_264),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_L g220 ( 
.A1(n_187),
.A2(n_121),
.B1(n_120),
.B2(n_102),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_220),
.A2(n_244),
.B1(n_263),
.B2(n_234),
.Y(n_311)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_221),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_222),
.Y(n_299)
);

INVx11_ASAP7_75t_L g225 ( 
.A(n_169),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g323 ( 
.A(n_225),
.Y(n_323)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_148),
.Y(n_227)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_227),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_164),
.B(n_4),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_139),
.B(n_7),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_230),
.B(n_258),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_134),
.A2(n_85),
.B1(n_83),
.B2(n_78),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_231),
.B(n_234),
.Y(n_333)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_153),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_232),
.B(n_235),
.Y(n_284)
);

AND2x2_ASAP7_75t_SL g234 ( 
.A(n_138),
.B(n_89),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_127),
.B(n_80),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_172),
.B(n_88),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_237),
.B(n_246),
.Y(n_319)
);

AND2x2_ASAP7_75t_SL g238 ( 
.A(n_142),
.B(n_100),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_238),
.B(n_255),
.Y(n_302)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_146),
.Y(n_239)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_239),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_177),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_240),
.Y(n_324)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_152),
.Y(n_242)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_242),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_243),
.Y(n_329)
);

OAI22xp33_ASAP7_75t_L g244 ( 
.A1(n_133),
.A2(n_131),
.B1(n_167),
.B2(n_126),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_170),
.Y(n_245)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_245),
.Y(n_336)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_174),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_137),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_154),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_251),
.B(n_252),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_150),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_198),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_253),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_160),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_254),
.B(n_257),
.Y(n_304)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_175),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_176),
.A2(n_91),
.B1(n_106),
.B2(n_100),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_256),
.A2(n_266),
.B1(n_280),
.B2(n_281),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_132),
.B(n_106),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_188),
.B(n_10),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_186),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_259),
.B(n_262),
.Y(n_325)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_165),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_260),
.B(n_265),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_192),
.B(n_11),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_261),
.B(n_264),
.Y(n_332)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_206),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_128),
.A2(n_211),
.B1(n_204),
.B2(n_143),
.Y(n_263)
);

A2O1A1Ixp33_ASAP7_75t_L g264 ( 
.A1(n_136),
.A2(n_207),
.B(n_158),
.C(n_159),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_159),
.B(n_190),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_176),
.A2(n_155),
.B1(n_191),
.B2(n_162),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_140),
.A2(n_198),
.B1(n_204),
.B2(n_128),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_267),
.A2(n_269),
.B1(n_271),
.B2(n_231),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_159),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_268),
.B(n_276),
.Y(n_330)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_199),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_270),
.B(n_273),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_205),
.A2(n_197),
.B1(n_208),
.B2(n_130),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_205),
.A2(n_130),
.B1(n_208),
.B2(n_179),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_180),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_189),
.B(n_194),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_274),
.B(n_279),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_147),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_275),
.Y(n_294)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_179),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_193),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_277),
.Y(n_307)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_171),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_278),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_193),
.B(n_191),
.Y(n_279)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_162),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_158),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_210),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_282),
.A2(n_268),
.B1(n_253),
.B2(n_275),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_182),
.B(n_178),
.Y(n_283)
);

OAI21xp33_ASAP7_75t_L g316 ( 
.A1(n_283),
.A2(n_221),
.B(n_238),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_219),
.A2(n_147),
.B1(n_151),
.B2(n_183),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_287),
.A2(n_305),
.B1(n_318),
.B2(n_321),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_269),
.A2(n_151),
.B1(n_183),
.B2(n_210),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_288),
.A2(n_290),
.B1(n_292),
.B2(n_317),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_229),
.A2(n_241),
.B1(n_216),
.B2(n_250),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_241),
.B(n_214),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_291),
.B(n_297),
.C(n_298),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_230),
.B(n_228),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_226),
.B(n_233),
.C(n_274),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_301),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_226),
.B(n_251),
.C(n_224),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_303),
.B(n_308),
.C(n_327),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_219),
.A2(n_244),
.B1(n_263),
.B2(n_247),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g355 ( 
.A(n_306),
.B(n_311),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_258),
.B(n_261),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_316),
.B(n_333),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_229),
.A2(n_249),
.B1(n_236),
.B2(n_273),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_234),
.A2(n_238),
.B1(n_270),
.B2(n_245),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_227),
.A2(n_242),
.B1(n_255),
.B2(n_218),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_326),
.A2(n_331),
.B1(n_294),
.B2(n_325),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_223),
.B(n_213),
.C(n_262),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g328 ( 
.A1(n_259),
.A2(n_246),
.B1(n_239),
.B2(n_243),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_328),
.A2(n_335),
.B1(n_326),
.B2(n_318),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_277),
.A2(n_225),
.B(n_280),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_334),
.A2(n_295),
.B(n_302),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_222),
.A2(n_250),
.B1(n_244),
.B2(n_217),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_212),
.A2(n_250),
.B1(n_241),
.B2(n_251),
.Y(n_337)
);

AOI31xp33_ASAP7_75t_SL g375 ( 
.A1(n_337),
.A2(n_294),
.A3(n_327),
.B(n_309),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_310),
.B(n_308),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_338),
.B(n_340),
.Y(n_386)
);

BUFx24_ASAP7_75t_SL g339 ( 
.A(n_293),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_339),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_310),
.B(n_290),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_343),
.A2(n_345),
.B(n_364),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_317),
.A2(n_288),
.B1(n_292),
.B2(n_335),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_344),
.A2(n_360),
.B1(n_321),
.B2(n_323),
.Y(n_384)
);

XOR2x2_ASAP7_75t_SL g346 ( 
.A(n_337),
.B(n_297),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_346),
.B(n_359),
.C(n_376),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_315),
.B(n_319),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_347),
.B(n_354),
.Y(n_400)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_296),
.Y(n_348)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_348),
.Y(n_381)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_296),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_286),
.Y(n_351)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_351),
.Y(n_398)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_320),
.Y(n_352)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_352),
.Y(n_401)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_320),
.Y(n_353)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_353),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_315),
.B(n_319),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_320),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_356),
.B(n_365),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_291),
.B(n_300),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_332),
.A2(n_305),
.B1(n_311),
.B2(n_302),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_286),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_362),
.A2(n_366),
.B1(n_331),
.B2(n_323),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_332),
.B(n_284),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_363),
.B(n_377),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_302),
.A2(n_333),
.B(n_334),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_314),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_284),
.A2(n_298),
.B1(n_303),
.B2(n_300),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_325),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_367),
.B(n_368),
.Y(n_389)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_314),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_336),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_369),
.B(n_371),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_304),
.B(n_322),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_370),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_325),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_372),
.A2(n_375),
.B(n_307),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_330),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_373),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_285),
.B(n_309),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_374),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_324),
.B(n_336),
.C(n_313),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_312),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_313),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_378),
.B(n_307),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_379),
.A2(n_390),
.B1(n_397),
.B2(n_383),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_352),
.B(n_353),
.Y(n_383)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_383),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_384),
.A2(n_408),
.B1(n_341),
.B2(n_348),
.Y(n_429)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_387),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_338),
.B(n_324),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_388),
.B(n_349),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g390 ( 
.A(n_360),
.B(n_289),
.Y(n_390)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_390),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_391),
.A2(n_394),
.B(n_395),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_364),
.A2(n_323),
.B(n_312),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_343),
.A2(n_329),
.B(n_289),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_355),
.A2(n_329),
.B(n_299),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_396),
.B(n_410),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_376),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_397),
.B(n_407),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_355),
.A2(n_299),
.B(n_340),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_405),
.B(n_356),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_359),
.B(n_349),
.C(n_346),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_406),
.B(n_357),
.C(n_366),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_351),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_342),
.A2(n_344),
.B1(n_372),
.B2(n_375),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_367),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_411),
.B(n_380),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_412),
.A2(n_416),
.B(n_419),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_387),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_414),
.B(n_415),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_379),
.A2(n_342),
.B1(n_347),
.B2(n_354),
.Y(n_415)
);

OAI22x1_ASAP7_75t_L g416 ( 
.A1(n_390),
.A2(n_341),
.B1(n_362),
.B2(n_358),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_387),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_417),
.B(n_418),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_387),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_399),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_399),
.Y(n_420)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_420),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_406),
.B(n_357),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_422),
.B(n_423),
.C(n_427),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_400),
.B(n_363),
.Y(n_424)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_424),
.Y(n_451)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_398),
.Y(n_425)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_425),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_406),
.B(n_358),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_429),
.A2(n_435),
.B1(n_438),
.B2(n_383),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_400),
.B(n_350),
.Y(n_430)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_430),
.Y(n_455)
);

OA21x2_ASAP7_75t_L g431 ( 
.A1(n_408),
.A2(n_378),
.B(n_361),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_431),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_392),
.B(n_377),
.Y(n_434)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_434),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_384),
.A2(n_408),
.B1(n_405),
.B2(n_403),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_389),
.Y(n_436)
);

INVxp33_ASAP7_75t_SL g461 ( 
.A(n_436),
.Y(n_461)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_381),
.Y(n_437)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_437),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_379),
.A2(n_390),
.B1(n_405),
.B2(n_404),
.Y(n_438)
);

FAx1_ASAP7_75t_SL g439 ( 
.A(n_386),
.B(n_380),
.CI(n_404),
.CON(n_439),
.SN(n_439)
);

NOR2xp67_ASAP7_75t_L g458 ( 
.A(n_439),
.B(n_403),
.Y(n_458)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_440),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_441),
.B(n_445),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_443),
.A2(n_444),
.B1(n_467),
.B2(n_431),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_435),
.A2(n_395),
.B1(n_386),
.B2(n_383),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_422),
.B(n_380),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_423),
.B(n_388),
.C(n_382),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_447),
.B(n_448),
.C(n_449),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_411),
.B(n_388),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_427),
.B(n_382),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_413),
.B(n_391),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_450),
.B(n_452),
.C(n_463),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_415),
.B(n_385),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_458),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_419),
.A2(n_409),
.B1(n_392),
.B2(n_402),
.Y(n_459)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_459),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_424),
.B(n_430),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_421),
.B(n_385),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_466),
.B(n_426),
.C(n_389),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_429),
.A2(n_395),
.B1(n_401),
.B2(n_384),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_456),
.B(n_393),
.Y(n_470)
);

CKINVDCx14_ASAP7_75t_R g502 ( 
.A(n_470),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_461),
.B(n_420),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_471),
.B(n_472),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_450),
.B(n_436),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_460),
.Y(n_473)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_473),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_453),
.A2(n_438),
.B1(n_433),
.B2(n_432),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_474),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_476),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_477),
.B(n_490),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_442),
.B(n_445),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_478),
.B(n_484),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_446),
.A2(n_428),
.B(n_433),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_479),
.B(n_481),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_442),
.B(n_432),
.C(n_418),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_480),
.B(n_486),
.C(n_452),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_464),
.A2(n_431),
.B1(n_412),
.B2(n_421),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_463),
.B(n_437),
.Y(n_483)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_483),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_455),
.B(n_417),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_SL g485 ( 
.A(n_448),
.B(n_439),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_485),
.B(n_466),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_441),
.B(n_447),
.C(n_449),
.Y(n_486)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_460),
.Y(n_488)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_488),
.Y(n_500)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_460),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_489),
.B(n_407),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_453),
.A2(n_401),
.B1(n_414),
.B2(n_416),
.Y(n_490)
);

BUFx24_ASAP7_75t_SL g494 ( 
.A(n_487),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_494),
.B(n_468),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_495),
.B(n_480),
.Y(n_519)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_497),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_487),
.B(n_451),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_501),
.B(n_503),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_478),
.B(n_465),
.C(n_462),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_477),
.B(n_439),
.Y(n_504)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_504),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_507),
.B(n_482),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_509),
.B(n_517),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_493),
.B(n_484),
.Y(n_510)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_510),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_505),
.A2(n_479),
.B(n_446),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_511),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_491),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g533 ( 
.A(n_512),
.B(n_513),
.Y(n_533)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_496),
.B(n_428),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_514),
.B(n_515),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g515 ( 
.A(n_503),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_500),
.B(n_454),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_519),
.B(n_506),
.C(n_482),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_495),
.B(n_475),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_520),
.B(n_521),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_502),
.B(n_475),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_522),
.B(n_523),
.Y(n_535)
);

BUFx24_ASAP7_75t_SL g523 ( 
.A(n_516),
.Y(n_523)
);

INVx6_ASAP7_75t_L g527 ( 
.A(n_518),
.Y(n_527)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_527),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_520),
.B(n_499),
.C(n_506),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_529),
.B(n_530),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_519),
.B(n_486),
.C(n_469),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_509),
.B(n_469),
.C(n_505),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_532),
.B(n_485),
.Y(n_538)
);

INVxp33_ASAP7_75t_L g534 ( 
.A(n_531),
.Y(n_534)
);

AOI21xp33_ASAP7_75t_L g547 ( 
.A1(n_534),
.A2(n_525),
.B(n_536),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_SL g543 ( 
.A(n_538),
.B(n_539),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_527),
.B(n_508),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_528),
.B(n_511),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_540),
.Y(n_546)
);

NOR2xp67_ASAP7_75t_SL g541 ( 
.A(n_524),
.B(n_507),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_541),
.A2(n_528),
.B(n_514),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_526),
.A2(n_492),
.B1(n_498),
.B2(n_500),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_542),
.B(n_510),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g554 ( 
.A1(n_544),
.A2(n_547),
.B(n_517),
.Y(n_554)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_545),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_535),
.B(n_525),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_548),
.B(n_549),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_537),
.B(n_533),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_546),
.B(n_534),
.C(n_540),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_550),
.B(n_552),
.Y(n_556)
);

INVxp33_ASAP7_75t_L g552 ( 
.A(n_543),
.Y(n_552)
);

A2O1A1O1Ixp25_ASAP7_75t_L g555 ( 
.A1(n_554),
.A2(n_546),
.B(n_553),
.C(n_551),
.D(n_396),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g559 ( 
.A1(n_555),
.A2(n_557),
.B(n_492),
.Y(n_559)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_551),
.Y(n_557)
);

OAI31xp33_ASAP7_75t_SL g558 ( 
.A1(n_556),
.A2(n_474),
.A3(n_481),
.B(n_444),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_558),
.A2(n_559),
.B1(n_467),
.B2(n_457),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_560),
.B(n_476),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_561),
.B(n_394),
.Y(n_562)
);


endmodule