module fake_netlist_6_2760_n_1805 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_442, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_67, n_15, n_443, n_246, n_38, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_397, n_155, n_109, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_414, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_363, n_395, n_323, n_393, n_411, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_102, n_204, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_433, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_328, n_429, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_64, n_288, n_427, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1805);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_397;
input n_155;
input n_109;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_102;
input n_204;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_433;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_328;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_64;
input n_288;
input n_427;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1805;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_1380;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_830;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_564;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_932;
wire n_1697;
wire n_979;
wire n_905;
wire n_1680;
wire n_993;
wire n_689;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_1386;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_811;
wire n_527;
wire n_683;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_1466;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_1060;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_1681;
wire n_520;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_1745;
wire n_914;
wire n_759;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_607;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1095;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_621;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_1361;
wire n_1491;
wire n_662;
wire n_1152;
wire n_1705;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_1222;
wire n_599;
wire n_776;
wire n_1720;
wire n_934;
wire n_482;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_799;
wire n_1548;
wire n_1155;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_1047;
wire n_1385;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_1276;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_1582;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1525;
wire n_1585;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_570;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1632;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_456),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_408),
.Y(n_464)
);

BUFx10_ASAP7_75t_L g465 ( 
.A(n_4),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_178),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_270),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_441),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_453),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_101),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_366),
.Y(n_471)
);

CKINVDCx14_ASAP7_75t_R g472 ( 
.A(n_401),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_172),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_341),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_36),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_403),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_49),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_340),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_30),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_156),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_82),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_255),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_232),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_84),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_244),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_33),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_123),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_254),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_182),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_225),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_445),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_47),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_356),
.Y(n_493)
);

BUFx10_ASAP7_75t_L g494 ( 
.A(n_457),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_234),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_189),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_450),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_425),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_387),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_91),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_253),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_167),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_302),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_337),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_301),
.Y(n_505)
);

BUFx10_ASAP7_75t_L g506 ( 
.A(n_368),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_396),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_295),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_306),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_446),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_311),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_93),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_398),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_364),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_280),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_31),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_404),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_386),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_266),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_179),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_336),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_352),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_71),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_134),
.Y(n_524)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_44),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_77),
.Y(n_526)
);

BUFx10_ASAP7_75t_L g527 ( 
.A(n_36),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_191),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_433),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_414),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_346),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_113),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_185),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_13),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_98),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_201),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_154),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_60),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_140),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_330),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_95),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_419),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_209),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_357),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_16),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_94),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_411),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_62),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_197),
.Y(n_549)
);

BUFx2_ASAP7_75t_SL g550 ( 
.A(n_233),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_130),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_444),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_328),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_360),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_451),
.Y(n_555)
);

CKINVDCx16_ASAP7_75t_R g556 ( 
.A(n_315),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_23),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_63),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_429),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_53),
.Y(n_560)
);

CKINVDCx16_ASAP7_75t_R g561 ( 
.A(n_460),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_43),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_314),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_384),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_442),
.Y(n_565)
);

BUFx8_ASAP7_75t_SL g566 ( 
.A(n_84),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_64),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_417),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_213),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_392),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_89),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_344),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_80),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_407),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_138),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_436),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_40),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_200),
.Y(n_578)
);

CKINVDCx16_ASAP7_75t_R g579 ( 
.A(n_153),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_348),
.Y(n_580)
);

BUFx10_ASAP7_75t_L g581 ( 
.A(n_265),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_281),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_219),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_420),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_402),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_124),
.Y(n_586)
);

BUFx10_ASAP7_75t_L g587 ( 
.A(n_30),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_13),
.Y(n_588)
);

CKINVDCx16_ASAP7_75t_R g589 ( 
.A(n_52),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_114),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_347),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_167),
.Y(n_592)
);

INVx2_ASAP7_75t_R g593 ( 
.A(n_210),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_106),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_262),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_55),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_100),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_247),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_79),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_6),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_141),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_440),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_351),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_173),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_145),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_197),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_293),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_195),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_125),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_145),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_251),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_69),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_355),
.Y(n_613)
);

BUFx10_ASAP7_75t_L g614 ( 
.A(n_89),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_19),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_220),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_54),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_305),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_109),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_16),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_210),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_421),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_192),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_376),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_454),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_447),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_202),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_128),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_264),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_430),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_354),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_313),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_359),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_182),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_102),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_62),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_148),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_458),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_452),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_246),
.Y(n_640)
);

INVx1_ASAP7_75t_SL g641 ( 
.A(n_34),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_431),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_105),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_162),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_79),
.Y(n_645)
);

BUFx10_ASAP7_75t_L g646 ( 
.A(n_199),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_276),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_395),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_325),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_415),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_335),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_400),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_233),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_95),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_110),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_223),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_92),
.Y(n_657)
);

CKINVDCx14_ASAP7_75t_R g658 ( 
.A(n_242),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_405),
.Y(n_659)
);

INVx1_ASAP7_75t_SL g660 ( 
.A(n_31),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_363),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_150),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_56),
.Y(n_663)
);

INVx1_ASAP7_75t_SL g664 ( 
.A(n_55),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_171),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_10),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_339),
.Y(n_667)
);

BUFx10_ASAP7_75t_L g668 ( 
.A(n_39),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_100),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_263),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_377),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_350),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_334),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_367),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_443),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_256),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_297),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_252),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_257),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_232),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_123),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_455),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_136),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_358),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_388),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_240),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_137),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_164),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_413),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_207),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_94),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_143),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_307),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_112),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_184),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_373),
.Y(n_696)
);

INVxp67_ASAP7_75t_L g697 ( 
.A(n_379),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_432),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_382),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_560),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g701 ( 
.A(n_566),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_560),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_493),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_493),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_635),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_463),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_464),
.Y(n_707)
);

INVxp67_ASAP7_75t_SL g708 ( 
.A(n_471),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_469),
.Y(n_709)
);

INVxp33_ASAP7_75t_SL g710 ( 
.A(n_492),
.Y(n_710)
);

CKINVDCx20_ASAP7_75t_R g711 ( 
.A(n_481),
.Y(n_711)
);

BUFx10_ASAP7_75t_L g712 ( 
.A(n_470),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_635),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_535),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_519),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_535),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_579),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_535),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_535),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_680),
.Y(n_720)
);

INVxp67_ASAP7_75t_SL g721 ( 
.A(n_478),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_680),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_466),
.Y(n_723)
);

BUFx10_ASAP7_75t_L g724 ( 
.A(n_473),
.Y(n_724)
);

CKINVDCx20_ASAP7_75t_R g725 ( 
.A(n_486),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_477),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_538),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_658),
.B(n_0),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_496),
.Y(n_729)
);

CKINVDCx14_ASAP7_75t_R g730 ( 
.A(n_472),
.Y(n_730)
);

INVxp67_ASAP7_75t_SL g731 ( 
.A(n_649),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_516),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_533),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_474),
.Y(n_734)
);

INVxp67_ASAP7_75t_SL g735 ( 
.A(n_671),
.Y(n_735)
);

INVxp67_ASAP7_75t_SL g736 ( 
.A(n_498),
.Y(n_736)
);

CKINVDCx14_ASAP7_75t_R g737 ( 
.A(n_472),
.Y(n_737)
);

INVxp67_ASAP7_75t_SL g738 ( 
.A(n_498),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_476),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_490),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_534),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_539),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_543),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_549),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_562),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_482),
.Y(n_746)
);

INVxp67_ASAP7_75t_SL g747 ( 
.A(n_499),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_512),
.Y(n_748)
);

INVxp67_ASAP7_75t_SL g749 ( 
.A(n_499),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_567),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_569),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_573),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_578),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_583),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_597),
.Y(n_755)
);

INVxp67_ASAP7_75t_SL g756 ( 
.A(n_510),
.Y(n_756)
);

INVxp67_ASAP7_75t_L g757 ( 
.A(n_620),
.Y(n_757)
);

INVxp67_ASAP7_75t_SL g758 ( 
.A(n_510),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_600),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_601),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_605),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_504),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_629),
.Y(n_763)
);

INVxp67_ASAP7_75t_L g764 ( 
.A(n_623),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_520),
.Y(n_765)
);

INVxp33_ASAP7_75t_L g766 ( 
.A(n_637),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_609),
.Y(n_767)
);

CKINVDCx16_ASAP7_75t_R g768 ( 
.A(n_589),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_612),
.Y(n_769)
);

NOR2xp67_ASAP7_75t_L g770 ( 
.A(n_528),
.B(n_0),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_519),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_488),
.Y(n_772)
);

CKINVDCx16_ASAP7_75t_R g773 ( 
.A(n_556),
.Y(n_773)
);

INVxp33_ASAP7_75t_SL g774 ( 
.A(n_475),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_628),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_629),
.Y(n_776)
);

INVxp67_ASAP7_75t_SL g777 ( 
.A(n_639),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_644),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_654),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_663),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_491),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_SL g782 ( 
.A1(n_710),
.A2(n_658),
.B1(n_526),
.B2(n_590),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_716),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_706),
.B(n_707),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_715),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_715),
.Y(n_786)
);

INVxp67_ASAP7_75t_L g787 ( 
.A(n_717),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_709),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_714),
.Y(n_789)
);

INVx6_ASAP7_75t_L g790 ( 
.A(n_715),
.Y(n_790)
);

INVx6_ASAP7_75t_L g791 ( 
.A(n_715),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_703),
.Y(n_792)
);

AND2x4_ASAP7_75t_L g793 ( 
.A(n_736),
.B(n_639),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_738),
.B(n_480),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_734),
.B(n_632),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_720),
.Y(n_796)
);

OA21x2_ASAP7_75t_L g797 ( 
.A1(n_720),
.A2(n_595),
.B(n_542),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_718),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_703),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_719),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_774),
.B(n_561),
.Y(n_801)
);

AND2x6_ASAP7_75t_L g802 ( 
.A(n_771),
.B(n_519),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_771),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_739),
.B(n_468),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_771),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_722),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_723),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_746),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_728),
.B(n_494),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_726),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_729),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_732),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_733),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_768),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_772),
.B(n_647),
.Y(n_815)
);

BUFx8_ASAP7_75t_L g816 ( 
.A(n_704),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_704),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_741),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_742),
.Y(n_819)
);

BUFx2_ASAP7_75t_L g820 ( 
.A(n_763),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_781),
.B(n_685),
.Y(n_821)
);

INVx4_ASAP7_75t_L g822 ( 
.A(n_763),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_743),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_747),
.B(n_542),
.Y(n_824)
);

INVx4_ASAP7_75t_L g825 ( 
.A(n_776),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_749),
.B(n_595),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_776),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_756),
.B(n_480),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_758),
.B(n_652),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_700),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_744),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_SL g832 ( 
.A1(n_711),
.A2(n_592),
.B1(n_604),
.B2(n_571),
.Y(n_832)
);

HB1xp67_ASAP7_75t_L g833 ( 
.A(n_727),
.Y(n_833)
);

AND2x6_ASAP7_75t_L g834 ( 
.A(n_728),
.B(n_519),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_745),
.Y(n_835)
);

OAI22xp33_ASAP7_75t_L g836 ( 
.A1(n_766),
.A2(n_764),
.B1(n_757),
.B2(n_721),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_702),
.Y(n_837)
);

CKINVDCx20_ASAP7_75t_R g838 ( 
.A(n_788),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_R g839 ( 
.A(n_788),
.B(n_762),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_808),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_808),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_820),
.B(n_792),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_804),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_784),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_823),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_830),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_816),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_803),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_814),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_827),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_837),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_837),
.Y(n_852)
);

AND2x6_ASAP7_75t_L g853 ( 
.A(n_826),
.B(n_652),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_785),
.Y(n_854)
);

CKINVDCx20_ASAP7_75t_R g855 ( 
.A(n_816),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_816),
.Y(n_856)
);

NAND2xp33_ASAP7_75t_R g857 ( 
.A(n_793),
.B(n_479),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_803),
.Y(n_858)
);

NAND2xp33_ASAP7_75t_R g859 ( 
.A(n_793),
.B(n_794),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_801),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_799),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_832),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_799),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_795),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_815),
.Y(n_865)
);

CKINVDCx16_ASAP7_75t_R g866 ( 
.A(n_833),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_807),
.Y(n_867)
);

BUFx10_ASAP7_75t_L g868 ( 
.A(n_793),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_785),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_821),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_792),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_807),
.Y(n_872)
);

CKINVDCx20_ASAP7_75t_R g873 ( 
.A(n_787),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_817),
.Y(n_874)
);

NOR2xp67_ASAP7_75t_L g875 ( 
.A(n_822),
.B(n_697),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_817),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_834),
.B(n_730),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_822),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_794),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_825),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_807),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_785),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_807),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_825),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_828),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_809),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_R g887 ( 
.A(n_834),
.B(n_730),
.Y(n_887)
);

CKINVDCx20_ASAP7_75t_R g888 ( 
.A(n_809),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_826),
.B(n_773),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_810),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_782),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_836),
.B(n_737),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_826),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_824),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_810),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_829),
.B(n_731),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_834),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_834),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_834),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_810),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_834),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_810),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_818),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_818),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_818),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_818),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_813),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_785),
.Y(n_908)
);

CKINVDCx20_ASAP7_75t_R g909 ( 
.A(n_811),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_813),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_866),
.B(n_735),
.Y(n_911)
);

INVx4_ASAP7_75t_L g912 ( 
.A(n_902),
.Y(n_912)
);

OR2x2_ASAP7_75t_L g913 ( 
.A(n_879),
.B(n_708),
.Y(n_913)
);

INVxp33_ASAP7_75t_L g914 ( 
.A(n_839),
.Y(n_914)
);

NAND2xp33_ASAP7_75t_L g915 ( 
.A(n_897),
.B(n_802),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_868),
.Y(n_916)
);

INVx4_ASAP7_75t_L g917 ( 
.A(n_903),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_868),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_894),
.B(n_712),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_848),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_893),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_858),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_845),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_889),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_896),
.B(n_797),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_854),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_910),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_846),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_842),
.B(n_766),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_909),
.Y(n_930)
);

AND3x1_ASAP7_75t_L g931 ( 
.A(n_892),
.B(n_879),
.C(n_850),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_861),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_863),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_854),
.Y(n_934)
);

CKINVDCx20_ASAP7_75t_R g935 ( 
.A(n_838),
.Y(n_935)
);

INVx5_ASAP7_75t_L g936 ( 
.A(n_853),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_854),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_885),
.B(n_777),
.Y(n_938)
);

BUFx3_ASAP7_75t_L g939 ( 
.A(n_851),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_843),
.B(n_724),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_852),
.B(n_904),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_854),
.Y(n_942)
);

INVxp33_ASAP7_75t_L g943 ( 
.A(n_875),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_867),
.B(n_872),
.Y(n_944)
);

INVxp67_ASAP7_75t_L g945 ( 
.A(n_857),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_869),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_853),
.B(n_831),
.Y(n_947)
);

BUFx10_ASAP7_75t_L g948 ( 
.A(n_840),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_841),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_907),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_871),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_881),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_883),
.B(n_812),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_859),
.A2(n_544),
.B1(n_613),
.B2(n_585),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_864),
.B(n_865),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_890),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_869),
.Y(n_957)
);

AND2x2_ASAP7_75t_SL g958 ( 
.A(n_862),
.B(n_523),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_844),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_882),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_870),
.B(n_624),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_895),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_900),
.B(n_812),
.Y(n_963)
);

OAI22xp33_ASAP7_75t_L g964 ( 
.A1(n_860),
.A2(n_770),
.B1(n_661),
.B2(n_525),
.Y(n_964)
);

INVxp67_ASAP7_75t_L g965 ( 
.A(n_874),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_882),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_876),
.B(n_737),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_905),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_906),
.B(n_501),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_878),
.B(n_711),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_849),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_882),
.Y(n_972)
);

OR2x6_ASAP7_75t_L g973 ( 
.A(n_855),
.B(n_550),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_908),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_908),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_891),
.B(n_705),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_853),
.B(n_831),
.Y(n_977)
);

AOI22xp5_ASAP7_75t_L g978 ( 
.A1(n_886),
.A2(n_669),
.B1(n_695),
.B2(n_643),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_898),
.B(n_831),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_899),
.B(n_783),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_873),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_880),
.B(n_725),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_901),
.B(n_783),
.Y(n_983)
);

INVx4_ASAP7_75t_SL g984 ( 
.A(n_908),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_908),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_888),
.A2(n_593),
.B1(n_659),
.B2(n_467),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_884),
.Y(n_987)
);

INVx8_ASAP7_75t_L g988 ( 
.A(n_847),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_856),
.Y(n_989)
);

INVx1_ASAP7_75t_SL g990 ( 
.A(n_887),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_877),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_843),
.B(n_725),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_909),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_893),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_893),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_868),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_893),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_893),
.Y(n_998)
);

OR2x2_ASAP7_75t_L g999 ( 
.A(n_866),
.B(n_713),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_894),
.B(n_805),
.Y(n_1000)
);

BUFx10_ASAP7_75t_L g1001 ( 
.A(n_892),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_842),
.B(n_819),
.Y(n_1002)
);

BUFx2_ASAP7_75t_L g1003 ( 
.A(n_849),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_848),
.Y(n_1004)
);

INVx6_ASAP7_75t_L g1005 ( 
.A(n_866),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_848),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_893),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_L g1008 ( 
.A1(n_853),
.A2(n_517),
.B1(n_518),
.B2(n_508),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_893),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_893),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_894),
.B(n_497),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_893),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_894),
.B(n_796),
.Y(n_1013)
);

AND2x4_ASAP7_75t_L g1014 ( 
.A(n_846),
.B(n_835),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_842),
.B(n_835),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_893),
.Y(n_1016)
);

BUFx10_ASAP7_75t_L g1017 ( 
.A(n_892),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_843),
.B(n_740),
.Y(n_1018)
);

BUFx10_ASAP7_75t_L g1019 ( 
.A(n_892),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_893),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_1002),
.B(n_540),
.Y(n_1021)
);

NOR2x1p5_ASAP7_75t_L g1022 ( 
.A(n_916),
.B(n_701),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_1015),
.B(n_554),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_931),
.A2(n_576),
.B1(n_580),
.B2(n_574),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_986),
.A2(n_607),
.B(n_622),
.C(n_603),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_925),
.A2(n_633),
.B(n_642),
.C(n_630),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_944),
.Y(n_1027)
);

AND2x6_ASAP7_75t_SL g1028 ( 
.A(n_992),
.B(n_686),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_923),
.Y(n_1029)
);

OR2x6_ASAP7_75t_L g1030 ( 
.A(n_1005),
.B(n_988),
.Y(n_1030)
);

AOI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_991),
.A2(n_675),
.B1(n_676),
.B2(n_667),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_945),
.B(n_503),
.Y(n_1032)
);

AND2x6_ASAP7_75t_L g1033 ( 
.A(n_979),
.B(n_677),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_955),
.B(n_740),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_959),
.B(n_748),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_929),
.B(n_748),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_953),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_912),
.B(n_505),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_961),
.B(n_765),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_1014),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1013),
.B(n_806),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1013),
.B(n_806),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_938),
.B(n_789),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_1000),
.B(n_798),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_963),
.Y(n_1045)
);

AND2x2_ASAP7_75t_SL g1046 ( 
.A(n_958),
.B(n_765),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_979),
.B(n_800),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_917),
.B(n_507),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_927),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_965),
.B(n_701),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_917),
.B(n_509),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_931),
.A2(n_513),
.B1(n_514),
.B2(n_511),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_913),
.B(n_465),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_951),
.B(n_515),
.Y(n_1054)
);

BUFx8_ASAP7_75t_L g1055 ( 
.A(n_1003),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_916),
.B(n_521),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_921),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_940),
.B(n_465),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_SL g1059 ( 
.A(n_949),
.B(n_494),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_980),
.B(n_522),
.Y(n_1060)
);

INVx1_ASAP7_75t_SL g1061 ( 
.A(n_1005),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_916),
.B(n_529),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_SL g1063 ( 
.A(n_948),
.B(n_494),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_983),
.B(n_530),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_994),
.Y(n_1065)
);

OR2x6_ASAP7_75t_L g1066 ( 
.A(n_988),
.B(n_523),
.Y(n_1066)
);

NOR2x1p5_ASAP7_75t_L g1067 ( 
.A(n_918),
.B(n_483),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_983),
.B(n_531),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_954),
.B(n_928),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_976),
.B(n_465),
.Y(n_1070)
);

INVx4_ASAP7_75t_L g1071 ( 
.A(n_918),
.Y(n_1071)
);

INVx2_ASAP7_75t_SL g1072 ( 
.A(n_999),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_995),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_935),
.Y(n_1074)
);

INVxp67_ASAP7_75t_L g1075 ( 
.A(n_911),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_918),
.Y(n_1076)
);

OAI22xp33_ASAP7_75t_L g1077 ( 
.A1(n_943),
.A2(n_641),
.B1(n_660),
.B2(n_545),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_950),
.B(n_547),
.Y(n_1078)
);

INVx2_ASAP7_75t_SL g1079 ( 
.A(n_930),
.Y(n_1079)
);

OR2x6_ASAP7_75t_L g1080 ( 
.A(n_988),
.B(n_588),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_941),
.B(n_968),
.Y(n_1081)
);

AOI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_997),
.A2(n_553),
.B1(n_555),
.B2(n_552),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_998),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_SL g1084 ( 
.A1(n_978),
.A2(n_664),
.B1(n_485),
.B2(n_487),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_1007),
.A2(n_570),
.B1(n_673),
.B2(n_602),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_964),
.B(n_484),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1009),
.B(n_559),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_914),
.B(n_489),
.Y(n_1088)
);

INVxp67_ASAP7_75t_L g1089 ( 
.A(n_924),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1010),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_1012),
.A2(n_570),
.B1(n_673),
.B2(n_602),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_1004),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1016),
.B(n_563),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1020),
.B(n_564),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_SL g1095 ( 
.A(n_948),
.B(n_506),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_987),
.B(n_565),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_952),
.B(n_568),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1006),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_993),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_920),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_920),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_922),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_919),
.B(n_495),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_956),
.B(n_572),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_970),
.B(n_500),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_947),
.A2(n_570),
.B1(n_673),
.B2(n_602),
.Y(n_1106)
);

NOR2xp67_ASAP7_75t_L g1107 ( 
.A(n_996),
.B(n_750),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_982),
.B(n_1018),
.Y(n_1108)
);

INVxp67_ASAP7_75t_L g1109 ( 
.A(n_981),
.Y(n_1109)
);

AOI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_947),
.A2(n_582),
.B1(n_591),
.B2(n_584),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_962),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_977),
.A2(n_570),
.B1(n_674),
.B2(n_581),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_939),
.Y(n_1113)
);

INVx2_ASAP7_75t_SL g1114 ( 
.A(n_971),
.Y(n_1114)
);

INVx4_ASAP7_75t_L g1115 ( 
.A(n_984),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_926),
.Y(n_1116)
);

HB1xp67_ASAP7_75t_L g1117 ( 
.A(n_932),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_1011),
.B(n_502),
.Y(n_1118)
);

NAND2x1p5_ASAP7_75t_L g1119 ( 
.A(n_936),
.B(n_674),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_969),
.B(n_611),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_934),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_936),
.B(n_967),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_942),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_946),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_933),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_977),
.A2(n_674),
.B1(n_581),
.B2(n_506),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_1001),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_960),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1008),
.B(n_618),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_990),
.B(n_625),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_1001),
.A2(n_674),
.B1(n_581),
.B2(n_506),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1017),
.A2(n_631),
.B1(n_638),
.B2(n_626),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1019),
.A2(n_617),
.B1(n_662),
.B2(n_599),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_990),
.B(n_966),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_972),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1019),
.A2(n_972),
.B1(n_985),
.B2(n_975),
.Y(n_1136)
);

INVxp67_ASAP7_75t_L g1137 ( 
.A(n_978),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_985),
.Y(n_1138)
);

AOI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_915),
.A2(n_650),
.B1(n_651),
.B2(n_648),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_937),
.B(n_957),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_937),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_984),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_989),
.B(n_524),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_937),
.Y(n_1144)
);

INVx2_ASAP7_75t_SL g1145 ( 
.A(n_973),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_973),
.B(n_532),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_974),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_SL g1148 ( 
.A(n_973),
.B(n_527),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1002),
.B(n_670),
.Y(n_1149)
);

HB1xp67_ASAP7_75t_L g1150 ( 
.A(n_924),
.Y(n_1150)
);

NOR3xp33_ASAP7_75t_L g1151 ( 
.A(n_961),
.B(n_767),
.C(n_761),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1002),
.B(n_672),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_944),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_945),
.B(n_536),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1002),
.B(n_678),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_945),
.B(n_537),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1002),
.B(n_679),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_945),
.B(n_541),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_1005),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1002),
.B(n_682),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1029),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_1046),
.B(n_684),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1140),
.A2(n_786),
.B(n_689),
.Y(n_1163)
);

INVx4_ASAP7_75t_L g1164 ( 
.A(n_1071),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_1141),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1044),
.B(n_693),
.Y(n_1166)
);

NOR2x1_ASAP7_75t_L g1167 ( 
.A(n_1071),
.B(n_751),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_1086),
.A2(n_698),
.B1(n_699),
.B2(n_696),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1049),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1021),
.B(n_1023),
.Y(n_1170)
);

AO21x1_ASAP7_75t_L g1171 ( 
.A1(n_1024),
.A2(n_690),
.B(n_688),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1041),
.A2(n_1042),
.B(n_1043),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1108),
.B(n_546),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1118),
.A2(n_692),
.B(n_617),
.C(n_662),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1075),
.B(n_548),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1069),
.A2(n_557),
.B1(n_558),
.B2(n_551),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1060),
.B(n_575),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1105),
.B(n_577),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1047),
.A2(n_802),
.B(n_753),
.Y(n_1179)
);

BUFx8_ASAP7_75t_SL g1180 ( 
.A(n_1030),
.Y(n_1180)
);

AOI33xp33_ASAP7_75t_L g1181 ( 
.A1(n_1077),
.A2(n_755),
.A3(n_752),
.B1(n_760),
.B2(n_759),
.B3(n_754),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1064),
.B(n_586),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1068),
.B(n_594),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_1027),
.B(n_1153),
.Y(n_1184)
);

INVx4_ASAP7_75t_L g1185 ( 
.A(n_1076),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1149),
.B(n_596),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_1137),
.B(n_1089),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_1125),
.Y(n_1188)
);

BUFx4f_ASAP7_75t_L g1189 ( 
.A(n_1030),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1154),
.A2(n_599),
.B(n_775),
.C(n_769),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1156),
.B(n_598),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1152),
.B(n_606),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1155),
.A2(n_779),
.B(n_778),
.Y(n_1193)
);

OAI321xp33_ASAP7_75t_L g1194 ( 
.A1(n_1084),
.A2(n_780),
.A3(n_646),
.B1(n_587),
.B2(n_668),
.C(n_614),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_1030),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1037),
.Y(n_1196)
);

INVx4_ASAP7_75t_L g1197 ( 
.A(n_1076),
.Y(n_1197)
);

O2A1O1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1158),
.A2(n_587),
.B(n_614),
.C(n_527),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1027),
.B(n_608),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1157),
.A2(n_791),
.B(n_790),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1160),
.B(n_610),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1113),
.B(n_250),
.Y(n_1202)
);

INVxp67_ASAP7_75t_L g1203 ( 
.A(n_1150),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1153),
.B(n_615),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1053),
.B(n_527),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1026),
.A2(n_619),
.B(n_616),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1070),
.B(n_587),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1092),
.Y(n_1208)
);

OAI21xp33_ASAP7_75t_L g1209 ( 
.A1(n_1059),
.A2(n_627),
.B(n_621),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1098),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1134),
.B(n_634),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1103),
.A2(n_636),
.B(n_645),
.C(n_640),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_1141),
.Y(n_1213)
);

NOR3xp33_ASAP7_75t_L g1214 ( 
.A(n_1035),
.B(n_655),
.C(n_653),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1036),
.B(n_1072),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1058),
.B(n_1039),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_1117),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_1141),
.Y(n_1218)
);

AO21x1_ASAP7_75t_L g1219 ( 
.A1(n_1024),
.A2(n_1),
.B(n_2),
.Y(n_1219)
);

O2A1O1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1025),
.A2(n_668),
.B(n_646),
.C(n_657),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1111),
.B(n_656),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1033),
.B(n_665),
.Y(n_1222)
);

INVx11_ASAP7_75t_L g1223 ( 
.A(n_1055),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1033),
.B(n_666),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1033),
.B(n_681),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_1081),
.B(n_683),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1040),
.B(n_687),
.Y(n_1227)
);

OAI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1110),
.A2(n_694),
.B(n_691),
.Y(n_1228)
);

AOI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1034),
.A2(n_668),
.B1(n_646),
.B2(n_259),
.Y(n_1229)
);

AOI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1107),
.A2(n_260),
.B1(n_261),
.B2(n_258),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1045),
.B(n_1),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1088),
.B(n_2),
.Y(n_1232)
);

INVx5_ASAP7_75t_L g1233 ( 
.A(n_1115),
.Y(n_1233)
);

NOR3xp33_ASAP7_75t_L g1234 ( 
.A(n_1084),
.B(n_3),
.C(n_4),
.Y(n_1234)
);

NAND3xp33_ASAP7_75t_L g1235 ( 
.A(n_1131),
.B(n_3),
.C(n_5),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1099),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1057),
.B(n_7),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1110),
.A2(n_268),
.B(n_267),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1109),
.B(n_7),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1119),
.A2(n_271),
.B(n_269),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1130),
.B(n_8),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1050),
.B(n_1096),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1065),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1073),
.B(n_8),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1116),
.A2(n_273),
.B(n_272),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1055),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1136),
.A2(n_275),
.B1(n_277),
.B2(n_274),
.Y(n_1247)
);

NAND2x1p5_ASAP7_75t_L g1248 ( 
.A(n_1115),
.B(n_278),
.Y(n_1248)
);

NAND2x1p5_ASAP7_75t_L g1249 ( 
.A(n_1159),
.B(n_279),
.Y(n_1249)
);

AOI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1121),
.A2(n_283),
.B(n_282),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1116),
.A2(n_285),
.B(n_284),
.Y(n_1251)
);

NOR3xp33_ASAP7_75t_L g1252 ( 
.A(n_1143),
.B(n_9),
.C(n_10),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_1052),
.B(n_286),
.Y(n_1253)
);

AND2x4_ASAP7_75t_L g1254 ( 
.A(n_1083),
.B(n_287),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1031),
.A2(n_289),
.B1(n_290),
.B2(n_288),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1142),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1090),
.Y(n_1257)
);

BUFx4f_ASAP7_75t_L g1258 ( 
.A(n_1127),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1147),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1100),
.B(n_9),
.Y(n_1260)
);

INVx1_ASAP7_75t_SL g1261 ( 
.A(n_1061),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1124),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1135),
.A2(n_292),
.B(n_291),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1101),
.B(n_11),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1135),
.A2(n_296),
.B(n_294),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1102),
.B(n_11),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1133),
.B(n_12),
.Y(n_1267)
);

HB1xp67_ASAP7_75t_L g1268 ( 
.A(n_1079),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_SL g1269 ( 
.A(n_1074),
.B(n_298),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_1114),
.B(n_12),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1122),
.A2(n_300),
.B(n_299),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1097),
.B(n_14),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1129),
.A2(n_1104),
.B(n_1144),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1078),
.A2(n_304),
.B(n_303),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1056),
.A2(n_309),
.B(n_308),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_R g1276 ( 
.A(n_1148),
.B(n_310),
.Y(n_1276)
);

INVx1_ASAP7_75t_SL g1277 ( 
.A(n_1066),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1123),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1062),
.A2(n_316),
.B(n_312),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_1138),
.Y(n_1280)
);

INVx8_ASAP7_75t_L g1281 ( 
.A(n_1066),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1120),
.B(n_15),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_1082),
.B(n_317),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1032),
.B(n_17),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_1128),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1087),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1093),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1066),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1132),
.B(n_18),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1082),
.B(n_19),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1094),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1106),
.A2(n_319),
.B(n_318),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1112),
.A2(n_321),
.B1(n_322),
.B2(n_320),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1151),
.B(n_20),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1139),
.Y(n_1295)
);

NOR3xp33_ASAP7_75t_L g1296 ( 
.A(n_1146),
.B(n_20),
.C(n_21),
.Y(n_1296)
);

A2O1A1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1126),
.A2(n_23),
.B(n_21),
.C(n_22),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1038),
.B(n_24),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1054),
.B(n_25),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1048),
.A2(n_324),
.B(n_323),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1051),
.B(n_26),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1216),
.B(n_1080),
.Y(n_1302)
);

O2A1O1Ixp5_ASAP7_75t_L g1303 ( 
.A1(n_1178),
.A2(n_1095),
.B(n_1063),
.C(n_1139),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1242),
.B(n_1028),
.Y(n_1304)
);

AO21x1_ASAP7_75t_L g1305 ( 
.A1(n_1238),
.A2(n_1091),
.B(n_1085),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1170),
.A2(n_1145),
.B1(n_1080),
.B2(n_1067),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_R g1307 ( 
.A(n_1188),
.B(n_1028),
.Y(n_1307)
);

NAND2x1p5_ASAP7_75t_L g1308 ( 
.A(n_1233),
.B(n_1022),
.Y(n_1308)
);

OR2x6_ASAP7_75t_L g1309 ( 
.A(n_1281),
.B(n_326),
.Y(n_1309)
);

INVx3_ASAP7_75t_L g1310 ( 
.A(n_1180),
.Y(n_1310)
);

A2O1A1Ixp33_ASAP7_75t_SL g1311 ( 
.A1(n_1232),
.A2(n_1191),
.B(n_1241),
.C(n_1299),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1286),
.B(n_27),
.Y(n_1312)
);

BUFx10_ASAP7_75t_L g1313 ( 
.A(n_1215),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1243),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1236),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1172),
.A2(n_329),
.B(n_327),
.Y(n_1316)
);

BUFx6f_ASAP7_75t_L g1317 ( 
.A(n_1218),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1273),
.A2(n_332),
.B(n_331),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1217),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_SL g1320 ( 
.A(n_1189),
.B(n_1269),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1195),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1257),
.Y(n_1322)
);

O2A1O1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1198),
.A2(n_29),
.B(n_27),
.C(n_28),
.Y(n_1323)
);

INVx2_ASAP7_75t_SL g1324 ( 
.A(n_1268),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1289),
.A2(n_32),
.B1(n_28),
.B2(n_29),
.Y(n_1325)
);

O2A1O1Ixp33_ASAP7_75t_L g1326 ( 
.A1(n_1234),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1205),
.B(n_35),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1223),
.Y(n_1328)
);

A2O1A1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1287),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_1329)
);

INVxp67_ASAP7_75t_L g1330 ( 
.A(n_1187),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1173),
.B(n_41),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1161),
.Y(n_1332)
);

A2O1A1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1291),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_1333)
);

AND2x6_ASAP7_75t_L g1334 ( 
.A(n_1295),
.B(n_333),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_1203),
.Y(n_1335)
);

CKINVDCx20_ASAP7_75t_R g1336 ( 
.A(n_1246),
.Y(n_1336)
);

BUFx4f_ASAP7_75t_L g1337 ( 
.A(n_1288),
.Y(n_1337)
);

BUFx12f_ASAP7_75t_L g1338 ( 
.A(n_1288),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1166),
.B(n_1211),
.Y(n_1339)
);

AND2x4_ASAP7_75t_SL g1340 ( 
.A(n_1164),
.B(n_338),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1169),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1262),
.Y(n_1342)
);

BUFx12f_ASAP7_75t_L g1343 ( 
.A(n_1288),
.Y(n_1343)
);

NOR2xp67_ASAP7_75t_SL g1344 ( 
.A(n_1233),
.B(n_1194),
.Y(n_1344)
);

INVx1_ASAP7_75t_SL g1345 ( 
.A(n_1261),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1259),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1177),
.B(n_45),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1182),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_1348)
);

AOI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1214),
.A2(n_1162),
.B1(n_1283),
.B2(n_1253),
.Y(n_1349)
);

OA22x2_ASAP7_75t_L g1350 ( 
.A1(n_1229),
.A2(n_1290),
.B1(n_1294),
.B2(n_1228),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_1218),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1272),
.A2(n_343),
.B(n_342),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1207),
.B(n_49),
.Y(n_1353)
);

O2A1O1Ixp33_ASAP7_75t_SL g1354 ( 
.A1(n_1297),
.A2(n_349),
.B(n_353),
.C(n_345),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1183),
.B(n_50),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_SL g1356 ( 
.A(n_1254),
.B(n_50),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1237),
.B(n_51),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1186),
.B(n_51),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_SL g1359 ( 
.A(n_1254),
.B(n_52),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1192),
.B(n_53),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1235),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_1361)
);

O2A1O1Ixp5_ASAP7_75t_L g1362 ( 
.A1(n_1282),
.A2(n_60),
.B(n_58),
.C(n_59),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_1258),
.B(n_61),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_SL g1364 ( 
.A1(n_1277),
.A2(n_64),
.B1(n_61),
.B2(n_63),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1292),
.A2(n_362),
.B(n_361),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1201),
.B(n_65),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1196),
.B(n_66),
.Y(n_1367)
);

AOI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1175),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_1368)
);

AOI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1226),
.A2(n_1199),
.B1(n_1301),
.B2(n_1298),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1221),
.B(n_70),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1296),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_1371)
);

INVx4_ASAP7_75t_L g1372 ( 
.A(n_1164),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1209),
.B(n_72),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1208),
.B(n_73),
.Y(n_1374)
);

NAND2x1p5_ASAP7_75t_L g1375 ( 
.A(n_1185),
.B(n_365),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1210),
.B(n_74),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1193),
.B(n_74),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1259),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1204),
.B(n_1212),
.Y(n_1379)
);

O2A1O1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1252),
.A2(n_78),
.B(n_75),
.C(n_76),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1244),
.B(n_78),
.Y(n_1381)
);

NAND2x1p5_ASAP7_75t_L g1382 ( 
.A(n_1185),
.B(n_369),
.Y(n_1382)
);

A2O1A1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1220),
.A2(n_83),
.B(n_81),
.C(n_82),
.Y(n_1383)
);

INVx5_ASAP7_75t_L g1384 ( 
.A(n_1197),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1278),
.Y(n_1385)
);

INVx4_ASAP7_75t_L g1386 ( 
.A(n_1197),
.Y(n_1386)
);

AO21x2_ASAP7_75t_L g1387 ( 
.A1(n_1200),
.A2(n_371),
.B(n_370),
.Y(n_1387)
);

OAI21xp33_ASAP7_75t_L g1388 ( 
.A1(n_1181),
.A2(n_85),
.B(n_86),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1256),
.Y(n_1389)
);

NAND3xp33_ASAP7_75t_L g1390 ( 
.A(n_1168),
.B(n_1174),
.C(n_1206),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_L g1391 ( 
.A(n_1284),
.B(n_86),
.Y(n_1391)
);

AOI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1202),
.A2(n_90),
.B1(n_87),
.B2(n_88),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_1276),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1260),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1227),
.B(n_87),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1256),
.B(n_372),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1231),
.B(n_88),
.Y(n_1397)
);

AND2x6_ASAP7_75t_L g1398 ( 
.A(n_1165),
.B(n_374),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1264),
.Y(n_1399)
);

BUFx12f_ASAP7_75t_L g1400 ( 
.A(n_1270),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_1256),
.Y(n_1401)
);

AOI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1163),
.A2(n_462),
.B(n_375),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1266),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_L g1404 ( 
.A(n_1176),
.B(n_90),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1281),
.Y(n_1405)
);

NOR2xp67_ASAP7_75t_R g1406 ( 
.A(n_1259),
.B(n_91),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_R g1407 ( 
.A(n_1165),
.B(n_378),
.Y(n_1407)
);

INVx4_ASAP7_75t_L g1408 ( 
.A(n_1213),
.Y(n_1408)
);

INVx2_ASAP7_75t_SL g1409 ( 
.A(n_1285),
.Y(n_1409)
);

NOR3xp33_ASAP7_75t_SL g1410 ( 
.A(n_1239),
.B(n_92),
.C(n_93),
.Y(n_1410)
);

OR2x6_ASAP7_75t_SL g1411 ( 
.A(n_1222),
.B(n_96),
.Y(n_1411)
);

BUFx6f_ASAP7_75t_L g1412 ( 
.A(n_1280),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1285),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1224),
.B(n_96),
.Y(n_1414)
);

O2A1O1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1190),
.A2(n_99),
.B(n_97),
.C(n_98),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1250),
.A2(n_381),
.B(n_380),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_SL g1417 ( 
.A(n_1280),
.B(n_97),
.Y(n_1417)
);

O2A1O1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1225),
.A2(n_102),
.B(n_99),
.C(n_101),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1167),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1341),
.Y(n_1420)
);

NAND3x1_ASAP7_75t_L g1421 ( 
.A(n_1304),
.B(n_1230),
.C(n_1267),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1311),
.A2(n_1300),
.B(n_1179),
.Y(n_1422)
);

OAI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1390),
.A2(n_1184),
.B(n_1275),
.Y(n_1423)
);

INVxp67_ASAP7_75t_L g1424 ( 
.A(n_1319),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1339),
.B(n_1171),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1330),
.B(n_1219),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1350),
.A2(n_1247),
.B1(n_1293),
.B2(n_1255),
.Y(n_1427)
);

NAND3xp33_ASAP7_75t_L g1428 ( 
.A(n_1404),
.B(n_1355),
.C(n_1347),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1345),
.B(n_1249),
.Y(n_1429)
);

INVxp67_ASAP7_75t_SL g1430 ( 
.A(n_1335),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1365),
.A2(n_1251),
.B(n_1245),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1379),
.A2(n_1265),
.B(n_1263),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1369),
.A2(n_1248),
.B1(n_1271),
.B2(n_1279),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_1320),
.B(n_1274),
.Y(n_1434)
);

AOI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1402),
.A2(n_1240),
.B(n_383),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1314),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1331),
.B(n_103),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1322),
.Y(n_1438)
);

AOI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1318),
.A2(n_461),
.B(n_385),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1416),
.A2(n_390),
.B(n_389),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1394),
.B(n_103),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1399),
.B(n_104),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1403),
.B(n_104),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_R g1444 ( 
.A(n_1413),
.B(n_391),
.Y(n_1444)
);

AO31x2_ASAP7_75t_L g1445 ( 
.A1(n_1305),
.A2(n_108),
.A3(n_106),
.B(n_107),
.Y(n_1445)
);

OA21x2_ASAP7_75t_L g1446 ( 
.A1(n_1316),
.A2(n_394),
.B(n_393),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1393),
.B(n_1356),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1352),
.A2(n_459),
.B(n_397),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1303),
.A2(n_107),
.B(n_108),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1359),
.B(n_399),
.Y(n_1450)
);

NOR4xp25_ASAP7_75t_L g1451 ( 
.A(n_1326),
.B(n_113),
.C(n_111),
.D(n_112),
.Y(n_1451)
);

AO31x2_ASAP7_75t_L g1452 ( 
.A1(n_1383),
.A2(n_116),
.A3(n_114),
.B(n_115),
.Y(n_1452)
);

AOI211x1_ASAP7_75t_L g1453 ( 
.A1(n_1348),
.A2(n_117),
.B(n_115),
.C(n_116),
.Y(n_1453)
);

INVx3_ASAP7_75t_L g1454 ( 
.A(n_1412),
.Y(n_1454)
);

INVx1_ASAP7_75t_SL g1455 ( 
.A(n_1315),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_1324),
.Y(n_1456)
);

BUFx12f_ASAP7_75t_L g1457 ( 
.A(n_1328),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1358),
.B(n_117),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1366),
.B(n_118),
.Y(n_1459)
);

OAI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1349),
.A2(n_1360),
.B(n_1373),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1302),
.B(n_119),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1397),
.B(n_120),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1357),
.B(n_121),
.Y(n_1463)
);

A2O1A1Ixp33_ASAP7_75t_L g1464 ( 
.A1(n_1391),
.A2(n_122),
.B(n_124),
.C(n_125),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1370),
.B(n_122),
.Y(n_1465)
);

NOR2xp67_ASAP7_75t_SL g1466 ( 
.A(n_1384),
.B(n_126),
.Y(n_1466)
);

OAI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1395),
.A2(n_126),
.B(n_127),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_SL g1468 ( 
.A1(n_1415),
.A2(n_127),
.B(n_128),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1312),
.B(n_129),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1332),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1313),
.B(n_406),
.Y(n_1471)
);

A2O1A1Ixp33_ASAP7_75t_L g1472 ( 
.A1(n_1414),
.A2(n_130),
.B(n_131),
.C(n_132),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1377),
.A2(n_131),
.B(n_132),
.Y(n_1473)
);

AO22x2_ASAP7_75t_L g1474 ( 
.A1(n_1306),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1342),
.Y(n_1475)
);

AOI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1354),
.A2(n_1406),
.B(n_1387),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1388),
.B(n_137),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_1412),
.Y(n_1478)
);

NOR2xp67_ASAP7_75t_L g1479 ( 
.A(n_1372),
.B(n_409),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_SL g1480 ( 
.A(n_1313),
.B(n_139),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1384),
.A2(n_412),
.B(n_410),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1385),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1374),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1317),
.Y(n_1484)
);

OAI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1362),
.A2(n_418),
.B(n_416),
.Y(n_1485)
);

O2A1O1Ixp33_ASAP7_75t_SL g1486 ( 
.A1(n_1329),
.A2(n_140),
.B(n_141),
.C(n_142),
.Y(n_1486)
);

INVx3_ASAP7_75t_L g1487 ( 
.A(n_1412),
.Y(n_1487)
);

CKINVDCx6p67_ASAP7_75t_R g1488 ( 
.A(n_1338),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1419),
.B(n_422),
.Y(n_1489)
);

AOI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1344),
.A2(n_424),
.B(n_423),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_SL g1491 ( 
.A(n_1337),
.B(n_426),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1376),
.Y(n_1492)
);

AOI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1375),
.A2(n_428),
.B(n_427),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1381),
.B(n_142),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1327),
.B(n_143),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1382),
.A2(n_435),
.B(n_434),
.Y(n_1496)
);

NAND2xp33_ASAP7_75t_L g1497 ( 
.A(n_1389),
.B(n_144),
.Y(n_1497)
);

AO31x2_ASAP7_75t_L g1498 ( 
.A1(n_1333),
.A2(n_144),
.A3(n_146),
.B(n_147),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1353),
.B(n_146),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1371),
.B(n_147),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1361),
.B(n_148),
.Y(n_1501)
);

A2O1A1Ixp33_ASAP7_75t_L g1502 ( 
.A1(n_1428),
.A2(n_1323),
.B(n_1380),
.C(n_1392),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1426),
.B(n_1367),
.Y(n_1503)
);

OA21x2_ASAP7_75t_L g1504 ( 
.A1(n_1476),
.A2(n_1417),
.B(n_1325),
.Y(n_1504)
);

OA21x2_ASAP7_75t_L g1505 ( 
.A1(n_1422),
.A2(n_1485),
.B(n_1432),
.Y(n_1505)
);

AO21x2_ASAP7_75t_L g1506 ( 
.A1(n_1460),
.A2(n_1418),
.B(n_1407),
.Y(n_1506)
);

OAI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1449),
.A2(n_1368),
.B(n_1410),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1430),
.B(n_1378),
.Y(n_1508)
);

INVx5_ASAP7_75t_L g1509 ( 
.A(n_1484),
.Y(n_1509)
);

O2A1O1Ixp33_ASAP7_75t_L g1510 ( 
.A1(n_1464),
.A2(n_1363),
.B(n_1308),
.C(n_1309),
.Y(n_1510)
);

A2O1A1Ixp33_ASAP7_75t_L g1511 ( 
.A1(n_1448),
.A2(n_1473),
.B(n_1467),
.C(n_1427),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1469),
.A2(n_1364),
.B1(n_1411),
.B2(n_1309),
.Y(n_1512)
);

AO21x2_ASAP7_75t_L g1513 ( 
.A1(n_1431),
.A2(n_1396),
.B(n_1307),
.Y(n_1513)
);

OR2x6_ASAP7_75t_L g1514 ( 
.A(n_1493),
.B(n_1343),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1483),
.B(n_1346),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1461),
.B(n_1409),
.Y(n_1516)
);

OAI21x1_ASAP7_75t_L g1517 ( 
.A1(n_1435),
.A2(n_1334),
.B(n_1310),
.Y(n_1517)
);

OAI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1458),
.A2(n_1400),
.B1(n_1405),
.B2(n_1321),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1492),
.B(n_1396),
.Y(n_1519)
);

AND2x4_ASAP7_75t_L g1520 ( 
.A(n_1454),
.B(n_1478),
.Y(n_1520)
);

AO31x2_ASAP7_75t_L g1521 ( 
.A1(n_1433),
.A2(n_1408),
.A3(n_1334),
.B(n_1386),
.Y(n_1521)
);

AOI21xp33_ASAP7_75t_L g1522 ( 
.A1(n_1425),
.A2(n_1401),
.B(n_1389),
.Y(n_1522)
);

NAND2x1_ASAP7_75t_L g1523 ( 
.A(n_1438),
.B(n_1398),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1438),
.B(n_1389),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1424),
.B(n_1401),
.Y(n_1525)
);

INVx2_ASAP7_75t_SL g1526 ( 
.A(n_1484),
.Y(n_1526)
);

NAND2x1p5_ASAP7_75t_L g1527 ( 
.A(n_1454),
.B(n_1317),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1478),
.Y(n_1528)
);

INVxp67_ASAP7_75t_L g1529 ( 
.A(n_1456),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1436),
.B(n_1340),
.Y(n_1530)
);

OA21x2_ASAP7_75t_L g1531 ( 
.A1(n_1423),
.A2(n_1351),
.B(n_1317),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1487),
.B(n_1351),
.Y(n_1532)
);

O2A1O1Ixp33_ASAP7_75t_SL g1533 ( 
.A1(n_1472),
.A2(n_1336),
.B(n_150),
.C(n_151),
.Y(n_1533)
);

BUFx2_ASAP7_75t_L g1534 ( 
.A(n_1487),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_1457),
.Y(n_1535)
);

OA21x2_ASAP7_75t_L g1536 ( 
.A1(n_1440),
.A2(n_149),
.B(n_152),
.Y(n_1536)
);

INVx5_ASAP7_75t_L g1537 ( 
.A(n_1484),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1420),
.B(n_149),
.Y(n_1538)
);

AND2x4_ASAP7_75t_L g1539 ( 
.A(n_1470),
.B(n_437),
.Y(n_1539)
);

OAI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_1421),
.A2(n_152),
.B(n_153),
.Y(n_1540)
);

AOI21xp5_ASAP7_75t_L g1541 ( 
.A1(n_1434),
.A2(n_449),
.B(n_448),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1445),
.Y(n_1542)
);

NAND3xp33_ASAP7_75t_L g1543 ( 
.A(n_1459),
.B(n_154),
.C(n_155),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1455),
.B(n_438),
.Y(n_1544)
);

AND2x2_ASAP7_75t_SL g1545 ( 
.A(n_1451),
.B(n_155),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1475),
.B(n_1482),
.Y(n_1546)
);

OAI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1500),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_1547)
);

OA21x2_ASAP7_75t_L g1548 ( 
.A1(n_1490),
.A2(n_157),
.B(n_158),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1498),
.Y(n_1549)
);

OAI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1512),
.A2(n_1501),
.B1(n_1491),
.B2(n_1477),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1549),
.B(n_1452),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1503),
.B(n_1441),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_SL g1553 ( 
.A1(n_1540),
.A2(n_1468),
.B(n_1481),
.Y(n_1553)
);

OAI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1511),
.A2(n_1450),
.B(n_1439),
.Y(n_1554)
);

BUFx3_ASAP7_75t_L g1555 ( 
.A(n_1523),
.Y(n_1555)
);

AOI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1506),
.A2(n_1446),
.B(n_1497),
.Y(n_1556)
);

AOI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1506),
.A2(n_1446),
.B(n_1486),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1549),
.B(n_1474),
.Y(n_1558)
);

AOI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1542),
.A2(n_1466),
.B(n_1474),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1546),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1546),
.Y(n_1561)
);

BUFx6f_ASAP7_75t_L g1562 ( 
.A(n_1514),
.Y(n_1562)
);

BUFx2_ASAP7_75t_L g1563 ( 
.A(n_1531),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1508),
.B(n_1442),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1505),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1531),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1513),
.A2(n_1496),
.B(n_1443),
.Y(n_1567)
);

OAI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1502),
.A2(n_1480),
.B(n_1447),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_SL g1569 ( 
.A(n_1507),
.B(n_1471),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1505),
.Y(n_1570)
);

OA21x2_ASAP7_75t_L g1571 ( 
.A1(n_1565),
.A2(n_1507),
.B(n_1517),
.Y(n_1571)
);

BUFx2_ASAP7_75t_L g1572 ( 
.A(n_1563),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1563),
.B(n_1524),
.Y(n_1573)
);

INVxp67_ASAP7_75t_L g1574 ( 
.A(n_1560),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1560),
.B(n_1521),
.Y(n_1575)
);

AOI21x1_ASAP7_75t_L g1576 ( 
.A1(n_1569),
.A2(n_1548),
.B(n_1536),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1561),
.Y(n_1577)
);

INVx3_ASAP7_75t_L g1578 ( 
.A(n_1565),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1561),
.B(n_1545),
.Y(n_1579)
);

AO21x2_ASAP7_75t_L g1580 ( 
.A1(n_1557),
.A2(n_1522),
.B(n_1543),
.Y(n_1580)
);

BUFx6f_ASAP7_75t_L g1581 ( 
.A(n_1562),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1566),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1551),
.B(n_1521),
.Y(n_1583)
);

AO21x2_ASAP7_75t_L g1584 ( 
.A1(n_1570),
.A2(n_1522),
.B(n_1543),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1582),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1572),
.B(n_1566),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1572),
.B(n_1558),
.Y(n_1587)
);

OAI222xp33_ASAP7_75t_L g1588 ( 
.A1(n_1579),
.A2(n_1512),
.B1(n_1550),
.B2(n_1556),
.C1(n_1559),
.C2(n_1552),
.Y(n_1588)
);

NAND3xp33_ASAP7_75t_L g1589 ( 
.A(n_1571),
.B(n_1568),
.C(n_1554),
.Y(n_1589)
);

OAI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1576),
.A2(n_1567),
.B(n_1518),
.Y(n_1590)
);

AOI21xp33_ASAP7_75t_L g1591 ( 
.A1(n_1580),
.A2(n_1553),
.B(n_1465),
.Y(n_1591)
);

A2O1A1Ixp33_ASAP7_75t_L g1592 ( 
.A1(n_1583),
.A2(n_1510),
.B(n_1544),
.C(n_1489),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1581),
.B(n_1575),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1582),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1573),
.Y(n_1595)
);

OAI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1581),
.A2(n_1562),
.B1(n_1559),
.B2(n_1555),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1577),
.B(n_1558),
.Y(n_1597)
);

OAI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1581),
.A2(n_1562),
.B1(n_1555),
.B2(n_1504),
.Y(n_1598)
);

INVx3_ASAP7_75t_L g1599 ( 
.A(n_1578),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1597),
.B(n_1581),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1595),
.B(n_1573),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1597),
.B(n_1587),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1587),
.B(n_1574),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1585),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1585),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1589),
.B(n_1583),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1594),
.Y(n_1607)
);

INVxp67_ASAP7_75t_SL g1608 ( 
.A(n_1606),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1600),
.B(n_1593),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1602),
.B(n_1593),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1603),
.B(n_1593),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1601),
.B(n_1581),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1608),
.A2(n_1590),
.B1(n_1591),
.B2(n_1580),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1608),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1611),
.B(n_1610),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1612),
.Y(n_1616)
);

OAI21xp33_ASAP7_75t_L g1617 ( 
.A1(n_1609),
.A2(n_1592),
.B(n_1564),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1609),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1614),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1615),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1616),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1620),
.B(n_1618),
.Y(n_1622)
);

OAI32xp33_ASAP7_75t_L g1623 ( 
.A1(n_1619),
.A2(n_1613),
.A3(n_1617),
.B1(n_1588),
.B2(n_1605),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1622),
.A2(n_1613),
.B1(n_1621),
.B2(n_1596),
.Y(n_1624)
);

OAI21xp33_ASAP7_75t_L g1625 ( 
.A1(n_1624),
.A2(n_1623),
.B(n_1499),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1625),
.B(n_1535),
.Y(n_1626)
);

AOI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1625),
.A2(n_1562),
.B1(n_1598),
.B2(n_1580),
.Y(n_1627)
);

AOI222xp33_ASAP7_75t_L g1628 ( 
.A1(n_1626),
.A2(n_1547),
.B1(n_1463),
.B2(n_1494),
.C1(n_1495),
.C2(n_1553),
.Y(n_1628)
);

OAI21xp5_ASAP7_75t_SL g1629 ( 
.A1(n_1627),
.A2(n_1529),
.B(n_1562),
.Y(n_1629)
);

AOI221xp5_ASAP7_75t_L g1630 ( 
.A1(n_1629),
.A2(n_1533),
.B1(n_1437),
.B2(n_1453),
.C(n_1462),
.Y(n_1630)
);

NAND2x1_ASAP7_75t_SL g1631 ( 
.A(n_1628),
.B(n_1429),
.Y(n_1631)
);

AOI322xp5_ASAP7_75t_L g1632 ( 
.A1(n_1629),
.A2(n_1586),
.A3(n_1516),
.B1(n_1607),
.B2(n_1604),
.C1(n_1525),
.C2(n_1539),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1631),
.B(n_1488),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1630),
.Y(n_1634)
);

INVx3_ASAP7_75t_SL g1635 ( 
.A(n_1632),
.Y(n_1635)
);

AOI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1633),
.A2(n_1586),
.B1(n_1538),
.B2(n_1539),
.Y(n_1636)
);

O2A1O1Ixp33_ASAP7_75t_L g1637 ( 
.A1(n_1635),
.A2(n_1541),
.B(n_1479),
.C(n_161),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1634),
.Y(n_1638)
);

AOI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1633),
.A2(n_1526),
.B1(n_1584),
.B2(n_1532),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1635),
.B(n_1584),
.Y(n_1640)
);

INVxp67_ASAP7_75t_SL g1641 ( 
.A(n_1633),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1633),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1641),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1638),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1642),
.B(n_1555),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1637),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1640),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1636),
.B(n_1599),
.Y(n_1648)
);

INVxp33_ASAP7_75t_L g1649 ( 
.A(n_1639),
.Y(n_1649)
);

AND3x2_ASAP7_75t_L g1650 ( 
.A(n_1641),
.B(n_1444),
.C(n_159),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1641),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1640),
.B(n_159),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_L g1653 ( 
.A(n_1650),
.B(n_160),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1652),
.Y(n_1654)
);

AO22x2_ASAP7_75t_L g1655 ( 
.A1(n_1644),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1645),
.Y(n_1656)
);

NOR2x1_ASAP7_75t_L g1657 ( 
.A(n_1643),
.B(n_163),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1651),
.B(n_1599),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1646),
.Y(n_1659)
);

NOR2x1_ASAP7_75t_L g1660 ( 
.A(n_1647),
.B(n_163),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1648),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1649),
.B(n_164),
.Y(n_1662)
);

AND2x4_ASAP7_75t_L g1663 ( 
.A(n_1643),
.B(n_1520),
.Y(n_1663)
);

NOR4xp75_ASAP7_75t_L g1664 ( 
.A(n_1645),
.B(n_165),
.C(n_166),
.D(n_168),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1650),
.B(n_165),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1643),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1643),
.B(n_1520),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_SL g1668 ( 
.A(n_1643),
.Y(n_1668)
);

NOR2xp67_ASAP7_75t_L g1669 ( 
.A(n_1652),
.B(n_166),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1650),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1650),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1645),
.B(n_1599),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1652),
.B(n_168),
.Y(n_1673)
);

NOR2x1_ASAP7_75t_L g1674 ( 
.A(n_1652),
.B(n_169),
.Y(n_1674)
);

INVxp33_ASAP7_75t_SL g1675 ( 
.A(n_1643),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1650),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1650),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1650),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1669),
.B(n_1509),
.Y(n_1679)
);

AOI211xp5_ASAP7_75t_L g1680 ( 
.A1(n_1653),
.A2(n_169),
.B(n_170),
.C(n_171),
.Y(n_1680)
);

AOI211xp5_ASAP7_75t_L g1681 ( 
.A1(n_1665),
.A2(n_170),
.B(n_172),
.C(n_173),
.Y(n_1681)
);

NAND4xp25_ASAP7_75t_SL g1682 ( 
.A(n_1670),
.B(n_1678),
.C(n_1677),
.D(n_1676),
.Y(n_1682)
);

NAND4xp25_ASAP7_75t_L g1683 ( 
.A(n_1659),
.B(n_174),
.C(n_175),
.D(n_176),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_SL g1684 ( 
.A(n_1671),
.B(n_1509),
.Y(n_1684)
);

O2A1O1Ixp33_ASAP7_75t_L g1685 ( 
.A1(n_1662),
.A2(n_174),
.B(n_175),
.C(n_176),
.Y(n_1685)
);

AOI221xp5_ASAP7_75t_L g1686 ( 
.A1(n_1675),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.C(n_180),
.Y(n_1686)
);

AOI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1666),
.A2(n_1515),
.B1(n_1584),
.B2(n_1532),
.Y(n_1687)
);

AOI211xp5_ASAP7_75t_L g1688 ( 
.A1(n_1673),
.A2(n_177),
.B(n_180),
.C(n_181),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1657),
.Y(n_1689)
);

AOI221xp5_ASAP7_75t_L g1690 ( 
.A1(n_1658),
.A2(n_181),
.B1(n_183),
.B2(n_184),
.C(n_185),
.Y(n_1690)
);

BUFx2_ASAP7_75t_L g1691 ( 
.A(n_1674),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1668),
.A2(n_1661),
.B1(n_1656),
.B2(n_1654),
.Y(n_1692)
);

AOI221x1_ASAP7_75t_L g1693 ( 
.A1(n_1655),
.A2(n_183),
.B1(n_186),
.B2(n_187),
.C(n_188),
.Y(n_1693)
);

NOR3xp33_ASAP7_75t_L g1694 ( 
.A(n_1660),
.B(n_186),
.C(n_187),
.Y(n_1694)
);

NAND4xp25_ASAP7_75t_SL g1695 ( 
.A(n_1672),
.B(n_1530),
.C(n_1519),
.D(n_190),
.Y(n_1695)
);

AO22x2_ASAP7_75t_L g1696 ( 
.A1(n_1663),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_1696)
);

NOR3xp33_ASAP7_75t_SL g1697 ( 
.A(n_1664),
.B(n_191),
.C(n_192),
.Y(n_1697)
);

OAI311xp33_ASAP7_75t_L g1698 ( 
.A1(n_1667),
.A2(n_1530),
.A3(n_194),
.B1(n_195),
.C1(n_196),
.Y(n_1698)
);

OAI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1655),
.A2(n_1537),
.B1(n_1509),
.B2(n_1594),
.Y(n_1699)
);

AOI221xp5_ASAP7_75t_L g1700 ( 
.A1(n_1670),
.A2(n_193),
.B1(n_194),
.B2(n_196),
.C(n_198),
.Y(n_1700)
);

OAI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1670),
.A2(n_1537),
.B1(n_1528),
.B2(n_1548),
.Y(n_1701)
);

NOR3x2_ASAP7_75t_L g1702 ( 
.A(n_1662),
.B(n_193),
.C(n_198),
.Y(n_1702)
);

O2A1O1Ixp33_ASAP7_75t_L g1703 ( 
.A1(n_1670),
.A2(n_199),
.B(n_200),
.C(n_201),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1655),
.Y(n_1704)
);

XNOR2xp5_ASAP7_75t_L g1705 ( 
.A(n_1664),
.B(n_202),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1675),
.A2(n_1534),
.B1(n_1571),
.B2(n_1537),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1653),
.B(n_203),
.Y(n_1707)
);

OAI211xp5_ASAP7_75t_L g1708 ( 
.A1(n_1670),
.A2(n_203),
.B(n_204),
.C(n_205),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1670),
.B(n_204),
.Y(n_1709)
);

INVxp67_ASAP7_75t_L g1710 ( 
.A(n_1653),
.Y(n_1710)
);

AOI211xp5_ASAP7_75t_L g1711 ( 
.A1(n_1653),
.A2(n_205),
.B(n_206),
.C(n_207),
.Y(n_1711)
);

XNOR2x1_ASAP7_75t_L g1712 ( 
.A(n_1705),
.B(n_206),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1702),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1696),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1683),
.B(n_208),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1691),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1704),
.Y(n_1717)
);

NAND2xp33_ASAP7_75t_L g1718 ( 
.A(n_1697),
.B(n_208),
.Y(n_1718)
);

OR3x2_ASAP7_75t_L g1719 ( 
.A(n_1689),
.B(n_209),
.C(n_211),
.Y(n_1719)
);

NOR2x1_ASAP7_75t_L g1720 ( 
.A(n_1708),
.B(n_1682),
.Y(n_1720)
);

NAND2xp33_ASAP7_75t_L g1721 ( 
.A(n_1694),
.B(n_212),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1709),
.Y(n_1722)
);

AND3x4_ASAP7_75t_L g1723 ( 
.A(n_1698),
.B(n_212),
.C(n_213),
.Y(n_1723)
);

OAI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1692),
.A2(n_1710),
.B(n_1684),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_L g1725 ( 
.A(n_1707),
.B(n_214),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1696),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1703),
.Y(n_1727)
);

NAND4xp75_ASAP7_75t_L g1728 ( 
.A(n_1693),
.B(n_214),
.C(n_215),
.D(n_216),
.Y(n_1728)
);

AO21x2_ASAP7_75t_L g1729 ( 
.A1(n_1679),
.A2(n_215),
.B(n_216),
.Y(n_1729)
);

NOR3xp33_ASAP7_75t_SL g1730 ( 
.A(n_1700),
.B(n_217),
.C(n_218),
.Y(n_1730)
);

NAND3xp33_ASAP7_75t_SL g1731 ( 
.A(n_1680),
.B(n_1711),
.C(n_1681),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1688),
.B(n_217),
.Y(n_1732)
);

NOR3xp33_ASAP7_75t_L g1733 ( 
.A(n_1685),
.B(n_218),
.C(n_219),
.Y(n_1733)
);

XNOR2xp5_ASAP7_75t_L g1734 ( 
.A(n_1686),
.B(n_220),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1699),
.Y(n_1735)
);

XNOR2x1_ASAP7_75t_L g1736 ( 
.A(n_1695),
.B(n_221),
.Y(n_1736)
);

INVx2_ASAP7_75t_SL g1737 ( 
.A(n_1690),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1687),
.B(n_221),
.Y(n_1738)
);

XNOR2x1_ASAP7_75t_L g1739 ( 
.A(n_1701),
.B(n_222),
.Y(n_1739)
);

BUFx2_ASAP7_75t_L g1740 ( 
.A(n_1706),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1709),
.B(n_222),
.Y(n_1741)
);

XNOR2x1_ASAP7_75t_L g1742 ( 
.A(n_1705),
.B(n_223),
.Y(n_1742)
);

NAND2x1p5_ASAP7_75t_L g1743 ( 
.A(n_1691),
.B(n_1528),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1707),
.B(n_224),
.Y(n_1744)
);

AND3x4_ASAP7_75t_L g1745 ( 
.A(n_1697),
.B(n_224),
.C(n_225),
.Y(n_1745)
);

NOR3xp33_ASAP7_75t_SL g1746 ( 
.A(n_1682),
.B(n_226),
.C(n_227),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1696),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1728),
.Y(n_1748)
);

NOR3xp33_ASAP7_75t_SL g1749 ( 
.A(n_1724),
.B(n_226),
.C(n_227),
.Y(n_1749)
);

XNOR2xp5_ASAP7_75t_L g1750 ( 
.A(n_1723),
.B(n_228),
.Y(n_1750)
);

INVx2_ASAP7_75t_SL g1751 ( 
.A(n_1729),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1719),
.Y(n_1752)
);

OAI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1745),
.A2(n_1527),
.B1(n_1571),
.B2(n_1536),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1717),
.B(n_228),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1726),
.B(n_229),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1714),
.Y(n_1756)
);

INVx3_ASAP7_75t_L g1757 ( 
.A(n_1743),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_L g1758 ( 
.A(n_1744),
.B(n_229),
.Y(n_1758)
);

INVx2_ASAP7_75t_SL g1759 ( 
.A(n_1713),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1747),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1736),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1712),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1742),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1746),
.B(n_230),
.Y(n_1764)
);

NAND2x1p5_ASAP7_75t_L g1765 ( 
.A(n_1720),
.B(n_230),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1715),
.B(n_231),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1741),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1765),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1751),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1750),
.Y(n_1770)
);

NAND3xp33_ASAP7_75t_L g1771 ( 
.A(n_1749),
.B(n_1718),
.C(n_1716),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1755),
.Y(n_1772)
);

OAI21x1_ASAP7_75t_L g1773 ( 
.A1(n_1764),
.A2(n_1734),
.B(n_1727),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1754),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1756),
.A2(n_1737),
.B1(n_1725),
.B2(n_1722),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1748),
.B(n_1732),
.Y(n_1776)
);

OAI22x1_ASAP7_75t_L g1777 ( 
.A1(n_1752),
.A2(n_1740),
.B1(n_1735),
.B2(n_1738),
.Y(n_1777)
);

AOI222xp33_ASAP7_75t_L g1778 ( 
.A1(n_1760),
.A2(n_1721),
.B1(n_1731),
.B2(n_1740),
.C1(n_1730),
.C2(n_1739),
.Y(n_1778)
);

INVxp67_ASAP7_75t_L g1779 ( 
.A(n_1758),
.Y(n_1779)
);

OAI21xp33_ASAP7_75t_L g1780 ( 
.A1(n_1778),
.A2(n_1759),
.B(n_1761),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_SL g1781 ( 
.A(n_1768),
.B(n_1733),
.Y(n_1781)
);

XNOR2xp5_ASAP7_75t_L g1782 ( 
.A(n_1777),
.B(n_1763),
.Y(n_1782)
);

AO22x2_ASAP7_75t_L g1783 ( 
.A1(n_1775),
.A2(n_1762),
.B1(n_1767),
.B2(n_1766),
.Y(n_1783)
);

XNOR2x1_ASAP7_75t_L g1784 ( 
.A(n_1776),
.B(n_1757),
.Y(n_1784)
);

AOI21xp5_ASAP7_75t_L g1785 ( 
.A1(n_1769),
.A2(n_1753),
.B(n_234),
.Y(n_1785)
);

AOI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1771),
.A2(n_1770),
.B(n_1772),
.Y(n_1786)
);

AOI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1779),
.A2(n_231),
.B(n_235),
.Y(n_1787)
);

CKINVDCx20_ASAP7_75t_R g1788 ( 
.A(n_1782),
.Y(n_1788)
);

AOI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1780),
.A2(n_1774),
.B1(n_1773),
.B2(n_237),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_SL g1790 ( 
.A1(n_1784),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_1790)
);

OAI22x1_ASAP7_75t_L g1791 ( 
.A1(n_1781),
.A2(n_236),
.B1(n_238),
.B2(n_239),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1783),
.A2(n_1571),
.B1(n_239),
.B2(n_240),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1787),
.Y(n_1793)
);

OAI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1788),
.A2(n_1783),
.B1(n_1786),
.B2(n_1785),
.Y(n_1794)
);

INVx2_ASAP7_75t_SL g1795 ( 
.A(n_1791),
.Y(n_1795)
);

INVxp33_ASAP7_75t_SL g1796 ( 
.A(n_1789),
.Y(n_1796)
);

INVx3_ASAP7_75t_L g1797 ( 
.A(n_1790),
.Y(n_1797)
);

OAI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1796),
.A2(n_1792),
.B1(n_1793),
.B2(n_242),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1797),
.Y(n_1799)
);

OAI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1795),
.A2(n_238),
.B1(n_241),
.B2(n_243),
.Y(n_1800)
);

AOI22x1_ASAP7_75t_L g1801 ( 
.A1(n_1799),
.A2(n_1794),
.B1(n_1798),
.B2(n_1800),
.Y(n_1801)
);

AOI22xp33_ASAP7_75t_L g1802 ( 
.A1(n_1801),
.A2(n_241),
.B1(n_243),
.B2(n_244),
.Y(n_1802)
);

OAI22xp5_ASAP7_75t_SL g1803 ( 
.A1(n_1802),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1803),
.A2(n_245),
.B(n_248),
.Y(n_1804)
);

AOI211xp5_ASAP7_75t_L g1805 ( 
.A1(n_1804),
.A2(n_248),
.B(n_249),
.C(n_439),
.Y(n_1805)
);


endmodule