module fake_jpeg_3160_n_539 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_539);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_539;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_26),
.B(n_10),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_52),
.B(n_69),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_54),
.Y(n_143)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_55),
.Y(n_131)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_57),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_61),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_62),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_32),
.A2(n_10),
.B1(n_17),
.B2(n_2),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_63),
.A2(n_22),
.B1(n_50),
.B2(n_33),
.Y(n_111)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_67),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_11),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_73),
.Y(n_148)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_74),
.Y(n_156)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_31),
.Y(n_81)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_24),
.B(n_11),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_82),
.B(n_83),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_24),
.B(n_11),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_86),
.Y(n_163)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_89),
.Y(n_141)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_94),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_23),
.Y(n_95)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_25),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_100),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_98),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_101),
.Y(n_107)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_103),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_58),
.B(n_50),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_109),
.B(n_114),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_111),
.A2(n_33),
.B1(n_49),
.B2(n_35),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_41),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_87),
.A2(n_28),
.B1(n_43),
.B2(n_45),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_119),
.A2(n_150),
.B1(n_159),
.B2(n_160),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_22),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_122),
.B(n_132),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_95),
.C(n_91),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_124),
.B(n_149),
.C(n_89),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_64),
.B(n_41),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_74),
.B(n_36),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_137),
.B(n_147),
.Y(n_198)
);

AOI21xp33_ASAP7_75t_L g147 ( 
.A1(n_60),
.A2(n_29),
.B(n_49),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_94),
.B(n_103),
.C(n_102),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_85),
.A2(n_43),
.B1(n_45),
.B2(n_30),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_76),
.B(n_51),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_154),
.Y(n_172)
);

OA22x2_ASAP7_75t_L g157 ( 
.A1(n_53),
.A2(n_23),
.B1(n_45),
.B2(n_43),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_157),
.A2(n_46),
.B1(n_40),
.B2(n_35),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_54),
.A2(n_43),
.B1(n_45),
.B2(n_37),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_57),
.A2(n_49),
.B1(n_34),
.B2(n_42),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_86),
.B(n_36),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_104),
.Y(n_168)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_113),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_166),
.Y(n_229)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_167),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_168),
.B(n_175),
.Y(n_255)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_169),
.Y(n_232)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_170),
.Y(n_228)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_173),
.Y(n_252)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_174),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_121),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_176),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_121),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_177),
.Y(n_260)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_178),
.Y(n_238)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_136),
.Y(n_179)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_179),
.Y(n_240)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_128),
.Y(n_180)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_180),
.Y(n_242)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_117),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_181),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_108),
.Y(n_183)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_183),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_184),
.A2(n_193),
.B1(n_212),
.B2(n_223),
.Y(n_272)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_185),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_106),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_186),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_30),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_187),
.B(n_197),
.Y(n_239)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_188),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_116),
.A2(n_30),
.B1(n_34),
.B2(n_42),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_190),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_116),
.A2(n_34),
.B1(n_42),
.B2(n_40),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_191),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_108),
.Y(n_192)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_192),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_157),
.A2(n_62),
.B1(n_99),
.B2(n_98),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_194),
.B(n_201),
.Y(n_262)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_128),
.Y(n_195)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_195),
.Y(n_250)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_196),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_153),
.B(n_23),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_159),
.A2(n_61),
.B1(n_79),
.B2(n_73),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_199),
.A2(n_129),
.B1(n_164),
.B2(n_145),
.Y(n_230)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_112),
.Y(n_200)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_200),
.Y(n_261)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_117),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_110),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_202),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_115),
.B(n_125),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_203),
.B(n_208),
.Y(n_258)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_127),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_204),
.Y(n_241)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_131),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_205),
.Y(n_234)
);

INVx4_ASAP7_75t_SL g206 ( 
.A(n_120),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_206),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_110),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_207),
.Y(n_277)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_131),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_135),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_209),
.B(n_211),
.Y(n_249)
);

OA22x2_ASAP7_75t_L g246 ( 
.A1(n_210),
.A2(n_118),
.B1(n_46),
.B2(n_39),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_135),
.B(n_40),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_119),
.A2(n_67),
.B1(n_101),
.B2(n_35),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_163),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_213),
.B(n_216),
.Y(n_263)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_118),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_214),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_257)
);

FAx1_ASAP7_75t_SL g215 ( 
.A(n_130),
.B(n_60),
.CI(n_66),
.CON(n_215),
.SN(n_215)
);

A2O1A1Ixp33_ASAP7_75t_L g271 ( 
.A1(n_215),
.A2(n_21),
.B(n_11),
.C(n_3),
.Y(n_271)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_146),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_162),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_133),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_133),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_220),
.A2(n_222),
.B1(n_226),
.B2(n_156),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_154),
.B(n_37),
.Y(n_221)
);

NOR2xp67_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_225),
.Y(n_233)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_105),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_150),
.A2(n_101),
.B1(n_39),
.B2(n_37),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_107),
.A2(n_39),
.B(n_46),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_224),
.B(n_0),
.Y(n_276)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_142),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_105),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_210),
.A2(n_160),
.B1(n_157),
.B2(n_142),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_227),
.A2(n_265),
.B1(n_273),
.B2(n_275),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_230),
.A2(n_248),
.B1(n_254),
.B2(n_268),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_194),
.B(n_172),
.C(n_198),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_235),
.B(n_267),
.C(n_278),
.Y(n_302)
);

OA21x2_ASAP7_75t_L g307 ( 
.A1(n_246),
.A2(n_271),
.B(n_4),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_189),
.A2(n_129),
.B1(n_107),
.B2(n_158),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_199),
.A2(n_164),
.B1(n_158),
.B2(n_143),
.Y(n_254)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_259),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_184),
.A2(n_145),
.B1(n_143),
.B2(n_148),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_200),
.B(n_123),
.C(n_120),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_188),
.A2(n_148),
.B1(n_123),
.B2(n_139),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_182),
.A2(n_139),
.B1(n_120),
.B2(n_21),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_270),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_171),
.A2(n_9),
.B1(n_17),
.B2(n_3),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_185),
.A2(n_204),
.B1(n_174),
.B2(n_173),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_218),
.Y(n_291)
);

AND2x2_ASAP7_75t_SL g278 ( 
.A(n_215),
.B(n_0),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_215),
.A2(n_0),
.B(n_1),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_279),
.A2(n_202),
.B(n_217),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_280),
.A2(n_316),
.B(n_307),
.Y(n_328)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_282),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_248),
.A2(n_262),
.B1(n_230),
.B2(n_254),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_283),
.A2(n_292),
.B1(n_295),
.B2(n_299),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_239),
.B(n_258),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_284),
.B(n_286),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_239),
.B(n_167),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_263),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_288),
.B(n_296),
.Y(n_339)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_229),
.Y(n_289)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_289),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_255),
.B(n_170),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_290),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_291),
.B(n_323),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_262),
.A2(n_183),
.B1(n_192),
.B2(n_226),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_213),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_293),
.B(n_294),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_249),
.B(n_181),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_278),
.A2(n_222),
.B1(n_201),
.B2(n_220),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_231),
.B(n_214),
.Y(n_296)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_235),
.B(n_216),
.C(n_195),
.Y(n_297)
);

MAJx2_ASAP7_75t_L g363 ( 
.A(n_297),
.B(n_300),
.C(n_247),
.Y(n_363)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_229),
.Y(n_298)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_298),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_278),
.A2(n_272),
.B1(n_249),
.B2(n_256),
.Y(n_299)
);

MAJx2_ASAP7_75t_L g300 ( 
.A(n_233),
.B(n_180),
.C(n_206),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_276),
.B(n_0),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_301),
.B(n_306),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_256),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_303),
.A2(n_314),
.B1(n_315),
.B2(n_318),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_304),
.A2(n_253),
.B1(n_247),
.B2(n_252),
.Y(n_362)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_229),
.Y(n_305)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_305),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_258),
.B(n_1),
.Y(n_306)
);

OAI21xp33_ASAP7_75t_SL g351 ( 
.A1(n_307),
.A2(n_250),
.B(n_242),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_231),
.B(n_5),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_308),
.B(n_310),
.Y(n_360)
);

INVx6_ASAP7_75t_L g309 ( 
.A(n_264),
.Y(n_309)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_309),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_263),
.B(n_6),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_232),
.B(n_7),
.C(n_9),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_311),
.B(n_261),
.C(n_244),
.Y(n_345)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_245),
.Y(n_312)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_312),
.Y(n_336)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_232),
.Y(n_313)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_313),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_266),
.A2(n_7),
.B1(n_9),
.B2(n_12),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_266),
.A2(n_7),
.B1(n_12),
.B2(n_13),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_279),
.B(n_13),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_316),
.B(n_317),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_234),
.B(n_13),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_270),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_246),
.A2(n_18),
.B1(n_14),
.B2(n_16),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_319),
.A2(n_275),
.B1(n_241),
.B2(n_261),
.Y(n_347)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_245),
.Y(n_320)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_320),
.Y(n_356)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_251),
.Y(n_321)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_321),
.Y(n_367)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_251),
.Y(n_322)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_322),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_246),
.B(n_14),
.Y(n_323)
);

NAND3xp33_ASAP7_75t_L g324 ( 
.A(n_243),
.B(n_236),
.C(n_277),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_324),
.B(n_325),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_237),
.B(n_16),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_246),
.B(n_277),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_326),
.B(n_327),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_237),
.B(n_238),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_328),
.A2(n_343),
.B(n_349),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_281),
.A2(n_265),
.B1(n_259),
.B2(n_271),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_331),
.A2(n_348),
.B1(n_318),
.B2(n_304),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_326),
.A2(n_267),
.B1(n_260),
.B2(n_257),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_332),
.A2(n_335),
.B1(n_362),
.B2(n_298),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_294),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_333),
.B(n_337),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_281),
.A2(n_257),
.B1(n_269),
.B2(n_243),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_308),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_288),
.A2(n_236),
.B(n_238),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_345),
.B(n_274),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_347),
.B(n_351),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_323),
.A2(n_269),
.B1(n_241),
.B2(n_244),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_280),
.A2(n_250),
.B(n_242),
.Y(n_349)
);

OA21x2_ASAP7_75t_L g352 ( 
.A1(n_287),
.A2(n_228),
.B(n_240),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_352),
.B(n_305),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_287),
.A2(n_293),
.B(n_299),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_354),
.A2(n_358),
.B(n_319),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_297),
.B(n_240),
.C(n_253),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_357),
.B(n_330),
.C(n_334),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_295),
.A2(n_283),
.B(n_307),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_363),
.B(n_369),
.Y(n_401)
);

AO21x2_ASAP7_75t_SL g364 ( 
.A1(n_285),
.A2(n_228),
.B(n_252),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_364),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_300),
.A2(n_302),
.B(n_306),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_365),
.A2(n_291),
.B(n_301),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_358),
.A2(n_310),
.B1(n_302),
.B2(n_289),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_370),
.A2(n_375),
.B1(n_389),
.B2(n_352),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_343),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_371),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_372),
.A2(n_392),
.B(n_405),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_L g427 ( 
.A1(n_374),
.A2(n_385),
.B1(n_395),
.B2(n_396),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_340),
.A2(n_292),
.B1(n_313),
.B2(n_321),
.Y(n_375)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_367),
.Y(n_377)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_377),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_378),
.A2(n_386),
.B1(n_399),
.B2(n_347),
.Y(n_406)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_367),
.Y(n_379)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_379),
.Y(n_430)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_368),
.Y(n_380)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_380),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_382),
.B(n_388),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_384),
.B(n_344),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_340),
.A2(n_303),
.B1(n_322),
.B2(n_315),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_368),
.Y(n_387)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_387),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_337),
.B(n_274),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_354),
.A2(n_312),
.B1(n_320),
.B2(n_282),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_336),
.Y(n_390)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_390),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_369),
.B(n_365),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_391),
.B(n_401),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_350),
.A2(n_314),
.B(n_309),
.Y(n_392)
);

INVx5_ASAP7_75t_L g393 ( 
.A(n_364),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_393),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_333),
.A2(n_311),
.B1(n_364),
.B2(n_335),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_394),
.A2(n_362),
.B1(n_352),
.B2(n_342),
.Y(n_410)
);

INVxp33_ASAP7_75t_L g395 ( 
.A(n_346),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_336),
.Y(n_396)
);

OAI32xp33_ASAP7_75t_L g397 ( 
.A1(n_339),
.A2(n_359),
.A3(n_364),
.B1(n_357),
.B2(n_363),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_397),
.B(n_398),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_339),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_331),
.A2(n_332),
.B1(n_364),
.B2(n_348),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_359),
.B(n_341),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_400),
.B(n_329),
.Y(n_436)
);

OR2x2_ASAP7_75t_L g402 ( 
.A(n_352),
.B(n_363),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_402),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_341),
.B(n_345),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_403),
.B(n_404),
.C(n_360),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_349),
.A2(n_328),
.B(n_353),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_406),
.A2(n_415),
.B1(n_394),
.B2(n_375),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_389),
.Y(n_409)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_409),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_410),
.A2(n_414),
.B1(n_417),
.B2(n_419),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_399),
.A2(n_342),
.B1(n_330),
.B2(n_334),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_372),
.A2(n_356),
.B1(n_338),
.B2(n_366),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_381),
.A2(n_356),
.B1(n_338),
.B2(n_366),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_371),
.B(n_360),
.Y(n_420)
);

OR2x2_ASAP7_75t_L g453 ( 
.A(n_420),
.B(n_429),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_391),
.B(n_361),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_421),
.B(n_422),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_401),
.B(n_361),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_398),
.B(n_355),
.Y(n_423)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_423),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_424),
.B(n_434),
.C(n_370),
.Y(n_440)
);

BUFx5_ASAP7_75t_L g425 ( 
.A(n_405),
.Y(n_425)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_425),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_403),
.B(n_355),
.Y(n_426)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_426),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_376),
.B(n_344),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_384),
.B(n_404),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_435),
.B(n_373),
.Y(n_442)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_436),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_429),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_438),
.B(n_418),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_440),
.B(n_446),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_441),
.A2(n_449),
.B1(n_461),
.B2(n_414),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_442),
.B(n_416),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_434),
.B(n_402),
.C(n_373),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_445),
.B(n_447),
.C(n_455),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_421),
.B(n_424),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_408),
.B(n_402),
.C(n_400),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_422),
.B(n_376),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_448),
.B(n_457),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_406),
.A2(n_374),
.B1(n_378),
.B2(n_392),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_411),
.B(n_329),
.Y(n_452)
);

CKINVDCx14_ASAP7_75t_R g476 ( 
.A(n_452),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_407),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_454),
.B(n_433),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_408),
.B(n_383),
.C(n_379),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_412),
.B(n_420),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_456),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_435),
.B(n_383),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_412),
.B(n_377),
.C(n_380),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_458),
.B(n_459),
.C(n_433),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_409),
.B(n_390),
.C(n_396),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_415),
.A2(n_386),
.B1(n_385),
.B2(n_381),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_427),
.B(n_397),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_462),
.B(n_410),
.Y(n_477)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_454),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_463),
.A2(n_468),
.B1(n_471),
.B2(n_481),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_459),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_465),
.Y(n_492)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_453),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_466),
.B(n_469),
.Y(n_494)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_453),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_470),
.B(n_472),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_437),
.A2(n_428),
.B1(n_431),
.B2(n_393),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_458),
.A2(n_416),
.B(n_428),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_475),
.B(n_477),
.Y(n_493)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_439),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_478),
.B(n_479),
.Y(n_491)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_451),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_480),
.B(n_484),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_460),
.A2(n_431),
.B1(n_436),
.B2(n_425),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_444),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_482),
.A2(n_483),
.B1(n_463),
.B2(n_476),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_448),
.B(n_419),
.Y(n_484)
);

BUFx24_ASAP7_75t_SL g485 ( 
.A(n_474),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_485),
.B(n_499),
.Y(n_512)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_487),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_464),
.B(n_446),
.C(n_440),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_488),
.B(n_490),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_464),
.B(n_467),
.C(n_465),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_467),
.B(n_443),
.C(n_455),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_495),
.B(n_498),
.Y(n_511)
);

XNOR2x1_ASAP7_75t_L g496 ( 
.A(n_472),
.B(n_442),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_496),
.B(n_489),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_470),
.B(n_443),
.C(n_445),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_473),
.B(n_475),
.C(n_484),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_481),
.A2(n_450),
.B1(n_462),
.B2(n_417),
.Y(n_500)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_500),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_480),
.A2(n_418),
.B1(n_430),
.B2(n_432),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_501),
.B(n_471),
.Y(n_503)
);

AO21x1_ASAP7_75t_L g502 ( 
.A1(n_492),
.A2(n_457),
.B(n_477),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_502),
.B(n_503),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_494),
.A2(n_447),
.B(n_473),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_506),
.A2(n_509),
.B(n_498),
.Y(n_518)
);

INVx11_ASAP7_75t_L g507 ( 
.A(n_492),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_507),
.A2(n_513),
.B1(n_510),
.B2(n_504),
.Y(n_522)
);

FAx1_ASAP7_75t_SL g508 ( 
.A(n_499),
.B(n_430),
.CI(n_432),
.CON(n_508),
.SN(n_508)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_508),
.B(n_493),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_486),
.A2(n_413),
.B(n_387),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_493),
.A2(n_413),
.B1(n_491),
.B2(n_497),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_514),
.B(n_496),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_505),
.B(n_490),
.C(n_511),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_515),
.B(n_516),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_512),
.B(n_495),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_517),
.A2(n_502),
.B(n_514),
.Y(n_526)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_518),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_510),
.B(n_488),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_520),
.B(n_521),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_522),
.A2(n_504),
.B1(n_507),
.B2(n_509),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_506),
.B(n_513),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_523),
.A2(n_503),
.B(n_508),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_525),
.B(n_526),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_528),
.B(n_519),
.Y(n_531)
);

NOR2xp67_ASAP7_75t_SL g534 ( 
.A(n_531),
.B(n_532),
.Y(n_534)
);

NOR2xp67_ASAP7_75t_L g532 ( 
.A(n_529),
.B(n_515),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_530),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_533),
.B(n_523),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_535),
.B(n_527),
.C(n_524),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_536),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_537),
.A2(n_534),
.B(n_526),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_538),
.A2(n_521),
.B(n_508),
.Y(n_539)
);


endmodule