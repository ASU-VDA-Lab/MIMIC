module fake_jpeg_17411_n_81 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_81);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_81;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_25),
.Y(n_30)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_26),
.B(n_29),
.Y(n_39)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_27),
.B(n_28),
.Y(n_36)
);

INVx5_ASAP7_75t_SL g28 ( 
.A(n_18),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_10),
.B(n_1),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_12),
.B1(n_11),
.B2(n_14),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_31),
.A2(n_11),
.B1(n_12),
.B2(n_19),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_27),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_21),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_18),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_17),
.C(n_19),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_1),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_45),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_47),
.C(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_10),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_46),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_20),
.B1(n_16),
.B2(n_5),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_21),
.C(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_50),
.A2(n_38),
.B1(n_32),
.B2(n_20),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_SL g60 ( 
.A(n_51),
.B(n_55),
.Y(n_60)
);

AOI32xp33_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_36),
.A3(n_22),
.B1(n_38),
.B2(n_39),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_54),
.B(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_36),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_57),
.A2(n_16),
.B1(n_44),
.B2(n_46),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_42),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_65),
.C(n_60),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_49),
.B1(n_41),
.B2(n_33),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_62),
.A2(n_63),
.B1(n_57),
.B2(n_56),
.Y(n_66)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_34),
.C(n_33),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_68),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_70),
.B(n_9),
.Y(n_72)
);

MAJx2_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_34),
.C(n_8),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_73),
.A2(n_2),
.B(n_3),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_68),
.C(n_65),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_74),
.A2(n_75),
.B(n_76),
.Y(n_77)
);

INVxp33_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_70),
.B(n_63),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_77),
.C(n_34),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_2),
.Y(n_81)
);


endmodule