module fake_jpeg_29381_n_159 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_159);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_159;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_54;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_7),
.B(n_27),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_24),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_0),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_1),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_46),
.B(n_2),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_69),
.Y(n_83)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_2),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_73),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_49),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_48),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_55),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_72),
.A2(n_64),
.B1(n_57),
.B2(n_59),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_65),
.C(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_86),
.B(n_64),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_87),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_61),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_88),
.B(n_93),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_92),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_83),
.B(n_63),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_56),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_62),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_102),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_55),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_78),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_101),
.B(n_103),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_54),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_51),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_99),
.A2(n_77),
.B1(n_64),
.B2(n_52),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_106),
.A2(n_122),
.B1(n_30),
.B2(n_31),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_103),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_108),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_89),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_97),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_115),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_121),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_50),
.B(n_59),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_51),
.C(n_52),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_17),
.C(n_19),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_120),
.B1(n_32),
.B2(n_34),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_91),
.B(n_98),
.C(n_89),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_116),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_3),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_118),
.B(n_119),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_5),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_10),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g124 ( 
.A1(n_105),
.A2(n_15),
.B(n_16),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_124),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_129),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_116),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_132),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_135),
.B1(n_137),
.B2(n_138),
.Y(n_144)
);

XNOR2x1_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_28),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_111),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_136),
.Y(n_142)
);

AO22x1_ASAP7_75t_SL g138 ( 
.A1(n_106),
.A2(n_104),
.B1(n_121),
.B2(n_41),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_126),
.A2(n_37),
.B(n_38),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_134),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_146),
.B(n_149),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_144),
.A2(n_123),
.B1(n_125),
.B2(n_132),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_148),
.Y(n_151)
);

HAxp5_ASAP7_75t_SL g149 ( 
.A(n_143),
.B(n_125),
.CON(n_149),
.SN(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_140),
.Y(n_153)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_149),
.C(n_141),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_150),
.Y(n_155)
);

AO21x1_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_142),
.B(n_147),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_139),
.C(n_141),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_157),
.A2(n_138),
.B(n_127),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_145),
.Y(n_159)
);


endmodule