module real_jpeg_21552_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_0),
.A2(n_40),
.B1(n_41),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_0),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_0),
.A2(n_48),
.B1(n_49),
.B2(n_65),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_0),
.A2(n_3),
.B1(n_32),
.B2(n_65),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_0),
.A2(n_5),
.B1(n_27),
.B2(n_65),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_1),
.A2(n_5),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_1),
.A2(n_28),
.B1(n_48),
.B2(n_49),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_2),
.A2(n_3),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_2),
.A2(n_33),
.B1(n_48),
.B2(n_49),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_2),
.A2(n_33),
.B1(n_40),
.B2(n_41),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_2),
.A2(n_5),
.B1(n_27),
.B2(n_33),
.Y(n_120)
);

AOI21xp33_ASAP7_75t_SL g132 ( 
.A1(n_2),
.A2(n_37),
.B(n_41),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_2),
.B(n_80),
.Y(n_145)
);

AOI21xp33_ASAP7_75t_L g160 ( 
.A1(n_2),
.A2(n_5),
.B(n_10),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_2),
.B(n_82),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_SL g183 ( 
.A1(n_2),
.A2(n_49),
.B(n_59),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_3),
.A2(n_33),
.B(n_38),
.C(n_132),
.Y(n_131)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_5),
.B(n_24),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_5),
.A2(n_10),
.B1(n_27),
.B2(n_46),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_5),
.A2(n_7),
.B1(n_27),
.B2(n_50),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_7),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_7),
.A2(n_40),
.B1(n_41),
.B2(n_50),
.Y(n_97)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_9),
.A2(n_32),
.B(n_36),
.C(n_39),
.Y(n_35)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_9),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_10),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_10),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_105),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_104),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_84),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_16),
.B(n_84),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_56),
.C(n_70),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_17),
.B(n_56),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_43),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_29),
.B2(n_42),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_19),
.A2(n_20),
.B1(n_44),
.B2(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_44),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_20),
.A2(n_29),
.B(n_43),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_26),
.Y(n_20)
);

INVxp33_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_22),
.B(n_119),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_25),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_23),
.A2(n_25),
.B1(n_26),
.B2(n_74),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_23),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_23),
.A2(n_24),
.B1(n_120),
.B2(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_25),
.A2(n_74),
.B(n_118),
.Y(n_117)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_25),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_25),
.B(n_33),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_27),
.B(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_34),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_30),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_31),
.B(n_35),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_37),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_33),
.A2(n_46),
.B(n_49),
.C(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_33),
.B(n_45),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_33),
.A2(n_41),
.B(n_60),
.C(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_39),
.Y(n_34)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_59),
.B(n_61),
.C(n_62),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_59),
.Y(n_61)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_44),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B(n_51),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_47),
.B1(n_54),
.B2(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_53),
.B1(n_54),
.B2(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_45),
.B(n_54),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_45),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_49),
.B1(n_59),
.B2(n_60),
.Y(n_62)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_52),
.A2(n_114),
.B(n_115),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_67),
.B(n_69),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_67),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_57),
.A2(n_77),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_57),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_57),
.B(n_144),
.C(n_146),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_57),
.A2(n_128),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_62),
.B1(n_63),
.B2(n_66),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_58),
.Y(n_222)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_62),
.A2(n_96),
.B(n_98),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_82),
.B(n_83),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_66),
.B(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_68),
.B(n_93),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_86),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_70),
.A2(n_71),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_77),
.C(n_81),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_72),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_73),
.A2(n_75),
.B1(n_176),
.B2(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_73),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_75),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_75),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_75),
.B(n_133),
.C(n_174),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_75),
.A2(n_176),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_75),
.B(n_192),
.C(n_199),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_77),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_77),
.B(n_128),
.C(n_129),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_77),
.A2(n_81),
.B1(n_127),
.B2(n_139),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_80),
.B(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_87),
.C(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_81),
.A2(n_123),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_81),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_81),
.A2(n_112),
.B1(n_113),
.B2(n_139),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_81),
.B(n_113),
.C(n_181),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_82),
.B(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_84)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_89),
.B1(n_90),
.B2(n_100),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_87),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_87),
.A2(n_100),
.B1(n_137),
.B2(n_140),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_87),
.A2(n_100),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_87),
.B(n_217),
.C(n_219),
.Y(n_236)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_95),
.B2(n_99),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_95),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_238),
.B(n_243),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_226),
.B(n_237),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_149),
.B(n_207),
.C(n_225),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_135),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_109),
.B(n_135),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_125),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_122),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_111),
.B(n_122),
.C(n_125),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_116),
.B2(n_117),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_112),
.A2(n_113),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_112),
.B(n_117),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_113),
.B(n_159),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_134),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_123),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_130),
.A2(n_131),
.B1(n_133),
.B2(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_166),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_133),
.A2(n_142),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_141),
.C(n_143),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_136),
.B(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_137),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_141),
.B(n_143),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_156),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_146),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_206),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_201),
.B(n_205),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_189),
.B(n_200),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_178),
.B(n_188),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_169),
.B(n_177),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_161),
.B(n_168),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_157),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_165),
.B(n_167),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_171),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_180),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_187),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_182),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_184),
.B(n_186),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_190),
.B(n_191),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_196),
.B2(n_197),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_194),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_198),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_203),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_208),
.B(n_209),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_223),
.B2(n_224),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_216),
.C(n_224),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_223),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_227),
.B(n_228),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_236),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_233),
.B2(n_234),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_234),
.C(n_236),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_240),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);


endmodule