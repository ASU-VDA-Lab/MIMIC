module fake_netlist_5_855_n_2353 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_237, n_90, n_127, n_75, n_101, n_180, n_184, n_226, n_235, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_229, n_108, n_231, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_236, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_46, n_233, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_234, n_17, n_92, n_19, n_149, n_120, n_232, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_225, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_223, n_188, n_190, n_8, n_201, n_158, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_230, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2353);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_237;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_235;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_236;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_46;
input n_233;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_234;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_232;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2353;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2076;
wire n_2031;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_2323;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_291;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_2249;
wire n_344;
wire n_1218;
wire n_1931;
wire n_2276;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_2300;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_283;
wire n_1403;
wire n_2248;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_310;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2324;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_407;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_857;
wire n_832;
wire n_2305;
wire n_561;
wire n_1319;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_604;
wire n_433;
wire n_368;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2320;
wire n_2339;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_2299;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_2346;
wire n_662;
wire n_459;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_1574;
wire n_473;
wire n_2048;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_2277;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_1982;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_860;
wire n_441;
wire n_450;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1205;
wire n_1044;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_2198;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_2266;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_2333;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_378;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_2289;
wire n_302;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_321;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_2269;
wire n_2309;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_2310;
wire n_323;
wire n_2287;
wire n_356;
wire n_2291;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_1735;
wire n_1575;
wire n_1697;
wire n_833;
wire n_2318;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2282;
wire n_2002;
wire n_510;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2340;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2148;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1726;
wire n_665;
wire n_1584;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1543;
wire n_1399;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_2286;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_2136;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_2332;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2183;
wire n_328;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_2278;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_1654;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1956;
wire n_1936;
wire n_437;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_2273;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;
wire n_2268;

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_156),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_47),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_15),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_110),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_187),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_98),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_56),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_103),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_38),
.Y(n_246)
);

BUFx5_ASAP7_75t_L g247 ( 
.A(n_85),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_213),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_203),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_158),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_96),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_232),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_1),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_66),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_182),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_72),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_25),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_129),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_202),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_4),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_86),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_150),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_32),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_55),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_91),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_231),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_141),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_70),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_120),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_113),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_169),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_128),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_37),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_41),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_76),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_60),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_135),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_27),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_210),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_11),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_176),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_57),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_217),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_145),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_188),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_45),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_130),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_180),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_173),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_208),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_229),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_40),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_237),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_172),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_147),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_171),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_3),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_78),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_24),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_72),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_64),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_4),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_207),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_228),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_152),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_148),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_11),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_52),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_68),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_95),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_167),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_127),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_206),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_100),
.Y(n_314)
);

BUFx5_ASAP7_75t_L g315 ( 
.A(n_7),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_183),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_193),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_14),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_219),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_107),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_174),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_149),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_64),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_104),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_119),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_77),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_51),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_27),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_200),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_197),
.Y(n_330)
);

BUFx10_ASAP7_75t_L g331 ( 
.A(n_83),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_51),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_94),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_137),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_136),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_29),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_61),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_170),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_74),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_23),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_47),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_19),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_65),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_84),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_31),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_30),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_185),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_92),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_218),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_142),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_175),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_163),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_82),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_223),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_10),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_70),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_190),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_57),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_144),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_125),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_162),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_40),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_124),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_121),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_56),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_78),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_224),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_134),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_133),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_76),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_75),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_75),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_186),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_17),
.Y(n_374)
);

BUFx10_ASAP7_75t_L g375 ( 
.A(n_26),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_28),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_77),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_89),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_37),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_25),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_230),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_53),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_235),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_181),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_55),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_204),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_184),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_14),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_71),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_165),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_109),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_221),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_234),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_17),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_79),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_216),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_20),
.Y(n_397)
);

BUFx10_ASAP7_75t_L g398 ( 
.A(n_24),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_44),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_32),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_117),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_225),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_222),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_168),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_49),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_153),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_22),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_90),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_122),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_192),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_23),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_66),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_10),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_73),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_99),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_106),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_79),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_138),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_54),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_43),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_236),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_16),
.Y(n_422)
);

BUFx10_ASAP7_75t_L g423 ( 
.A(n_140),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_199),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_46),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_215),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_97),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_179),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_81),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_26),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_30),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_44),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_233),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_114),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_205),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_45),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_31),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_220),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_194),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_191),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_93),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_166),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_155),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_131),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_43),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_39),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_226),
.Y(n_447)
);

INVxp67_ASAP7_75t_SL g448 ( 
.A(n_198),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_6),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_42),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_7),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_116),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_5),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_1),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_112),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_69),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_49),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_33),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_108),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_67),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_214),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_5),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_161),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_105),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_87),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_299),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_315),
.B(n_0),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_446),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_315),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_300),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_315),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_315),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_307),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_315),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_258),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_308),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_315),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_265),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_361),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_315),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_309),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_318),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_267),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_315),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_240),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_282),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_283),
.Y(n_487)
);

INVxp67_ASAP7_75t_SL g488 ( 
.A(n_421),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_297),
.Y(n_489)
);

NOR2xp67_ASAP7_75t_L g490 ( 
.A(n_292),
.B(n_0),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_297),
.Y(n_491)
);

INVxp67_ASAP7_75t_SL g492 ( 
.A(n_434),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_297),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_334),
.B(n_2),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_297),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_297),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_302),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_338),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_386),
.Y(n_499)
);

INVxp67_ASAP7_75t_SL g500 ( 
.A(n_243),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_282),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_343),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_387),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_243),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_438),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_343),
.Y(n_506)
);

INVxp67_ASAP7_75t_SL g507 ( 
.A(n_302),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_334),
.B(n_2),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_345),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_250),
.B(n_3),
.Y(n_510)
);

INVxp67_ASAP7_75t_SL g511 ( 
.A(n_302),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_455),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_345),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_R g514 ( 
.A(n_304),
.B(n_88),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_327),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_436),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_328),
.Y(n_517)
);

CKINVDCx16_ASAP7_75t_R g518 ( 
.A(n_249),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_250),
.B(n_6),
.Y(n_519)
);

CKINVDCx16_ASAP7_75t_R g520 ( 
.A(n_364),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_331),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_332),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_302),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_426),
.Y(n_524)
);

INVxp33_ASAP7_75t_SL g525 ( 
.A(n_240),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_436),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_302),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_291),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_293),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_246),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_244),
.Y(n_531)
);

NOR2xp67_ASAP7_75t_L g532 ( 
.A(n_292),
.B(n_8),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_294),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_247),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_337),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_257),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_296),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_303),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_339),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_273),
.Y(n_540)
);

INVxp33_ASAP7_75t_SL g541 ( 
.A(n_246),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_276),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_278),
.Y(n_543)
);

INVxp67_ASAP7_75t_SL g544 ( 
.A(n_248),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_346),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_305),
.Y(n_546)
);

OR2x2_ASAP7_75t_L g547 ( 
.A(n_298),
.B(n_8),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_306),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_301),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_323),
.Y(n_550)
);

CKINVDCx16_ASAP7_75t_R g551 ( 
.A(n_331),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_262),
.B(n_9),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_353),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_326),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_336),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_311),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_314),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_355),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_341),
.Y(n_559)
);

INVxp67_ASAP7_75t_SL g560 ( 
.A(n_255),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_331),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_262),
.B(n_9),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_344),
.Y(n_563)
);

CKINVDCx16_ASAP7_75t_R g564 ( 
.A(n_375),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_356),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_317),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_358),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_288),
.B(n_12),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_319),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_370),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_371),
.Y(n_571)
);

INVxp33_ASAP7_75t_SL g572 ( 
.A(n_253),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_374),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_320),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_321),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_385),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_286),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_362),
.Y(n_578)
);

INVxp67_ASAP7_75t_SL g579 ( 
.A(n_266),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_361),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_324),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_253),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_397),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_286),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_414),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_423),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_365),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_366),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_417),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_419),
.Y(n_590)
);

NOR2xp67_ASAP7_75t_L g591 ( 
.A(n_411),
.B(n_12),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_420),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_372),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_485),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_472),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_466),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_490),
.B(n_423),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_507),
.B(n_238),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_479),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_544),
.B(n_288),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_489),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_489),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_479),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_491),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_511),
.B(n_391),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_479),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_491),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_560),
.B(n_391),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_579),
.B(n_408),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_SL g610 ( 
.A1(n_475),
.A2(n_239),
.B1(n_394),
.B2(n_340),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_523),
.B(n_408),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_472),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_493),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_479),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_479),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_493),
.B(n_427),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_495),
.Y(n_617)
);

OA21x2_ASAP7_75t_L g618 ( 
.A1(n_467),
.A2(n_432),
.B(n_430),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_530),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_466),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_500),
.B(n_427),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_495),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_580),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_496),
.B(n_452),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_527),
.B(n_494),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_580),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_496),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_497),
.Y(n_628)
);

AND3x2_ASAP7_75t_L g629 ( 
.A(n_519),
.B(n_452),
.C(n_445),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g630 ( 
.A(n_582),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_508),
.B(n_238),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_580),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_580),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_497),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_580),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_478),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_469),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_471),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_534),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_474),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_477),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_480),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_484),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_470),
.Y(n_644)
);

NAND2xp33_ASAP7_75t_SL g645 ( 
.A(n_547),
.B(n_411),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_534),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_577),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_510),
.B(n_270),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_577),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_483),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_584),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_562),
.B(n_241),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_584),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_552),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_568),
.B(n_241),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_531),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_536),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_540),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_504),
.B(n_242),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_582),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_542),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_543),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_549),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_532),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_550),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_554),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_504),
.B(n_242),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_555),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_559),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_563),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_470),
.Y(n_671)
);

AND2x2_ASAP7_75t_SL g672 ( 
.A(n_547),
.B(n_361),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_567),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_591),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_570),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_486),
.B(n_245),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_571),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_573),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_576),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_583),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_501),
.B(n_462),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_585),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_589),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_502),
.B(n_506),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_514),
.B(n_423),
.Y(n_685)
);

OAI22xp5_ASAP7_75t_L g686 ( 
.A1(n_468),
.A2(n_456),
.B1(n_342),
.B2(n_453),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_590),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_592),
.Y(n_688)
);

HB1xp67_ASAP7_75t_L g689 ( 
.A(n_473),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_518),
.B(n_375),
.Y(n_690)
);

OA21x2_ASAP7_75t_L g691 ( 
.A1(n_509),
.A2(n_449),
.B(n_437),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_631),
.B(n_520),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_638),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_685),
.B(n_551),
.Y(n_694)
);

NOR3xp33_ASAP7_75t_L g695 ( 
.A(n_686),
.B(n_564),
.C(n_492),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_638),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_595),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_672),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_595),
.Y(n_699)
);

INVx1_ASAP7_75t_SL g700 ( 
.A(n_636),
.Y(n_700)
);

OR2x2_ASAP7_75t_L g701 ( 
.A(n_598),
.B(n_488),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_654),
.B(n_473),
.Y(n_702)
);

BUFx4f_ASAP7_75t_L g703 ( 
.A(n_618),
.Y(n_703)
);

AO22x2_ASAP7_75t_L g704 ( 
.A1(n_686),
.A2(n_462),
.B1(n_460),
.B2(n_458),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_672),
.Y(n_705)
);

INVxp33_ASAP7_75t_L g706 ( 
.A(n_660),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_618),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_595),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_685),
.B(n_476),
.Y(n_709)
);

INVx4_ASAP7_75t_L g710 ( 
.A(n_642),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_640),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_640),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_612),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_643),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_643),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_612),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_612),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_646),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_618),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_646),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_605),
.B(n_448),
.Y(n_721)
);

OR2x2_ASAP7_75t_L g722 ( 
.A(n_598),
.B(n_521),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_646),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_637),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_637),
.Y(n_725)
);

NOR3xp33_ASAP7_75t_L g726 ( 
.A(n_610),
.B(n_561),
.C(n_481),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_637),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_641),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_641),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_641),
.Y(n_730)
);

BUFx10_ASAP7_75t_L g731 ( 
.A(n_672),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_SL g732 ( 
.A(n_672),
.B(n_524),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_661),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_631),
.B(n_525),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_SL g735 ( 
.A(n_597),
.B(n_476),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_629),
.Y(n_736)
);

INVx5_ASAP7_75t_L g737 ( 
.A(n_642),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_661),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_601),
.Y(n_739)
);

BUFx2_ASAP7_75t_L g740 ( 
.A(n_664),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_654),
.B(n_481),
.Y(n_741)
);

INVxp67_ASAP7_75t_SL g742 ( 
.A(n_603),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_654),
.B(n_482),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_601),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_599),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_605),
.B(n_272),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_618),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_599),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_654),
.B(n_482),
.Y(n_749)
);

INVx5_ASAP7_75t_L g750 ( 
.A(n_642),
.Y(n_750)
);

OR2x6_ASAP7_75t_L g751 ( 
.A(n_659),
.B(n_277),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_661),
.Y(n_752)
);

INVxp33_ASAP7_75t_SL g753 ( 
.A(n_610),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_602),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_602),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_661),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_652),
.B(n_525),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_661),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_621),
.B(n_600),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_652),
.B(n_541),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_599),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_687),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_599),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_599),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_654),
.B(n_515),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_604),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_655),
.B(n_541),
.Y(n_767)
);

INVx5_ASAP7_75t_L g768 ( 
.A(n_642),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_664),
.B(n_515),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_687),
.Y(n_770)
);

INVx4_ASAP7_75t_L g771 ( 
.A(n_642),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_655),
.B(n_572),
.Y(n_772)
);

AND2x6_ASAP7_75t_L g773 ( 
.A(n_654),
.B(n_361),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_599),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_636),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_604),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_674),
.B(n_517),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_607),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_687),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_674),
.B(n_517),
.Y(n_780)
);

NAND3xp33_ASAP7_75t_L g781 ( 
.A(n_618),
.B(n_516),
.C(n_513),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_687),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_607),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_613),
.Y(n_784)
);

NAND2xp33_ASAP7_75t_L g785 ( 
.A(n_654),
.B(n_522),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_687),
.Y(n_786)
);

INVx5_ASAP7_75t_L g787 ( 
.A(n_642),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_613),
.Y(n_788)
);

BUFx2_ASAP7_75t_L g789 ( 
.A(n_660),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_654),
.B(n_522),
.Y(n_790)
);

INVx5_ASAP7_75t_L g791 ( 
.A(n_642),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_621),
.B(n_535),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_605),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_648),
.A2(n_572),
.B1(n_526),
.B2(n_361),
.Y(n_794)
);

INVx4_ASAP7_75t_L g795 ( 
.A(n_639),
.Y(n_795)
);

INVx1_ASAP7_75t_SL g796 ( 
.A(n_650),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_617),
.Y(n_797)
);

AND2x6_ASAP7_75t_L g798 ( 
.A(n_648),
.B(n_281),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_617),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_621),
.B(n_586),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_599),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_622),
.Y(n_802)
);

NAND2xp33_ASAP7_75t_L g803 ( 
.A(n_659),
.B(n_593),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_605),
.B(n_535),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_600),
.B(n_586),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_622),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_615),
.Y(n_807)
);

NAND2xp33_ASAP7_75t_SL g808 ( 
.A(n_597),
.B(n_539),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_627),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_627),
.Y(n_810)
);

CKINVDCx6p67_ASAP7_75t_R g811 ( 
.A(n_650),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_628),
.Y(n_812)
);

BUFx2_ASAP7_75t_L g813 ( 
.A(n_630),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_605),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_611),
.B(n_287),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_667),
.B(n_528),
.Y(n_816)
);

OR2x6_ASAP7_75t_L g817 ( 
.A(n_667),
.B(n_295),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_596),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_628),
.Y(n_819)
);

INVx3_ASAP7_75t_L g820 ( 
.A(n_615),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_619),
.B(n_529),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_615),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_634),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_615),
.Y(n_824)
);

BUFx10_ASAP7_75t_L g825 ( 
.A(n_648),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_634),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_611),
.B(n_539),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_619),
.B(n_533),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_611),
.B(n_600),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_611),
.B(n_608),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_608),
.B(n_545),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_639),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_611),
.B(n_310),
.Y(n_833)
);

INVxp33_ASAP7_75t_L g834 ( 
.A(n_594),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_615),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_625),
.B(n_537),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_616),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_615),
.Y(n_838)
);

NOR2x1p5_ASAP7_75t_L g839 ( 
.A(n_676),
.B(n_254),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_608),
.B(n_545),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_616),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_639),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_629),
.Y(n_843)
);

NAND2xp33_ASAP7_75t_SL g844 ( 
.A(n_594),
.B(n_553),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_648),
.A2(n_313),
.B1(n_316),
.B2(n_312),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_609),
.B(n_684),
.Y(n_846)
);

OAI22xp33_ASAP7_75t_L g847 ( 
.A1(n_630),
.A2(n_377),
.B1(n_379),
.B2(n_376),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_596),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_639),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_639),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_615),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_616),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_649),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_793),
.Y(n_854)
);

INVx1_ASAP7_75t_SL g855 ( 
.A(n_789),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_698),
.B(n_648),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_739),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_698),
.A2(n_645),
.B1(n_691),
.B2(n_609),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_705),
.B(n_759),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_800),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_793),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_731),
.B(n_596),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_705),
.B(n_609),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_759),
.B(n_625),
.Y(n_864)
);

NAND2x1p5_ASAP7_75t_L g865 ( 
.A(n_793),
.B(n_691),
.Y(n_865)
);

AOI22xp5_ASAP7_75t_L g866 ( 
.A1(n_757),
.A2(n_689),
.B1(n_644),
.B2(n_671),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_829),
.B(n_691),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_814),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_805),
.B(n_620),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_739),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_814),
.Y(n_871)
);

NAND2xp33_ASAP7_75t_L g872 ( 
.A(n_798),
.B(n_689),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_744),
.Y(n_873)
);

AOI221xp5_ASAP7_75t_L g874 ( 
.A1(n_704),
.A2(n_645),
.B1(n_451),
.B2(n_457),
.C(n_254),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_731),
.B(n_620),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_830),
.B(n_691),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_814),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_837),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_731),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_837),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_734),
.B(n_721),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_721),
.B(n_691),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_721),
.B(n_676),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_744),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_707),
.A2(n_681),
.B1(n_624),
.B2(n_616),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_721),
.B(n_666),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_754),
.Y(n_887)
);

XNOR2xp5_ASAP7_75t_L g888 ( 
.A(n_775),
.B(n_487),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_841),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_841),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_731),
.B(n_620),
.Y(n_891)
);

INVx5_ASAP7_75t_L g892 ( 
.A(n_773),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_702),
.B(n_666),
.Y(n_893)
);

AND2x4_ASAP7_75t_SL g894 ( 
.A(n_811),
.B(n_498),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_741),
.B(n_666),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_825),
.B(n_644),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_805),
.B(n_644),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_743),
.B(n_666),
.Y(n_898)
);

AOI21x1_ASAP7_75t_L g899 ( 
.A1(n_693),
.A2(n_623),
.B(n_614),
.Y(n_899)
);

INVxp67_ASAP7_75t_L g900 ( 
.A(n_740),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_800),
.B(n_671),
.Y(n_901)
);

NAND2xp33_ASAP7_75t_L g902 ( 
.A(n_798),
.B(n_247),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_825),
.B(n_671),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_852),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_749),
.B(n_666),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_754),
.Y(n_906)
);

AOI21x1_ASAP7_75t_L g907 ( 
.A1(n_693),
.A2(n_623),
.B(n_614),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_825),
.B(n_247),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_755),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_825),
.B(n_247),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_765),
.B(n_247),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_852),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_790),
.B(n_247),
.Y(n_913)
);

AO22x1_ASAP7_75t_L g914 ( 
.A1(n_760),
.A2(n_558),
.B1(n_565),
.B2(n_553),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_767),
.B(n_772),
.Y(n_915)
);

NOR2xp67_ASAP7_75t_L g916 ( 
.A(n_821),
.B(n_558),
.Y(n_916)
);

OR2x2_ASAP7_75t_L g917 ( 
.A(n_722),
.B(n_565),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_696),
.B(n_666),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_696),
.B(n_666),
.Y(n_919)
);

NOR2xp67_ASAP7_75t_L g920 ( 
.A(n_828),
.B(n_578),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_755),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_722),
.B(n_578),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_766),
.Y(n_923)
);

OR2x2_ASAP7_75t_L g924 ( 
.A(n_789),
.B(n_587),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_701),
.B(n_690),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_740),
.Y(n_926)
);

BUFx6f_ASAP7_75t_SL g927 ( 
.A(n_736),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_711),
.B(n_678),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_703),
.B(n_247),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_701),
.B(n_690),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_711),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_836),
.B(n_538),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_822),
.Y(n_933)
);

INVxp67_ASAP7_75t_L g934 ( 
.A(n_813),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_766),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_792),
.B(n_840),
.Y(n_936)
);

AOI22xp5_ASAP7_75t_L g937 ( 
.A1(n_732),
.A2(n_548),
.B1(n_556),
.B2(n_546),
.Y(n_937)
);

NAND3xp33_ASAP7_75t_L g938 ( 
.A(n_794),
.B(n_588),
.C(n_587),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_712),
.B(n_678),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_703),
.B(n_247),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_703),
.B(n_657),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_712),
.B(n_678),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_714),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_714),
.B(n_678),
.Y(n_944)
);

AOI22xp33_ASAP7_75t_L g945 ( 
.A1(n_707),
.A2(n_681),
.B1(n_624),
.B2(n_616),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_715),
.B(n_678),
.Y(n_946)
);

NOR3xp33_ASAP7_75t_L g947 ( 
.A(n_844),
.B(n_593),
.C(n_588),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_715),
.B(n_678),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_692),
.A2(n_566),
.B1(n_569),
.B2(n_557),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_846),
.B(n_678),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_707),
.B(n_657),
.Y(n_951)
);

NOR3xp33_ASAP7_75t_L g952 ( 
.A(n_694),
.B(n_816),
.C(n_709),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_797),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_719),
.B(n_657),
.Y(n_954)
);

BUFx6f_ASAP7_75t_SL g955 ( 
.A(n_736),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_776),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_846),
.B(n_657),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_804),
.B(n_657),
.Y(n_958)
);

AOI22xp33_ASAP7_75t_L g959 ( 
.A1(n_719),
.A2(n_681),
.B1(n_624),
.B2(n_325),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_719),
.B(n_657),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_827),
.B(n_657),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_831),
.B(n_684),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_746),
.B(n_657),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_797),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_799),
.Y(n_965)
);

AOI22xp33_ASAP7_75t_L g966 ( 
.A1(n_747),
.A2(n_624),
.B1(n_330),
.B2(n_333),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_776),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_778),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_778),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_747),
.B(n_673),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_L g971 ( 
.A1(n_747),
.A2(n_624),
.B1(n_335),
.B2(n_350),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_799),
.Y(n_972)
);

NOR3xp33_ASAP7_75t_L g973 ( 
.A(n_843),
.B(n_684),
.C(n_663),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_843),
.B(n_662),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_806),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_783),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_746),
.B(n_673),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_746),
.B(n_673),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_806),
.Y(n_979)
);

INVxp67_ASAP7_75t_L g980 ( 
.A(n_813),
.Y(n_980)
);

AND2x6_ASAP7_75t_L g981 ( 
.A(n_733),
.B(n_322),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_706),
.B(n_831),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_783),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_746),
.B(n_673),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_815),
.B(n_673),
.Y(n_985)
);

NAND2xp33_ASAP7_75t_L g986 ( 
.A(n_798),
.B(n_329),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_784),
.Y(n_987)
);

INVx2_ASAP7_75t_SL g988 ( 
.A(n_839),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_819),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_815),
.B(n_673),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_815),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_815),
.B(n_673),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_834),
.B(n_848),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_742),
.A2(n_626),
.B(n_615),
.Y(n_994)
);

INVxp67_ASAP7_75t_L g995 ( 
.A(n_769),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_785),
.A2(n_575),
.B1(n_581),
.B2(n_574),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_833),
.B(n_673),
.Y(n_997)
);

OR2x6_ASAP7_75t_L g998 ( 
.A(n_751),
.B(n_662),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_781),
.B(n_680),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_833),
.B(n_680),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_819),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_781),
.B(n_680),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_833),
.B(n_680),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_848),
.B(n_499),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_833),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_823),
.B(n_680),
.Y(n_1006)
);

OR2x6_ASAP7_75t_L g1007 ( 
.A(n_751),
.B(n_663),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_777),
.B(n_392),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_823),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_826),
.B(n_751),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_780),
.B(n_669),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_826),
.Y(n_1012)
);

INVx2_ASAP7_75t_SL g1013 ( 
.A(n_839),
.Y(n_1013)
);

NAND2xp33_ASAP7_75t_L g1014 ( 
.A(n_798),
.B(n_347),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_784),
.Y(n_1015)
);

OAI22xp33_ASAP7_75t_SL g1016 ( 
.A1(n_753),
.A2(n_413),
.B1(n_256),
.B2(n_260),
.Y(n_1016)
);

INVx2_ASAP7_75t_SL g1017 ( 
.A(n_751),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_795),
.Y(n_1018)
);

INVxp67_ASAP7_75t_L g1019 ( 
.A(n_700),
.Y(n_1019)
);

NAND3x1_ASAP7_75t_L g1020 ( 
.A(n_726),
.B(n_363),
.C(n_354),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_795),
.B(n_680),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_751),
.B(n_680),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_798),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_817),
.B(n_680),
.Y(n_1024)
);

NAND2xp33_ASAP7_75t_L g1025 ( 
.A(n_798),
.B(n_773),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_795),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_882),
.A2(n_795),
.B(n_738),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_915),
.B(n_817),
.Y(n_1028)
);

OAI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_929),
.A2(n_738),
.B(n_733),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_857),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_932),
.B(n_503),
.Y(n_1031)
);

AOI21x1_ASAP7_75t_L g1032 ( 
.A1(n_941),
.A2(n_756),
.B(n_752),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_881),
.A2(n_756),
.B(n_752),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_878),
.Y(n_1034)
);

INVx4_ASAP7_75t_L g1035 ( 
.A(n_879),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_991),
.Y(n_1036)
);

AO21x1_ASAP7_75t_L g1037 ( 
.A1(n_929),
.A2(n_808),
.B(n_735),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_936),
.B(n_864),
.Y(n_1038)
);

INVxp67_ASAP7_75t_L g1039 ( 
.A(n_993),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_880),
.Y(n_1040)
);

OAI321xp33_ASAP7_75t_L g1041 ( 
.A1(n_925),
.A2(n_847),
.A3(n_817),
.B1(n_845),
.B2(n_428),
.C(n_410),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_936),
.A2(n_803),
.B1(n_817),
.B2(n_512),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_856),
.A2(n_762),
.B(n_758),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_886),
.A2(n_762),
.B(n_758),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_932),
.B(n_505),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_883),
.B(n_817),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_925),
.A2(n_770),
.B(n_782),
.C(n_779),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_867),
.A2(n_779),
.B(n_770),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_876),
.A2(n_786),
.B(n_782),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_940),
.A2(n_786),
.B(n_727),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_859),
.A2(n_788),
.B(n_809),
.C(n_802),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_1018),
.A2(n_771),
.B(n_710),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_861),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_863),
.B(n_798),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_930),
.A2(n_788),
.B(n_809),
.C(n_802),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_930),
.A2(n_695),
.B1(n_773),
.B2(n_810),
.Y(n_1056)
);

OAI21xp33_ASAP7_75t_L g1057 ( 
.A1(n_1008),
.A2(n_704),
.B(n_753),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_855),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_931),
.B(n_943),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_940),
.A2(n_727),
.B(n_725),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_889),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_1018),
.A2(n_1026),
.B(n_895),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_SL g1063 ( 
.A(n_1004),
.B(n_796),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_1026),
.A2(n_771),
.B(n_710),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_SL g1065 ( 
.A(n_1019),
.B(n_811),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_953),
.B(n_964),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_893),
.A2(n_771),
.B(n_710),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_899),
.A2(n_820),
.B(n_807),
.Y(n_1068)
);

O2A1O1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_1010),
.A2(n_812),
.B(n_810),
.C(n_725),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_898),
.A2(n_771),
.B(n_710),
.Y(n_1070)
);

AO21x1_ASAP7_75t_L g1071 ( 
.A1(n_911),
.A2(n_373),
.B(n_369),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_934),
.B(n_818),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_965),
.B(n_972),
.Y(n_1073)
);

O2A1O1Ixp5_ASAP7_75t_L g1074 ( 
.A1(n_911),
.A2(n_853),
.B(n_728),
.C(n_730),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_991),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_926),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_980),
.B(n_245),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_975),
.B(n_853),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_979),
.B(n_729),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_860),
.B(n_669),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_989),
.B(n_729),
.Y(n_1081)
);

AOI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_952),
.A2(n_1008),
.B1(n_1017),
.B2(n_901),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_857),
.Y(n_1083)
);

AOI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_897),
.A2(n_773),
.B1(n_724),
.B2(n_730),
.Y(n_1084)
);

NAND2xp33_ASAP7_75t_SL g1085 ( 
.A(n_927),
.B(n_251),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_905),
.A2(n_824),
.B(n_822),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_890),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_958),
.A2(n_824),
.B(n_822),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1001),
.B(n_1009),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_870),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_904),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_862),
.A2(n_728),
.B(n_724),
.C(n_679),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_917),
.B(n_251),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_900),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_996),
.B(n_962),
.Y(n_1095)
);

INVxp67_ASAP7_75t_L g1096 ( 
.A(n_982),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_961),
.A2(n_824),
.B(n_822),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_862),
.A2(n_891),
.B(n_875),
.C(n_896),
.Y(n_1098)
);

OAI21xp33_ASAP7_75t_SL g1099 ( 
.A1(n_858),
.A2(n_396),
.B(n_384),
.Y(n_1099)
);

OR2x2_ASAP7_75t_L g1100 ( 
.A(n_922),
.B(n_677),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_941),
.A2(n_824),
.B(n_822),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1012),
.B(n_861),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_966),
.B(n_807),
.Y(n_1103)
);

INVx2_ASAP7_75t_SL g1104 ( 
.A(n_924),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_SL g1105 ( 
.A(n_894),
.B(n_252),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_916),
.B(n_252),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_870),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_894),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_1011),
.A2(n_403),
.B(n_404),
.C(n_402),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_966),
.B(n_807),
.Y(n_1110)
);

INVx1_ASAP7_75t_SL g1111 ( 
.A(n_888),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_995),
.B(n_259),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_1005),
.B(n_677),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_912),
.Y(n_1114)
);

AOI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_854),
.A2(n_773),
.B1(n_704),
.B2(n_832),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_951),
.A2(n_699),
.B(n_697),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_950),
.A2(n_842),
.B(n_832),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_957),
.A2(n_849),
.B(n_842),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_1011),
.A2(n_442),
.B(n_461),
.C(n_435),
.Y(n_1119)
);

AOI22x1_ASAP7_75t_L g1120 ( 
.A1(n_865),
.A2(n_704),
.B1(n_851),
.B2(n_820),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_866),
.B(n_259),
.Y(n_1121)
);

OR2x2_ASAP7_75t_L g1122 ( 
.A(n_949),
.B(n_679),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_971),
.B(n_820),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_954),
.A2(n_850),
.B(n_849),
.Y(n_1124)
);

AO21x1_ASAP7_75t_L g1125 ( 
.A1(n_913),
.A2(n_850),
.B(n_713),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_954),
.A2(n_713),
.B(n_708),
.Y(n_1126)
);

INVx4_ASAP7_75t_L g1127 ( 
.A(n_879),
.Y(n_1127)
);

O2A1O1Ixp5_ASAP7_75t_L g1128 ( 
.A1(n_913),
.A2(n_851),
.B(n_838),
.C(n_835),
.Y(n_1128)
);

OAI21xp33_ASAP7_75t_L g1129 ( 
.A1(n_974),
.A2(n_260),
.B(n_256),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_873),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_1005),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_937),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_971),
.B(n_835),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_959),
.B(n_835),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_873),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_960),
.A2(n_716),
.B(n_708),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_884),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_960),
.A2(n_717),
.B(n_716),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_959),
.B(n_838),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_970),
.A2(n_718),
.B(n_717),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_858),
.B(n_838),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_879),
.A2(n_440),
.B1(n_269),
.B2(n_271),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_887),
.Y(n_1143)
);

INVx4_ASAP7_75t_L g1144 ( 
.A(n_879),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_914),
.B(n_261),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_970),
.A2(n_720),
.B(n_718),
.Y(n_1146)
);

INVx4_ASAP7_75t_L g1147 ( 
.A(n_933),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_906),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_974),
.B(n_851),
.Y(n_1149)
);

BUFx2_ASAP7_75t_SL g1150 ( 
.A(n_927),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_906),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_999),
.A2(n_723),
.B(n_720),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_920),
.B(n_973),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_909),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_999),
.A2(n_723),
.B(n_745),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_868),
.B(n_745),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_998),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1002),
.A2(n_773),
.B(n_748),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_875),
.B(n_261),
.Y(n_1159)
);

AOI21xp33_ASAP7_75t_L g1160 ( 
.A1(n_938),
.A2(n_382),
.B(n_380),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_891),
.B(n_269),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1002),
.A2(n_748),
.B(n_745),
.Y(n_1162)
);

OR2x4_ASAP7_75t_L g1163 ( 
.A(n_1016),
.B(n_683),
.Y(n_1163)
);

NOR2x1_ASAP7_75t_L g1164 ( 
.A(n_896),
.B(n_683),
.Y(n_1164)
);

BUFx4f_ASAP7_75t_L g1165 ( 
.A(n_998),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_909),
.Y(n_1166)
);

INVx11_ASAP7_75t_L g1167 ( 
.A(n_981),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_865),
.A2(n_773),
.B(n_761),
.Y(n_1168)
);

INVx2_ASAP7_75t_SL g1169 ( 
.A(n_988),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_885),
.A2(n_409),
.B1(n_279),
.B2(n_284),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_872),
.A2(n_977),
.B(n_963),
.Y(n_1171)
);

AND2x2_ASAP7_75t_SL g1172 ( 
.A(n_947),
.B(n_688),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_871),
.B(n_877),
.Y(n_1173)
);

AOI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_903),
.A2(n_748),
.B1(n_801),
.B2(n_774),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_885),
.A2(n_688),
.B(n_649),
.C(n_774),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_903),
.B(n_271),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_945),
.B(n_761),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_892),
.B(n_945),
.Y(n_1178)
);

NOR2x1p5_ASAP7_75t_SL g1179 ( 
.A(n_907),
.B(n_614),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_921),
.B(n_761),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_978),
.A2(n_774),
.B(n_763),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_892),
.B(n_279),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_923),
.B(n_763),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1022),
.A2(n_658),
.B(n_656),
.C(n_682),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_923),
.B(n_801),
.Y(n_1185)
);

BUFx4f_ASAP7_75t_L g1186 ( 
.A(n_998),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_935),
.B(n_801),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1013),
.B(n_656),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_892),
.B(n_284),
.Y(n_1189)
);

AOI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1021),
.A2(n_632),
.B(n_623),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_935),
.B(n_956),
.Y(n_1191)
);

AOI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1021),
.A2(n_633),
.B(n_632),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_955),
.B(n_285),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_956),
.B(n_824),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_955),
.B(n_285),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1007),
.B(n_1023),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_967),
.B(n_764),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_1007),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1007),
.B(n_289),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1024),
.A2(n_658),
.B(n_682),
.C(n_675),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_967),
.Y(n_1201)
);

AO21x1_ASAP7_75t_L g1202 ( 
.A1(n_908),
.A2(n_651),
.B(n_647),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_968),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_984),
.A2(n_764),
.B(n_750),
.Y(n_1204)
);

OR2x2_ASAP7_75t_L g1205 ( 
.A(n_968),
.B(n_656),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_969),
.B(n_764),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_985),
.A2(n_764),
.B(n_750),
.Y(n_1207)
);

OAI21xp33_ASAP7_75t_L g1208 ( 
.A1(n_874),
.A2(n_264),
.B(n_263),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1023),
.B(n_658),
.Y(n_1209)
);

O2A1O1Ixp5_ASAP7_75t_L g1210 ( 
.A1(n_908),
.A2(n_910),
.B(n_969),
.C(n_1015),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_910),
.A2(n_750),
.B(n_737),
.Y(n_1211)
);

INVx1_ASAP7_75t_SL g1212 ( 
.A(n_1020),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_976),
.B(n_983),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_990),
.A2(n_764),
.B(n_750),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_976),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_992),
.A2(n_750),
.B(n_737),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1038),
.B(n_983),
.Y(n_1217)
);

AOI21xp33_ASAP7_75t_L g1218 ( 
.A1(n_1041),
.A2(n_1015),
.B(n_987),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_R g1219 ( 
.A(n_1132),
.B(n_1025),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1095),
.A2(n_1014),
.B1(n_986),
.B2(n_1003),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1028),
.B(n_987),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1042),
.A2(n_997),
.B1(n_1000),
.B2(n_944),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_R g1223 ( 
.A(n_1058),
.B(n_981),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1148),
.Y(n_1224)
);

O2A1O1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1160),
.A2(n_928),
.B(n_918),
.C(n_919),
.Y(n_1225)
);

O2A1O1Ixp5_ASAP7_75t_L g1226 ( 
.A1(n_1037),
.A2(n_946),
.B(n_939),
.C(n_942),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1096),
.B(n_948),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_1036),
.Y(n_1228)
);

INVx2_ASAP7_75t_SL g1229 ( 
.A(n_1076),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1198),
.B(n_933),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1046),
.B(n_1034),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1057),
.A2(n_1006),
.B(n_902),
.C(n_668),
.Y(n_1232)
);

CKINVDCx14_ASAP7_75t_R g1233 ( 
.A(n_1072),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1082),
.A2(n_1059),
.B1(n_1073),
.B2(n_1066),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1062),
.A2(n_933),
.B(n_892),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1148),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1040),
.B(n_981),
.Y(n_1237)
);

O2A1O1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1098),
.A2(n_1161),
.B(n_1159),
.C(n_1119),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1052),
.A2(n_933),
.B(n_994),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1166),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_1111),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1153),
.B(n_289),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1036),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1031),
.B(n_388),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1061),
.B(n_1087),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_1150),
.Y(n_1246)
);

AOI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1045),
.A2(n_1176),
.B1(n_1039),
.B2(n_1172),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1166),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1201),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1215),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_SL g1251 ( 
.A1(n_1121),
.A2(n_275),
.B1(n_263),
.B2(n_264),
.Y(n_1251)
);

INVx4_ASAP7_75t_L g1252 ( 
.A(n_1036),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1048),
.A2(n_981),
.B(n_633),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1091),
.B(n_981),
.Y(n_1254)
);

A2O1A1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1056),
.A2(n_424),
.B(n_409),
.C(n_415),
.Y(n_1255)
);

OAI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1122),
.A2(n_275),
.B1(n_268),
.B2(n_274),
.Y(n_1256)
);

NOR3xp33_ASAP7_75t_L g1257 ( 
.A(n_1145),
.B(n_1093),
.C(n_1193),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1064),
.A2(n_750),
.B(n_737),
.Y(n_1258)
);

O2A1O1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1109),
.A2(n_668),
.B(n_682),
.C(n_675),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1030),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1083),
.Y(n_1261)
);

O2A1O1Ixp5_ASAP7_75t_L g1262 ( 
.A1(n_1202),
.A2(n_651),
.B(n_647),
.C(n_653),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1114),
.B(n_665),
.Y(n_1263)
);

BUFx10_ASAP7_75t_L g1264 ( 
.A(n_1195),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1094),
.B(n_389),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1075),
.B(n_290),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1112),
.A2(n_424),
.B(n_290),
.C(n_415),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1089),
.B(n_665),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1210),
.A2(n_416),
.B(n_418),
.C(n_433),
.Y(n_1269)
);

AOI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1063),
.A2(n_348),
.B1(n_349),
.B2(n_351),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_SL g1271 ( 
.A(n_1075),
.B(n_416),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1090),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1134),
.A2(n_268),
.B1(n_274),
.B2(n_280),
.Y(n_1273)
);

OAI21xp33_ASAP7_75t_SL g1274 ( 
.A1(n_1178),
.A2(n_653),
.B(n_670),
.Y(n_1274)
);

AO21x1_ASAP7_75t_L g1275 ( 
.A1(n_1171),
.A2(n_668),
.B(n_670),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1205),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1080),
.B(n_670),
.Y(n_1277)
);

INVx1_ASAP7_75t_SL g1278 ( 
.A(n_1100),
.Y(n_1278)
);

NOR3xp33_ASAP7_75t_SL g1279 ( 
.A(n_1208),
.B(n_422),
.C(n_454),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1171),
.A2(n_791),
.B(n_787),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1104),
.B(n_395),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1048),
.A2(n_632),
.B(n_633),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1107),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_R g1284 ( 
.A(n_1065),
.B(n_418),
.Y(n_1284)
);

O2A1O1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1106),
.A2(n_675),
.B(n_649),
.C(n_635),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1067),
.A2(n_791),
.B(n_787),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1108),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1135),
.Y(n_1288)
);

O2A1O1Ixp5_ASAP7_75t_L g1289 ( 
.A1(n_1071),
.A2(n_649),
.B(n_603),
.C(n_635),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1075),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_SL g1291 ( 
.A(n_1131),
.B(n_433),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1139),
.A2(n_431),
.B1(n_412),
.B2(n_413),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1130),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1080),
.B(n_1113),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1077),
.B(n_375),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1188),
.B(n_398),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1151),
.Y(n_1297)
);

A2O1A1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1099),
.A2(n_439),
.B(n_440),
.C(n_441),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1213),
.B(n_649),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1070),
.A2(n_791),
.B(n_787),
.Y(n_1300)
);

INVxp67_ASAP7_75t_L g1301 ( 
.A(n_1169),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1131),
.B(n_439),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1105),
.B(n_399),
.Y(n_1303)
);

OR2x6_ASAP7_75t_L g1304 ( 
.A(n_1196),
.B(n_1131),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1137),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1054),
.A2(n_791),
.B(n_787),
.Y(n_1306)
);

BUFx6f_ASAP7_75t_L g1307 ( 
.A(n_1196),
.Y(n_1307)
);

O2A1O1Ixp33_ASAP7_75t_SL g1308 ( 
.A1(n_1047),
.A2(n_603),
.B(n_635),
.C(n_606),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1113),
.B(n_441),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1115),
.A2(n_429),
.B1(n_412),
.B2(n_422),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1102),
.B(n_443),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1053),
.B(n_443),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_1212),
.B(n_400),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_1157),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1203),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1053),
.B(n_444),
.Y(n_1316)
);

AOI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1032),
.A2(n_791),
.B(n_787),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1143),
.Y(n_1318)
);

INVxp67_ASAP7_75t_L g1319 ( 
.A(n_1199),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1129),
.B(n_405),
.Y(n_1320)
);

INVxp67_ASAP7_75t_L g1321 ( 
.A(n_1085),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1165),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1164),
.B(n_444),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1163),
.B(n_407),
.Y(n_1324)
);

NOR2xp67_ASAP7_75t_L g1325 ( 
.A(n_1142),
.B(n_352),
.Y(n_1325)
);

OA21x2_ASAP7_75t_L g1326 ( 
.A1(n_1060),
.A2(n_406),
.B(n_357),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1086),
.A2(n_791),
.B(n_787),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1165),
.Y(n_1328)
);

INVx4_ASAP7_75t_L g1329 ( 
.A(n_1035),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1103),
.A2(n_280),
.B1(n_425),
.B2(n_429),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1163),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1170),
.B(n_425),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_SL g1333 ( 
.A(n_1186),
.B(n_447),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1173),
.B(n_431),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1110),
.A2(n_451),
.B1(n_457),
.B2(n_450),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1209),
.B(n_447),
.Y(n_1336)
);

NAND3xp33_ASAP7_75t_SL g1337 ( 
.A(n_1055),
.B(n_454),
.C(n_450),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1088),
.A2(n_768),
.B(n_737),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1097),
.A2(n_768),
.B(n_737),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1154),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1209),
.B(n_459),
.Y(n_1341)
);

NOR2x1_ASAP7_75t_L g1342 ( 
.A(n_1035),
.B(n_603),
.Y(n_1342)
);

BUFx6f_ASAP7_75t_L g1343 ( 
.A(n_1186),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_1167),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_L g1345 ( 
.A(n_1149),
.B(n_459),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1079),
.B(n_463),
.Y(n_1346)
);

INVx2_ASAP7_75t_SL g1347 ( 
.A(n_1081),
.Y(n_1347)
);

OAI21xp33_ASAP7_75t_L g1348 ( 
.A1(n_1177),
.A2(n_465),
.B(n_464),
.Y(n_1348)
);

AOI222xp33_ASAP7_75t_L g1349 ( 
.A1(n_1141),
.A2(n_398),
.B1(n_465),
.B2(n_464),
.C1(n_463),
.C2(n_378),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1123),
.A2(n_393),
.B1(n_360),
.B2(n_367),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1120),
.A2(n_401),
.B1(n_368),
.B2(n_381),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1191),
.B(n_359),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1078),
.B(n_398),
.Y(n_1353)
);

OR2x6_ASAP7_75t_SL g1354 ( 
.A(n_1156),
.B(n_383),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1033),
.B(n_390),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1133),
.A2(n_768),
.B(n_737),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1175),
.B(n_13),
.Y(n_1357)
);

NAND2x1p5_ASAP7_75t_L g1358 ( 
.A(n_1127),
.B(n_768),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1027),
.A2(n_768),
.B(n_626),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_1182),
.Y(n_1360)
);

INVxp67_ASAP7_75t_L g1361 ( 
.A(n_1189),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1127),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_L g1363 ( 
.A(n_1144),
.B(n_13),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1027),
.A2(n_768),
.B(n_626),
.Y(n_1364)
);

OR2x6_ASAP7_75t_SL g1365 ( 
.A(n_1180),
.B(n_15),
.Y(n_1365)
);

BUFx6f_ASAP7_75t_L g1366 ( 
.A(n_1147),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1033),
.B(n_603),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1049),
.B(n_606),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1051),
.Y(n_1369)
);

OR2x6_ASAP7_75t_SL g1370 ( 
.A(n_1183),
.B(n_16),
.Y(n_1370)
);

O2A1O1Ixp33_ASAP7_75t_L g1371 ( 
.A1(n_1092),
.A2(n_635),
.B(n_606),
.C(n_20),
.Y(n_1371)
);

INVx8_ASAP7_75t_L g1372 ( 
.A(n_1147),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1049),
.A2(n_635),
.B(n_606),
.Y(n_1373)
);

O2A1O1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1069),
.A2(n_606),
.B(n_19),
.C(n_21),
.Y(n_1374)
);

INVx2_ASAP7_75t_SL g1375 ( 
.A(n_1144),
.Y(n_1375)
);

A2O1A1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1044),
.A2(n_626),
.B(n_21),
.C(n_22),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1174),
.B(n_227),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1185),
.Y(n_1378)
);

AOI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1190),
.A2(n_626),
.B(n_212),
.Y(n_1379)
);

AOI222xp33_ASAP7_75t_L g1380 ( 
.A1(n_1029),
.A2(n_18),
.B1(n_28),
.B2(n_29),
.C1(n_33),
.C2(n_34),
.Y(n_1380)
);

A2O1A1Ixp33_ASAP7_75t_L g1381 ( 
.A1(n_1044),
.A2(n_626),
.B(n_34),
.C(n_35),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1084),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1318),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1238),
.A2(n_1168),
.B(n_1101),
.Y(n_1384)
);

AOI221x1_ASAP7_75t_L g1385 ( 
.A1(n_1257),
.A2(n_1043),
.B1(n_1117),
.B2(n_1118),
.C(n_1050),
.Y(n_1385)
);

AOI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1221),
.A2(n_1117),
.B(n_1118),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1239),
.A2(n_1158),
.B(n_1194),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_1314),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1217),
.A2(n_1197),
.B(n_1206),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1220),
.A2(n_1204),
.B(n_1214),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1366),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1317),
.A2(n_1192),
.B(n_1068),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1226),
.A2(n_1043),
.B(n_1074),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1347),
.B(n_1187),
.Y(n_1394)
);

NAND3xp33_ASAP7_75t_SL g1395 ( 
.A(n_1244),
.B(n_1184),
.C(n_1200),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1332),
.A2(n_1125),
.B1(n_1181),
.B2(n_1124),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1234),
.A2(n_1214),
.B(n_1207),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1231),
.B(n_1152),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1280),
.A2(n_1379),
.B(n_1364),
.Y(n_1399)
);

OAI22x1_ASAP7_75t_L g1400 ( 
.A1(n_1247),
.A2(n_18),
.B1(n_35),
.B2(n_36),
.Y(n_1400)
);

A2O1A1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1320),
.A2(n_1377),
.B(n_1303),
.C(n_1234),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1382),
.A2(n_1377),
.B1(n_1231),
.B2(n_1245),
.Y(n_1402)
);

INVx4_ASAP7_75t_L g1403 ( 
.A(n_1372),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1227),
.B(n_1378),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1288),
.Y(n_1405)
);

O2A1O1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1267),
.A2(n_1128),
.B(n_1181),
.C(n_1116),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1268),
.B(n_1152),
.Y(n_1407)
);

NAND3xp33_ASAP7_75t_SL g1408 ( 
.A(n_1349),
.B(n_1124),
.C(n_1146),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1225),
.A2(n_1207),
.B(n_1204),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1235),
.A2(n_1162),
.B(n_1155),
.Y(n_1410)
);

BUFx2_ASAP7_75t_L g1411 ( 
.A(n_1287),
.Y(n_1411)
);

A2O1A1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1255),
.A2(n_1162),
.B(n_1155),
.C(n_1179),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1241),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1276),
.B(n_1146),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1304),
.B(n_1328),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1278),
.B(n_1140),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1359),
.A2(n_1140),
.B(n_1138),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1299),
.A2(n_1138),
.B(n_1136),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1282),
.A2(n_1126),
.B(n_1216),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1282),
.A2(n_1126),
.B(n_1216),
.Y(n_1420)
);

BUFx2_ASAP7_75t_R g1421 ( 
.A(n_1246),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1262),
.A2(n_1211),
.B(n_211),
.Y(n_1422)
);

AOI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1369),
.A2(n_626),
.B(n_209),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_1233),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1319),
.B(n_36),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1299),
.A2(n_626),
.B(n_201),
.Y(n_1426)
);

OAI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1222),
.A2(n_1232),
.B(n_1269),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1286),
.A2(n_196),
.B(n_195),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_1328),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1355),
.A2(n_189),
.B(n_178),
.Y(n_1430)
);

AO31x2_ASAP7_75t_L g1431 ( 
.A1(n_1275),
.A2(n_38),
.A3(n_39),
.B(n_41),
.Y(n_1431)
);

AOI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1380),
.A2(n_42),
.B1(n_46),
.B2(n_48),
.Y(n_1432)
);

INVxp67_ASAP7_75t_L g1433 ( 
.A(n_1331),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1300),
.A2(n_177),
.B(n_164),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_1229),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1356),
.A2(n_1373),
.B(n_1339),
.Y(n_1436)
);

AO21x1_ASAP7_75t_L g1437 ( 
.A1(n_1374),
.A2(n_48),
.B(n_50),
.Y(n_1437)
);

OAI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1294),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1301),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1328),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1305),
.Y(n_1441)
);

OAI22x1_ASAP7_75t_L g1442 ( 
.A1(n_1242),
.A2(n_54),
.B1(n_58),
.B2(n_59),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1340),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1249),
.B(n_58),
.Y(n_1444)
);

AOI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1380),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_1445)
);

OAI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1222),
.A2(n_102),
.B(n_159),
.Y(n_1446)
);

A2O1A1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1295),
.A2(n_62),
.B(n_63),
.C(n_65),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_SL g1448 ( 
.A(n_1264),
.B(n_62),
.Y(n_1448)
);

CKINVDCx11_ASAP7_75t_R g1449 ( 
.A(n_1264),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1373),
.A2(n_111),
.B(n_157),
.Y(n_1450)
);

NAND3xp33_ASAP7_75t_L g1451 ( 
.A(n_1349),
.B(n_63),
.C(n_67),
.Y(n_1451)
);

BUFx10_ASAP7_75t_L g1452 ( 
.A(n_1324),
.Y(n_1452)
);

INVx3_ASAP7_75t_SL g1453 ( 
.A(n_1322),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1334),
.B(n_68),
.Y(n_1454)
);

BUFx6f_ASAP7_75t_L g1455 ( 
.A(n_1343),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1260),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1261),
.Y(n_1457)
);

A2O1A1Ixp33_ASAP7_75t_L g1458 ( 
.A1(n_1279),
.A2(n_69),
.B(n_71),
.C(n_73),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1272),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1277),
.B(n_74),
.Y(n_1460)
);

BUFx10_ASAP7_75t_L g1461 ( 
.A(n_1265),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1304),
.B(n_1343),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1343),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1368),
.A2(n_123),
.B(n_154),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1338),
.A2(n_118),
.B(n_151),
.Y(n_1465)
);

OAI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1253),
.A2(n_160),
.B(n_115),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1283),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1293),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1367),
.A2(n_101),
.B(n_143),
.Y(n_1469)
);

AOI31xp67_ASAP7_75t_L g1470 ( 
.A1(n_1237),
.A2(n_146),
.A3(n_139),
.B(n_132),
.Y(n_1470)
);

INVx2_ASAP7_75t_SL g1471 ( 
.A(n_1228),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1357),
.B(n_80),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1251),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1296),
.B(n_1353),
.Y(n_1474)
);

OAI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1253),
.A2(n_126),
.B(n_83),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1327),
.A2(n_84),
.B(n_1258),
.Y(n_1476)
);

AO31x2_ASAP7_75t_L g1477 ( 
.A1(n_1376),
.A2(n_1381),
.A3(n_1298),
.B(n_1310),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1297),
.B(n_1315),
.Y(n_1478)
);

NAND2x1p5_ASAP7_75t_L g1479 ( 
.A(n_1362),
.B(n_1329),
.Y(n_1479)
);

OA21x2_ASAP7_75t_L g1480 ( 
.A1(n_1289),
.A2(n_1218),
.B(n_1351),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1224),
.B(n_1236),
.Y(n_1481)
);

INVxp67_ASAP7_75t_SL g1482 ( 
.A(n_1250),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1218),
.A2(n_1254),
.B(n_1306),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1313),
.B(n_1281),
.Y(n_1484)
);

INVx2_ASAP7_75t_SL g1485 ( 
.A(n_1228),
.Y(n_1485)
);

A2O1A1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1371),
.A2(n_1361),
.B(n_1345),
.C(n_1348),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1263),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1309),
.B(n_1360),
.Y(n_1488)
);

NOR2xp67_ASAP7_75t_L g1489 ( 
.A(n_1321),
.B(n_1344),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1352),
.A2(n_1308),
.B(n_1326),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1365),
.B(n_1370),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1285),
.A2(n_1342),
.B(n_1259),
.Y(n_1492)
);

AOI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1326),
.A2(n_1346),
.B(n_1311),
.Y(n_1493)
);

INVx2_ASAP7_75t_SL g1494 ( 
.A(n_1228),
.Y(n_1494)
);

INVx3_ASAP7_75t_L g1495 ( 
.A(n_1366),
.Y(n_1495)
);

AO31x2_ASAP7_75t_L g1496 ( 
.A1(n_1310),
.A2(n_1350),
.A3(n_1363),
.B(n_1330),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1240),
.Y(n_1497)
);

AO31x2_ASAP7_75t_L g1498 ( 
.A1(n_1350),
.A2(n_1335),
.A3(n_1330),
.B(n_1273),
.Y(n_1498)
);

O2A1O1Ixp33_ASAP7_75t_SL g1499 ( 
.A1(n_1333),
.A2(n_1337),
.B(n_1271),
.C(n_1291),
.Y(n_1499)
);

OAI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1274),
.A2(n_1323),
.B(n_1325),
.Y(n_1500)
);

AOI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1335),
.A2(n_1292),
.B1(n_1273),
.B2(n_1256),
.Y(n_1501)
);

AO31x2_ASAP7_75t_L g1502 ( 
.A1(n_1292),
.A2(n_1248),
.A3(n_1316),
.B(n_1312),
.Y(n_1502)
);

AOI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1362),
.A2(n_1341),
.B(n_1336),
.Y(n_1503)
);

OAI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1304),
.A2(n_1307),
.B1(n_1354),
.B2(n_1230),
.Y(n_1504)
);

NOR2xp67_ASAP7_75t_L g1505 ( 
.A(n_1252),
.B(n_1270),
.Y(n_1505)
);

AO31x2_ASAP7_75t_L g1506 ( 
.A1(n_1252),
.A2(n_1329),
.A3(n_1223),
.B(n_1358),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1358),
.A2(n_1266),
.B(n_1302),
.Y(n_1507)
);

INVx3_ASAP7_75t_SL g1508 ( 
.A(n_1307),
.Y(n_1508)
);

BUFx2_ASAP7_75t_R g1509 ( 
.A(n_1219),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_SL g1510 ( 
.A(n_1307),
.B(n_1284),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1230),
.B(n_1243),
.Y(n_1511)
);

OAI21x1_ASAP7_75t_L g1512 ( 
.A1(n_1372),
.A2(n_1375),
.B(n_1366),
.Y(n_1512)
);

OAI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1372),
.A2(n_1243),
.B(n_1290),
.Y(n_1513)
);

A2O1A1Ixp33_ASAP7_75t_L g1514 ( 
.A1(n_1290),
.A2(n_915),
.B(n_1238),
.C(n_930),
.Y(n_1514)
);

A2O1A1Ixp33_ASAP7_75t_L g1515 ( 
.A1(n_1290),
.A2(n_915),
.B(n_1238),
.C(n_930),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1318),
.Y(n_1516)
);

OAI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1226),
.A2(n_915),
.B(n_1038),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1245),
.Y(n_1518)
);

INVx4_ASAP7_75t_L g1519 ( 
.A(n_1372),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1347),
.B(n_1038),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1347),
.B(n_1038),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1347),
.B(n_1038),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_1366),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1245),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1328),
.Y(n_1525)
);

AOI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1238),
.A2(n_1026),
.B(n_1018),
.Y(n_1526)
);

NAND2xp33_ASAP7_75t_SL g1527 ( 
.A(n_1219),
.B(n_1328),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1238),
.A2(n_1026),
.B(n_1018),
.Y(n_1528)
);

OR2x6_ASAP7_75t_L g1529 ( 
.A(n_1304),
.B(n_1372),
.Y(n_1529)
);

BUFx6f_ASAP7_75t_L g1530 ( 
.A(n_1328),
.Y(n_1530)
);

INVx5_ASAP7_75t_L g1531 ( 
.A(n_1372),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1245),
.Y(n_1532)
);

OAI21x1_ASAP7_75t_L g1533 ( 
.A1(n_1239),
.A2(n_1317),
.B(n_1280),
.Y(n_1533)
);

BUFx10_ASAP7_75t_L g1534 ( 
.A(n_1324),
.Y(n_1534)
);

AOI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1238),
.A2(n_1026),
.B(n_1018),
.Y(n_1535)
);

INVxp67_ASAP7_75t_L g1536 ( 
.A(n_1331),
.Y(n_1536)
);

NOR2xp67_ASAP7_75t_L g1537 ( 
.A(n_1301),
.B(n_1058),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1245),
.Y(n_1538)
);

OAI21x1_ASAP7_75t_SL g1539 ( 
.A1(n_1231),
.A2(n_1037),
.B(n_1238),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1245),
.Y(n_1540)
);

BUFx2_ASAP7_75t_R g1541 ( 
.A(n_1246),
.Y(n_1541)
);

OAI21x1_ASAP7_75t_L g1542 ( 
.A1(n_1239),
.A2(n_1317),
.B(n_1280),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_1229),
.Y(n_1543)
);

NOR2xp67_ASAP7_75t_L g1544 ( 
.A(n_1301),
.B(n_1058),
.Y(n_1544)
);

A2O1A1Ixp33_ASAP7_75t_L g1545 ( 
.A1(n_1238),
.A2(n_915),
.B(n_930),
.C(n_925),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_SL g1546 ( 
.A(n_1278),
.B(n_937),
.Y(n_1546)
);

OAI21x1_ASAP7_75t_L g1547 ( 
.A1(n_1239),
.A2(n_1317),
.B(n_1280),
.Y(n_1547)
);

AOI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1221),
.A2(n_1379),
.B(n_913),
.Y(n_1548)
);

AO21x1_ASAP7_75t_L g1549 ( 
.A1(n_1238),
.A2(n_915),
.B(n_1234),
.Y(n_1549)
);

OAI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1226),
.A2(n_915),
.B(n_1038),
.Y(n_1550)
);

AO31x2_ASAP7_75t_L g1551 ( 
.A1(n_1275),
.A2(n_1269),
.A3(n_1369),
.B(n_1202),
.Y(n_1551)
);

BUFx3_ASAP7_75t_L g1552 ( 
.A(n_1229),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1382),
.A2(n_915),
.B1(n_1038),
.B2(n_971),
.Y(n_1553)
);

OAI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1226),
.A2(n_915),
.B(n_1038),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1278),
.B(n_869),
.Y(n_1555)
);

OAI21x1_ASAP7_75t_L g1556 ( 
.A1(n_1239),
.A2(n_1317),
.B(n_1280),
.Y(n_1556)
);

AOI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1238),
.A2(n_1026),
.B(n_1018),
.Y(n_1557)
);

OAI22x1_ASAP7_75t_L g1558 ( 
.A1(n_1247),
.A2(n_866),
.B1(n_1042),
.B2(n_930),
.Y(n_1558)
);

O2A1O1Ixp33_ASAP7_75t_SL g1559 ( 
.A1(n_1238),
.A2(n_915),
.B(n_1298),
.C(n_1255),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_SL g1560 ( 
.A1(n_1238),
.A2(n_879),
.B(n_705),
.Y(n_1560)
);

OAI21x1_ASAP7_75t_L g1561 ( 
.A1(n_1239),
.A2(n_1317),
.B(n_1280),
.Y(n_1561)
);

AOI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1238),
.A2(n_1026),
.B(n_1018),
.Y(n_1562)
);

CKINVDCx6p67_ASAP7_75t_R g1563 ( 
.A(n_1453),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1383),
.Y(n_1564)
);

AOI21xp5_ASAP7_75t_SL g1565 ( 
.A1(n_1401),
.A2(n_1545),
.B(n_1475),
.Y(n_1565)
);

INVx1_ASAP7_75t_SL g1566 ( 
.A(n_1439),
.Y(n_1566)
);

BUFx8_ASAP7_75t_L g1567 ( 
.A(n_1429),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1484),
.B(n_1404),
.Y(n_1568)
);

CKINVDCx20_ASAP7_75t_R g1569 ( 
.A(n_1413),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_1543),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1451),
.A2(n_1445),
.B1(n_1432),
.B2(n_1558),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1552),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1449),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1411),
.Y(n_1574)
);

BUFx3_ASAP7_75t_L g1575 ( 
.A(n_1435),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1516),
.Y(n_1576)
);

INVx2_ASAP7_75t_SL g1577 ( 
.A(n_1429),
.Y(n_1577)
);

CKINVDCx20_ASAP7_75t_R g1578 ( 
.A(n_1424),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1451),
.A2(n_1432),
.B1(n_1445),
.B2(n_1501),
.Y(n_1579)
);

BUFx12f_ASAP7_75t_L g1580 ( 
.A(n_1452),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1553),
.A2(n_1402),
.B1(n_1501),
.B2(n_1404),
.Y(n_1581)
);

INVx6_ASAP7_75t_L g1582 ( 
.A(n_1531),
.Y(n_1582)
);

INVx6_ASAP7_75t_L g1583 ( 
.A(n_1531),
.Y(n_1583)
);

INVx8_ASAP7_75t_L g1584 ( 
.A(n_1531),
.Y(n_1584)
);

OAI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1454),
.A2(n_1553),
.B1(n_1475),
.B2(n_1472),
.Y(n_1585)
);

BUFx12f_ASAP7_75t_L g1586 ( 
.A(n_1452),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1456),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1549),
.A2(n_1400),
.B1(n_1473),
.B2(n_1402),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1441),
.Y(n_1589)
);

CKINVDCx11_ASAP7_75t_R g1590 ( 
.A(n_1534),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1457),
.Y(n_1591)
);

CKINVDCx20_ASAP7_75t_R g1592 ( 
.A(n_1527),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1467),
.Y(n_1593)
);

BUFx2_ASAP7_75t_SL g1594 ( 
.A(n_1537),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_L g1595 ( 
.A1(n_1446),
.A2(n_1437),
.B1(n_1472),
.B2(n_1438),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_SL g1596 ( 
.A1(n_1491),
.A2(n_1446),
.B1(n_1466),
.B2(n_1425),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1518),
.B(n_1524),
.Y(n_1597)
);

INVx4_ASAP7_75t_SL g1598 ( 
.A(n_1529),
.Y(n_1598)
);

BUFx12f_ASAP7_75t_L g1599 ( 
.A(n_1534),
.Y(n_1599)
);

INVx6_ASAP7_75t_L g1600 ( 
.A(n_1403),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1443),
.Y(n_1601)
);

CKINVDCx11_ASAP7_75t_R g1602 ( 
.A(n_1461),
.Y(n_1602)
);

BUFx3_ASAP7_75t_L g1603 ( 
.A(n_1388),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1474),
.A2(n_1546),
.B1(n_1466),
.B2(n_1408),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1520),
.B(n_1521),
.Y(n_1605)
);

INVx6_ASAP7_75t_L g1606 ( 
.A(n_1519),
.Y(n_1606)
);

AOI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1488),
.A2(n_1504),
.B1(n_1461),
.B2(n_1510),
.Y(n_1607)
);

BUFx5_ASAP7_75t_L g1608 ( 
.A(n_1487),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1459),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1468),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1497),
.Y(n_1611)
);

OAI21xp5_ASAP7_75t_SL g1612 ( 
.A1(n_1447),
.A2(n_1458),
.B(n_1448),
.Y(n_1612)
);

INVx1_ASAP7_75t_SL g1613 ( 
.A(n_1509),
.Y(n_1613)
);

BUFx12f_ASAP7_75t_L g1614 ( 
.A(n_1429),
.Y(n_1614)
);

CKINVDCx20_ASAP7_75t_R g1615 ( 
.A(n_1508),
.Y(n_1615)
);

INVx2_ASAP7_75t_SL g1616 ( 
.A(n_1440),
.Y(n_1616)
);

OAI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1522),
.A2(n_1532),
.B1(n_1538),
.B2(n_1540),
.Y(n_1617)
);

BUFx3_ASAP7_75t_L g1618 ( 
.A(n_1440),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1394),
.B(n_1514),
.Y(n_1619)
);

OAI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1442),
.A2(n_1416),
.B1(n_1444),
.B2(n_1460),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1478),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_SL g1622 ( 
.A1(n_1427),
.A2(n_1422),
.B1(n_1539),
.B2(n_1482),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_SL g1623 ( 
.A1(n_1427),
.A2(n_1422),
.B1(n_1554),
.B2(n_1550),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1481),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1515),
.A2(n_1486),
.B1(n_1536),
.B2(n_1433),
.Y(n_1625)
);

BUFx2_ASAP7_75t_SL g1626 ( 
.A(n_1544),
.Y(n_1626)
);

OAI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1460),
.A2(n_1517),
.B1(n_1554),
.B2(n_1550),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1517),
.A2(n_1395),
.B1(n_1414),
.B2(n_1398),
.Y(n_1628)
);

INVx6_ASAP7_75t_L g1629 ( 
.A(n_1519),
.Y(n_1629)
);

BUFx3_ASAP7_75t_L g1630 ( 
.A(n_1455),
.Y(n_1630)
);

OAI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1493),
.A2(n_1503),
.B(n_1500),
.Y(n_1631)
);

CKINVDCx8_ASAP7_75t_R g1632 ( 
.A(n_1455),
.Y(n_1632)
);

CKINVDCx11_ASAP7_75t_R g1633 ( 
.A(n_1463),
.Y(n_1633)
);

CKINVDCx6p67_ASAP7_75t_R g1634 ( 
.A(n_1463),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_SL g1635 ( 
.A1(n_1504),
.A2(n_1498),
.B1(n_1500),
.B2(n_1415),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1398),
.A2(n_1384),
.B1(n_1505),
.B2(n_1430),
.Y(n_1636)
);

INVx1_ASAP7_75t_SL g1637 ( 
.A(n_1421),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1407),
.A2(n_1480),
.B1(n_1462),
.B2(n_1415),
.Y(n_1638)
);

INVx4_ASAP7_75t_L g1639 ( 
.A(n_1463),
.Y(n_1639)
);

AOI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1499),
.A2(n_1489),
.B1(n_1462),
.B2(n_1559),
.Y(n_1640)
);

OAI21xp33_ASAP7_75t_SL g1641 ( 
.A1(n_1560),
.A2(n_1507),
.B(n_1450),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_1511),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_SL g1643 ( 
.A1(n_1498),
.A2(n_1496),
.B1(n_1480),
.B2(n_1525),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_SL g1644 ( 
.A1(n_1496),
.A2(n_1525),
.B1(n_1530),
.B2(n_1469),
.Y(n_1644)
);

CKINVDCx11_ASAP7_75t_R g1645 ( 
.A(n_1530),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1431),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1407),
.A2(n_1464),
.B1(n_1396),
.B2(n_1529),
.Y(n_1647)
);

BUFx3_ASAP7_75t_L g1648 ( 
.A(n_1530),
.Y(n_1648)
);

CKINVDCx6p67_ASAP7_75t_R g1649 ( 
.A(n_1529),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1397),
.A2(n_1426),
.B1(n_1393),
.B2(n_1389),
.Y(n_1650)
);

INVx2_ASAP7_75t_SL g1651 ( 
.A(n_1471),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_SL g1652 ( 
.A1(n_1485),
.A2(n_1494),
.B1(n_1479),
.B2(n_1541),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1431),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1479),
.A2(n_1562),
.B1(n_1528),
.B2(n_1557),
.Y(n_1654)
);

BUFx3_ASAP7_75t_L g1655 ( 
.A(n_1391),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1495),
.B(n_1523),
.Y(n_1656)
);

INVx3_ASAP7_75t_SL g1657 ( 
.A(n_1495),
.Y(n_1657)
);

OAI21xp5_ASAP7_75t_SL g1658 ( 
.A1(n_1385),
.A2(n_1490),
.B(n_1406),
.Y(n_1658)
);

INVx2_ASAP7_75t_R g1659 ( 
.A(n_1470),
.Y(n_1659)
);

BUFx2_ASAP7_75t_L g1660 ( 
.A(n_1523),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1502),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1393),
.A2(n_1483),
.B1(n_1535),
.B2(n_1526),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1390),
.A2(n_1409),
.B1(n_1387),
.B2(n_1418),
.Y(n_1663)
);

OAI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1386),
.A2(n_1423),
.B1(n_1548),
.B2(n_1477),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1431),
.Y(n_1665)
);

OAI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1412),
.A2(n_1410),
.B(n_1436),
.Y(n_1666)
);

BUFx3_ASAP7_75t_L g1667 ( 
.A(n_1513),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1502),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_SL g1669 ( 
.A1(n_1477),
.A2(n_1428),
.B1(n_1434),
.B2(n_1465),
.Y(n_1669)
);

INVx4_ASAP7_75t_L g1670 ( 
.A(n_1506),
.Y(n_1670)
);

OAI21xp5_ASAP7_75t_SL g1671 ( 
.A1(n_1477),
.A2(n_1502),
.B(n_1551),
.Y(n_1671)
);

OAI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1551),
.A2(n_1506),
.B1(n_1512),
.B2(n_1492),
.Y(n_1672)
);

OAI22x1_ASAP7_75t_L g1673 ( 
.A1(n_1551),
.A2(n_1476),
.B1(n_1506),
.B2(n_1419),
.Y(n_1673)
);

BUFx3_ASAP7_75t_L g1674 ( 
.A(n_1420),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1417),
.Y(n_1675)
);

BUFx4f_ASAP7_75t_SL g1676 ( 
.A(n_1399),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_1533),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1542),
.A2(n_1547),
.B1(n_1556),
.B2(n_1561),
.Y(n_1678)
);

CKINVDCx20_ASAP7_75t_R g1679 ( 
.A(n_1392),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1405),
.Y(n_1680)
);

INVx3_ASAP7_75t_L g1681 ( 
.A(n_1403),
.Y(n_1681)
);

CKINVDCx20_ASAP7_75t_R g1682 ( 
.A(n_1413),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1451),
.A2(n_1445),
.B1(n_1432),
.B2(n_1380),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1405),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1555),
.B(n_1474),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1451),
.A2(n_1445),
.B1(n_1432),
.B2(n_1380),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1405),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1484),
.A2(n_1451),
.B1(n_1244),
.B2(n_1257),
.Y(n_1688)
);

BUFx2_ASAP7_75t_SL g1689 ( 
.A(n_1537),
.Y(n_1689)
);

INVx2_ASAP7_75t_SL g1690 ( 
.A(n_1543),
.Y(n_1690)
);

CKINVDCx20_ASAP7_75t_R g1691 ( 
.A(n_1413),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1405),
.Y(n_1692)
);

INVx4_ASAP7_75t_L g1693 ( 
.A(n_1531),
.Y(n_1693)
);

OAI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1484),
.A2(n_915),
.B1(n_932),
.B2(n_1257),
.C(n_1244),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1555),
.B(n_1474),
.Y(n_1695)
);

BUFx4_ASAP7_75t_R g1696 ( 
.A(n_1461),
.Y(n_1696)
);

BUFx12f_ASAP7_75t_L g1697 ( 
.A(n_1413),
.Y(n_1697)
);

NAND2x1p5_ASAP7_75t_L g1698 ( 
.A(n_1531),
.B(n_1403),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1451),
.A2(n_1445),
.B1(n_1432),
.B2(n_1380),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1451),
.A2(n_1445),
.B1(n_1432),
.B2(n_1380),
.Y(n_1700)
);

BUFx2_ASAP7_75t_L g1701 ( 
.A(n_1543),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1555),
.B(n_1474),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1484),
.A2(n_915),
.B1(n_1401),
.B2(n_932),
.Y(n_1703)
);

CKINVDCx11_ASAP7_75t_R g1704 ( 
.A(n_1453),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1484),
.A2(n_915),
.B1(n_1401),
.B2(n_932),
.Y(n_1705)
);

BUFx4f_ASAP7_75t_L g1706 ( 
.A(n_1429),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1451),
.A2(n_1445),
.B1(n_1432),
.B2(n_1380),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_SL g1708 ( 
.A1(n_1451),
.A2(n_915),
.B1(n_1484),
.B2(n_930),
.Y(n_1708)
);

BUFx3_ASAP7_75t_L g1709 ( 
.A(n_1543),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1383),
.Y(n_1710)
);

BUFx3_ASAP7_75t_L g1711 ( 
.A(n_1543),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1484),
.B(n_1038),
.Y(n_1712)
);

INVx3_ASAP7_75t_L g1713 ( 
.A(n_1403),
.Y(n_1713)
);

INVx5_ASAP7_75t_L g1714 ( 
.A(n_1529),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1415),
.B(n_1462),
.Y(n_1715)
);

INVx1_ASAP7_75t_SL g1716 ( 
.A(n_1439),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1383),
.Y(n_1717)
);

CKINVDCx11_ASAP7_75t_R g1718 ( 
.A(n_1453),
.Y(n_1718)
);

AOI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1451),
.A2(n_1445),
.B1(n_1432),
.B2(n_1380),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1484),
.B(n_1038),
.Y(n_1720)
);

OAI21xp33_ASAP7_75t_L g1721 ( 
.A1(n_1484),
.A2(n_915),
.B(n_925),
.Y(n_1721)
);

BUFx3_ASAP7_75t_L g1722 ( 
.A(n_1543),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1402),
.Y(n_1723)
);

INVx3_ASAP7_75t_SL g1724 ( 
.A(n_1413),
.Y(n_1724)
);

INVx5_ASAP7_75t_L g1725 ( 
.A(n_1529),
.Y(n_1725)
);

AOI22xp33_ASAP7_75t_L g1726 ( 
.A1(n_1451),
.A2(n_1445),
.B1(n_1432),
.B2(n_1380),
.Y(n_1726)
);

NAND2x1p5_ASAP7_75t_L g1727 ( 
.A(n_1531),
.B(n_1403),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_1413),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_L g1729 ( 
.A1(n_1451),
.A2(n_1445),
.B1(n_1432),
.B2(n_1380),
.Y(n_1729)
);

BUFx6f_ASAP7_75t_L g1730 ( 
.A(n_1429),
.Y(n_1730)
);

INVx4_ASAP7_75t_SL g1731 ( 
.A(n_1529),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_1413),
.Y(n_1732)
);

AOI22xp33_ASAP7_75t_L g1733 ( 
.A1(n_1451),
.A2(n_1445),
.B1(n_1432),
.B2(n_1380),
.Y(n_1733)
);

OAI22xp5_ASAP7_75t_L g1734 ( 
.A1(n_1484),
.A2(n_915),
.B1(n_1401),
.B2(n_932),
.Y(n_1734)
);

AOI22xp33_ASAP7_75t_SL g1735 ( 
.A1(n_1451),
.A2(n_915),
.B1(n_1484),
.B2(n_930),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_1413),
.Y(n_1736)
);

INVx6_ASAP7_75t_L g1737 ( 
.A(n_1531),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1451),
.A2(n_1445),
.B1(n_1432),
.B2(n_1380),
.Y(n_1738)
);

BUFx10_ASAP7_75t_L g1739 ( 
.A(n_1413),
.Y(n_1739)
);

AOI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1451),
.A2(n_1445),
.B1(n_1432),
.B2(n_1380),
.Y(n_1740)
);

BUFx12f_ASAP7_75t_L g1741 ( 
.A(n_1413),
.Y(n_1741)
);

INVx5_ASAP7_75t_L g1742 ( 
.A(n_1529),
.Y(n_1742)
);

OAI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1484),
.A2(n_915),
.B1(n_1401),
.B2(n_932),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_1413),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1405),
.Y(n_1745)
);

AOI22xp33_ASAP7_75t_SL g1746 ( 
.A1(n_1451),
.A2(n_915),
.B1(n_1484),
.B2(n_930),
.Y(n_1746)
);

INVx4_ASAP7_75t_SL g1747 ( 
.A(n_1529),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_SL g1748 ( 
.A1(n_1451),
.A2(n_915),
.B1(n_1484),
.B2(n_930),
.Y(n_1748)
);

AOI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1451),
.A2(n_1445),
.B1(n_1432),
.B2(n_1380),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1608),
.Y(n_1750)
);

NAND3xp33_ASAP7_75t_L g1751 ( 
.A(n_1688),
.B(n_1705),
.C(n_1703),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_L g1752 ( 
.A1(n_1683),
.A2(n_1699),
.B1(n_1700),
.B2(n_1686),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1668),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1646),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1608),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1653),
.Y(n_1756)
);

OA21x2_ASAP7_75t_L g1757 ( 
.A1(n_1658),
.A2(n_1631),
.B(n_1671),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1608),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1608),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1723),
.B(n_1643),
.Y(n_1760)
);

OAI21x1_ASAP7_75t_L g1761 ( 
.A1(n_1666),
.A2(n_1678),
.B(n_1654),
.Y(n_1761)
);

AOI21x1_ASAP7_75t_L g1762 ( 
.A1(n_1673),
.A2(n_1675),
.B(n_1665),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1642),
.Y(n_1763)
);

HB1xp67_ASAP7_75t_L g1764 ( 
.A(n_1625),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1598),
.B(n_1731),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1643),
.B(n_1635),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1661),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1683),
.A2(n_1749),
.B1(n_1686),
.B2(n_1699),
.Y(n_1768)
);

INVx3_ASAP7_75t_L g1769 ( 
.A(n_1670),
.Y(n_1769)
);

OAI21x1_ASAP7_75t_L g1770 ( 
.A1(n_1678),
.A2(n_1663),
.B(n_1662),
.Y(n_1770)
);

OAI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1694),
.A2(n_1743),
.B(n_1734),
.Y(n_1771)
);

INVx3_ASAP7_75t_L g1772 ( 
.A(n_1674),
.Y(n_1772)
);

NOR2x1_ASAP7_75t_L g1773 ( 
.A(n_1617),
.B(n_1693),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1568),
.B(n_1712),
.Y(n_1774)
);

INVxp33_ASAP7_75t_L g1775 ( 
.A(n_1685),
.Y(n_1775)
);

AOI21x1_ASAP7_75t_L g1776 ( 
.A1(n_1581),
.A2(n_1619),
.B(n_1601),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1589),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1720),
.B(n_1605),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1680),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1684),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1687),
.Y(n_1781)
);

HB1xp67_ASAP7_75t_L g1782 ( 
.A(n_1692),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1597),
.B(n_1721),
.Y(n_1783)
);

INVx1_ASAP7_75t_SL g1784 ( 
.A(n_1566),
.Y(n_1784)
);

OAI21x1_ASAP7_75t_L g1785 ( 
.A1(n_1663),
.A2(n_1662),
.B(n_1650),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1574),
.B(n_1695),
.Y(n_1786)
);

AO31x2_ASAP7_75t_L g1787 ( 
.A1(n_1623),
.A2(n_1565),
.A3(n_1659),
.B(n_1664),
.Y(n_1787)
);

INVx2_ASAP7_75t_SL g1788 ( 
.A(n_1714),
.Y(n_1788)
);

HB1xp67_ASAP7_75t_L g1789 ( 
.A(n_1745),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1672),
.Y(n_1790)
);

INVx3_ASAP7_75t_L g1791 ( 
.A(n_1667),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1672),
.Y(n_1792)
);

BUFx6f_ASAP7_75t_L g1793 ( 
.A(n_1714),
.Y(n_1793)
);

NOR2xp33_ASAP7_75t_L g1794 ( 
.A(n_1702),
.B(n_1716),
.Y(n_1794)
);

OA21x2_ASAP7_75t_L g1795 ( 
.A1(n_1650),
.A2(n_1628),
.B(n_1638),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1635),
.B(n_1623),
.Y(n_1796)
);

OAI21x1_ASAP7_75t_L g1797 ( 
.A1(n_1636),
.A2(n_1647),
.B(n_1604),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1610),
.Y(n_1798)
);

INVx2_ASAP7_75t_SL g1799 ( 
.A(n_1714),
.Y(n_1799)
);

INVx3_ASAP7_75t_L g1800 ( 
.A(n_1676),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1708),
.B(n_1735),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1624),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1660),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1622),
.B(n_1609),
.Y(n_1804)
);

BUFx3_ASAP7_75t_L g1805 ( 
.A(n_1567),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1677),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1621),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1596),
.B(n_1564),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1708),
.B(n_1735),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1664),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1596),
.B(n_1576),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1627),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1710),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1587),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1717),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1591),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1593),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1611),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1620),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1676),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1679),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1714),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1585),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1725),
.Y(n_1824)
);

OAI21x1_ASAP7_75t_L g1825 ( 
.A1(n_1636),
.A2(n_1647),
.B(n_1640),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1725),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1725),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_SL g1828 ( 
.A1(n_1700),
.A2(n_1749),
.B1(n_1738),
.B2(n_1707),
.Y(n_1828)
);

AOI21x1_ASAP7_75t_L g1829 ( 
.A1(n_1659),
.A2(n_1656),
.B(n_1715),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1585),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1571),
.B(n_1579),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1644),
.Y(n_1832)
);

BUFx6f_ASAP7_75t_L g1833 ( 
.A(n_1742),
.Y(n_1833)
);

AOI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1707),
.A2(n_1726),
.B(n_1719),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1644),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1620),
.B(n_1571),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_L g1837 ( 
.A(n_1613),
.B(n_1607),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1641),
.Y(n_1838)
);

CKINVDCx5p33_ASAP7_75t_R g1839 ( 
.A(n_1704),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1579),
.B(n_1588),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1746),
.B(n_1748),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1747),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1669),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1669),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1649),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1746),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1748),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1588),
.B(n_1595),
.Y(n_1848)
);

OAI31xp33_ASAP7_75t_L g1849 ( 
.A1(n_1719),
.A2(n_1738),
.A3(n_1733),
.B(n_1729),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1612),
.B(n_1726),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1595),
.Y(n_1851)
);

INVx2_ASAP7_75t_SL g1852 ( 
.A(n_1582),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1729),
.A2(n_1733),
.B1(n_1740),
.B2(n_1603),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1582),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1656),
.Y(n_1855)
);

HB1xp67_ASAP7_75t_L g1856 ( 
.A(n_1575),
.Y(n_1856)
);

HB1xp67_ASAP7_75t_L g1857 ( 
.A(n_1655),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1583),
.Y(n_1858)
);

OAI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1740),
.A2(n_1592),
.B1(n_1652),
.B2(n_1689),
.Y(n_1859)
);

BUFx2_ASAP7_75t_L g1860 ( 
.A(n_1570),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1737),
.Y(n_1861)
);

OA21x2_ASAP7_75t_L g1862 ( 
.A1(n_1715),
.A2(n_1616),
.B(n_1577),
.Y(n_1862)
);

HB1xp67_ASAP7_75t_L g1863 ( 
.A(n_1701),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1698),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1690),
.B(n_1657),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1698),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1727),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1618),
.Y(n_1868)
);

HB1xp67_ASAP7_75t_L g1869 ( 
.A(n_1630),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1730),
.B(n_1648),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1727),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1584),
.Y(n_1872)
);

INVxp67_ASAP7_75t_L g1873 ( 
.A(n_1572),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1730),
.B(n_1639),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1584),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1584),
.Y(n_1876)
);

OAI21x1_ASAP7_75t_L g1877 ( 
.A1(n_1681),
.A2(n_1713),
.B(n_1606),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1681),
.Y(n_1878)
);

HB1xp67_ASAP7_75t_L g1879 ( 
.A(n_1651),
.Y(n_1879)
);

OAI21x1_ASAP7_75t_L g1880 ( 
.A1(n_1713),
.A2(n_1606),
.B(n_1600),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_1718),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1594),
.B(n_1626),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1724),
.B(n_1744),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1600),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1634),
.B(n_1637),
.Y(n_1885)
);

INVx2_ASAP7_75t_SL g1886 ( 
.A(n_1629),
.Y(n_1886)
);

BUFx6f_ASAP7_75t_L g1887 ( 
.A(n_1633),
.Y(n_1887)
);

AO21x1_ASAP7_75t_SL g1888 ( 
.A1(n_1696),
.A2(n_1567),
.B(n_1632),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1706),
.Y(n_1889)
);

HB1xp67_ASAP7_75t_L g1890 ( 
.A(n_1709),
.Y(n_1890)
);

INVx2_ASAP7_75t_SL g1891 ( 
.A(n_1706),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1614),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1711),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1645),
.B(n_1722),
.Y(n_1894)
);

HB1xp67_ASAP7_75t_L g1895 ( 
.A(n_1580),
.Y(n_1895)
);

OAI22xp33_ASAP7_75t_L g1896 ( 
.A1(n_1586),
.A2(n_1599),
.B1(n_1724),
.B2(n_1563),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1615),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1821),
.B(n_1739),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1828),
.A2(n_1573),
.B1(n_1569),
.B2(n_1682),
.Y(n_1899)
);

INVxp67_ASAP7_75t_L g1900 ( 
.A(n_1782),
.Y(n_1900)
);

AND2x4_ASAP7_75t_L g1901 ( 
.A(n_1820),
.B(n_1691),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1789),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1779),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1779),
.Y(n_1904)
);

AND2x6_ASAP7_75t_L g1905 ( 
.A(n_1765),
.B(n_1590),
.Y(n_1905)
);

OA21x2_ASAP7_75t_L g1906 ( 
.A1(n_1770),
.A2(n_1732),
.B(n_1728),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1780),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1821),
.B(n_1739),
.Y(n_1908)
);

NOR2xp67_ASAP7_75t_SL g1909 ( 
.A(n_1751),
.B(n_1697),
.Y(n_1909)
);

OAI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1771),
.A2(n_1736),
.B(n_1578),
.Y(n_1910)
);

CKINVDCx5p33_ASAP7_75t_R g1911 ( 
.A(n_1839),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1775),
.B(n_1602),
.Y(n_1912)
);

O2A1O1Ixp33_ASAP7_75t_SL g1913 ( 
.A1(n_1850),
.A2(n_1741),
.B(n_1834),
.C(n_1764),
.Y(n_1913)
);

OAI21x1_ASAP7_75t_SL g1914 ( 
.A1(n_1752),
.A2(n_1768),
.B(n_1776),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1808),
.B(n_1811),
.Y(n_1915)
);

AND2x4_ASAP7_75t_SL g1916 ( 
.A(n_1887),
.B(n_1894),
.Y(n_1916)
);

OAI21x1_ASAP7_75t_SL g1917 ( 
.A1(n_1776),
.A2(n_1783),
.B(n_1801),
.Y(n_1917)
);

A2O1A1Ixp33_ASAP7_75t_L g1918 ( 
.A1(n_1849),
.A2(n_1853),
.B(n_1797),
.C(n_1825),
.Y(n_1918)
);

AOI21xp5_ASAP7_75t_L g1919 ( 
.A1(n_1785),
.A2(n_1757),
.B(n_1795),
.Y(n_1919)
);

A2O1A1Ixp33_ASAP7_75t_L g1920 ( 
.A1(n_1836),
.A2(n_1848),
.B(n_1831),
.C(n_1840),
.Y(n_1920)
);

OAI21x1_ASAP7_75t_SL g1921 ( 
.A1(n_1809),
.A2(n_1841),
.B(n_1773),
.Y(n_1921)
);

OAI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1785),
.A2(n_1848),
.B(n_1830),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1763),
.B(n_1804),
.Y(n_1923)
);

O2A1O1Ixp33_ASAP7_75t_L g1924 ( 
.A1(n_1840),
.A2(n_1831),
.B(n_1859),
.C(n_1851),
.Y(n_1924)
);

NOR2xp33_ASAP7_75t_L g1925 ( 
.A(n_1774),
.B(n_1778),
.Y(n_1925)
);

NOR2x1_ASAP7_75t_SL g1926 ( 
.A(n_1888),
.B(n_1793),
.Y(n_1926)
);

AND2x4_ASAP7_75t_L g1927 ( 
.A(n_1820),
.B(n_1765),
.Y(n_1927)
);

O2A1O1Ixp33_ASAP7_75t_SL g1928 ( 
.A1(n_1896),
.A2(n_1882),
.B(n_1891),
.C(n_1889),
.Y(n_1928)
);

BUFx3_ASAP7_75t_L g1929 ( 
.A(n_1887),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1796),
.B(n_1806),
.Y(n_1930)
);

HB1xp67_ASAP7_75t_L g1931 ( 
.A(n_1862),
.Y(n_1931)
);

BUFx3_ASAP7_75t_L g1932 ( 
.A(n_1887),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1786),
.B(n_1855),
.Y(n_1933)
);

A2O1A1Ixp33_ASAP7_75t_L g1934 ( 
.A1(n_1837),
.A2(n_1819),
.B(n_1851),
.C(n_1846),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1855),
.B(n_1794),
.Y(n_1935)
);

NOR3xp33_ASAP7_75t_L g1936 ( 
.A(n_1823),
.B(n_1830),
.C(n_1846),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1777),
.B(n_1781),
.Y(n_1937)
);

OAI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1823),
.A2(n_1847),
.B(n_1812),
.Y(n_1938)
);

AOI221xp5_ASAP7_75t_L g1939 ( 
.A1(n_1847),
.A2(n_1812),
.B1(n_1766),
.B2(n_1832),
.C(n_1835),
.Y(n_1939)
);

CKINVDCx11_ASAP7_75t_R g1940 ( 
.A(n_1887),
.Y(n_1940)
);

BUFx3_ASAP7_75t_L g1941 ( 
.A(n_1887),
.Y(n_1941)
);

OA21x2_ASAP7_75t_L g1942 ( 
.A1(n_1761),
.A2(n_1810),
.B(n_1838),
.Y(n_1942)
);

AO32x2_ASAP7_75t_L g1943 ( 
.A1(n_1788),
.A2(n_1799),
.A3(n_1852),
.B1(n_1886),
.B2(n_1760),
.Y(n_1943)
);

BUFx3_ASAP7_75t_L g1944 ( 
.A(n_1860),
.Y(n_1944)
);

OAI31xp33_ASAP7_75t_SL g1945 ( 
.A1(n_1766),
.A2(n_1835),
.A3(n_1832),
.B(n_1760),
.Y(n_1945)
);

AOI22xp5_ASAP7_75t_L g1946 ( 
.A1(n_1897),
.A2(n_1845),
.B1(n_1873),
.B2(n_1784),
.Y(n_1946)
);

INVx3_ASAP7_75t_L g1947 ( 
.A(n_1862),
.Y(n_1947)
);

OAI21x1_ASAP7_75t_L g1948 ( 
.A1(n_1762),
.A2(n_1877),
.B(n_1880),
.Y(n_1948)
);

A2O1A1Ixp33_ASAP7_75t_L g1949 ( 
.A1(n_1882),
.A2(n_1843),
.B(n_1844),
.C(n_1845),
.Y(n_1949)
);

OAI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1795),
.A2(n_1757),
.B(n_1844),
.Y(n_1950)
);

CKINVDCx20_ASAP7_75t_R g1951 ( 
.A(n_1839),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1881),
.Y(n_1952)
);

OR2x2_ASAP7_75t_L g1953 ( 
.A(n_1798),
.B(n_1757),
.Y(n_1953)
);

NOR2xp33_ASAP7_75t_L g1954 ( 
.A(n_1897),
.B(n_1890),
.Y(n_1954)
);

AOI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1893),
.A2(n_1895),
.B1(n_1795),
.B2(n_1885),
.Y(n_1955)
);

AOI21xp5_ASAP7_75t_L g1956 ( 
.A1(n_1757),
.A2(n_1795),
.B(n_1838),
.Y(n_1956)
);

OAI21xp5_ASAP7_75t_L g1957 ( 
.A1(n_1843),
.A2(n_1880),
.B(n_1877),
.Y(n_1957)
);

BUFx6f_ASAP7_75t_L g1958 ( 
.A(n_1888),
.Y(n_1958)
);

OAI21xp5_ASAP7_75t_SL g1959 ( 
.A1(n_1894),
.A2(n_1885),
.B(n_1883),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1803),
.B(n_1860),
.Y(n_1960)
);

AND2x4_ASAP7_75t_L g1961 ( 
.A(n_1842),
.B(n_1791),
.Y(n_1961)
);

AOI22xp5_ASAP7_75t_L g1962 ( 
.A1(n_1893),
.A2(n_1881),
.B1(n_1856),
.B2(n_1892),
.Y(n_1962)
);

CKINVDCx20_ASAP7_75t_R g1963 ( 
.A(n_1863),
.Y(n_1963)
);

NAND3xp33_ASAP7_75t_L g1964 ( 
.A(n_1790),
.B(n_1792),
.C(n_1879),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1862),
.B(n_1870),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1862),
.B(n_1870),
.Y(n_1966)
);

NAND2xp33_ASAP7_75t_L g1967 ( 
.A(n_1793),
.B(n_1833),
.Y(n_1967)
);

INVxp33_ASAP7_75t_L g1968 ( 
.A(n_1865),
.Y(n_1968)
);

AND2x4_ASAP7_75t_L g1969 ( 
.A(n_1791),
.B(n_1800),
.Y(n_1969)
);

AO32x2_ASAP7_75t_L g1970 ( 
.A1(n_1788),
.A2(n_1799),
.A3(n_1852),
.B1(n_1886),
.B2(n_1787),
.Y(n_1970)
);

AOI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1750),
.A2(n_1759),
.B(n_1755),
.Y(n_1971)
);

AOI221xp5_ASAP7_75t_L g1972 ( 
.A1(n_1790),
.A2(n_1792),
.B1(n_1802),
.B2(n_1817),
.C(n_1813),
.Y(n_1972)
);

OR2x2_ASAP7_75t_L g1973 ( 
.A(n_1754),
.B(n_1756),
.Y(n_1973)
);

NOR2xp33_ASAP7_75t_L g1974 ( 
.A(n_1857),
.B(n_1868),
.Y(n_1974)
);

NAND3xp33_ASAP7_75t_L g1975 ( 
.A(n_1815),
.B(n_1818),
.C(n_1869),
.Y(n_1975)
);

AO21x2_ASAP7_75t_L g1976 ( 
.A1(n_1762),
.A2(n_1753),
.B(n_1767),
.Y(n_1976)
);

OR2x6_ASAP7_75t_L g1977 ( 
.A(n_1800),
.B(n_1793),
.Y(n_1977)
);

OAI22xp5_ASAP7_75t_L g1978 ( 
.A1(n_1805),
.A2(n_1892),
.B1(n_1807),
.B2(n_1889),
.Y(n_1978)
);

INVxp67_ASAP7_75t_L g1979 ( 
.A(n_1814),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1791),
.B(n_1814),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1816),
.B(n_1874),
.Y(n_1981)
);

OR2x2_ASAP7_75t_L g1982 ( 
.A(n_1772),
.B(n_1767),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1772),
.Y(n_1983)
);

OR2x6_ASAP7_75t_L g1984 ( 
.A(n_1800),
.B(n_1793),
.Y(n_1984)
);

OAI21xp5_ASAP7_75t_L g1985 ( 
.A1(n_1864),
.A2(n_1866),
.B(n_1867),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1878),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1903),
.Y(n_1987)
);

HB1xp67_ASAP7_75t_L g1988 ( 
.A(n_1931),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1950),
.B(n_1787),
.Y(n_1989)
);

AND2x4_ASAP7_75t_L g1990 ( 
.A(n_1947),
.B(n_1787),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1950),
.B(n_1787),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1965),
.B(n_1787),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1904),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1966),
.B(n_1750),
.Y(n_1994)
);

INVx1_ASAP7_75t_SL g1995 ( 
.A(n_1960),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1953),
.Y(n_1996)
);

NOR2x1_ASAP7_75t_L g1997 ( 
.A(n_1975),
.B(n_1769),
.Y(n_1997)
);

INVxp67_ASAP7_75t_SL g1998 ( 
.A(n_1964),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1907),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1976),
.Y(n_2000)
);

OAI221xp5_ASAP7_75t_SL g2001 ( 
.A1(n_1918),
.A2(n_1805),
.B1(n_1871),
.B2(n_1867),
.C(n_1866),
.Y(n_2001)
);

INVx3_ASAP7_75t_L g2002 ( 
.A(n_1948),
.Y(n_2002)
);

INVxp67_ASAP7_75t_L g2003 ( 
.A(n_1964),
.Y(n_2003)
);

INVx3_ASAP7_75t_L g2004 ( 
.A(n_1942),
.Y(n_2004)
);

BUFx2_ASAP7_75t_L g2005 ( 
.A(n_1943),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1942),
.B(n_1758),
.Y(n_2006)
);

BUFx12f_ASAP7_75t_L g2007 ( 
.A(n_1940),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1943),
.B(n_1758),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1919),
.B(n_1956),
.Y(n_2009)
);

INVxp67_ASAP7_75t_SL g2010 ( 
.A(n_1900),
.Y(n_2010)
);

AND2x4_ASAP7_75t_L g2011 ( 
.A(n_1971),
.B(n_1769),
.Y(n_2011)
);

HB1xp67_ASAP7_75t_L g2012 ( 
.A(n_1900),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1973),
.Y(n_2013)
);

HB1xp67_ASAP7_75t_L g2014 ( 
.A(n_1980),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1922),
.B(n_1829),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1922),
.B(n_1829),
.Y(n_2016)
);

BUFx3_ASAP7_75t_L g2017 ( 
.A(n_1905),
.Y(n_2017)
);

AOI21xp5_ASAP7_75t_L g2018 ( 
.A1(n_1967),
.A2(n_1793),
.B(n_1833),
.Y(n_2018)
);

HB1xp67_ASAP7_75t_L g2019 ( 
.A(n_1980),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1902),
.B(n_1822),
.Y(n_2020)
);

AND2x4_ASAP7_75t_L g2021 ( 
.A(n_1957),
.B(n_1824),
.Y(n_2021)
);

BUFx3_ASAP7_75t_L g2022 ( 
.A(n_1905),
.Y(n_2022)
);

NOR2xp33_ASAP7_75t_L g2023 ( 
.A(n_1968),
.B(n_1884),
.Y(n_2023)
);

HB1xp67_ASAP7_75t_L g2024 ( 
.A(n_1979),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1930),
.B(n_1970),
.Y(n_2025)
);

HB1xp67_ASAP7_75t_L g2026 ( 
.A(n_1979),
.Y(n_2026)
);

AOI22xp33_ASAP7_75t_L g2027 ( 
.A1(n_1914),
.A2(n_1861),
.B1(n_1858),
.B2(n_1854),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_1970),
.B(n_1826),
.Y(n_2028)
);

NOR2xp33_ASAP7_75t_L g2029 ( 
.A(n_1925),
.B(n_1959),
.Y(n_2029)
);

BUFx3_ASAP7_75t_L g2030 ( 
.A(n_1905),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1970),
.B(n_1827),
.Y(n_2031)
);

BUFx2_ASAP7_75t_L g2032 ( 
.A(n_2021),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_2025),
.B(n_1923),
.Y(n_2033)
);

OAI22xp5_ASAP7_75t_L g2034 ( 
.A1(n_2001),
.A2(n_1920),
.B1(n_1899),
.B2(n_1959),
.Y(n_2034)
);

AOI221xp5_ASAP7_75t_L g2035 ( 
.A1(n_2003),
.A2(n_1899),
.B1(n_1921),
.B2(n_1917),
.C(n_1934),
.Y(n_2035)
);

AOI33xp33_ASAP7_75t_L g2036 ( 
.A1(n_1989),
.A2(n_1991),
.A3(n_2009),
.B1(n_1939),
.B2(n_2027),
.B3(n_2015),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_2025),
.B(n_1955),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_2025),
.B(n_1915),
.Y(n_2038)
);

NAND3xp33_ASAP7_75t_L g2039 ( 
.A(n_2003),
.B(n_1949),
.C(n_1945),
.Y(n_2039)
);

OAI21xp33_ASAP7_75t_SL g2040 ( 
.A1(n_1998),
.A2(n_1945),
.B(n_1939),
.Y(n_2040)
);

AOI22xp33_ASAP7_75t_L g2041 ( 
.A1(n_2029),
.A2(n_1909),
.B1(n_1936),
.B2(n_1908),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_2014),
.Y(n_2042)
);

AO21x2_ASAP7_75t_L g2043 ( 
.A1(n_2000),
.A2(n_1985),
.B(n_1938),
.Y(n_2043)
);

AND2x4_ASAP7_75t_L g2044 ( 
.A(n_2021),
.B(n_1969),
.Y(n_2044)
);

OAI221xp5_ASAP7_75t_L g2045 ( 
.A1(n_1998),
.A2(n_1910),
.B1(n_1962),
.B2(n_1928),
.C(n_1946),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2014),
.Y(n_2046)
);

AND2x4_ASAP7_75t_L g2047 ( 
.A(n_2021),
.B(n_1961),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2019),
.Y(n_2048)
);

OAI22xp5_ASAP7_75t_SL g2049 ( 
.A1(n_2007),
.A2(n_1910),
.B1(n_1963),
.B2(n_1951),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_2019),
.Y(n_2050)
);

HB1xp67_ASAP7_75t_L g2051 ( 
.A(n_2024),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1988),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_1992),
.B(n_1944),
.Y(n_2053)
);

AOI22xp33_ASAP7_75t_L g2054 ( 
.A1(n_2017),
.A2(n_1898),
.B1(n_1912),
.B2(n_1905),
.Y(n_2054)
);

INVxp67_ASAP7_75t_SL g2055 ( 
.A(n_1997),
.Y(n_2055)
);

AND2x4_ASAP7_75t_L g2056 ( 
.A(n_2021),
.B(n_1961),
.Y(n_2056)
);

OAI221xp5_ASAP7_75t_L g2057 ( 
.A1(n_2001),
.A2(n_1913),
.B1(n_1924),
.B2(n_1938),
.C(n_1954),
.Y(n_2057)
);

BUFx6f_ASAP7_75t_L g2058 ( 
.A(n_2007),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1988),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1987),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1987),
.Y(n_2061)
);

AOI322xp5_ASAP7_75t_L g2062 ( 
.A1(n_1989),
.A2(n_1972),
.A3(n_1901),
.B1(n_1924),
.B2(n_1958),
.C1(n_1941),
.C2(n_1929),
.Y(n_2062)
);

AOI21xp5_ASAP7_75t_L g2063 ( 
.A1(n_1997),
.A2(n_1926),
.B(n_1906),
.Y(n_2063)
);

AOI22xp33_ASAP7_75t_L g2064 ( 
.A1(n_2017),
.A2(n_1927),
.B1(n_1958),
.B2(n_1901),
.Y(n_2064)
);

OAI33xp33_ASAP7_75t_L g2065 ( 
.A1(n_2020),
.A2(n_1978),
.A3(n_1975),
.B1(n_1982),
.B2(n_1983),
.B3(n_1986),
.Y(n_2065)
);

AOI21xp5_ASAP7_75t_SL g2066 ( 
.A1(n_2017),
.A2(n_1906),
.B(n_1958),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1993),
.Y(n_2067)
);

BUFx2_ASAP7_75t_L g2068 ( 
.A(n_2021),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_2006),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1993),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1999),
.Y(n_2071)
);

BUFx3_ASAP7_75t_L g2072 ( 
.A(n_2007),
.Y(n_2072)
);

AOI22xp33_ASAP7_75t_L g2073 ( 
.A1(n_2022),
.A2(n_1927),
.B1(n_1933),
.B2(n_1935),
.Y(n_2073)
);

INVx5_ASAP7_75t_L g2074 ( 
.A(n_2004),
.Y(n_2074)
);

OAI221xp5_ASAP7_75t_SL g2075 ( 
.A1(n_1989),
.A2(n_1972),
.B1(n_1974),
.B2(n_1984),
.C(n_1977),
.Y(n_2075)
);

HB1xp67_ASAP7_75t_L g2076 ( 
.A(n_2026),
.Y(n_2076)
);

AND2x4_ASAP7_75t_L g2077 ( 
.A(n_1990),
.B(n_1977),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_1992),
.B(n_1981),
.Y(n_2078)
);

OAI31xp33_ASAP7_75t_L g2079 ( 
.A1(n_1991),
.A2(n_1978),
.A3(n_1916),
.B(n_1932),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1999),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_1994),
.B(n_1937),
.Y(n_2081)
);

INVx2_ASAP7_75t_SL g2082 ( 
.A(n_2074),
.Y(n_2082)
);

INVxp67_ASAP7_75t_SL g2083 ( 
.A(n_2051),
.Y(n_2083)
);

AND2x4_ASAP7_75t_L g2084 ( 
.A(n_2032),
.B(n_1990),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2042),
.B(n_2010),
.Y(n_2085)
);

BUFx3_ASAP7_75t_L g2086 ( 
.A(n_2058),
.Y(n_2086)
);

AOI21xp33_ASAP7_75t_L g2087 ( 
.A1(n_2040),
.A2(n_1991),
.B(n_2009),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_2032),
.B(n_2005),
.Y(n_2088)
);

INVx3_ASAP7_75t_L g2089 ( 
.A(n_2074),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_2042),
.B(n_2010),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_2046),
.B(n_2012),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_2046),
.B(n_2012),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_2068),
.B(n_2005),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_2048),
.B(n_1996),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2060),
.Y(n_2095)
);

BUFx2_ASAP7_75t_L g2096 ( 
.A(n_2055),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2060),
.Y(n_2097)
);

HB1xp67_ASAP7_75t_L g2098 ( 
.A(n_2076),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2061),
.Y(n_2099)
);

AOI22xp5_ASAP7_75t_L g2100 ( 
.A1(n_2034),
.A2(n_2023),
.B1(n_2022),
.B2(n_2030),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2068),
.B(n_2028),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_2037),
.B(n_2028),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2061),
.Y(n_2103)
);

INVx3_ASAP7_75t_L g2104 ( 
.A(n_2074),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_2037),
.B(n_2028),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_2038),
.B(n_2031),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2038),
.B(n_2031),
.Y(n_2107)
);

OR2x2_ASAP7_75t_L g2108 ( 
.A(n_2069),
.B(n_2031),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2067),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2067),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2070),
.Y(n_2111)
);

OR2x2_ASAP7_75t_L g2112 ( 
.A(n_2052),
.B(n_2000),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_2033),
.B(n_2015),
.Y(n_2113)
);

AND2x4_ASAP7_75t_L g2114 ( 
.A(n_2077),
.B(n_1990),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2033),
.B(n_2015),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_2078),
.B(n_2016),
.Y(n_2116)
);

AOI22xp5_ASAP7_75t_L g2117 ( 
.A1(n_2040),
.A2(n_2030),
.B1(n_2016),
.B2(n_2009),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_2078),
.B(n_2016),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_2050),
.B(n_2013),
.Y(n_2119)
);

AND2x4_ASAP7_75t_L g2120 ( 
.A(n_2077),
.B(n_2011),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2070),
.Y(n_2121)
);

BUFx2_ASAP7_75t_L g2122 ( 
.A(n_2077),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_2077),
.B(n_2008),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2071),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2080),
.Y(n_2125)
);

OR2x2_ASAP7_75t_L g2126 ( 
.A(n_2083),
.B(n_2050),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2095),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2095),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2102),
.B(n_2105),
.Y(n_2129)
);

NOR2xp33_ASAP7_75t_L g2130 ( 
.A(n_2086),
.B(n_2058),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_2102),
.B(n_2044),
.Y(n_2131)
);

INVxp67_ASAP7_75t_L g2132 ( 
.A(n_2098),
.Y(n_2132)
);

AND2x4_ASAP7_75t_L g2133 ( 
.A(n_2122),
.B(n_2044),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2097),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_2108),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2102),
.B(n_2044),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2097),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_2105),
.B(n_2044),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2105),
.B(n_2047),
.Y(n_2139)
);

AOI211xp5_ASAP7_75t_L g2140 ( 
.A1(n_2087),
.A2(n_2045),
.B(n_2039),
.C(n_2049),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2122),
.B(n_2047),
.Y(n_2141)
);

NOR2xp33_ASAP7_75t_L g2142 ( 
.A(n_2086),
.B(n_2058),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_2122),
.B(n_2047),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2099),
.Y(n_2144)
);

HB1xp67_ASAP7_75t_L g2145 ( 
.A(n_2098),
.Y(n_2145)
);

OR2x2_ASAP7_75t_L g2146 ( 
.A(n_2083),
.B(n_2052),
.Y(n_2146)
);

NOR2xp33_ASAP7_75t_L g2147 ( 
.A(n_2086),
.B(n_2058),
.Y(n_2147)
);

AND2x2_ASAP7_75t_L g2148 ( 
.A(n_2116),
.B(n_2047),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2116),
.B(n_2056),
.Y(n_2149)
);

NOR2x1_ASAP7_75t_R g2150 ( 
.A(n_2086),
.B(n_2058),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2116),
.B(n_2056),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2099),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2118),
.B(n_2056),
.Y(n_2153)
);

OAI211xp5_ASAP7_75t_SL g2154 ( 
.A1(n_2117),
.A2(n_2062),
.B(n_2035),
.C(n_2036),
.Y(n_2154)
);

INVxp67_ASAP7_75t_L g2155 ( 
.A(n_2100),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_2118),
.B(n_2123),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2103),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2100),
.B(n_2062),
.Y(n_2158)
);

NAND3x1_ASAP7_75t_L g2159 ( 
.A(n_2117),
.B(n_2063),
.C(n_2079),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2103),
.Y(n_2160)
);

INVx4_ASAP7_75t_L g2161 ( 
.A(n_2089),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2109),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_2118),
.B(n_2056),
.Y(n_2163)
);

OR2x2_ASAP7_75t_L g2164 ( 
.A(n_2085),
.B(n_2059),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2109),
.Y(n_2165)
);

AOI22xp5_ASAP7_75t_L g2166 ( 
.A1(n_2087),
.A2(n_2057),
.B1(n_2049),
.B2(n_2065),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2110),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2091),
.B(n_1995),
.Y(n_2168)
);

OR2x2_ASAP7_75t_L g2169 ( 
.A(n_2085),
.B(n_2059),
.Y(n_2169)
);

AND2x4_ASAP7_75t_L g2170 ( 
.A(n_2123),
.B(n_2030),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2110),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2111),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2123),
.B(n_2081),
.Y(n_2173)
);

HB1xp67_ASAP7_75t_L g2174 ( 
.A(n_2096),
.Y(n_2174)
);

INVxp67_ASAP7_75t_SL g2175 ( 
.A(n_2096),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2111),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_2113),
.B(n_2081),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2121),
.Y(n_2178)
);

INVxp67_ASAP7_75t_SL g2179 ( 
.A(n_2096),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_2113),
.B(n_2053),
.Y(n_2180)
);

INVx5_ASAP7_75t_L g2181 ( 
.A(n_2089),
.Y(n_2181)
);

OR2x2_ASAP7_75t_L g2182 ( 
.A(n_2090),
.B(n_2091),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2127),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_2129),
.B(n_2113),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2166),
.B(n_2115),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2127),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_2129),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2180),
.B(n_2115),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_2180),
.B(n_2115),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_2131),
.B(n_2114),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_2155),
.B(n_2092),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2134),
.Y(n_2192)
);

AOI21xp5_ASAP7_75t_L g2193 ( 
.A1(n_2140),
.A2(n_2075),
.B(n_2041),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_2156),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2134),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2158),
.B(n_2092),
.Y(n_2196)
);

INVx1_ASAP7_75t_SL g2197 ( 
.A(n_2145),
.Y(n_2197)
);

INVx1_ASAP7_75t_SL g2198 ( 
.A(n_2130),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2137),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2137),
.Y(n_2200)
);

OR2x2_ASAP7_75t_L g2201 ( 
.A(n_2182),
.B(n_2164),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_2131),
.B(n_2114),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_2136),
.B(n_2114),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_2136),
.B(n_2114),
.Y(n_2204)
);

OAI21xp33_ASAP7_75t_L g2205 ( 
.A1(n_2154),
.A2(n_2093),
.B(n_2088),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2144),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2132),
.B(n_2090),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2144),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_2142),
.B(n_2119),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2147),
.B(n_2173),
.Y(n_2210)
);

AND2x4_ASAP7_75t_L g2211 ( 
.A(n_2170),
.B(n_2082),
.Y(n_2211)
);

AND2x2_ASAP7_75t_L g2212 ( 
.A(n_2138),
.B(n_2156),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_2173),
.B(n_2119),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_2182),
.B(n_2088),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2152),
.Y(n_2215)
);

AOI21xp33_ASAP7_75t_SL g2216 ( 
.A1(n_2174),
.A2(n_1952),
.B(n_1911),
.Y(n_2216)
);

OR2x2_ASAP7_75t_L g2217 ( 
.A(n_2164),
.B(n_2094),
.Y(n_2217)
);

INVx2_ASAP7_75t_SL g2218 ( 
.A(n_2181),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2152),
.Y(n_2219)
);

HB1xp67_ASAP7_75t_L g2220 ( 
.A(n_2175),
.Y(n_2220)
);

OR2x2_ASAP7_75t_L g2221 ( 
.A(n_2169),
.B(n_2146),
.Y(n_2221)
);

AND2x2_ASAP7_75t_SL g2222 ( 
.A(n_2161),
.B(n_2054),
.Y(n_2222)
);

OR2x2_ASAP7_75t_L g2223 ( 
.A(n_2169),
.B(n_2094),
.Y(n_2223)
);

INVx1_ASAP7_75t_SL g2224 ( 
.A(n_2170),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_2138),
.B(n_2114),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_2212),
.B(n_2170),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_2218),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_2218),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2220),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_2197),
.B(n_2177),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_SL g2231 ( 
.A(n_2216),
.B(n_2072),
.Y(n_2231)
);

NOR2xp33_ASAP7_75t_L g2232 ( 
.A(n_2198),
.B(n_2072),
.Y(n_2232)
);

O2A1O1Ixp33_ASAP7_75t_L g2233 ( 
.A1(n_2193),
.A2(n_2179),
.B(n_2082),
.C(n_2159),
.Y(n_2233)
);

OR2x2_ASAP7_75t_L g2234 ( 
.A(n_2221),
.B(n_2146),
.Y(n_2234)
);

AOI322xp5_ASAP7_75t_L g2235 ( 
.A1(n_2205),
.A2(n_2093),
.A3(n_2088),
.B1(n_2101),
.B2(n_2177),
.C1(n_2106),
.C2(n_2107),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_2212),
.B(n_2139),
.Y(n_2236)
);

OAI21xp33_ASAP7_75t_L g2237 ( 
.A1(n_2196),
.A2(n_2185),
.B(n_2191),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2183),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2183),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2186),
.Y(n_2240)
);

OAI21xp33_ASAP7_75t_L g2241 ( 
.A1(n_2210),
.A2(n_2143),
.B(n_2141),
.Y(n_2241)
);

AOI21xp33_ASAP7_75t_L g2242 ( 
.A1(n_2222),
.A2(n_2150),
.B(n_2159),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_2190),
.B(n_2139),
.Y(n_2243)
);

INVxp67_ASAP7_75t_SL g2244 ( 
.A(n_2211),
.Y(n_2244)
);

AOI31xp33_ASAP7_75t_L g2245 ( 
.A1(n_2224),
.A2(n_2209),
.A3(n_2207),
.B(n_2201),
.Y(n_2245)
);

NOR2xp67_ASAP7_75t_SL g2246 ( 
.A(n_2221),
.B(n_2066),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2190),
.B(n_2141),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2186),
.Y(n_2248)
);

OAI221xp5_ASAP7_75t_L g2249 ( 
.A1(n_2214),
.A2(n_2082),
.B1(n_2089),
.B2(n_2104),
.C(n_2161),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_2184),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2188),
.B(n_2143),
.Y(n_2251)
);

AOI221xp5_ASAP7_75t_L g2252 ( 
.A1(n_2194),
.A2(n_2135),
.B1(n_2133),
.B2(n_2176),
.C(n_2172),
.Y(n_2252)
);

OAI22xp33_ASAP7_75t_SL g2253 ( 
.A1(n_2201),
.A2(n_2181),
.B1(n_2161),
.B2(n_2104),
.Y(n_2253)
);

OAI31xp33_ASAP7_75t_L g2254 ( 
.A1(n_2211),
.A2(n_2133),
.A3(n_2089),
.B(n_2104),
.Y(n_2254)
);

OAI21xp5_ASAP7_75t_L g2255 ( 
.A1(n_2222),
.A2(n_2181),
.B(n_2126),
.Y(n_2255)
);

OAI221xp5_ASAP7_75t_L g2256 ( 
.A1(n_2233),
.A2(n_2194),
.B1(n_2187),
.B2(n_2213),
.C(n_2217),
.Y(n_2256)
);

OR2x2_ASAP7_75t_L g2257 ( 
.A(n_2234),
.B(n_2187),
.Y(n_2257)
);

AOI22xp33_ASAP7_75t_L g2258 ( 
.A1(n_2242),
.A2(n_2237),
.B1(n_2241),
.B2(n_2222),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2238),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2238),
.Y(n_2260)
);

NOR2xp33_ASAP7_75t_SL g2261 ( 
.A(n_2232),
.B(n_2181),
.Y(n_2261)
);

NAND4xp75_ASAP7_75t_L g2262 ( 
.A(n_2255),
.B(n_2200),
.C(n_2199),
.D(n_2195),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2226),
.B(n_2211),
.Y(n_2263)
);

AND2x2_ASAP7_75t_SL g2264 ( 
.A(n_2229),
.B(n_2133),
.Y(n_2264)
);

OAI221xp5_ASAP7_75t_L g2265 ( 
.A1(n_2245),
.A2(n_2223),
.B1(n_2217),
.B2(n_2089),
.C(n_2104),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2244),
.B(n_2188),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_2226),
.B(n_2202),
.Y(n_2267)
);

AOI22xp5_ASAP7_75t_L g2268 ( 
.A1(n_2231),
.A2(n_2225),
.B1(n_2202),
.B2(n_2203),
.Y(n_2268)
);

AOI22xp33_ASAP7_75t_L g2269 ( 
.A1(n_2250),
.A2(n_2225),
.B1(n_2203),
.B2(n_2204),
.Y(n_2269)
);

OR2x2_ASAP7_75t_L g2270 ( 
.A(n_2234),
.B(n_2223),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_2247),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_2247),
.Y(n_2272)
);

AOI221xp5_ASAP7_75t_L g2273 ( 
.A1(n_2229),
.A2(n_2219),
.B1(n_2215),
.B2(n_2208),
.C(n_2206),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2239),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2227),
.B(n_2189),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2239),
.Y(n_2276)
);

HB1xp67_ASAP7_75t_L g2277 ( 
.A(n_2227),
.Y(n_2277)
);

AND2x4_ASAP7_75t_SL g2278 ( 
.A(n_2228),
.B(n_2104),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2277),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2257),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_2258),
.B(n_2228),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2257),
.Y(n_2282)
);

INVx1_ASAP7_75t_SL g2283 ( 
.A(n_2264),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2271),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2271),
.Y(n_2285)
);

BUFx2_ASAP7_75t_L g2286 ( 
.A(n_2264),
.Y(n_2286)
);

OAI21xp5_ASAP7_75t_L g2287 ( 
.A1(n_2262),
.A2(n_2235),
.B(n_2253),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2272),
.Y(n_2288)
);

INVx1_ASAP7_75t_SL g2289 ( 
.A(n_2263),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2272),
.Y(n_2290)
);

AND3x1_ASAP7_75t_L g2291 ( 
.A(n_2261),
.B(n_2254),
.C(n_2252),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2263),
.Y(n_2292)
);

INVxp67_ASAP7_75t_L g2293 ( 
.A(n_2266),
.Y(n_2293)
);

AOI22xp5_ASAP7_75t_L g2294 ( 
.A1(n_2268),
.A2(n_2250),
.B1(n_2230),
.B2(n_2246),
.Y(n_2294)
);

AOI21xp5_ASAP7_75t_L g2295 ( 
.A1(n_2287),
.A2(n_2265),
.B(n_2256),
.Y(n_2295)
);

HB1xp67_ASAP7_75t_L g2296 ( 
.A(n_2286),
.Y(n_2296)
);

NOR3xp33_ASAP7_75t_L g2297 ( 
.A(n_2281),
.B(n_2262),
.C(n_2273),
.Y(n_2297)
);

INVxp67_ASAP7_75t_L g2298 ( 
.A(n_2286),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2280),
.Y(n_2299)
);

BUFx2_ASAP7_75t_L g2300 ( 
.A(n_2280),
.Y(n_2300)
);

NOR4xp25_ASAP7_75t_L g2301 ( 
.A(n_2283),
.B(n_2259),
.C(n_2274),
.D(n_2260),
.Y(n_2301)
);

NOR2xp67_ASAP7_75t_L g2302 ( 
.A(n_2282),
.B(n_2270),
.Y(n_2302)
);

AOI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_2291),
.A2(n_2267),
.B1(n_2275),
.B2(n_2246),
.Y(n_2303)
);

NOR2xp33_ASAP7_75t_L g2304 ( 
.A(n_2293),
.B(n_2270),
.Y(n_2304)
);

OAI21xp5_ASAP7_75t_L g2305 ( 
.A1(n_2294),
.A2(n_2289),
.B(n_2282),
.Y(n_2305)
);

NOR2xp33_ASAP7_75t_L g2306 ( 
.A(n_2292),
.B(n_2267),
.Y(n_2306)
);

NOR4xp25_ASAP7_75t_L g2307 ( 
.A(n_2279),
.B(n_2276),
.C(n_2248),
.D(n_2240),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2292),
.B(n_2269),
.Y(n_2308)
);

AOI221xp5_ASAP7_75t_L g2309 ( 
.A1(n_2297),
.A2(n_2290),
.B1(n_2288),
.B2(n_2285),
.C(n_2284),
.Y(n_2309)
);

XOR2xp5_ASAP7_75t_L g2310 ( 
.A(n_2303),
.B(n_2251),
.Y(n_2310)
);

OAI21xp33_ASAP7_75t_L g2311 ( 
.A1(n_2306),
.A2(n_2278),
.B(n_2249),
.Y(n_2311)
);

AOI221xp5_ASAP7_75t_L g2312 ( 
.A1(n_2301),
.A2(n_2276),
.B1(n_2248),
.B2(n_2240),
.C(n_2278),
.Y(n_2312)
);

AOI22xp5_ASAP7_75t_L g2313 ( 
.A1(n_2295),
.A2(n_2236),
.B1(n_2243),
.B2(n_2219),
.Y(n_2313)
);

NOR2x1_ASAP7_75t_L g2314 ( 
.A(n_2302),
.B(n_2192),
.Y(n_2314)
);

O2A1O1Ixp33_ASAP7_75t_L g2315 ( 
.A1(n_2296),
.A2(n_2199),
.B(n_2215),
.C(n_2192),
.Y(n_2315)
);

AND3x4_ASAP7_75t_L g2316 ( 
.A(n_2307),
.B(n_2120),
.C(n_2084),
.Y(n_2316)
);

AO221x1_ASAP7_75t_L g2317 ( 
.A1(n_2298),
.A2(n_2195),
.B1(n_2208),
.B2(n_2206),
.C(n_2200),
.Y(n_2317)
);

O2A1O1Ixp33_ASAP7_75t_L g2318 ( 
.A1(n_2298),
.A2(n_2236),
.B(n_2126),
.C(n_2243),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2300),
.B(n_2189),
.Y(n_2319)
);

OAI221xp5_ASAP7_75t_SL g2320 ( 
.A1(n_2311),
.A2(n_2308),
.B1(n_2304),
.B2(n_2299),
.C(n_2305),
.Y(n_2320)
);

XNOR2x2_ASAP7_75t_L g2321 ( 
.A(n_2314),
.B(n_2184),
.Y(n_2321)
);

AOI221xp5_ASAP7_75t_L g2322 ( 
.A1(n_2309),
.A2(n_2181),
.B1(n_2135),
.B2(n_2204),
.C(n_2157),
.Y(n_2322)
);

AOI21xp33_ASAP7_75t_R g2323 ( 
.A1(n_2319),
.A2(n_2157),
.B(n_2128),
.Y(n_2323)
);

AOI321xp33_ASAP7_75t_L g2324 ( 
.A1(n_2318),
.A2(n_2313),
.A3(n_2312),
.B1(n_2315),
.B2(n_2310),
.C(n_2316),
.Y(n_2324)
);

OAI21xp33_ASAP7_75t_L g2325 ( 
.A1(n_2317),
.A2(n_2162),
.B(n_2160),
.Y(n_2325)
);

AOI32xp33_ASAP7_75t_L g2326 ( 
.A1(n_2314),
.A2(n_2093),
.A3(n_2151),
.B1(n_2153),
.B2(n_2149),
.Y(n_2326)
);

AOI32xp33_ASAP7_75t_L g2327 ( 
.A1(n_2314),
.A2(n_2163),
.A3(n_2149),
.B1(n_2148),
.B2(n_2153),
.Y(n_2327)
);

XNOR2x1_ASAP7_75t_L g2328 ( 
.A(n_2310),
.B(n_2148),
.Y(n_2328)
);

XOR2xp5_ASAP7_75t_L g2329 ( 
.A(n_2328),
.B(n_2064),
.Y(n_2329)
);

NOR2x1_ASAP7_75t_L g2330 ( 
.A(n_2325),
.B(n_2165),
.Y(n_2330)
);

NOR2xp67_ASAP7_75t_SL g2331 ( 
.A(n_2320),
.B(n_2066),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2321),
.Y(n_2332)
);

AO22x2_ASAP7_75t_L g2333 ( 
.A1(n_2324),
.A2(n_2178),
.B1(n_2171),
.B2(n_2167),
.Y(n_2333)
);

AOI22xp5_ASAP7_75t_L g2334 ( 
.A1(n_2322),
.A2(n_2163),
.B1(n_2151),
.B2(n_2084),
.Y(n_2334)
);

OAI22xp5_ASAP7_75t_L g2335 ( 
.A1(n_2326),
.A2(n_2168),
.B1(n_2084),
.B2(n_2112),
.Y(n_2335)
);

NOR2x1p5_ASAP7_75t_L g2336 ( 
.A(n_2332),
.B(n_2323),
.Y(n_2336)
);

AOI22xp33_ASAP7_75t_L g2337 ( 
.A1(n_2333),
.A2(n_2327),
.B1(n_2002),
.B2(n_2043),
.Y(n_2337)
);

OAI22xp5_ASAP7_75t_L g2338 ( 
.A1(n_2334),
.A2(n_2112),
.B1(n_2101),
.B2(n_2084),
.Y(n_2338)
);

OAI211xp5_ASAP7_75t_SL g2339 ( 
.A1(n_2330),
.A2(n_2018),
.B(n_2073),
.C(n_1875),
.Y(n_2339)
);

AND3x2_ASAP7_75t_L g2340 ( 
.A(n_2336),
.B(n_2331),
.C(n_2329),
.Y(n_2340)
);

OAI22xp5_ASAP7_75t_SL g2341 ( 
.A1(n_2337),
.A2(n_2335),
.B1(n_1891),
.B2(n_2084),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2340),
.B(n_2338),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2342),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2342),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_2343),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2344),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2345),
.Y(n_2347)
);

INVxp67_ASAP7_75t_SL g2348 ( 
.A(n_2346),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_2347),
.Y(n_2349)
);

XNOR2xp5_ASAP7_75t_L g2350 ( 
.A(n_2349),
.B(n_2348),
.Y(n_2350)
);

NOR2xp67_ASAP7_75t_L g2351 ( 
.A(n_2350),
.B(n_2341),
.Y(n_2351)
);

AOI221xp5_ASAP7_75t_L g2352 ( 
.A1(n_2351),
.A2(n_2339),
.B1(n_2121),
.B2(n_2125),
.C(n_2124),
.Y(n_2352)
);

AOI211xp5_ASAP7_75t_L g2353 ( 
.A1(n_2352),
.A2(n_1872),
.B(n_1875),
.C(n_1876),
.Y(n_2353)
);


endmodule