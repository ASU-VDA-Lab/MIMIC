module real_jpeg_26358_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_206;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_1),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_1),
.A2(n_27),
.B1(n_53),
.B2(n_54),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_1),
.A2(n_27),
.B1(n_67),
.B2(n_68),
.Y(n_221)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_2),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_2),
.B(n_30),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_L g195 ( 
.A1(n_2),
.A2(n_53),
.B1(n_54),
.B2(n_61),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_2),
.B(n_68),
.C(n_82),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_2),
.B(n_52),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_2),
.A2(n_105),
.B1(n_214),
.B2(n_221),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_3),
.A2(n_67),
.B1(n_68),
.B2(n_73),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_3),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_3),
.A2(n_53),
.B1(n_54),
.B2(n_73),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_4),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_5),
.A2(n_46),
.B1(n_96),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_5),
.A2(n_46),
.B1(n_53),
.B2(n_54),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_5),
.A2(n_46),
.B1(n_67),
.B2(n_68),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

INVx8_ASAP7_75t_SL g36 ( 
.A(n_7),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_8),
.A2(n_25),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_40),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_8),
.A2(n_40),
.B1(n_53),
.B2(n_54),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_8),
.A2(n_40),
.B1(n_67),
.B2(n_68),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_9),
.A2(n_67),
.B1(n_68),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_9),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_9),
.A2(n_53),
.B1(n_54),
.B2(n_75),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_10),
.A2(n_53),
.B1(n_54),
.B2(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_10),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_10),
.A2(n_67),
.B1(n_68),
.B2(n_89),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_89),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_12),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_12),
.A2(n_53),
.B1(n_54),
.B2(n_57),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_12),
.A2(n_57),
.B1(n_67),
.B2(n_68),
.Y(n_119)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_15),
.Y(n_110)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_15),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_142),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_140),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_111),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_19),
.B(n_111),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_76),
.C(n_99),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_20),
.B(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_58),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_43),
.B2(n_44),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_23),
.B(n_43),
.C(n_58),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B1(n_30),
.B2(n_39),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_24),
.Y(n_98)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_28),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_28),
.A2(n_30),
.B1(n_39),
.B2(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_37),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_29),
.A2(n_94),
.B1(n_95),
.B2(n_98),
.Y(n_93)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_31),
.A2(n_32),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_31),
.A2(n_35),
.B(n_60),
.C(n_63),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g169 ( 
.A(n_31),
.B(n_61),
.CON(n_169),
.SN(n_169)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_32),
.B(n_34),
.C(n_42),
.Y(n_63)
);

OAI32xp33_ASAP7_75t_L g168 ( 
.A1(n_32),
.A2(n_51),
.A3(n_54),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp33_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B(n_55),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_45),
.A2(n_47),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_47),
.A2(n_134),
.B(n_135),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_47),
.A2(n_91),
.B1(n_92),
.B2(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_48),
.A2(n_52),
.B1(n_159),
.B2(n_169),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

AO22x1_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_50),
.B(n_53),
.Y(n_170)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_52),
.B(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_52),
.B(n_136),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_53),
.A2(n_54),
.B1(n_82),
.B2(n_84),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_54),
.B(n_198),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_56),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_64),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_59),
.A2(n_64),
.B1(n_65),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_59),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_60),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_61),
.B(n_85),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_61),
.B(n_222),
.Y(n_227)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_69),
.B1(n_71),
.B2(n_74),
.Y(n_65)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_66),
.B(n_108),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_66),
.A2(n_210),
.B1(n_212),
.B2(n_213),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_67),
.A2(n_68),
.B1(n_82),
.B2(n_84),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_67),
.B(n_227),
.Y(n_226)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_69),
.Y(n_154)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_70),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_72),
.A2(n_120),
.B(n_154),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_76),
.A2(n_77),
.B1(n_99),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_90),
.C(n_93),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_78),
.A2(n_79),
.B1(n_90),
.B2(n_149),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_86),
.B(n_87),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_80),
.B(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_80),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_80),
.A2(n_123),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_80),
.A2(n_176),
.B(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_80),
.A2(n_123),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_80),
.A2(n_123),
.B1(n_175),
.B2(n_196),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.Y(n_80)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

BUFx24_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_101),
.B(n_102),
.Y(n_100)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_85),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_86),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_93),
.B(n_148),
.Y(n_147)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_99),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_104),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B(n_107),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_105),
.A2(n_107),
.B(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_105),
.A2(n_117),
.B(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_105),
.A2(n_211),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_SL g118 ( 
.A(n_110),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_138),
.B2(n_139),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_126),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_121),
.B2(n_125),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_119),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_121),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_137),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_132),
.B2(n_133),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_138),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_242),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_163),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_160),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_146),
.B(n_160),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.C(n_152),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_147),
.B(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_150),
.B(n_152),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.C(n_157),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_155),
.B1(n_156),
.B2(n_181),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_153),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_237),
.B(n_241),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_190),
.B(n_236),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_177),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_166),
.B(n_177),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_173),
.C(n_174),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_167),
.B(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_171),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_173),
.B(n_174),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_182),
.B2(n_183),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_178),
.B(n_185),
.C(n_189),
.Y(n_238)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_189),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_184),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_231),
.B(n_235),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_207),
.B(n_230),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_199),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_193),
.B(n_199),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_197),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_205),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_204),
.C(n_205),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_203),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_206),
.Y(n_212)
);

AOI21xp33_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_217),
.B(n_229),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_216),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_216),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_224),
.B(n_228),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_219),
.B(n_220),
.Y(n_228)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_232),
.B(n_233),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_238),
.B(n_239),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);


endmodule