module fake_netlist_1_3576_n_541 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_541);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_541;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_10), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_16), .Y(n_79) );
INVxp33_ASAP7_75t_SL g80 ( .A(n_1), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_42), .Y(n_81) );
INVx1_ASAP7_75t_SL g82 ( .A(n_4), .Y(n_82) );
INVxp33_ASAP7_75t_SL g83 ( .A(n_58), .Y(n_83) );
INVxp33_ASAP7_75t_SL g84 ( .A(n_8), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_44), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_29), .Y(n_86) );
BUFx10_ASAP7_75t_L g87 ( .A(n_68), .Y(n_87) );
BUFx3_ASAP7_75t_L g88 ( .A(n_16), .Y(n_88) );
CKINVDCx16_ASAP7_75t_R g89 ( .A(n_75), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_55), .Y(n_90) );
CKINVDCx20_ASAP7_75t_R g91 ( .A(n_56), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_4), .Y(n_92) );
INVxp33_ASAP7_75t_L g93 ( .A(n_3), .Y(n_93) );
INVxp33_ASAP7_75t_L g94 ( .A(n_51), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_38), .Y(n_95) );
INVx1_ASAP7_75t_SL g96 ( .A(n_34), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_22), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_36), .Y(n_98) );
CKINVDCx16_ASAP7_75t_R g99 ( .A(n_10), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_71), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_19), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g102 ( .A(n_8), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_53), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_7), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_9), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_67), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_70), .Y(n_107) );
CKINVDCx14_ASAP7_75t_R g108 ( .A(n_27), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_63), .Y(n_109) );
INVx1_ASAP7_75t_SL g110 ( .A(n_19), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_28), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_72), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_11), .Y(n_113) );
BUFx2_ASAP7_75t_L g114 ( .A(n_88), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_88), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_89), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_99), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_99), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_79), .B(n_0), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_98), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_88), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_89), .Y(n_122) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_93), .B(n_0), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_98), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_91), .Y(n_125) );
BUFx2_ASAP7_75t_L g126 ( .A(n_102), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_102), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_109), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_87), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_81), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_79), .B(n_1), .Y(n_131) );
BUFx2_ASAP7_75t_L g132 ( .A(n_108), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_81), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_92), .B(n_2), .Y(n_134) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_92), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_85), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_130), .Y(n_137) );
INVxp67_ASAP7_75t_L g138 ( .A(n_126), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_114), .B(n_85), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_117), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_124), .Y(n_141) );
INVx5_ASAP7_75t_L g142 ( .A(n_130), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_129), .B(n_94), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_130), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_130), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_132), .B(n_87), .Y(n_146) );
AOI22xp5_ASAP7_75t_L g147 ( .A1(n_123), .A2(n_80), .B1(n_84), .B2(n_112), .Y(n_147) );
INVx4_ASAP7_75t_L g148 ( .A(n_129), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_130), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_124), .Y(n_150) );
CKINVDCx16_ASAP7_75t_R g151 ( .A(n_126), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_124), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_114), .B(n_86), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_130), .Y(n_154) );
AND2x6_ASAP7_75t_L g155 ( .A(n_129), .B(n_86), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_130), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_132), .B(n_87), .Y(n_157) );
INVxp67_ASAP7_75t_L g158 ( .A(n_132), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_124), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_124), .Y(n_160) );
AOI22xp5_ASAP7_75t_L g161 ( .A1(n_123), .A2(n_113), .B1(n_82), .B2(n_110), .Y(n_161) );
AND2x2_ASAP7_75t_L g162 ( .A(n_135), .B(n_87), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_148), .Y(n_163) );
NOR2x1_ASAP7_75t_L g164 ( .A(n_139), .B(n_129), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_162), .B(n_129), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_162), .B(n_135), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_151), .Y(n_167) );
OR2x6_ASAP7_75t_L g168 ( .A(n_158), .B(n_119), .Y(n_168) );
BUFx4_ASAP7_75t_SL g169 ( .A(n_140), .Y(n_169) );
INVxp67_ASAP7_75t_L g170 ( .A(n_157), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_148), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_143), .B(n_133), .Y(n_172) );
BUFx2_ASAP7_75t_L g173 ( .A(n_138), .Y(n_173) );
INVx4_ASAP7_75t_L g174 ( .A(n_155), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_158), .B(n_116), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_148), .Y(n_176) );
AND2x6_ASAP7_75t_SL g177 ( .A(n_157), .B(n_119), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_148), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_L g179 ( .A1(n_139), .A2(n_134), .B(n_131), .C(n_133), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_153), .B(n_122), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_151), .Y(n_181) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_153), .Y(n_182) );
BUFx8_ASAP7_75t_SL g183 ( .A(n_149), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_155), .A2(n_136), .B1(n_134), .B2(n_131), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_155), .B(n_136), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_161), .B(n_97), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_155), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_155), .B(n_115), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_155), .Y(n_189) );
AND2x4_ASAP7_75t_L g190 ( .A(n_146), .B(n_97), .Y(n_190) );
XNOR2xp5_ASAP7_75t_L g191 ( .A(n_147), .B(n_117), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_147), .B(n_118), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_155), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_161), .B(n_83), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_155), .B(n_104), .Y(n_195) );
OAI21x1_ASAP7_75t_SL g196 ( .A1(n_184), .A2(n_95), .B(n_100), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_176), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_165), .B(n_125), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_174), .B(n_128), .Y(n_199) );
O2A1O1Ixp5_ASAP7_75t_L g200 ( .A1(n_172), .A2(n_149), .B(n_121), .C(n_115), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_184), .A2(n_121), .B1(n_120), .B2(n_127), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_182), .B(n_104), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_176), .Y(n_203) );
BUFx2_ASAP7_75t_L g204 ( .A(n_174), .Y(n_204) );
BUFx10_ASAP7_75t_L g205 ( .A(n_189), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_176), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_176), .Y(n_207) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_169), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_166), .B(n_105), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_176), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_176), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_189), .Y(n_212) );
INVx5_ASAP7_75t_L g213 ( .A(n_174), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_163), .A2(n_137), .B(n_144), .Y(n_214) );
BUFx3_ASAP7_75t_L g215 ( .A(n_189), .Y(n_215) );
INVx3_ASAP7_75t_L g216 ( .A(n_174), .Y(n_216) );
INVx2_ASAP7_75t_SL g217 ( .A(n_171), .Y(n_217) );
CKINVDCx16_ASAP7_75t_R g218 ( .A(n_181), .Y(n_218) );
OAI21xp5_ASAP7_75t_L g219 ( .A1(n_179), .A2(n_137), .B(n_144), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_171), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_189), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_171), .Y(n_222) );
NAND2x1p5_ASAP7_75t_L g223 ( .A(n_171), .B(n_95), .Y(n_223) );
INVx4_ASAP7_75t_L g224 ( .A(n_189), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_168), .B(n_118), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_195), .A2(n_120), .B1(n_127), .B2(n_105), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_163), .Y(n_227) );
AO32x2_ASAP7_75t_L g228 ( .A1(n_177), .A2(n_124), .A3(n_120), .B1(n_103), .B2(n_106), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_227), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_203), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_201), .A2(n_168), .B1(n_186), .B2(n_170), .Y(n_231) );
AND2x4_ASAP7_75t_L g232 ( .A(n_213), .B(n_168), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_227), .Y(n_233) );
NAND2xp33_ASAP7_75t_R g234 ( .A(n_225), .B(n_168), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_201), .B(n_168), .Y(n_235) );
CKINVDCx6p67_ASAP7_75t_R g236 ( .A(n_213), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_213), .B(n_165), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_196), .A2(n_186), .B1(n_165), .B2(n_190), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_225), .B(n_166), .Y(n_239) );
INVx2_ASAP7_75t_SL g240 ( .A(n_213), .Y(n_240) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_203), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_227), .B(n_165), .Y(n_242) );
INVx4_ASAP7_75t_L g243 ( .A(n_213), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_203), .Y(n_244) );
AO31x2_ASAP7_75t_L g245 ( .A1(n_209), .A2(n_103), .A3(n_106), .B(n_107), .Y(n_245) );
AND2x2_ASAP7_75t_SL g246 ( .A(n_204), .B(n_189), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_220), .Y(n_247) );
BUFx3_ASAP7_75t_L g248 ( .A(n_213), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_203), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_219), .A2(n_214), .B(n_200), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_196), .A2(n_190), .B1(n_195), .B2(n_164), .Y(n_251) );
OAI222xp33_ASAP7_75t_L g252 ( .A1(n_226), .A2(n_191), .B1(n_101), .B2(n_78), .C1(n_192), .C2(n_167), .Y(n_252) );
OR2x2_ASAP7_75t_L g253 ( .A(n_226), .B(n_173), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_223), .B(n_173), .Y(n_254) );
INVx2_ASAP7_75t_SL g255 ( .A(n_203), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g256 ( .A1(n_231), .A2(n_223), .B1(n_198), .B2(n_202), .Y(n_256) );
INVx4_ASAP7_75t_SL g257 ( .A(n_232), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_231), .A2(n_223), .B1(n_198), .B2(n_191), .Y(n_258) );
OAI221xp5_ASAP7_75t_L g259 ( .A1(n_253), .A2(n_175), .B1(n_180), .B2(n_194), .C(n_208), .Y(n_259) );
OAI221xp5_ASAP7_75t_L g260 ( .A1(n_253), .A2(n_180), .B1(n_164), .B2(n_219), .C(n_199), .Y(n_260) );
OAI22xp33_ASAP7_75t_L g261 ( .A1(n_253), .A2(n_218), .B1(n_198), .B2(n_204), .Y(n_261) );
OAI211xp5_ASAP7_75t_L g262 ( .A1(n_238), .A2(n_90), .B(n_111), .C(n_100), .Y(n_262) );
OAI21x1_ASAP7_75t_L g263 ( .A1(n_250), .A2(n_206), .B(n_197), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_235), .A2(n_198), .B1(n_190), .B2(n_218), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_239), .B(n_177), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_235), .A2(n_190), .B1(n_222), .B2(n_220), .Y(n_266) );
INVxp67_ASAP7_75t_L g267 ( .A(n_254), .Y(n_267) );
AOI22xp5_ASAP7_75t_L g268 ( .A1(n_234), .A2(n_217), .B1(n_216), .B2(n_222), .Y(n_268) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_238), .A2(n_207), .B1(n_210), .B2(n_211), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_229), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_229), .Y(n_271) );
AOI221xp5_ASAP7_75t_L g272 ( .A1(n_252), .A2(n_185), .B1(n_188), .B2(n_207), .C(n_210), .Y(n_272) );
OAI22xp5_ASAP7_75t_L g273 ( .A1(n_235), .A2(n_251), .B1(n_229), .B2(n_233), .Y(n_273) );
AO21x2_ASAP7_75t_L g274 ( .A1(n_250), .A2(n_197), .B(n_188), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_233), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g276 ( .A1(n_239), .A2(n_217), .B1(n_216), .B2(n_206), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_233), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_257), .B(n_232), .Y(n_278) );
OAI21x1_ASAP7_75t_L g279 ( .A1(n_263), .A2(n_244), .B(n_230), .Y(n_279) );
INVx8_ASAP7_75t_L g280 ( .A(n_257), .Y(n_280) );
INVx4_ASAP7_75t_L g281 ( .A(n_257), .Y(n_281) );
OAI31xp33_ASAP7_75t_L g282 ( .A1(n_258), .A2(n_252), .A3(n_254), .B(n_239), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_263), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_275), .Y(n_284) );
XNOR2xp5_ASAP7_75t_L g285 ( .A(n_264), .B(n_254), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_256), .A2(n_251), .B1(n_246), .B2(n_232), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_261), .A2(n_232), .B1(n_237), .B2(n_242), .Y(n_287) );
OAI22xp5_ASAP7_75t_L g288 ( .A1(n_272), .A2(n_232), .B1(n_246), .B2(n_236), .Y(n_288) );
OAI33xp33_ASAP7_75t_L g289 ( .A1(n_265), .A2(n_107), .A3(n_111), .B1(n_247), .B2(n_145), .B3(n_154), .Y(n_289) );
A2O1A1Ixp33_ASAP7_75t_L g290 ( .A1(n_260), .A2(n_232), .B(n_237), .C(n_240), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_267), .A2(n_246), .B1(n_236), .B2(n_234), .Y(n_291) );
AOI31xp33_ASAP7_75t_SL g292 ( .A1(n_257), .A2(n_228), .A3(n_236), .B(n_5), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_275), .B(n_242), .Y(n_293) );
AOI22xp33_ASAP7_75t_SL g294 ( .A1(n_273), .A2(n_246), .B1(n_243), .B2(n_248), .Y(n_294) );
AND2x4_ASAP7_75t_L g295 ( .A(n_277), .B(n_230), .Y(n_295) );
OAI33xp33_ASAP7_75t_L g296 ( .A1(n_277), .A2(n_247), .A3(n_154), .B1(n_145), .B2(n_156), .B3(n_228), .Y(n_296) );
OAI211xp5_ASAP7_75t_L g297 ( .A1(n_259), .A2(n_242), .B(n_247), .C(n_96), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_274), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_270), .Y(n_299) );
BUFx2_ASAP7_75t_L g300 ( .A(n_281), .Y(n_300) );
OAI33xp33_ASAP7_75t_L g301 ( .A1(n_299), .A2(n_269), .A3(n_271), .B1(n_156), .B2(n_6), .B3(n_7), .Y(n_301) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_284), .Y(n_302) );
NAND3xp33_ASAP7_75t_L g303 ( .A(n_282), .B(n_262), .C(n_124), .Y(n_303) );
INVx2_ASAP7_75t_SL g304 ( .A(n_280), .Y(n_304) );
NAND2x1p5_ASAP7_75t_L g305 ( .A(n_281), .B(n_243), .Y(n_305) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_284), .Y(n_306) );
AOI211xp5_ASAP7_75t_L g307 ( .A1(n_292), .A2(n_237), .B(n_268), .C(n_240), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_284), .B(n_274), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_299), .B(n_245), .Y(n_309) );
OAI221xp5_ASAP7_75t_SL g310 ( .A1(n_282), .A2(n_266), .B1(n_276), .B2(n_236), .C(n_228), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_293), .B(n_245), .Y(n_311) );
OR2x2_ASAP7_75t_L g312 ( .A(n_286), .B(n_245), .Y(n_312) );
AOI221xp5_ASAP7_75t_L g313 ( .A1(n_289), .A2(n_237), .B1(n_274), .B2(n_149), .C(n_141), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_283), .Y(n_314) );
AOI32xp33_ASAP7_75t_L g315 ( .A1(n_286), .A2(n_237), .A3(n_243), .B1(n_248), .B2(n_240), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_295), .Y(n_316) );
INVx1_ASAP7_75t_SL g317 ( .A(n_278), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_283), .Y(n_318) );
AOI33xp33_ASAP7_75t_L g319 ( .A1(n_287), .A2(n_237), .A3(n_150), .B1(n_152), .B2(n_159), .B3(n_160), .Y(n_319) );
NAND3xp33_ASAP7_75t_L g320 ( .A(n_297), .B(n_243), .C(n_249), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_295), .B(n_228), .Y(n_321) );
OR2x2_ASAP7_75t_L g322 ( .A(n_298), .B(n_245), .Y(n_322) );
INVx1_ASAP7_75t_SL g323 ( .A(n_278), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_298), .B(n_245), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_281), .B(n_230), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_298), .B(n_245), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_295), .B(n_228), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_295), .B(n_228), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_283), .Y(n_329) );
NOR2xp33_ASAP7_75t_R g330 ( .A(n_304), .B(n_280), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_302), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_306), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_311), .B(n_293), .Y(n_333) );
NAND2xp33_ASAP7_75t_R g334 ( .A(n_300), .B(n_278), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_311), .B(n_278), .Y(n_335) );
OR2x6_ASAP7_75t_L g336 ( .A(n_300), .B(n_280), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_316), .B(n_285), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_309), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_309), .B(n_245), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_321), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_321), .Y(n_341) );
AND2x2_ASAP7_75t_SL g342 ( .A(n_312), .B(n_281), .Y(n_342) );
AOI31xp67_ASAP7_75t_L g343 ( .A1(n_314), .A2(n_292), .A3(n_230), .B(n_249), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_317), .B(n_285), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_310), .B(n_288), .Y(n_345) );
AOI21xp33_ASAP7_75t_L g346 ( .A1(n_312), .A2(n_291), .B(n_280), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_322), .B(n_280), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_327), .B(n_245), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_327), .B(n_245), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_322), .B(n_290), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_317), .B(n_294), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_324), .B(n_279), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_301), .B(n_296), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_323), .B(n_2), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_324), .Y(n_355) );
NAND2xp33_ASAP7_75t_SL g356 ( .A(n_304), .B(n_243), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_303), .B(n_3), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_328), .B(n_308), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_328), .B(n_5), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_308), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_326), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_323), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_326), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_307), .B(n_6), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_314), .B(n_279), .Y(n_365) );
INVx3_ASAP7_75t_SL g366 ( .A(n_325), .Y(n_366) );
NAND2xp33_ASAP7_75t_SL g367 ( .A(n_319), .B(n_243), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_314), .Y(n_368) );
NAND2xp33_ASAP7_75t_SL g369 ( .A(n_315), .B(n_241), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_303), .B(n_9), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_318), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_307), .B(n_11), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_318), .B(n_12), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_325), .B(n_12), .Y(n_374) );
OAI21xp33_ASAP7_75t_L g375 ( .A1(n_345), .A2(n_315), .B(n_320), .Y(n_375) );
OAI221xp5_ASAP7_75t_L g376 ( .A1(n_372), .A2(n_320), .B1(n_305), .B2(n_313), .C(n_318), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_338), .B(n_329), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_364), .B(n_13), .Y(n_378) );
INVxp67_ASAP7_75t_SL g379 ( .A(n_334), .Y(n_379) );
AOI211xp5_ASAP7_75t_SL g380 ( .A1(n_345), .A2(n_325), .B(n_329), .C(n_305), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_371), .Y(n_381) );
XNOR2x2_ASAP7_75t_L g382 ( .A(n_339), .B(n_329), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_371), .Y(n_383) );
NAND3xp33_ASAP7_75t_L g384 ( .A(n_353), .B(n_325), .C(n_141), .Y(n_384) );
O2A1O1Ixp5_ASAP7_75t_L g385 ( .A1(n_356), .A2(n_160), .B(n_150), .C(n_152), .Y(n_385) );
OAI21xp5_ASAP7_75t_L g386 ( .A1(n_357), .A2(n_305), .B(n_255), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_360), .B(n_244), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_334), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_340), .B(n_244), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_336), .A2(n_248), .B1(n_255), .B2(n_249), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_341), .B(n_244), .Y(n_391) );
OAI21xp33_ASAP7_75t_SL g392 ( .A1(n_336), .A2(n_255), .B(n_249), .Y(n_392) );
AOI32xp33_ASAP7_75t_L g393 ( .A1(n_369), .A2(n_248), .A3(n_14), .B1(n_15), .B2(n_17), .Y(n_393) );
AO21x1_ASAP7_75t_L g394 ( .A1(n_356), .A2(n_13), .B(n_14), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_358), .B(n_15), .Y(n_395) );
INVx1_ASAP7_75t_SL g396 ( .A(n_366), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_336), .A2(n_255), .B1(n_241), .B2(n_224), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_357), .A2(n_241), .B1(n_197), .B2(n_206), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_331), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_370), .A2(n_241), .B1(n_206), .B2(n_203), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_342), .B(n_17), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_361), .B(n_18), .Y(n_402) );
INVxp67_ASAP7_75t_L g403 ( .A(n_367), .Y(n_403) );
O2A1O1Ixp33_ASAP7_75t_L g404 ( .A1(n_370), .A2(n_141), .B(n_150), .C(n_152), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_342), .A2(n_241), .B1(n_224), .B2(n_211), .Y(n_405) );
OAI211xp5_ASAP7_75t_L g406 ( .A1(n_330), .A2(n_159), .B(n_160), .C(n_224), .Y(n_406) );
INVxp67_ASAP7_75t_L g407 ( .A(n_367), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_332), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_363), .Y(n_409) );
INVxp67_ASAP7_75t_L g410 ( .A(n_374), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_366), .A2(n_241), .B1(n_224), .B2(n_211), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_347), .A2(n_241), .B1(n_211), .B2(n_216), .Y(n_412) );
OAI322xp33_ASAP7_75t_L g413 ( .A1(n_350), .A2(n_18), .A3(n_20), .B1(n_21), .B2(n_22), .C1(n_23), .C2(n_24), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_335), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_355), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_352), .B(n_20), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_333), .B(n_21), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_351), .B(n_23), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_348), .B(n_24), .Y(n_419) );
NAND3xp33_ASAP7_75t_L g420 ( .A(n_353), .B(n_159), .C(n_241), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_373), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_368), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_354), .Y(n_423) );
OAI21xp5_ASAP7_75t_SL g424 ( .A1(n_346), .A2(n_25), .B(n_241), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_365), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_349), .B(n_25), .Y(n_426) );
NAND2xp5_ASAP7_75t_SL g427 ( .A(n_369), .B(n_211), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_399), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_425), .B(n_362), .Y(n_429) );
INVxp33_ASAP7_75t_L g430 ( .A(n_388), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_414), .B(n_344), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_415), .B(n_359), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_379), .B(n_409), .Y(n_433) );
INVxp67_ASAP7_75t_L g434 ( .A(n_418), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_381), .B(n_337), .Y(n_435) );
NOR2x1_ASAP7_75t_L g436 ( .A(n_401), .B(n_330), .Y(n_436) );
AND4x1_ASAP7_75t_L g437 ( .A(n_380), .B(n_343), .C(n_183), .D(n_31), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_408), .Y(n_438) );
NOR3xp33_ASAP7_75t_L g439 ( .A(n_413), .B(n_149), .C(n_216), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_381), .B(n_26), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_426), .B(n_30), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_383), .B(n_32), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_383), .B(n_33), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_401), .A2(n_211), .B1(n_215), .B2(n_212), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_410), .B(n_35), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_426), .B(n_37), .Y(n_446) );
NOR3xp33_ASAP7_75t_SL g447 ( .A(n_375), .B(n_193), .C(n_187), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_423), .B(n_39), .Y(n_448) );
NOR2xp33_ASAP7_75t_R g449 ( .A(n_396), .B(n_40), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_418), .B(n_41), .Y(n_450) );
NAND2xp33_ASAP7_75t_SL g451 ( .A(n_427), .B(n_221), .Y(n_451) );
XOR2x2_ASAP7_75t_L g452 ( .A(n_378), .B(n_43), .Y(n_452) );
INVx1_ASAP7_75t_SL g453 ( .A(n_416), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_422), .B(n_45), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_416), .B(n_46), .Y(n_455) );
NAND2xp33_ASAP7_75t_SL g456 ( .A(n_427), .B(n_221), .Y(n_456) );
NOR4xp25_ASAP7_75t_SL g457 ( .A(n_424), .B(n_47), .C(n_48), .D(n_49), .Y(n_457) );
NAND3xp33_ASAP7_75t_L g458 ( .A(n_393), .B(n_142), .C(n_212), .Y(n_458) );
INVxp67_ASAP7_75t_L g459 ( .A(n_417), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_378), .A2(n_215), .B1(n_221), .B2(n_212), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_421), .B(n_50), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_387), .B(n_52), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_395), .B(n_54), .Y(n_463) );
NOR3xp33_ASAP7_75t_L g464 ( .A(n_384), .B(n_193), .C(n_187), .Y(n_464) );
AND2x4_ASAP7_75t_L g465 ( .A(n_377), .B(n_57), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_387), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_395), .B(n_59), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_402), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_417), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_389), .B(n_60), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_419), .B(n_61), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_389), .B(n_62), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_449), .Y(n_473) );
NOR3xp33_ASAP7_75t_L g474 ( .A(n_458), .B(n_407), .C(n_403), .Y(n_474) );
INVxp67_ASAP7_75t_L g475 ( .A(n_468), .Y(n_475) );
OAI211xp5_ASAP7_75t_L g476 ( .A1(n_436), .A2(n_392), .B(n_406), .C(n_386), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_435), .B(n_433), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_435), .B(n_391), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_451), .B(n_405), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_451), .A2(n_394), .B(n_385), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_433), .B(n_391), .Y(n_481) );
NOR2x1_ASAP7_75t_L g482 ( .A(n_453), .B(n_420), .Y(n_482) );
XNOR2x2_ASAP7_75t_L g483 ( .A(n_452), .B(n_382), .Y(n_483) );
OAI21xp33_ASAP7_75t_SL g484 ( .A1(n_430), .A2(n_382), .B(n_400), .Y(n_484) );
AOI31xp33_ASAP7_75t_L g485 ( .A1(n_430), .A2(n_390), .A3(n_397), .B(n_411), .Y(n_485) );
INVxp33_ASAP7_75t_L g486 ( .A(n_452), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_469), .B(n_376), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_431), .B(n_398), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_431), .B(n_412), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_466), .B(n_64), .Y(n_490) );
INVxp67_ASAP7_75t_SL g491 ( .A(n_434), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_459), .A2(n_404), .B1(n_215), .B2(n_221), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_432), .A2(n_142), .B1(n_212), .B2(n_221), .Y(n_493) );
OAI22xp33_ASAP7_75t_L g494 ( .A1(n_460), .A2(n_221), .B1(n_212), .B2(n_142), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_428), .Y(n_495) );
XOR2xp5_ASAP7_75t_L g496 ( .A(n_432), .B(n_65), .Y(n_496) );
INVx1_ASAP7_75t_SL g497 ( .A(n_429), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_429), .B(n_66), .Y(n_498) );
AOI211x1_ASAP7_75t_SL g499 ( .A1(n_463), .A2(n_69), .B(n_73), .C(n_74), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_438), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_450), .A2(n_212), .B1(n_205), .B2(n_142), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_466), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_495), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_500), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_475), .Y(n_505) );
INVx1_ASAP7_75t_SL g506 ( .A(n_473), .Y(n_506) );
AO22x2_ASAP7_75t_L g507 ( .A1(n_491), .A2(n_444), .B1(n_465), .B2(n_454), .Y(n_507) );
INVxp67_ASAP7_75t_L g508 ( .A(n_487), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_474), .B(n_454), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_478), .Y(n_510) );
NOR2xp33_ASAP7_75t_R g511 ( .A(n_473), .B(n_456), .Y(n_511) );
NOR2xp33_ASAP7_75t_R g512 ( .A(n_498), .B(n_456), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_483), .A2(n_448), .B1(n_445), .B2(n_446), .Y(n_513) );
OAI211xp5_ASAP7_75t_L g514 ( .A1(n_484), .A2(n_467), .B(n_441), .C(n_457), .Y(n_514) );
AOI32xp33_ASAP7_75t_L g515 ( .A1(n_486), .A2(n_462), .A3(n_470), .B1(n_464), .B2(n_455), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_486), .A2(n_470), .B1(n_462), .B2(n_465), .Y(n_516) );
AOI21xp33_ASAP7_75t_SL g517 ( .A1(n_485), .A2(n_465), .B(n_461), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_488), .A2(n_471), .B1(n_447), .B2(n_472), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_497), .B(n_437), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_481), .B(n_443), .Y(n_520) );
AOI222xp33_ASAP7_75t_L g521 ( .A1(n_483), .A2(n_443), .B1(n_442), .B2(n_440), .C1(n_439), .C2(n_142), .Y(n_521) );
OAI321xp33_ASAP7_75t_L g522 ( .A1(n_476), .A2(n_440), .A3(n_442), .B1(n_76), .B2(n_77), .C(n_178), .Y(n_522) );
NOR4xp25_ASAP7_75t_L g523 ( .A(n_479), .B(n_178), .C(n_142), .D(n_205), .Y(n_523) );
NOR3xp33_ASAP7_75t_L g524 ( .A(n_479), .B(n_205), .C(n_142), .Y(n_524) );
OAI211xp5_ASAP7_75t_SL g525 ( .A1(n_489), .A2(n_205), .B(n_482), .C(n_499), .Y(n_525) );
NOR4xp25_ASAP7_75t_L g526 ( .A(n_477), .B(n_493), .C(n_502), .D(n_490), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_480), .A2(n_496), .B(n_481), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_481), .A2(n_502), .B1(n_492), .B2(n_501), .Y(n_528) );
OAI322xp33_ASAP7_75t_L g529 ( .A1(n_508), .A2(n_527), .A3(n_517), .B1(n_505), .B2(n_506), .C1(n_509), .C2(n_528), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_507), .B(n_526), .Y(n_530) );
OAI211xp5_ASAP7_75t_SL g531 ( .A1(n_513), .A2(n_521), .B(n_515), .C(n_514), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_510), .B(n_503), .Y(n_532) );
OAI221xp5_ASAP7_75t_R g533 ( .A1(n_518), .A2(n_524), .B1(n_507), .B2(n_516), .C(n_512), .Y(n_533) );
NAND4xp25_ASAP7_75t_L g534 ( .A(n_531), .B(n_519), .C(n_525), .D(n_493), .Y(n_534) );
XNOR2xp5_ASAP7_75t_L g535 ( .A(n_530), .B(n_507), .Y(n_535) );
NAND4xp25_ASAP7_75t_L g536 ( .A(n_533), .B(n_522), .C(n_511), .D(n_523), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_534), .Y(n_537) );
AND2x4_ASAP7_75t_L g538 ( .A(n_535), .B(n_532), .Y(n_538) );
INVx2_ASAP7_75t_SL g539 ( .A(n_537), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_539), .A2(n_538), .B1(n_536), .B2(n_529), .Y(n_540) );
AOI221xp5_ASAP7_75t_L g541 ( .A1(n_540), .A2(n_538), .B1(n_504), .B2(n_520), .C(n_494), .Y(n_541) );
endmodule