module fake_jpeg_860_n_544 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_544);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_544;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_19;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx10_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_7),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_45),
.B(n_55),
.Y(n_105)
);

BUFx4f_ASAP7_75t_SL g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx4f_ASAP7_75t_SL g108 ( 
.A(n_46),
.Y(n_108)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_50),
.Y(n_127)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_25),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_39),
.B(n_7),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_58),
.B(n_62),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_18),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_64),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_23),
.B(n_0),
.Y(n_65)
);

AND2x2_ASAP7_75t_SL g138 ( 
.A(n_65),
.B(n_20),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_66),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_69),
.Y(n_130)
);

INVx6_ASAP7_75t_SL g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx16f_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_71),
.Y(n_143)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_38),
.B(n_8),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_73),
.B(n_76),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_74),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_36),
.B(n_8),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_25),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_77),
.B(n_79),
.Y(n_140)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_25),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_28),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_80),
.B(n_82),
.Y(n_146)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_28),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_83),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

BUFx24_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_44),
.B(n_8),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_87),
.B(n_6),
.Y(n_152)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

BUFx8_ASAP7_75t_L g89 ( 
.A(n_17),
.Y(n_89)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_89),
.Y(n_157)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_21),
.Y(n_90)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_15),
.Y(n_91)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

BUFx24_ASAP7_75t_L g92 ( 
.A(n_17),
.Y(n_92)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_70),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_99),
.B(n_104),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_85),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_84),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_117),
.B(n_135),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_65),
.A2(n_44),
.B1(n_43),
.B2(n_41),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_119),
.B(n_155),
.C(n_27),
.Y(n_173)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_123),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_52),
.A2(n_21),
.B1(n_20),
.B2(n_37),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_131),
.A2(n_153),
.B1(n_89),
.B2(n_92),
.Y(n_169)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_56),
.Y(n_134)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_86),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_63),
.Y(n_136)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_138),
.Y(n_166)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_L g147 ( 
.A1(n_96),
.A2(n_34),
.B1(n_28),
.B2(n_41),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_147),
.A2(n_43),
.B1(n_32),
.B2(n_33),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_152),
.B(n_12),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_89),
.A2(n_20),
.B1(n_33),
.B2(n_32),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_65),
.B(n_20),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_91),
.Y(n_156)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_90),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_46),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_160),
.A2(n_168),
.B1(n_133),
.B2(n_92),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_64),
.B1(n_61),
.B2(n_59),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_161),
.A2(n_196),
.B1(n_169),
.B2(n_178),
.Y(n_220)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_162),
.B(n_163),
.Y(n_211)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_165),
.Y(n_226)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_102),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_167),
.B(n_191),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_131),
.A2(n_74),
.B1(n_66),
.B2(n_67),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_169),
.A2(n_154),
.B(n_17),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_136),
.A2(n_94),
.B1(n_93),
.B2(n_88),
.Y(n_171)
);

BUFx24_ASAP7_75t_L g219 ( 
.A(n_171),
.Y(n_219)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_172),
.Y(n_209)
);

NAND3xp33_ASAP7_75t_L g239 ( 
.A(n_173),
.B(n_198),
.C(n_204),
.Y(n_239)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_101),
.Y(n_175)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_121),
.A2(n_20),
.B1(n_95),
.B2(n_60),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_118),
.Y(n_179)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_179),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_103),
.B(n_81),
.C(n_50),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_193),
.C(n_199),
.Y(n_207)
);

CKINVDCx12_ASAP7_75t_R g181 ( 
.A(n_129),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_181),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_118),
.Y(n_182)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_182),
.Y(n_237)
);

INVx3_ASAP7_75t_SL g183 ( 
.A(n_111),
.Y(n_183)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_109),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_185),
.Y(n_236)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_139),
.Y(n_186)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_186),
.Y(n_229)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_115),
.Y(n_187)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_115),
.Y(n_188)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_188),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_141),
.B(n_69),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_189),
.B(n_200),
.Y(n_210)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_127),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_194),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_105),
.B(n_49),
.C(n_48),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_126),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_140),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_197),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_L g196 ( 
.A1(n_153),
.A2(n_75),
.B1(n_54),
.B2(n_34),
.Y(n_196)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_113),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_106),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_203),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_132),
.B(n_57),
.C(n_47),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_130),
.B(n_46),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_202),
.B(n_13),
.Y(n_222)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_107),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_123),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_205),
.Y(n_235)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_129),
.Y(n_205)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_139),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_206),
.B(n_142),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_161),
.A2(n_138),
.B1(n_155),
.B2(n_125),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_217),
.A2(n_220),
.B1(n_223),
.B2(n_113),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_218),
.A2(n_171),
.B1(n_133),
.B2(n_122),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_9),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_168),
.A2(n_120),
.B1(n_150),
.B2(n_144),
.Y(n_223)
);

A2O1A1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_166),
.A2(n_112),
.B(n_98),
.C(n_151),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_227),
.B(n_115),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_196),
.A2(n_108),
.B(n_151),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

OAI21xp33_ASAP7_75t_L g231 ( 
.A1(n_190),
.A2(n_151),
.B(n_108),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_231),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_238),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_97),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_201),
.B(n_124),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_241),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_177),
.B(n_100),
.Y(n_241)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_242),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_243),
.A2(n_261),
.B1(n_263),
.B2(n_217),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_244),
.Y(n_297)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_213),
.Y(n_247)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_247),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_248),
.B(n_254),
.Y(n_293)
);

MAJx2_ASAP7_75t_L g250 ( 
.A(n_207),
.B(n_176),
.C(n_159),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_250),
.B(n_235),
.C(n_215),
.Y(n_301)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_208),
.Y(n_251)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_251),
.Y(n_280)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_212),
.Y(n_252)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_252),
.Y(n_300)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_212),
.Y(n_253)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_253),
.Y(n_306)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_256),
.Y(n_286)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_232),
.Y(n_256)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_228),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_257),
.B(n_260),
.Y(n_295)
);

INVx13_ASAP7_75t_L g258 ( 
.A(n_216),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_258),
.Y(n_298)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_232),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_203),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_264),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_220),
.A2(n_125),
.B1(n_142),
.B2(n_148),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_226),
.B(n_170),
.Y(n_264)
);

OA21x2_ASAP7_75t_L g265 ( 
.A1(n_228),
.A2(n_227),
.B(n_217),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_265),
.A2(n_219),
.B(n_241),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_170),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_272),
.Y(n_279)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_224),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_269),
.Y(n_302)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_224),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_211),
.B(n_205),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_270),
.B(n_274),
.Y(n_284)
);

OA22x2_ASAP7_75t_SL g271 ( 
.A1(n_227),
.A2(n_110),
.B1(n_120),
.B2(n_78),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_271),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_210),
.B(n_207),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_210),
.B(n_116),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_208),
.Y(n_292)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_221),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_244),
.A2(n_214),
.B(n_238),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_276),
.A2(n_283),
.B(n_288),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_243),
.A2(n_218),
.B1(n_219),
.B2(n_221),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_277),
.A2(n_291),
.B1(n_307),
.B2(n_271),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_278),
.A2(n_281),
.B1(n_290),
.B2(n_271),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_265),
.A2(n_239),
.B1(n_207),
.B2(n_219),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_245),
.A2(n_219),
.B(n_231),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_259),
.B(n_222),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_287),
.B(n_248),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_250),
.B(n_225),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_289),
.B(n_303),
.C(n_267),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_265),
.A2(n_219),
.B1(n_242),
.B2(n_229),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_272),
.A2(n_225),
.B1(n_229),
.B2(n_209),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_292),
.B(n_230),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_266),
.A2(n_235),
.B(n_233),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_294),
.A2(n_304),
.B(n_188),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_246),
.B(n_211),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_305),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_265),
.A2(n_213),
.B1(n_209),
.B2(n_237),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_299),
.A2(n_255),
.B1(n_263),
.B2(n_262),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_260),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_250),
.B(n_234),
.C(n_233),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_257),
.A2(n_234),
.B(n_215),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_246),
.B(n_213),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_255),
.A2(n_257),
.B1(n_259),
.B2(n_256),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_300),
.Y(n_308)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_308),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_309),
.A2(n_315),
.B1(n_327),
.B2(n_335),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_310),
.B(n_289),
.Y(n_343)
);

OAI21xp33_ASAP7_75t_L g312 ( 
.A1(n_283),
.A2(n_273),
.B(n_264),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_312),
.B(n_322),
.Y(n_351)
);

OAI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_313),
.A2(n_280),
.B1(n_298),
.B2(n_293),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_296),
.B(n_274),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_314),
.B(n_320),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_316),
.B(n_289),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_269),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_317),
.B(n_328),
.Y(n_349)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_300),
.Y(n_318)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_318),
.Y(n_344)
);

AO22x1_ASAP7_75t_L g319 ( 
.A1(n_307),
.A2(n_271),
.B1(n_268),
.B2(n_261),
.Y(n_319)
);

A2O1A1Ixp33_ASAP7_75t_SL g363 ( 
.A1(n_319),
.A2(n_313),
.B(n_329),
.C(n_332),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_302),
.B(n_284),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_306),
.Y(n_321)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_321),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_284),
.B(n_208),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_306),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_323),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_324),
.B(n_330),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_290),
.A2(n_281),
.B1(n_288),
.B2(n_277),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_325),
.A2(n_282),
.B1(n_295),
.B2(n_299),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_297),
.A2(n_249),
.B1(n_253),
.B2(n_252),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_326),
.B(n_336),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_278),
.A2(n_209),
.B1(n_247),
.B2(n_237),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_286),
.B(n_251),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_305),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_329),
.B(n_331),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_287),
.B(n_258),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_275),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_275),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_332),
.B(n_333),
.Y(n_373)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_285),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_288),
.A2(n_237),
.B1(n_230),
.B2(n_182),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_286),
.A2(n_230),
.B1(n_175),
.B2(n_186),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_285),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_337),
.B(n_338),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_304),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_339),
.A2(n_328),
.B(n_326),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_304),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_340),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_341),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_343),
.B(n_358),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_345),
.B(n_311),
.C(n_339),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_310),
.B(n_301),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_346),
.B(n_354),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_319),
.A2(n_295),
.B1(n_291),
.B2(n_282),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_348),
.B(n_362),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_350),
.A2(n_361),
.B1(n_365),
.B2(n_366),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_316),
.B(n_301),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_330),
.B(n_279),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_355),
.B(n_363),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_317),
.B(n_279),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_325),
.A2(n_299),
.B1(n_276),
.B2(n_292),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_319),
.A2(n_340),
.B1(n_338),
.B2(n_335),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_331),
.B(n_303),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_364),
.B(n_97),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_334),
.A2(n_294),
.B1(n_303),
.B2(n_280),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_324),
.B(n_298),
.Y(n_368)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_368),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_334),
.A2(n_293),
.B(n_184),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_369),
.A2(n_374),
.B(n_111),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_311),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_372),
.B(n_27),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_349),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_377),
.B(n_382),
.Y(n_422)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_349),
.Y(n_379)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_379),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_381),
.B(n_383),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_360),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_345),
.B(n_341),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_370),
.Y(n_384)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_384),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_348),
.A2(n_315),
.B1(n_308),
.B2(n_323),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_385),
.A2(n_352),
.B1(n_363),
.B2(n_356),
.Y(n_407)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_370),
.Y(n_386)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_386),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_350),
.A2(n_327),
.B1(n_318),
.B2(n_321),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_387),
.A2(n_390),
.B1(n_397),
.B2(n_403),
.Y(n_417)
);

FAx1_ASAP7_75t_SL g388 ( 
.A(n_358),
.B(n_258),
.CI(n_337),
.CON(n_388),
.SN(n_388)
);

NOR3xp33_ASAP7_75t_SL g431 ( 
.A(n_388),
.B(n_205),
.C(n_187),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_354),
.B(n_346),
.C(n_343),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_389),
.B(n_391),
.C(n_396),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_353),
.A2(n_333),
.B1(n_172),
.B2(n_206),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_164),
.C(n_236),
.Y(n_391)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_392),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_360),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_395),
.B(n_15),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_365),
.B(n_164),
.C(n_116),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_361),
.A2(n_359),
.B1(n_371),
.B2(n_374),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_347),
.B(n_197),
.Y(n_398)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_398),
.Y(n_429)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_373),
.Y(n_399)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_399),
.Y(n_430)
);

AND2x2_ASAP7_75t_SL g400 ( 
.A(n_356),
.B(n_97),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_400),
.Y(n_428)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_373),
.Y(n_401)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_401),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_402),
.A2(n_352),
.B(n_356),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_359),
.A2(n_352),
.B1(n_367),
.B2(n_363),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_342),
.Y(n_404)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_404),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_405),
.B(n_406),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_351),
.B(n_183),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_407),
.A2(n_402),
.B1(n_378),
.B2(n_380),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_394),
.B(n_369),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_408),
.B(n_375),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_409),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_400),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_410),
.B(n_412),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_400),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_394),
.B(n_362),
.C(n_357),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_414),
.B(n_420),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_393),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_389),
.B(n_344),
.C(n_363),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_421),
.B(n_425),
.C(n_405),
.Y(n_445)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_424),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_391),
.B(n_114),
.C(n_179),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_387),
.B(n_148),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_426),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_403),
.B(n_110),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_427),
.Y(n_452)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_431),
.Y(n_439)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_385),
.Y(n_433)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_433),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_417),
.A2(n_433),
.B1(n_422),
.B2(n_427),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_437),
.A2(n_457),
.B1(n_428),
.B2(n_409),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_438),
.B(n_451),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_415),
.B(n_381),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_440),
.B(n_445),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_429),
.B(n_376),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_441),
.B(n_443),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_430),
.A2(n_380),
.B1(n_397),
.B2(n_378),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_423),
.B(n_383),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_444),
.B(n_459),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_432),
.A2(n_378),
.B1(n_388),
.B2(n_406),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_SL g473 ( 
.A1(n_447),
.A2(n_449),
.B1(n_122),
.B2(n_83),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_407),
.A2(n_388),
.B1(n_396),
.B2(n_375),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_450),
.B(n_428),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_415),
.B(n_51),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_421),
.B(n_51),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_453),
.B(n_418),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_414),
.B(n_150),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_454),
.B(n_456),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_413),
.B(n_408),
.C(n_434),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_455),
.B(n_434),
.C(n_425),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_413),
.B(n_144),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_427),
.A2(n_114),
.B1(n_53),
.B2(n_71),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_416),
.B(n_149),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_436),
.Y(n_460)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_460),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_461),
.B(n_479),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_462),
.A2(n_471),
.B1(n_17),
.B2(n_29),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_465),
.B(n_473),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_446),
.A2(n_431),
.B(n_419),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_466),
.A2(n_472),
.B(n_10),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_440),
.B(n_456),
.C(n_455),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_469),
.B(n_475),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_470),
.B(n_477),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_437),
.A2(n_426),
.B1(n_411),
.B2(n_34),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_458),
.A2(n_426),
.B(n_411),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_445),
.B(n_78),
.C(n_19),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_454),
.B(n_19),
.C(n_30),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_476),
.B(n_478),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_453),
.B(n_19),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_446),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_442),
.B(n_19),
.C(n_30),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_451),
.C(n_448),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_480),
.B(n_481),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_463),
.B(n_448),
.C(n_452),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_469),
.B(n_461),
.C(n_470),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_482),
.B(n_484),
.Y(n_500)
);

NOR2x1_ASAP7_75t_L g483 ( 
.A(n_465),
.B(n_466),
.Y(n_483)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_483),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_474),
.B(n_435),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_468),
.A2(n_439),
.B(n_450),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_486),
.A2(n_492),
.B(n_475),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_471),
.A2(n_457),
.B1(n_19),
.B2(n_29),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_489),
.A2(n_496),
.B1(n_17),
.B2(n_479),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_464),
.B(n_19),
.C(n_30),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_490),
.B(n_0),
.C(n_1),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_491),
.B(n_477),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_467),
.B(n_9),
.Y(n_492)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_497),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_498),
.B(n_1),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_501),
.B(n_502),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_482),
.B(n_464),
.C(n_476),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_487),
.A2(n_29),
.B1(n_6),
.B2(n_12),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_503),
.B(n_507),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_483),
.A2(n_14),
.B(n_13),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_504),
.B(n_506),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_485),
.B(n_14),
.Y(n_506)
);

NOR3xp33_ASAP7_75t_SL g507 ( 
.A(n_495),
.B(n_14),
.C(n_13),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_508),
.B(n_509),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_481),
.B(n_6),
.Y(n_509)
);

BUFx24_ASAP7_75t_SL g510 ( 
.A(n_494),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_510),
.B(n_4),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_491),
.A2(n_13),
.B1(n_2),
.B2(n_3),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_511),
.A2(n_480),
.B1(n_488),
.B2(n_490),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_493),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_512),
.B(n_508),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_513),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_499),
.B(n_505),
.C(n_506),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_517),
.B(n_519),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_498),
.B(n_495),
.C(n_2),
.Y(n_519)
);

NOR2x1_ASAP7_75t_L g520 ( 
.A(n_507),
.B(n_1),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_520),
.A2(n_1),
.B(n_3),
.Y(n_525)
);

INVxp33_ASAP7_75t_L g526 ( 
.A(n_522),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_523),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_524),
.A2(n_531),
.B(n_518),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_525),
.B(n_3),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_514),
.B(n_4),
.C(n_1),
.Y(n_530)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_530),
.B(n_518),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_512),
.A2(n_3),
.B(n_515),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_532),
.Y(n_539)
);

INVxp33_ASAP7_75t_L g538 ( 
.A(n_533),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_534),
.A2(n_535),
.B(n_536),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_528),
.B(n_516),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_527),
.A2(n_521),
.B(n_3),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_538),
.B(n_524),
.C(n_529),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_540),
.B(n_541),
.C(n_537),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_539),
.B(n_526),
.Y(n_541)
);

BUFx24_ASAP7_75t_SL g543 ( 
.A(n_542),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_543),
.Y(n_544)
);


endmodule