module real_jpeg_6102_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g88 ( 
.A(n_0),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_1),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_60)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_1),
.A2(n_155),
.B1(n_157),
.B2(n_158),
.Y(n_154)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_1),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_1),
.A2(n_157),
.B1(n_211),
.B2(n_214),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_2),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_50)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_2),
.A2(n_53),
.B1(n_141),
.B2(n_143),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_2),
.A2(n_53),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_2),
.A2(n_53),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

O2A1O1Ixp33_ASAP7_75t_L g264 ( 
.A1(n_2),
.A2(n_265),
.B(n_268),
.C(n_271),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_2),
.B(n_220),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_2),
.B(n_106),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_2),
.B(n_305),
.C(n_308),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_2),
.B(n_96),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_2),
.B(n_302),
.C(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_2),
.B(n_32),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_3),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_3),
.A2(n_28),
.B1(n_38),
.B2(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_3),
.A2(n_28),
.B1(n_204),
.B2(n_206),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_3),
.A2(n_28),
.B1(n_275),
.B2(n_276),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_4),
.Y(n_110)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_4),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_4),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_5),
.Y(n_401)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_7),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_7),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_7),
.A2(n_98),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_7),
.A2(n_98),
.B1(n_167),
.B2(n_170),
.Y(n_166)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_8),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_8),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_8),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g293 ( 
.A(n_8),
.Y(n_293)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_9),
.Y(n_267)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_11),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_13),
.Y(n_108)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_13),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_396),
.B(n_399),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_191),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_190),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_146),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_19),
.B(n_146),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_135),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_133),
.B2(n_134),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_56),
.B2(n_57),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_23),
.A2(n_24),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_23),
.A2(n_24),
.B1(n_159),
.B2(n_349),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_24),
.B(n_199),
.C(n_223),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_24),
.B(n_159),
.C(n_263),
.Y(n_262)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_50),
.B2(n_55),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g133 ( 
.A1(n_25),
.A2(n_31),
.B1(n_50),
.B2(n_55),
.Y(n_133)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_31),
.A2(n_50),
.B(n_55),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_42),
.Y(n_31)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_36),
.B1(n_38),
.B2(n_40),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_34),
.Y(n_328)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_35),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_43),
.B1(n_45),
.B2(n_47),
.Y(n_42)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g269 ( 
.A(n_37),
.Y(n_269)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_43),
.Y(n_271)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_L g268 ( 
.A1(n_53),
.A2(n_269),
.B(n_270),
.Y(n_268)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_103),
.B2(n_132),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_68),
.B1(n_96),
.B2(n_97),
.Y(n_59)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_63),
.Y(n_142)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_67),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_68),
.B(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g159 ( 
.A1(n_69),
.A2(n_84),
.B1(n_140),
.B2(n_160),
.Y(n_159)
);

OA22x2_ASAP7_75t_L g223 ( 
.A1(n_69),
.A2(n_84),
.B1(n_140),
.B2(n_160),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_69),
.B(n_84),
.Y(n_240)
);

NAND2x1_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_84),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_75),
.B1(n_79),
.B2(n_81),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_78),
.Y(n_270)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_80),
.Y(n_333)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_84),
.A2(n_137),
.B(n_138),
.Y(n_136)
);

AOI22x1_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_89),
.B1(n_91),
.B2(n_93),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_86),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_88),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_88),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_103),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_133),
.C(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_103),
.A2(n_132),
.B1(n_136),
.B2(n_150),
.Y(n_149)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_127),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_104),
.B(n_186),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_116),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g201 ( 
.A1(n_105),
.A2(n_116),
.B1(n_202),
.B2(n_207),
.Y(n_201)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2x1_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_106),
.A2(n_117),
.B1(n_127),
.B2(n_154),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_106),
.A2(n_154),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_106),
.B(n_203),
.Y(n_238)
);

AO22x1_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_109),
.B1(n_111),
.B2(n_114),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_108),
.Y(n_307)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_109),
.Y(n_236)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_110),
.Y(n_176)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_112),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_113),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_113),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_117),
.B(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_120),
.Y(n_188)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_133),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_134),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_133),
.B(n_228),
.C(n_239),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_133),
.A2(n_134),
.B1(n_239),
.B2(n_259),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_133),
.A2(n_134),
.B1(n_357),
.B2(n_358),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_133),
.B(n_223),
.C(n_359),
.Y(n_376)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_139),
.B(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.C(n_163),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_147),
.A2(n_151),
.B1(n_152),
.B2(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_147),
.Y(n_393)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_152),
.A2(n_153),
.B(n_159),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_159),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_159),
.A2(n_345),
.B1(n_346),
.B2(n_349),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_159),
.Y(n_349)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_163),
.B(n_392),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B(n_189),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_164),
.B(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_183),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_165),
.A2(n_183),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_165),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_165),
.A2(n_189),
.B1(n_226),
.B2(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_172),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_169),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_172),
.B(n_233),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_181),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_173),
.A2(n_209),
.B1(n_216),
.B2(n_217),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_173),
.B(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_174),
.A2(n_233),
.B1(n_274),
.B2(n_277),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_174),
.A2(n_233),
.B1(n_274),
.B2(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_176),
.Y(n_276)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_180),
.Y(n_278)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_183),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

AND2x2_ASAP7_75t_SL g237 ( 
.A(n_185),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_189),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_390),
.B(n_395),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI211xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_279),
.B(n_384),
.C(n_389),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_252),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g384 ( 
.A1(n_196),
.A2(n_252),
.B(n_385),
.C(n_388),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_241),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g389 ( 
.A(n_197),
.B(n_241),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_224),
.C(n_227),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_198),
.B(n_224),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_221),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_208),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_200),
.A2(n_201),
.B1(n_208),
.B2(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_200),
.A2(n_201),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_200),
.A2(n_201),
.B1(n_341),
.B2(n_342),
.Y(n_340)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_201),
.B(n_273),
.C(n_316),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_201),
.B(n_341),
.C(n_343),
.Y(n_354)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_208),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_210),
.A2(n_218),
.B(n_231),
.Y(n_230)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_213),
.Y(n_309)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_222),
.A2(n_223),
.B1(n_237),
.B2(n_300),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_222),
.B(n_300),
.C(n_323),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_222),
.A2(n_223),
.B1(n_359),
.B2(n_360),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_254),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_258),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_237),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_230),
.A2(n_237),
.B1(n_300),
.B2(n_375),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_230),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_237),
.A2(n_300),
.B1(n_301),
.B2(n_310),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_237),
.Y(n_300)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_239),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_250),
.B2(n_251),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.Y(n_243)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_244),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_247),
.B(n_249),
.C(n_251),
.Y(n_394)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_250),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_253),
.B(n_255),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_260),
.C(n_262),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_256),
.A2(n_257),
.B1(n_260),
.B2(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_260),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_262),
.B(n_382),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_263),
.B(n_372),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_272),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_264),
.A2(n_272),
.B1(n_273),
.B2(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_264),
.Y(n_366)
);

INVx6_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_272),
.A2(n_273),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_295),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_295),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_276),
.Y(n_288)
);

INVx8_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_368),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_353),
.B(n_367),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_338),
.B(n_352),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_320),
.B(n_337),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_312),
.B(n_319),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_297),
.B(n_311),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_294),
.B(n_296),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_290),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_290),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_290),
.A2(n_298),
.B1(n_347),
.B2(n_348),
.Y(n_346)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_299),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_298),
.B(n_347),
.C(n_349),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_310),
.Y(n_318)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_301),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.Y(n_301)
);

INVx5_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_318),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_318),
.Y(n_319)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_316),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_321),
.B(n_322),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_336),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_325),
.B1(n_334),
.B2(n_335),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_324),
.B(n_335),
.Y(n_341)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_329),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx6_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_351),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_339),
.B(n_351),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_343),
.B1(n_344),
.B2(n_350),
.Y(n_339)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_340),
.Y(n_350)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_341),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_348),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_355),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_361),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_356),
.B(n_363),
.C(n_364),
.Y(n_377)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_359),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_362),
.A2(n_363),
.B1(n_364),
.B2(n_365),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

NOR2x1_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_378),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_370),
.B(n_377),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_370),
.B(n_377),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_373),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_371),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_376),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_374),
.B(n_376),
.C(n_380),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_378),
.A2(n_386),
.B(n_387),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_381),
.Y(n_378)
);

OR2x2_ASAP7_75t_L g387 ( 
.A(n_379),
.B(n_381),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_391),
.B(n_394),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_391),
.B(n_394),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx13_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx8_ASAP7_75t_L g400 ( 
.A(n_398),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_401),
.Y(n_399)
);


endmodule