module fake_jpeg_6237_n_44 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_44);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_44;

wire n_33;
wire n_23;
wire n_27;
wire n_40;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_SL g23 ( 
.A(n_0),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_0),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_22),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_8),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_10),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_1),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_36),
.C(n_25),
.Y(n_38)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_2),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_34),
.B1(n_35),
.B2(n_27),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_29),
.A2(n_12),
.B1(n_5),
.B2(n_6),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_2),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_38),
.B1(n_33),
.B2(n_30),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_38),
.Y(n_41)
);

AOI322xp5_ASAP7_75t_L g42 ( 
.A1(n_41),
.A2(n_30),
.A3(n_39),
.B1(n_15),
.B2(n_17),
.C1(n_7),
.C2(n_20),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_11),
.C(n_19),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_26),
.Y(n_44)
);


endmodule