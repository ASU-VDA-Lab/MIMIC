module fake_netlist_1_11414_n_1374 (n_117, n_44, n_361, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_348, n_252, n_152, n_113, n_353, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_351, n_83, n_28, n_48, n_100, n_305, n_228, n_345, n_360, n_236, n_340, n_150, n_373, n_3, n_18, n_301, n_66, n_222, n_234, n_366, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_367, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_354, n_32, n_235, n_243, n_331, n_352, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_369, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_362, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_370, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_357, n_260, n_78, n_197, n_201, n_317, n_4, n_374, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_365, n_179, n_315, n_363, n_86, n_143, n_295, n_263, n_166, n_186, n_364, n_75, n_376, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_349, n_51, n_225, n_220, n_358, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_378, n_359, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_377, n_343, n_127, n_291, n_170, n_356, n_281, n_341, n_58, n_122, n_187, n_375, n_138, n_371, n_323, n_347, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_368, n_355, n_226, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_372, n_194, n_287, n_110, n_261, n_332, n_350, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1374);
input n_117;
input n_44;
input n_361;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_348;
input n_252;
input n_152;
input n_113;
input n_353;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_351;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_360;
input n_236;
input n_340;
input n_150;
input n_373;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_366;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_367;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_354;
input n_32;
input n_235;
input n_243;
input n_331;
input n_352;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_369;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_362;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_370;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_357;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_374;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_365;
input n_179;
input n_315;
input n_363;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_364;
input n_75;
input n_376;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_349;
input n_51;
input n_225;
input n_220;
input n_358;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_378;
input n_359;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_377;
input n_343;
input n_127;
input n_291;
input n_170;
input n_356;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_375;
input n_138;
input n_371;
input n_323;
input n_347;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_368;
input n_355;
input n_226;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_372;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_350;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1374;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_1363;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_382;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1271;
wire n_708;
wire n_1062;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_733;
wire n_894;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_901;
wire n_834;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_688;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1372;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_1273;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_495;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_584;
wire n_1130;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_458;
wire n_1084;
wire n_618;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_1022;
wire n_802;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_401;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_1275;
wire n_955;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_653;
wire n_881;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1239;
wire n_1335;
wire n_924;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_600;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
wire n_1291;
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_237), .Y(n_379) );
INVx1_ASAP7_75t_SL g380 ( .A(n_154), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_344), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_18), .Y(n_382) );
INVxp33_ASAP7_75t_L g383 ( .A(n_293), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_359), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_365), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_48), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_324), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_91), .Y(n_388) );
BUFx3_ASAP7_75t_L g389 ( .A(n_303), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_361), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_74), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_348), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_242), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_302), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_106), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_325), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_357), .Y(n_397) );
CKINVDCx5p33_ASAP7_75t_R g398 ( .A(n_246), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_353), .Y(n_399) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_179), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_243), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_298), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_253), .Y(n_403) );
CKINVDCx16_ASAP7_75t_R g404 ( .A(n_143), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_99), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_276), .Y(n_406) );
BUFx3_ASAP7_75t_L g407 ( .A(n_45), .Y(n_407) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_345), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_285), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_3), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_326), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_356), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_272), .Y(n_413) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_89), .Y(n_414) );
CKINVDCx5p33_ASAP7_75t_R g415 ( .A(n_249), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_81), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_76), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_202), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_364), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_323), .B(n_196), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_85), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_172), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_352), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_266), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_209), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_80), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_156), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_314), .Y(n_428) );
CKINVDCx5p33_ASAP7_75t_R g429 ( .A(n_50), .Y(n_429) );
CKINVDCx5p33_ASAP7_75t_R g430 ( .A(n_316), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_227), .Y(n_431) );
CKINVDCx5p33_ASAP7_75t_R g432 ( .A(n_299), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_349), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_155), .Y(n_434) );
CKINVDCx5p33_ASAP7_75t_R g435 ( .A(n_49), .Y(n_435) );
INVxp67_ASAP7_75t_L g436 ( .A(n_319), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_373), .B(n_90), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_8), .Y(n_438) );
BUFx3_ASAP7_75t_L g439 ( .A(n_197), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_141), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_281), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_330), .Y(n_442) );
BUFx8_ASAP7_75t_SL g443 ( .A(n_150), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_247), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_346), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_358), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_354), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_308), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_283), .Y(n_449) );
CKINVDCx16_ASAP7_75t_R g450 ( .A(n_218), .Y(n_450) );
INVx1_ASAP7_75t_SL g451 ( .A(n_304), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_22), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_374), .Y(n_453) );
BUFx10_ASAP7_75t_L g454 ( .A(n_236), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_284), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g456 ( .A(n_166), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_273), .Y(n_457) );
CKINVDCx5p33_ASAP7_75t_R g458 ( .A(n_174), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_52), .Y(n_459) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_191), .Y(n_460) );
CKINVDCx5p33_ASAP7_75t_R g461 ( .A(n_109), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_100), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_238), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_61), .Y(n_464) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_208), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_287), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_369), .B(n_201), .Y(n_467) );
CKINVDCx5p33_ASAP7_75t_R g468 ( .A(n_25), .Y(n_468) );
BUFx3_ASAP7_75t_L g469 ( .A(n_355), .Y(n_469) );
BUFx5_ASAP7_75t_L g470 ( .A(n_248), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_267), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_198), .Y(n_472) );
CKINVDCx16_ASAP7_75t_R g473 ( .A(n_212), .Y(n_473) );
INVxp33_ASAP7_75t_SL g474 ( .A(n_171), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g475 ( .A(n_360), .Y(n_475) );
BUFx3_ASAP7_75t_L g476 ( .A(n_371), .Y(n_476) );
CKINVDCx5p33_ASAP7_75t_R g477 ( .A(n_87), .Y(n_477) );
CKINVDCx14_ASAP7_75t_R g478 ( .A(n_40), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_235), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_233), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_254), .Y(n_481) );
CKINVDCx5p33_ASAP7_75t_R g482 ( .A(n_5), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_301), .Y(n_483) );
CKINVDCx5p33_ASAP7_75t_R g484 ( .A(n_41), .Y(n_484) );
CKINVDCx5p33_ASAP7_75t_R g485 ( .A(n_135), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_363), .Y(n_486) );
CKINVDCx5p33_ASAP7_75t_R g487 ( .A(n_269), .Y(n_487) );
INVxp67_ASAP7_75t_SL g488 ( .A(n_97), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_189), .Y(n_489) );
BUFx3_ASAP7_75t_L g490 ( .A(n_126), .Y(n_490) );
CKINVDCx5p33_ASAP7_75t_R g491 ( .A(n_288), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_98), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_211), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_309), .Y(n_494) );
CKINVDCx5p33_ASAP7_75t_R g495 ( .A(n_351), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_315), .Y(n_496) );
INVx1_ASAP7_75t_SL g497 ( .A(n_334), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_12), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_72), .Y(n_499) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_129), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_350), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_30), .Y(n_502) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_103), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_219), .Y(n_504) );
CKINVDCx16_ASAP7_75t_R g505 ( .A(n_116), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_186), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_164), .Y(n_507) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_338), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_262), .Y(n_509) );
CKINVDCx5p33_ASAP7_75t_R g510 ( .A(n_278), .Y(n_510) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_264), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_327), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_216), .Y(n_513) );
CKINVDCx5p33_ASAP7_75t_R g514 ( .A(n_295), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g515 ( .A(n_124), .Y(n_515) );
CKINVDCx16_ASAP7_75t_R g516 ( .A(n_39), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_362), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_30), .Y(n_518) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_311), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_29), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_185), .Y(n_521) );
BUFx8_ASAP7_75t_SL g522 ( .A(n_378), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_297), .Y(n_523) );
CKINVDCx5p33_ASAP7_75t_R g524 ( .A(n_279), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_19), .Y(n_525) );
CKINVDCx5p33_ASAP7_75t_R g526 ( .A(n_34), .Y(n_526) );
INVx2_ASAP7_75t_SL g527 ( .A(n_332), .Y(n_527) );
CKINVDCx5p33_ASAP7_75t_R g528 ( .A(n_117), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_252), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_366), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_470), .Y(n_531) );
BUFx8_ASAP7_75t_SL g532 ( .A(n_443), .Y(n_532) );
BUFx2_ASAP7_75t_L g533 ( .A(n_478), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_503), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_470), .Y(n_535) );
AND2x4_ASAP7_75t_L g536 ( .A(n_410), .B(n_0), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_470), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_470), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_470), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_527), .B(n_516), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_438), .Y(n_541) );
NAND2xp33_ASAP7_75t_L g542 ( .A(n_420), .B(n_46), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_383), .B(n_0), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_385), .Y(n_544) );
BUFx2_ASAP7_75t_L g545 ( .A(n_382), .Y(n_545) );
AND2x4_ASAP7_75t_L g546 ( .A(n_452), .B(n_1), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_395), .B(n_418), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_468), .Y(n_548) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_400), .Y(n_549) );
OAI21x1_ASAP7_75t_L g550 ( .A1(n_431), .A2(n_51), .B(n_47), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_404), .B(n_1), .Y(n_551) );
INVx2_ASAP7_75t_SL g552 ( .A(n_454), .Y(n_552) );
INVx3_ASAP7_75t_L g553 ( .A(n_454), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_434), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_471), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_436), .B(n_2), .Y(n_556) );
INVx3_ASAP7_75t_L g557 ( .A(n_535), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_536), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_532), .Y(n_559) );
INVx3_ASAP7_75t_L g560 ( .A(n_531), .Y(n_560) );
NAND2xp33_ASAP7_75t_L g561 ( .A(n_543), .B(n_437), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_536), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_534), .A2(n_473), .B1(n_505), .B2(n_450), .Y(n_563) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_532), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_546), .Y(n_565) );
INVx4_ASAP7_75t_L g566 ( .A(n_546), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_531), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_537), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_548), .A2(n_482), .B1(n_520), .B2(n_484), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_533), .B(n_498), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_537), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_540), .B(n_526), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_538), .Y(n_573) );
BUFx3_ASAP7_75t_L g574 ( .A(n_550), .Y(n_574) );
INVx2_ASAP7_75t_SL g575 ( .A(n_545), .Y(n_575) );
OR2x6_ASAP7_75t_L g576 ( .A(n_552), .B(n_502), .Y(n_576) );
INVx3_ASAP7_75t_L g577 ( .A(n_538), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_553), .B(n_379), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_539), .Y(n_579) );
INVx2_ASAP7_75t_SL g580 ( .A(n_548), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_560), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_566), .B(n_553), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_558), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g584 ( .A1(n_562), .A2(n_541), .B1(n_462), .B2(n_388), .Y(n_584) );
INVx2_ASAP7_75t_SL g585 ( .A(n_576), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_572), .B(n_556), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_566), .B(n_551), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_560), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_565), .B(n_556), .Y(n_589) );
INVx3_ASAP7_75t_L g590 ( .A(n_566), .Y(n_590) );
O2A1O1Ixp33_ASAP7_75t_L g591 ( .A1(n_561), .A2(n_542), .B(n_547), .C(n_554), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_578), .B(n_474), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_560), .Y(n_593) );
NOR2xp67_ASAP7_75t_L g594 ( .A(n_563), .B(n_544), .Y(n_594) );
INVxp67_ASAP7_75t_SL g595 ( .A(n_561), .Y(n_595) );
BUFx3_ASAP7_75t_L g596 ( .A(n_576), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_580), .B(n_381), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_575), .B(n_384), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_570), .B(n_554), .Y(n_599) );
INVx8_ASAP7_75t_L g600 ( .A(n_576), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_557), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_571), .B(n_555), .Y(n_602) );
AO221x1_ASAP7_75t_L g603 ( .A1(n_569), .A2(n_522), .B1(n_465), .B2(n_511), .C(n_414), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_573), .B(n_542), .Y(n_604) );
NOR3xp33_ASAP7_75t_L g605 ( .A(n_559), .B(n_525), .C(n_518), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_577), .B(n_555), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_557), .Y(n_607) );
OAI21xp5_ASAP7_75t_L g608 ( .A1(n_574), .A2(n_539), .B(n_390), .Y(n_608) );
INVx2_ASAP7_75t_SL g609 ( .A(n_574), .Y(n_609) );
NAND2xp5_ASAP7_75t_SL g610 ( .A(n_557), .B(n_387), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_577), .Y(n_611) );
OAI22xp33_ASAP7_75t_L g612 ( .A1(n_559), .A2(n_386), .B1(n_392), .B2(n_391), .Y(n_612) );
O2A1O1Ixp5_ASAP7_75t_L g613 ( .A1(n_567), .A2(n_488), .B(n_393), .C(n_406), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_577), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_567), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_568), .B(n_380), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_564), .B(n_2), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_568), .B(n_380), .Y(n_618) );
NAND2x1p5_ASAP7_75t_L g619 ( .A(n_579), .B(n_467), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_579), .B(n_451), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_564), .Y(n_621) );
OAI221xp5_ASAP7_75t_L g622 ( .A1(n_569), .A2(n_497), .B1(n_451), .B2(n_411), .C(n_416), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_572), .B(n_497), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_595), .B(n_394), .Y(n_624) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_596), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g626 ( .A1(n_608), .A2(n_409), .B(n_401), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_583), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_619), .A2(n_419), .B1(n_421), .B2(n_417), .Y(n_628) );
OA22x2_ASAP7_75t_L g629 ( .A1(n_584), .A2(n_424), .B1(n_426), .B2(n_422), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_619), .A2(n_428), .B1(n_433), .B2(n_427), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_587), .B(n_396), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_586), .B(n_397), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_585), .B(n_398), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_589), .B(n_399), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_606), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_589), .B(n_402), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_608), .A2(n_447), .B(n_440), .Y(n_637) );
BUFx8_ASAP7_75t_SL g638 ( .A(n_621), .Y(n_638) );
BUFx8_ASAP7_75t_L g639 ( .A(n_617), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_584), .B(n_3), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_623), .B(n_403), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_599), .B(n_405), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_600), .B(n_408), .Y(n_643) );
NOR2xp67_ASAP7_75t_L g644 ( .A(n_590), .B(n_53), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_604), .A2(n_455), .B(n_453), .Y(n_645) );
INVx3_ASAP7_75t_L g646 ( .A(n_590), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_602), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_604), .A2(n_459), .B(n_457), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_620), .B(n_412), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_620), .B(n_413), .Y(n_650) );
OA22x2_ASAP7_75t_L g651 ( .A1(n_603), .A2(n_464), .B1(n_466), .B2(n_463), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_581), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_588), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_601), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_609), .A2(n_479), .B(n_472), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_607), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_600), .B(n_4), .Y(n_657) );
OAI321xp33_ASAP7_75t_L g658 ( .A1(n_591), .A2(n_549), .A3(n_483), .B1(n_489), .B2(n_494), .C(n_493), .Y(n_658) );
O2A1O1Ixp33_ASAP7_75t_SL g659 ( .A1(n_614), .A2(n_496), .B(n_499), .C(n_486), .Y(n_659) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_600), .Y(n_660) );
OR2x6_ASAP7_75t_L g661 ( .A(n_597), .B(n_501), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_582), .Y(n_662) );
O2A1O1Ixp33_ASAP7_75t_L g663 ( .A1(n_622), .A2(n_612), .B(n_613), .C(n_605), .Y(n_663) );
OAI21x1_ASAP7_75t_L g664 ( .A1(n_615), .A2(n_504), .B(n_492), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_593), .Y(n_665) );
BUFx4f_ASAP7_75t_L g666 ( .A(n_611), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_594), .B(n_415), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g668 ( .A(n_592), .B(n_423), .Y(n_668) );
O2A1O1Ixp33_ASAP7_75t_L g669 ( .A1(n_598), .A2(n_507), .B(n_512), .C(n_506), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_610), .A2(n_517), .B(n_513), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_616), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_618), .B(n_425), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_595), .B(n_429), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_595), .A2(n_523), .B1(n_529), .B2(n_521), .Y(n_674) );
AOI21xp5_ASAP7_75t_L g675 ( .A1(n_608), .A2(n_407), .B(n_389), .Y(n_675) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_645), .A2(n_432), .B(n_430), .Y(n_676) );
AO21x2_ASAP7_75t_L g677 ( .A1(n_658), .A2(n_664), .B(n_637), .Y(n_677) );
NAND3x1_ASAP7_75t_L g678 ( .A(n_640), .B(n_4), .C(n_5), .Y(n_678) );
INVx3_ASAP7_75t_L g679 ( .A(n_646), .Y(n_679) );
BUFx2_ASAP7_75t_R g680 ( .A(n_638), .Y(n_680) );
OAI21x1_ASAP7_75t_L g681 ( .A1(n_644), .A2(n_414), .B(n_400), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_647), .A2(n_441), .B1(n_442), .B2(n_435), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_648), .A2(n_445), .B(n_444), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_657), .B(n_446), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_627), .B(n_448), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_635), .A2(n_449), .B1(n_458), .B2(n_456), .Y(n_686) );
AO22x2_ASAP7_75t_L g687 ( .A1(n_628), .A2(n_469), .B1(n_476), .B2(n_439), .Y(n_687) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_649), .A2(n_461), .B(n_460), .Y(n_688) );
OAI21x1_ASAP7_75t_L g689 ( .A1(n_644), .A2(n_414), .B(n_400), .Y(n_689) );
OR2x2_ASAP7_75t_L g690 ( .A(n_660), .B(n_6), .Y(n_690) );
NAND2x1_ASAP7_75t_L g691 ( .A(n_646), .B(n_465), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g692 ( .A(n_663), .B(n_511), .C(n_465), .Y(n_692) );
AOI221x1_ASAP7_75t_L g693 ( .A1(n_675), .A2(n_549), .B1(n_519), .B2(n_511), .C(n_490), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_671), .B(n_475), .Y(n_694) );
OAI21xp5_ASAP7_75t_L g695 ( .A1(n_626), .A2(n_480), .B(n_477), .Y(n_695) );
BUFx3_ASAP7_75t_L g696 ( .A(n_625), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_630), .A2(n_485), .B1(n_487), .B2(n_481), .Y(n_697) );
INVx3_ASAP7_75t_SL g698 ( .A(n_651), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_629), .B(n_6), .Y(n_699) );
AOI21x1_ASAP7_75t_L g700 ( .A1(n_655), .A2(n_519), .B(n_549), .Y(n_700) );
AOI221xp5_ASAP7_75t_SL g701 ( .A1(n_674), .A2(n_519), .B1(n_549), .B2(n_9), .C(n_7), .Y(n_701) );
AOI21xp5_ASAP7_75t_L g702 ( .A1(n_650), .A2(n_495), .B(n_491), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_654), .Y(n_703) );
BUFx2_ASAP7_75t_L g704 ( .A(n_639), .Y(n_704) );
NAND3xp33_ASAP7_75t_L g705 ( .A(n_669), .B(n_508), .C(n_500), .Y(n_705) );
OAI21x1_ASAP7_75t_L g706 ( .A1(n_656), .A2(n_55), .B(n_54), .Y(n_706) );
BUFx6f_ASAP7_75t_L g707 ( .A(n_666), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_652), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_634), .A2(n_510), .B(n_509), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_636), .B(n_514), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_632), .B(n_515), .Y(n_711) );
BUFx6f_ASAP7_75t_L g712 ( .A(n_666), .Y(n_712) );
AND2x4_ASAP7_75t_L g713 ( .A(n_661), .B(n_662), .Y(n_713) );
NAND2xp5_ASAP7_75t_SL g714 ( .A(n_643), .B(n_524), .Y(n_714) );
INVx3_ASAP7_75t_SL g715 ( .A(n_661), .Y(n_715) );
AOI21x1_ASAP7_75t_L g716 ( .A1(n_670), .A2(n_672), .B(n_665), .Y(n_716) );
OAI21xp5_ASAP7_75t_L g717 ( .A1(n_658), .A2(n_530), .B(n_528), .Y(n_717) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_661), .Y(n_718) );
BUFx3_ASAP7_75t_L g719 ( .A(n_639), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g720 ( .A1(n_624), .A2(n_57), .B(n_56), .Y(n_720) );
AOI221x1_ASAP7_75t_L g721 ( .A1(n_667), .A2(n_9), .B1(n_7), .B2(n_8), .C(n_10), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_653), .Y(n_722) );
INVx2_ASAP7_75t_L g723 ( .A(n_673), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g724 ( .A1(n_631), .A2(n_59), .B(n_58), .Y(n_724) );
AO21x1_ASAP7_75t_L g725 ( .A1(n_641), .A2(n_62), .B(n_60), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_642), .B(n_10), .Y(n_726) );
OAI21xp5_ASAP7_75t_L g727 ( .A1(n_668), .A2(n_64), .B(n_63), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_659), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g729 ( .A1(n_633), .A2(n_66), .B(n_65), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_647), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_647), .B(n_11), .Y(n_731) );
INVx3_ASAP7_75t_L g732 ( .A(n_646), .Y(n_732) );
BUFx2_ASAP7_75t_L g733 ( .A(n_660), .Y(n_733) );
OAI21xp5_ASAP7_75t_L g734 ( .A1(n_645), .A2(n_68), .B(n_67), .Y(n_734) );
OAI21x1_ASAP7_75t_L g735 ( .A1(n_664), .A2(n_70), .B(n_69), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_730), .Y(n_736) );
BUFx8_ASAP7_75t_L g737 ( .A(n_704), .Y(n_737) );
OAI21x1_ASAP7_75t_L g738 ( .A1(n_681), .A2(n_73), .B(n_71), .Y(n_738) );
OA21x2_ASAP7_75t_L g739 ( .A1(n_693), .A2(n_77), .B(n_75), .Y(n_739) );
INVx6_ASAP7_75t_L g740 ( .A(n_719), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_730), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_703), .Y(n_742) );
OR2x2_ASAP7_75t_L g743 ( .A(n_715), .B(n_718), .Y(n_743) );
AO31x2_ASAP7_75t_L g744 ( .A1(n_725), .A2(n_13), .A3(n_11), .B(n_12), .Y(n_744) );
INVx3_ASAP7_75t_L g745 ( .A(n_707), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_703), .B(n_13), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_699), .Y(n_747) );
OAI21x1_ASAP7_75t_L g748 ( .A1(n_689), .A2(n_79), .B(n_78), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_708), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_731), .Y(n_750) );
OA21x2_ASAP7_75t_L g751 ( .A1(n_701), .A2(n_83), .B(n_82), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_722), .Y(n_752) );
OAI21x1_ASAP7_75t_SL g753 ( .A1(n_727), .A2(n_14), .B(n_15), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_716), .Y(n_754) );
OAI21x1_ASAP7_75t_L g755 ( .A1(n_735), .A2(n_86), .B(n_84), .Y(n_755) );
OR2x2_ASAP7_75t_L g756 ( .A(n_733), .B(n_14), .Y(n_756) );
OR2x2_ASAP7_75t_L g757 ( .A(n_690), .B(n_15), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_728), .Y(n_758) );
INVxp67_ASAP7_75t_SL g759 ( .A(n_696), .Y(n_759) );
OAI21x1_ASAP7_75t_L g760 ( .A1(n_706), .A2(n_92), .B(n_88), .Y(n_760) );
INVx2_ASAP7_75t_L g761 ( .A(n_723), .Y(n_761) );
INVx3_ASAP7_75t_L g762 ( .A(n_707), .Y(n_762) );
INVxp33_ASAP7_75t_L g763 ( .A(n_707), .Y(n_763) );
INVxp67_ASAP7_75t_SL g764 ( .A(n_713), .Y(n_764) );
OAI21x1_ASAP7_75t_L g765 ( .A1(n_700), .A2(n_94), .B(n_93), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_728), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_726), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_678), .Y(n_768) );
AO31x2_ASAP7_75t_L g769 ( .A1(n_721), .A2(n_18), .A3(n_16), .B(n_17), .Y(n_769) );
OA21x2_ASAP7_75t_L g770 ( .A1(n_692), .A2(n_96), .B(n_95), .Y(n_770) );
NOR2x1_ASAP7_75t_R g771 ( .A(n_680), .B(n_16), .Y(n_771) );
OAI21xp5_ASAP7_75t_L g772 ( .A1(n_695), .A2(n_17), .B(n_19), .Y(n_772) );
OAI21x1_ASAP7_75t_L g773 ( .A1(n_720), .A2(n_102), .B(n_101), .Y(n_773) );
CKINVDCx11_ASAP7_75t_R g774 ( .A(n_698), .Y(n_774) );
OAI21xp5_ASAP7_75t_L g775 ( .A1(n_705), .A2(n_20), .B(n_21), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_679), .Y(n_776) );
NOR2xp33_ASAP7_75t_L g777 ( .A(n_713), .B(n_20), .Y(n_777) );
INVx2_ASAP7_75t_SL g778 ( .A(n_712), .Y(n_778) );
INVx2_ASAP7_75t_L g779 ( .A(n_679), .Y(n_779) );
NOR2x1_ASAP7_75t_R g780 ( .A(n_712), .B(n_21), .Y(n_780) );
INVxp67_ASAP7_75t_L g781 ( .A(n_687), .Y(n_781) );
OAI21x1_ASAP7_75t_L g782 ( .A1(n_724), .A2(n_105), .B(n_104), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_694), .B(n_22), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_732), .Y(n_784) );
OAI21x1_ASAP7_75t_L g785 ( .A1(n_691), .A2(n_108), .B(n_107), .Y(n_785) );
INVx2_ASAP7_75t_SL g786 ( .A(n_712), .Y(n_786) );
OAI21x1_ASAP7_75t_L g787 ( .A1(n_734), .A2(n_111), .B(n_110), .Y(n_787) );
INVx2_ASAP7_75t_L g788 ( .A(n_732), .Y(n_788) );
OA21x2_ASAP7_75t_L g789 ( .A1(n_729), .A2(n_113), .B(n_112), .Y(n_789) );
NOR2xp67_ASAP7_75t_L g790 ( .A(n_684), .B(n_23), .Y(n_790) );
INVx2_ASAP7_75t_L g791 ( .A(n_677), .Y(n_791) );
AND2x2_ASAP7_75t_L g792 ( .A(n_687), .B(n_697), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_685), .Y(n_793) );
INVx3_ASAP7_75t_L g794 ( .A(n_710), .Y(n_794) );
BUFx3_ASAP7_75t_L g795 ( .A(n_682), .Y(n_795) );
OAI21x1_ASAP7_75t_L g796 ( .A1(n_688), .A2(n_115), .B(n_114), .Y(n_796) );
OAI21x1_ASAP7_75t_L g797 ( .A1(n_702), .A2(n_119), .B(n_118), .Y(n_797) );
OAI21x1_ASAP7_75t_L g798 ( .A1(n_709), .A2(n_121), .B(n_120), .Y(n_798) );
OA21x2_ASAP7_75t_L g799 ( .A1(n_717), .A2(n_123), .B(n_122), .Y(n_799) );
NAND2x1p5_ASAP7_75t_L g800 ( .A(n_714), .B(n_676), .Y(n_800) );
NAND2xp5_ASAP7_75t_SL g801 ( .A(n_686), .B(n_23), .Y(n_801) );
AND2x2_ASAP7_75t_L g802 ( .A(n_711), .B(n_24), .Y(n_802) );
AO21x1_ASAP7_75t_L g803 ( .A1(n_683), .A2(n_24), .B(n_25), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_730), .B(n_26), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_730), .B(n_26), .Y(n_805) );
NAND2xp5_ASAP7_75t_SL g806 ( .A(n_715), .B(n_27), .Y(n_806) );
INVxp67_ASAP7_75t_SL g807 ( .A(n_730), .Y(n_807) );
INVx2_ASAP7_75t_L g808 ( .A(n_730), .Y(n_808) );
AND2x4_ASAP7_75t_L g809 ( .A(n_730), .B(n_27), .Y(n_809) );
AO31x2_ASAP7_75t_L g810 ( .A1(n_725), .A2(n_31), .A3(n_28), .B(n_29), .Y(n_810) );
INVx2_ASAP7_75t_L g811 ( .A(n_736), .Y(n_811) );
INVx2_ASAP7_75t_L g812 ( .A(n_808), .Y(n_812) );
INVxp67_ASAP7_75t_L g813 ( .A(n_807), .Y(n_813) );
AO31x2_ASAP7_75t_L g814 ( .A1(n_754), .A2(n_244), .A3(n_376), .B(n_375), .Y(n_814) );
HB1xp67_ASAP7_75t_L g815 ( .A(n_741), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_761), .Y(n_816) );
BUFx6f_ASAP7_75t_L g817 ( .A(n_778), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_742), .Y(n_818) );
AND2x2_ASAP7_75t_L g819 ( .A(n_747), .B(n_759), .Y(n_819) );
HB1xp67_ASAP7_75t_L g820 ( .A(n_756), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_742), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_741), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_809), .Y(n_823) );
AO31x2_ASAP7_75t_L g824 ( .A1(n_754), .A2(n_241), .A3(n_372), .B(n_370), .Y(n_824) );
AND2x4_ASAP7_75t_SL g825 ( .A(n_809), .B(n_28), .Y(n_825) );
OAI22xp33_ASAP7_75t_SL g826 ( .A1(n_781), .A2(n_31), .B1(n_32), .B2(n_33), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_752), .Y(n_827) );
INVx2_ASAP7_75t_L g828 ( .A(n_752), .Y(n_828) );
HB1xp67_ASAP7_75t_L g829 ( .A(n_749), .Y(n_829) );
INVx1_ASAP7_75t_SL g830 ( .A(n_743), .Y(n_830) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_768), .B(n_32), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_804), .Y(n_832) );
HB1xp67_ASAP7_75t_L g833 ( .A(n_764), .Y(n_833) );
AOI21x1_ASAP7_75t_L g834 ( .A1(n_791), .A2(n_33), .B(n_34), .Y(n_834) );
INVx2_ASAP7_75t_SL g835 ( .A(n_737), .Y(n_835) );
INVx2_ASAP7_75t_L g836 ( .A(n_793), .Y(n_836) );
BUFx2_ASAP7_75t_L g837 ( .A(n_737), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_805), .Y(n_838) );
AND2x2_ASAP7_75t_L g839 ( .A(n_793), .B(n_35), .Y(n_839) );
AND2x2_ASAP7_75t_L g840 ( .A(n_757), .B(n_35), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_746), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_767), .B(n_36), .Y(n_842) );
HB1xp67_ASAP7_75t_L g843 ( .A(n_758), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_758), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_766), .Y(n_845) );
AND2x2_ASAP7_75t_L g846 ( .A(n_777), .B(n_36), .Y(n_846) );
INVxp67_ASAP7_75t_SL g847 ( .A(n_751), .Y(n_847) );
AND2x2_ASAP7_75t_L g848 ( .A(n_792), .B(n_37), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_766), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_790), .Y(n_850) );
INVx1_ASAP7_75t_SL g851 ( .A(n_745), .Y(n_851) );
BUFx2_ASAP7_75t_L g852 ( .A(n_745), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_803), .Y(n_853) );
INVx2_ASAP7_75t_L g854 ( .A(n_769), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_750), .Y(n_855) );
INVx2_ASAP7_75t_L g856 ( .A(n_769), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_767), .Y(n_857) );
INVxp67_ASAP7_75t_L g858 ( .A(n_780), .Y(n_858) );
INVx3_ASAP7_75t_L g859 ( .A(n_762), .Y(n_859) );
OR2x2_ASAP7_75t_L g860 ( .A(n_795), .B(n_37), .Y(n_860) );
HB1xp67_ASAP7_75t_L g861 ( .A(n_751), .Y(n_861) );
NOR2xp67_ASAP7_75t_SL g862 ( .A(n_740), .B(n_38), .Y(n_862) );
OAI21x1_ASAP7_75t_L g863 ( .A1(n_765), .A2(n_127), .B(n_125), .Y(n_863) );
INVx3_ASAP7_75t_L g864 ( .A(n_762), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_802), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_784), .B(n_38), .Y(n_866) );
INVx2_ASAP7_75t_L g867 ( .A(n_769), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_783), .Y(n_868) );
HB1xp67_ASAP7_75t_L g869 ( .A(n_784), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_794), .Y(n_870) );
INVx2_ASAP7_75t_L g871 ( .A(n_744), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_794), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_786), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_806), .Y(n_874) );
INVx2_ASAP7_75t_L g875 ( .A(n_810), .Y(n_875) );
OAI21x1_ASAP7_75t_L g876 ( .A1(n_760), .A2(n_130), .B(n_128), .Y(n_876) );
OA21x2_ASAP7_75t_L g877 ( .A1(n_787), .A2(n_132), .B(n_131), .Y(n_877) );
AO21x2_ASAP7_75t_L g878 ( .A1(n_753), .A2(n_39), .B(n_40), .Y(n_878) );
INVx2_ASAP7_75t_L g879 ( .A(n_744), .Y(n_879) );
INVxp67_ASAP7_75t_SL g880 ( .A(n_772), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_776), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_779), .Y(n_882) );
AND2x2_ASAP7_75t_L g883 ( .A(n_763), .B(n_774), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_788), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_801), .Y(n_885) );
BUFx3_ASAP7_75t_L g886 ( .A(n_740), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_744), .Y(n_887) );
INVx2_ASAP7_75t_L g888 ( .A(n_810), .Y(n_888) );
BUFx2_ASAP7_75t_L g889 ( .A(n_771), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_810), .Y(n_890) );
HB1xp67_ASAP7_75t_L g891 ( .A(n_799), .Y(n_891) );
HB1xp67_ASAP7_75t_L g892 ( .A(n_775), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_800), .Y(n_893) );
INVxp67_ASAP7_75t_L g894 ( .A(n_799), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_789), .B(n_41), .Y(n_895) );
INVx2_ASAP7_75t_L g896 ( .A(n_785), .Y(n_896) );
BUFx2_ASAP7_75t_L g897 ( .A(n_796), .Y(n_897) );
BUFx2_ASAP7_75t_L g898 ( .A(n_797), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_798), .Y(n_899) );
INVx2_ASAP7_75t_L g900 ( .A(n_755), .Y(n_900) );
HB1xp67_ASAP7_75t_L g901 ( .A(n_738), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_748), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_773), .Y(n_903) );
INVx2_ASAP7_75t_SL g904 ( .A(n_782), .Y(n_904) );
INVx2_ASAP7_75t_L g905 ( .A(n_789), .Y(n_905) );
AO31x2_ASAP7_75t_L g906 ( .A1(n_770), .A2(n_259), .A3(n_368), .B(n_367), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_739), .Y(n_907) );
BUFx6f_ASAP7_75t_L g908 ( .A(n_770), .Y(n_908) );
INVx2_ASAP7_75t_L g909 ( .A(n_739), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_761), .Y(n_910) );
CKINVDCx20_ASAP7_75t_R g911 ( .A(n_737), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_761), .Y(n_912) );
INVx2_ASAP7_75t_L g913 ( .A(n_736), .Y(n_913) );
INVx2_ASAP7_75t_L g914 ( .A(n_736), .Y(n_914) );
OAI21x1_ASAP7_75t_L g915 ( .A1(n_754), .A2(n_134), .B(n_133), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_761), .Y(n_916) );
INVx2_ASAP7_75t_L g917 ( .A(n_736), .Y(n_917) );
AND2x4_ASAP7_75t_L g918 ( .A(n_736), .B(n_42), .Y(n_918) );
AND2x2_ASAP7_75t_L g919 ( .A(n_819), .B(n_42), .Y(n_919) );
AND2x2_ASAP7_75t_L g920 ( .A(n_840), .B(n_43), .Y(n_920) );
NOR2xp67_ASAP7_75t_L g921 ( .A(n_858), .B(n_43), .Y(n_921) );
AND2x2_ASAP7_75t_L g922 ( .A(n_848), .B(n_44), .Y(n_922) );
BUFx3_ASAP7_75t_L g923 ( .A(n_911), .Y(n_923) );
INVx3_ASAP7_75t_L g924 ( .A(n_817), .Y(n_924) );
AND2x2_ASAP7_75t_L g925 ( .A(n_829), .B(n_44), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_818), .B(n_821), .Y(n_926) );
INVx2_ASAP7_75t_L g927 ( .A(n_828), .Y(n_927) );
AND2x2_ASAP7_75t_L g928 ( .A(n_865), .B(n_136), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_855), .Y(n_929) );
INVx2_ASAP7_75t_L g930 ( .A(n_811), .Y(n_930) );
INVx2_ASAP7_75t_L g931 ( .A(n_812), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_836), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_857), .Y(n_933) );
INVx2_ASAP7_75t_L g934 ( .A(n_913), .Y(n_934) );
HB1xp67_ASAP7_75t_L g935 ( .A(n_815), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_822), .B(n_137), .Y(n_936) );
INVx1_ASAP7_75t_SL g937 ( .A(n_833), .Y(n_937) );
AND2x2_ASAP7_75t_L g938 ( .A(n_830), .B(n_138), .Y(n_938) );
HB1xp67_ASAP7_75t_L g939 ( .A(n_815), .Y(n_939) );
HB1xp67_ASAP7_75t_L g940 ( .A(n_843), .Y(n_940) );
HB1xp67_ASAP7_75t_L g941 ( .A(n_843), .Y(n_941) );
OR2x2_ASAP7_75t_L g942 ( .A(n_830), .B(n_139), .Y(n_942) );
INVx3_ASAP7_75t_L g943 ( .A(n_817), .Y(n_943) );
BUFx2_ASAP7_75t_SL g944 ( .A(n_835), .Y(n_944) );
AND2x2_ASAP7_75t_L g945 ( .A(n_846), .B(n_839), .Y(n_945) );
HB1xp67_ASAP7_75t_L g946 ( .A(n_813), .Y(n_946) );
HB1xp67_ASAP7_75t_L g947 ( .A(n_813), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_827), .Y(n_948) );
AND2x4_ASAP7_75t_L g949 ( .A(n_833), .B(n_140), .Y(n_949) );
HB1xp67_ASAP7_75t_L g950 ( .A(n_869), .Y(n_950) );
INVx2_ASAP7_75t_L g951 ( .A(n_914), .Y(n_951) );
AND2x2_ASAP7_75t_L g952 ( .A(n_820), .B(n_142), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_816), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_910), .Y(n_954) );
HB1xp67_ASAP7_75t_L g955 ( .A(n_869), .Y(n_955) );
INVx2_ASAP7_75t_L g956 ( .A(n_917), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_825), .B(n_144), .Y(n_957) );
OR2x2_ASAP7_75t_L g958 ( .A(n_912), .B(n_145), .Y(n_958) );
HB1xp67_ASAP7_75t_L g959 ( .A(n_893), .Y(n_959) );
AND2x2_ASAP7_75t_L g960 ( .A(n_916), .B(n_146), .Y(n_960) );
AOI22xp5_ASAP7_75t_L g961 ( .A1(n_823), .A2(n_147), .B1(n_148), .B2(n_149), .Y(n_961) );
INVxp67_ASAP7_75t_SL g962 ( .A(n_901), .Y(n_962) );
INVx2_ASAP7_75t_L g963 ( .A(n_844), .Y(n_963) );
INVx2_ASAP7_75t_L g964 ( .A(n_845), .Y(n_964) );
INVx2_ASAP7_75t_R g965 ( .A(n_907), .Y(n_965) );
INVx3_ASAP7_75t_L g966 ( .A(n_817), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_849), .Y(n_967) );
INVx2_ASAP7_75t_L g968 ( .A(n_881), .Y(n_968) );
INVx2_ASAP7_75t_L g969 ( .A(n_882), .Y(n_969) );
AND2x2_ASAP7_75t_L g970 ( .A(n_831), .B(n_151), .Y(n_970) );
HB1xp67_ASAP7_75t_L g971 ( .A(n_854), .Y(n_971) );
INVx2_ASAP7_75t_L g972 ( .A(n_884), .Y(n_972) );
AND2x2_ASAP7_75t_L g973 ( .A(n_918), .B(n_152), .Y(n_973) );
INVx1_ASAP7_75t_L g974 ( .A(n_842), .Y(n_974) );
INVx2_ASAP7_75t_L g975 ( .A(n_918), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_842), .Y(n_976) );
AND2x2_ASAP7_75t_L g977 ( .A(n_860), .B(n_870), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_872), .B(n_153), .Y(n_978) );
INVx2_ASAP7_75t_L g979 ( .A(n_866), .Y(n_979) );
BUFx2_ASAP7_75t_L g980 ( .A(n_837), .Y(n_980) );
AND2x2_ASAP7_75t_L g981 ( .A(n_868), .B(n_157), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_866), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_832), .B(n_838), .Y(n_983) );
INVxp67_ASAP7_75t_R g984 ( .A(n_883), .Y(n_984) );
INVx2_ASAP7_75t_L g985 ( .A(n_834), .Y(n_985) );
AND2x2_ASAP7_75t_L g986 ( .A(n_873), .B(n_158), .Y(n_986) );
INVx1_ASAP7_75t_SL g987 ( .A(n_852), .Y(n_987) );
BUFx6f_ASAP7_75t_L g988 ( .A(n_886), .Y(n_988) );
AND2x2_ASAP7_75t_L g989 ( .A(n_850), .B(n_159), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_841), .B(n_160), .Y(n_990) );
AND2x2_ASAP7_75t_L g991 ( .A(n_874), .B(n_161), .Y(n_991) );
INVx2_ASAP7_75t_L g992 ( .A(n_856), .Y(n_992) );
INVx2_ASAP7_75t_L g993 ( .A(n_867), .Y(n_993) );
BUFx3_ASAP7_75t_L g994 ( .A(n_889), .Y(n_994) );
OAI21xp33_ASAP7_75t_L g995 ( .A1(n_826), .A2(n_162), .B(n_163), .Y(n_995) );
HB1xp67_ASAP7_75t_L g996 ( .A(n_890), .Y(n_996) );
HB1xp67_ASAP7_75t_L g997 ( .A(n_871), .Y(n_997) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_853), .B(n_165), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_885), .Y(n_999) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_858), .B(n_167), .Y(n_1000) );
INVx1_ASAP7_75t_L g1001 ( .A(n_878), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_859), .B(n_168), .Y(n_1002) );
NOR2xp67_ASAP7_75t_L g1003 ( .A(n_892), .B(n_169), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_878), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1005 ( .A(n_880), .B(n_875), .Y(n_1005) );
INVx2_ASAP7_75t_L g1006 ( .A(n_859), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_864), .Y(n_1007) );
INVx2_ASAP7_75t_L g1008 ( .A(n_864), .Y(n_1008) );
AND2x2_ASAP7_75t_L g1009 ( .A(n_851), .B(n_170), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_826), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_851), .B(n_173), .Y(n_1011) );
HB1xp67_ASAP7_75t_L g1012 ( .A(n_879), .Y(n_1012) );
OAI22xp5_ASAP7_75t_L g1013 ( .A1(n_880), .A2(n_175), .B1(n_176), .B2(n_177), .Y(n_1013) );
INVx2_ASAP7_75t_L g1014 ( .A(n_887), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_888), .B(n_178), .Y(n_1015) );
HB1xp67_ASAP7_75t_L g1016 ( .A(n_901), .Y(n_1016) );
NOR2x1_ASAP7_75t_L g1017 ( .A(n_895), .B(n_180), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_895), .Y(n_1018) );
HB1xp67_ASAP7_75t_L g1019 ( .A(n_902), .Y(n_1019) );
INVxp67_ASAP7_75t_L g1020 ( .A(n_862), .Y(n_1020) );
NOR2xp33_ASAP7_75t_L g1021 ( .A(n_897), .B(n_181), .Y(n_1021) );
INVx2_ASAP7_75t_L g1022 ( .A(n_814), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_814), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_861), .A2(n_182), .B1(n_183), .B2(n_184), .Y(n_1024) );
AND2x4_ASAP7_75t_L g1025 ( .A(n_814), .B(n_187), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_824), .B(n_188), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_824), .Y(n_1027) );
BUFx3_ASAP7_75t_L g1028 ( .A(n_915), .Y(n_1028) );
AND2x2_ASAP7_75t_L g1029 ( .A(n_824), .B(n_190), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_903), .Y(n_1030) );
INVx4_ASAP7_75t_L g1031 ( .A(n_877), .Y(n_1031) );
OR2x2_ASAP7_75t_L g1032 ( .A(n_899), .B(n_377), .Y(n_1032) );
BUFx3_ASAP7_75t_L g1033 ( .A(n_876), .Y(n_1033) );
BUFx6f_ASAP7_75t_L g1034 ( .A(n_863), .Y(n_1034) );
OR2x2_ASAP7_75t_L g1035 ( .A(n_898), .B(n_192), .Y(n_1035) );
HB1xp67_ASAP7_75t_L g1036 ( .A(n_861), .Y(n_1036) );
HB1xp67_ASAP7_75t_L g1037 ( .A(n_891), .Y(n_1037) );
INVx2_ASAP7_75t_L g1038 ( .A(n_896), .Y(n_1038) );
NAND2xp5_ASAP7_75t_L g1039 ( .A(n_891), .B(n_193), .Y(n_1039) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_906), .B(n_194), .Y(n_1040) );
INVx2_ASAP7_75t_L g1041 ( .A(n_904), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_894), .B(n_195), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_900), .Y(n_1043) );
INVx1_ASAP7_75t_SL g1044 ( .A(n_877), .Y(n_1044) );
BUFx3_ASAP7_75t_L g1045 ( .A(n_906), .Y(n_1045) );
INVx2_ASAP7_75t_L g1046 ( .A(n_906), .Y(n_1046) );
INVx2_ASAP7_75t_L g1047 ( .A(n_909), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_905), .Y(n_1048) );
HB1xp67_ASAP7_75t_L g1049 ( .A(n_894), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_847), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_847), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_908), .Y(n_1052) );
INVx2_ASAP7_75t_L g1053 ( .A(n_908), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_908), .B(n_199), .Y(n_1054) );
HB1xp67_ASAP7_75t_L g1055 ( .A(n_815), .Y(n_1055) );
BUFx3_ASAP7_75t_L g1056 ( .A(n_911), .Y(n_1056) );
OR2x2_ASAP7_75t_L g1057 ( .A(n_937), .B(n_200), .Y(n_1057) );
INVx3_ASAP7_75t_L g1058 ( .A(n_937), .Y(n_1058) );
NOR2xp33_ASAP7_75t_L g1059 ( .A(n_980), .B(n_203), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_945), .B(n_204), .Y(n_1060) );
AND2x2_ASAP7_75t_L g1061 ( .A(n_977), .B(n_205), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_919), .B(n_206), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_946), .B(n_207), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_946), .B(n_210), .Y(n_1064) );
AND2x2_ASAP7_75t_L g1065 ( .A(n_947), .B(n_213), .Y(n_1065) );
AND2x4_ASAP7_75t_L g1066 ( .A(n_947), .B(n_214), .Y(n_1066) );
OR2x2_ASAP7_75t_L g1067 ( .A(n_935), .B(n_215), .Y(n_1067) );
OR2x2_ASAP7_75t_L g1068 ( .A(n_935), .B(n_217), .Y(n_1068) );
INVx1_ASAP7_75t_L g1069 ( .A(n_929), .Y(n_1069) );
OR2x2_ASAP7_75t_L g1070 ( .A(n_939), .B(n_220), .Y(n_1070) );
OR2x2_ASAP7_75t_L g1071 ( .A(n_939), .B(n_221), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_948), .Y(n_1072) );
OR2x2_ASAP7_75t_L g1073 ( .A(n_940), .B(n_222), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_967), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_987), .B(n_223), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_953), .B(n_224), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_933), .Y(n_1077) );
INVx1_ASAP7_75t_L g1078 ( .A(n_954), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_987), .B(n_225), .Y(n_1079) );
BUFx2_ASAP7_75t_L g1080 ( .A(n_924), .Y(n_1080) );
INVx1_ASAP7_75t_L g1081 ( .A(n_963), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_968), .B(n_226), .Y(n_1082) );
BUFx3_ASAP7_75t_L g1083 ( .A(n_988), .Y(n_1083) );
BUFx2_ASAP7_75t_L g1084 ( .A(n_924), .Y(n_1084) );
INVx2_ASAP7_75t_L g1085 ( .A(n_930), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_964), .Y(n_1086) );
INVx1_ASAP7_75t_L g1087 ( .A(n_926), .Y(n_1087) );
BUFx3_ASAP7_75t_L g1088 ( .A(n_988), .Y(n_1088) );
INVx2_ASAP7_75t_L g1089 ( .A(n_931), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_926), .Y(n_1090) );
BUFx2_ASAP7_75t_L g1091 ( .A(n_943), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1030), .Y(n_1092) );
AND2x2_ASAP7_75t_SL g1093 ( .A(n_949), .B(n_228), .Y(n_1093) );
INVx1_ASAP7_75t_L g1094 ( .A(n_996), .Y(n_1094) );
OR2x2_ASAP7_75t_L g1095 ( .A(n_940), .B(n_229), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_969), .B(n_230), .Y(n_1096) );
INVx1_ASAP7_75t_L g1097 ( .A(n_996), .Y(n_1097) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1018), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_972), .B(n_231), .Y(n_1099) );
INVx2_ASAP7_75t_SL g1100 ( .A(n_988), .Y(n_1100) );
INVx1_ASAP7_75t_L g1101 ( .A(n_983), .Y(n_1101) );
OR2x2_ASAP7_75t_L g1102 ( .A(n_941), .B(n_232), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_983), .Y(n_1103) );
INVx1_ASAP7_75t_L g1104 ( .A(n_932), .Y(n_1104) );
AND2x4_ASAP7_75t_L g1105 ( .A(n_941), .B(n_234), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_959), .B(n_239), .Y(n_1106) );
NAND2xp5_ASAP7_75t_L g1107 ( .A(n_974), .B(n_240), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1019), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1019), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1048), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_959), .B(n_245), .Y(n_1111) );
HB1xp67_ASAP7_75t_L g1112 ( .A(n_950), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_922), .B(n_250), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1055), .Y(n_1114) );
INVx1_ASAP7_75t_SL g1115 ( .A(n_944), .Y(n_1115) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_976), .B(n_251), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1117 ( .A(n_934), .B(n_255), .Y(n_1117) );
OR2x2_ASAP7_75t_L g1118 ( .A(n_1055), .B(n_256), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_951), .B(n_257), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_927), .Y(n_1120) );
AOI21xp33_ASAP7_75t_L g1121 ( .A1(n_1020), .A2(n_258), .B(n_260), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_956), .B(n_261), .Y(n_1122) );
AND2x2_ASAP7_75t_L g1123 ( .A(n_920), .B(n_263), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1124 ( .A(n_925), .B(n_265), .Y(n_1124) );
OR2x2_ASAP7_75t_L g1125 ( .A(n_950), .B(n_268), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_955), .B(n_270), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_955), .B(n_271), .Y(n_1127) );
OR2x2_ASAP7_75t_L g1128 ( .A(n_979), .B(n_274), .Y(n_1128) );
OR2x2_ASAP7_75t_L g1129 ( .A(n_999), .B(n_275), .Y(n_1129) );
AND2x4_ASAP7_75t_SL g1130 ( .A(n_943), .B(n_277), .Y(n_1130) );
INVx1_ASAP7_75t_L g1131 ( .A(n_982), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_975), .B(n_280), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_984), .B(n_282), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1007), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_1010), .B(n_286), .Y(n_1135) );
OR2x2_ASAP7_75t_L g1136 ( .A(n_942), .B(n_289), .Y(n_1136) );
NAND2xp5_ASAP7_75t_SL g1137 ( .A(n_1020), .B(n_290), .Y(n_1137) );
AND2x4_ASAP7_75t_L g1138 ( .A(n_949), .B(n_291), .Y(n_1138) );
NAND2xp5_ASAP7_75t_L g1139 ( .A(n_1006), .B(n_292), .Y(n_1139) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1008), .B(n_294), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_938), .B(n_296), .Y(n_1141) );
INVxp67_ASAP7_75t_SL g1142 ( .A(n_1049), .Y(n_1142) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1049), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_998), .Y(n_1144) );
AND2x4_ASAP7_75t_L g1145 ( .A(n_966), .B(n_300), .Y(n_1145) );
OR2x2_ASAP7_75t_L g1146 ( .A(n_1005), .B(n_305), .Y(n_1146) );
HB1xp67_ASAP7_75t_L g1147 ( .A(n_966), .Y(n_1147) );
CKINVDCx20_ASAP7_75t_R g1148 ( .A(n_923), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_998), .Y(n_1149) );
HB1xp67_ASAP7_75t_L g1150 ( .A(n_1016), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_971), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g1152 ( .A(n_952), .B(n_306), .Y(n_1152) );
OR2x2_ASAP7_75t_L g1153 ( .A(n_1005), .B(n_307), .Y(n_1153) );
INVxp67_ASAP7_75t_SL g1154 ( .A(n_1037), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_971), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_992), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_928), .B(n_310), .Y(n_1157) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_973), .B(n_312), .Y(n_1158) );
INVx2_ASAP7_75t_L g1159 ( .A(n_1047), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_981), .B(n_313), .Y(n_1160) );
HB1xp67_ASAP7_75t_L g1161 ( .A(n_1016), .Y(n_1161) );
INVx2_ASAP7_75t_L g1162 ( .A(n_1050), .Y(n_1162) );
OR2x2_ASAP7_75t_L g1163 ( .A(n_1037), .B(n_958), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1164 ( .A(n_970), .B(n_317), .Y(n_1164) );
OR2x2_ASAP7_75t_L g1165 ( .A(n_994), .B(n_318), .Y(n_1165) );
INVx1_ASAP7_75t_L g1166 ( .A(n_993), .Y(n_1166) );
INVx2_ASAP7_75t_L g1167 ( .A(n_1051), .Y(n_1167) );
NAND2x1_ASAP7_75t_SL g1168 ( .A(n_1133), .B(n_921), .Y(n_1168) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1069), .Y(n_1169) );
INVx2_ASAP7_75t_L g1170 ( .A(n_1058), .Y(n_1170) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1078), .Y(n_1171) );
NAND2xp5_ASAP7_75t_L g1172 ( .A(n_1101), .B(n_1001), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1103), .B(n_1004), .Y(n_1173) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1072), .Y(n_1174) );
NAND2xp5_ASAP7_75t_L g1175 ( .A(n_1087), .B(n_1023), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1058), .B(n_1041), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1112), .B(n_965), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1090), .B(n_965), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1131), .B(n_962), .Y(n_1179) );
OR2x2_ASAP7_75t_L g1180 ( .A(n_1114), .B(n_1014), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1081), .B(n_962), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1074), .Y(n_1182) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1077), .Y(n_1183) );
OR2x2_ASAP7_75t_L g1184 ( .A(n_1142), .B(n_1036), .Y(n_1184) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1086), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1104), .B(n_1036), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1143), .B(n_997), .Y(n_1187) );
NAND2xp5_ASAP7_75t_L g1188 ( .A(n_1098), .B(n_1027), .Y(n_1188) );
INVx2_ASAP7_75t_L g1189 ( .A(n_1162), .Y(n_1189) );
NAND2xp5_ASAP7_75t_SL g1190 ( .A(n_1093), .B(n_1025), .Y(n_1190) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1098), .B(n_1022), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1092), .Y(n_1192) );
AND2x2_ASAP7_75t_SL g1193 ( .A(n_1138), .B(n_1025), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1147), .B(n_997), .Y(n_1194) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1150), .B(n_1012), .Y(n_1195) );
OR2x2_ASAP7_75t_L g1196 ( .A(n_1154), .B(n_1012), .Y(n_1196) );
NAND2xp5_ASAP7_75t_L g1197 ( .A(n_1110), .B(n_1043), .Y(n_1197) );
OR2x6_ASAP7_75t_L g1198 ( .A(n_1138), .B(n_1035), .Y(n_1198) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1110), .B(n_985), .Y(n_1199) );
INVxp67_ASAP7_75t_L g1200 ( .A(n_1161), .Y(n_1200) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1092), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1134), .Y(n_1202) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1167), .Y(n_1203) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1120), .Y(n_1204) );
INVx2_ASAP7_75t_L g1205 ( .A(n_1159), .Y(n_1205) );
INVx3_ASAP7_75t_L g1206 ( .A(n_1105), .Y(n_1206) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1085), .B(n_1052), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1089), .B(n_1053), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1120), .B(n_1009), .Y(n_1209) );
NOR2xp33_ASAP7_75t_SL g1210 ( .A(n_1115), .B(n_995), .Y(n_1210) );
NAND2xp5_ASAP7_75t_SL g1211 ( .A(n_1105), .B(n_1003), .Y(n_1211) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1094), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1213 ( .A(n_1094), .B(n_1046), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1080), .B(n_1011), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1084), .B(n_989), .Y(n_1215) );
NAND2xp5_ASAP7_75t_L g1216 ( .A(n_1097), .B(n_1038), .Y(n_1216) );
HB1xp67_ASAP7_75t_L g1217 ( .A(n_1151), .Y(n_1217) );
INVx2_ASAP7_75t_L g1218 ( .A(n_1156), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1091), .B(n_1039), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1097), .Y(n_1220) );
AND2x4_ASAP7_75t_L g1221 ( .A(n_1108), .B(n_1045), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1163), .B(n_1039), .Y(n_1222) );
INVx2_ASAP7_75t_SL g1223 ( .A(n_1083), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1108), .Y(n_1224) );
OR2x2_ASAP7_75t_L g1225 ( .A(n_1151), .B(n_1042), .Y(n_1225) );
OR2x2_ASAP7_75t_L g1226 ( .A(n_1155), .B(n_1042), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1088), .B(n_991), .Y(n_1227) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1109), .Y(n_1228) );
INVx2_ASAP7_75t_L g1229 ( .A(n_1156), .Y(n_1229) );
HB1xp67_ASAP7_75t_L g1230 ( .A(n_1155), .Y(n_1230) );
OR2x2_ASAP7_75t_L g1231 ( .A(n_1109), .B(n_1056), .Y(n_1231) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1166), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1100), .B(n_1054), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1144), .B(n_1017), .Y(n_1234) );
INVx2_ASAP7_75t_L g1235 ( .A(n_1166), .Y(n_1235) );
INVx2_ASAP7_75t_L g1236 ( .A(n_1196), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1169), .Y(n_1237) );
INVx2_ASAP7_75t_L g1238 ( .A(n_1184), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1200), .B(n_1149), .Y(n_1239) );
INVx3_ASAP7_75t_SL g1240 ( .A(n_1223), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1171), .Y(n_1241) );
NAND2xp5_ASAP7_75t_L g1242 ( .A(n_1186), .B(n_1135), .Y(n_1242) );
INVxp67_ASAP7_75t_L g1243 ( .A(n_1231), .Y(n_1243) );
OR2x2_ASAP7_75t_L g1244 ( .A(n_1200), .B(n_1067), .Y(n_1244) );
AOI22xp5_ASAP7_75t_L g1245 ( .A1(n_1190), .A2(n_1193), .B1(n_1198), .B2(n_1210), .Y(n_1245) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1174), .Y(n_1246) );
INVx2_ASAP7_75t_L g1247 ( .A(n_1194), .Y(n_1247) );
INVx2_ASAP7_75t_L g1248 ( .A(n_1195), .Y(n_1248) );
INVx2_ASAP7_75t_L g1249 ( .A(n_1218), .Y(n_1249) );
NOR2xp33_ASAP7_75t_L g1250 ( .A(n_1168), .B(n_1148), .Y(n_1250) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1182), .Y(n_1251) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1183), .Y(n_1252) );
OR2x2_ASAP7_75t_L g1253 ( .A(n_1217), .B(n_1068), .Y(n_1253) );
INVx2_ASAP7_75t_SL g1254 ( .A(n_1207), .Y(n_1254) );
INVxp67_ASAP7_75t_SL g1255 ( .A(n_1217), .Y(n_1255) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1202), .Y(n_1256) );
AND2x4_ASAP7_75t_L g1257 ( .A(n_1178), .B(n_1066), .Y(n_1257) );
NAND2xp5_ASAP7_75t_L g1258 ( .A(n_1230), .B(n_1146), .Y(n_1258) );
NAND2xp5_ASAP7_75t_L g1259 ( .A(n_1173), .B(n_1126), .Y(n_1259) );
OAI21xp5_ASAP7_75t_L g1260 ( .A1(n_1190), .A2(n_1066), .B(n_1059), .Y(n_1260) );
NAND2xp5_ASAP7_75t_L g1261 ( .A(n_1212), .B(n_1127), .Y(n_1261) );
NAND2xp5_ASAP7_75t_L g1262 ( .A(n_1220), .B(n_1153), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1230), .Y(n_1263) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1185), .Y(n_1264) );
AOI21xp5_ASAP7_75t_L g1265 ( .A1(n_1193), .A2(n_1137), .B(n_1013), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_1224), .B(n_1031), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1214), .B(n_1075), .Y(n_1267) );
NAND2xp5_ASAP7_75t_L g1268 ( .A(n_1228), .B(n_1031), .Y(n_1268) );
BUFx2_ASAP7_75t_L g1269 ( .A(n_1206), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1176), .B(n_1079), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g1271 ( .A(n_1203), .B(n_1063), .Y(n_1271) );
OR2x2_ASAP7_75t_L g1272 ( .A(n_1189), .B(n_1070), .Y(n_1272) );
OR2x2_ASAP7_75t_L g1273 ( .A(n_1205), .B(n_1071), .Y(n_1273) );
NAND2xp5_ASAP7_75t_L g1274 ( .A(n_1179), .B(n_1064), .Y(n_1274) );
NAND4xp25_ASAP7_75t_L g1275 ( .A(n_1210), .B(n_1060), .C(n_1113), .D(n_1123), .Y(n_1275) );
INVx2_ASAP7_75t_L g1276 ( .A(n_1218), .Y(n_1276) );
OAI22xp5_ASAP7_75t_L g1277 ( .A1(n_1245), .A2(n_1198), .B1(n_1206), .B2(n_1211), .Y(n_1277) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1239), .B(n_1181), .Y(n_1278) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1237), .Y(n_1279) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1241), .Y(n_1280) );
OAI21xp5_ASAP7_75t_SL g1281 ( .A1(n_1245), .A2(n_1211), .B(n_1215), .Y(n_1281) );
OAI22xp5_ASAP7_75t_L g1282 ( .A1(n_1240), .A2(n_1198), .B1(n_1125), .B2(n_1118), .Y(n_1282) );
NAND2xp5_ASAP7_75t_L g1283 ( .A(n_1263), .B(n_1187), .Y(n_1283) );
NAND2xp5_ASAP7_75t_L g1284 ( .A(n_1236), .B(n_1222), .Y(n_1284) );
AOI22xp33_ASAP7_75t_L g1285 ( .A1(n_1275), .A2(n_1234), .B1(n_1219), .B2(n_1221), .Y(n_1285) );
AOI22xp33_ASAP7_75t_L g1286 ( .A1(n_1275), .A2(n_1221), .B1(n_1227), .B2(n_1233), .Y(n_1286) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1246), .Y(n_1287) );
INVx1_ASAP7_75t_SL g1288 ( .A(n_1254), .Y(n_1288) );
NOR2x1p5_ASAP7_75t_L g1289 ( .A(n_1255), .B(n_1165), .Y(n_1289) );
INVx2_ASAP7_75t_L g1290 ( .A(n_1249), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1291 ( .A(n_1238), .B(n_1192), .Y(n_1291) );
OAI21xp33_ASAP7_75t_L g1292 ( .A1(n_1250), .A2(n_1177), .B(n_1172), .Y(n_1292) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1251), .Y(n_1293) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1252), .Y(n_1294) );
OAI22xp33_ASAP7_75t_L g1295 ( .A1(n_1260), .A2(n_1095), .B1(n_1073), .B2(n_1102), .Y(n_1295) );
AOI22xp5_ASAP7_75t_L g1296 ( .A1(n_1260), .A2(n_1209), .B1(n_1201), .B2(n_1172), .Y(n_1296) );
O2A1O1Ixp33_ASAP7_75t_L g1297 ( .A1(n_1265), .A2(n_1013), .B(n_957), .C(n_1000), .Y(n_1297) );
INVx2_ASAP7_75t_L g1298 ( .A(n_1276), .Y(n_1298) );
OAI21xp33_ASAP7_75t_L g1299 ( .A1(n_1247), .A2(n_1175), .B(n_1170), .Y(n_1299) );
O2A1O1Ixp5_ASAP7_75t_L g1300 ( .A1(n_1258), .A2(n_1175), .B(n_1188), .C(n_1199), .Y(n_1300) );
OAI211xp5_ASAP7_75t_SL g1301 ( .A1(n_1243), .A2(n_1199), .B(n_1164), .C(n_1226), .Y(n_1301) );
NOR2xp67_ASAP7_75t_L g1302 ( .A(n_1257), .B(n_1229), .Y(n_1302) );
AOI221x1_ASAP7_75t_L g1303 ( .A1(n_1277), .A2(n_1256), .B1(n_1264), .B2(n_1258), .C(n_1266), .Y(n_1303) );
NOR3xp33_ASAP7_75t_L g1304 ( .A(n_1277), .B(n_1121), .C(n_1116), .Y(n_1304) );
OAI22xp5_ASAP7_75t_L g1305 ( .A1(n_1285), .A2(n_1269), .B1(n_1257), .B2(n_1248), .Y(n_1305) );
AOI22xp33_ASAP7_75t_SL g1306 ( .A1(n_1288), .A2(n_1267), .B1(n_1270), .B2(n_1242), .Y(n_1306) );
AOI22xp5_ASAP7_75t_L g1307 ( .A1(n_1281), .A2(n_1259), .B1(n_1274), .B2(n_1271), .Y(n_1307) );
OAI22xp33_ASAP7_75t_L g1308 ( .A1(n_1302), .A2(n_1253), .B1(n_1244), .B2(n_1272), .Y(n_1308) );
OAI22xp5_ASAP7_75t_L g1309 ( .A1(n_1286), .A2(n_1261), .B1(n_1273), .B2(n_1262), .Y(n_1309) );
OAI221xp5_ASAP7_75t_L g1310 ( .A1(n_1292), .A2(n_1268), .B1(n_1266), .B2(n_1225), .C(n_1188), .Y(n_1310) );
AOI222xp33_ASAP7_75t_L g1311 ( .A1(n_1282), .A2(n_1232), .B1(n_1204), .B2(n_1268), .C1(n_1197), .C2(n_1235), .Y(n_1311) );
O2A1O1Ixp33_ASAP7_75t_L g1312 ( .A1(n_1297), .A2(n_990), .B(n_1062), .C(n_1107), .Y(n_1312) );
OR2x2_ASAP7_75t_L g1313 ( .A(n_1291), .B(n_1180), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1296), .B(n_1208), .Y(n_1314) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1279), .Y(n_1315) );
A2O1A1Ixp33_ASAP7_75t_L g1316 ( .A1(n_1300), .A2(n_1158), .B(n_1061), .C(n_1130), .Y(n_1316) );
AOI221xp5_ASAP7_75t_L g1317 ( .A1(n_1301), .A2(n_1197), .B1(n_1213), .B2(n_1191), .C(n_1216), .Y(n_1317) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1280), .Y(n_1318) );
INVx2_ASAP7_75t_L g1319 ( .A(n_1290), .Y(n_1319) );
AO21x1_ASAP7_75t_L g1320 ( .A1(n_1305), .A2(n_1282), .B(n_1295), .Y(n_1320) );
AOI21xp5_ASAP7_75t_L g1321 ( .A1(n_1303), .A2(n_1299), .B(n_1294), .Y(n_1321) );
NOR2xp33_ASAP7_75t_R g1322 ( .A(n_1313), .B(n_1124), .Y(n_1322) );
NAND4xp25_ASAP7_75t_L g1323 ( .A(n_1304), .B(n_1152), .C(n_1111), .D(n_1106), .Y(n_1323) );
AOI21xp5_ASAP7_75t_L g1324 ( .A1(n_1316), .A2(n_1293), .B(n_1287), .Y(n_1324) );
OAI22xp5_ASAP7_75t_L g1325 ( .A1(n_1306), .A2(n_1289), .B1(n_1278), .B2(n_1284), .Y(n_1325) );
OAI21xp33_ASAP7_75t_L g1326 ( .A1(n_1311), .A2(n_1283), .B(n_1298), .Y(n_1326) );
AOI222xp33_ASAP7_75t_L g1327 ( .A1(n_1309), .A2(n_1213), .B1(n_1191), .B2(n_1216), .C1(n_1065), .C2(n_1229), .Y(n_1327) );
AOI21xp5_ASAP7_75t_L g1328 ( .A1(n_1312), .A2(n_1145), .B(n_1057), .Y(n_1328) );
AOI211xp5_ASAP7_75t_L g1329 ( .A1(n_1308), .A2(n_1141), .B(n_1136), .C(n_1160), .Y(n_1329) );
NOR2xp33_ASAP7_75t_L g1330 ( .A(n_1307), .B(n_990), .Y(n_1330) );
AOI221xp5_ASAP7_75t_SL g1331 ( .A1(n_1310), .A2(n_1157), .B1(n_1076), .B2(n_1029), .C(n_1026), .Y(n_1331) );
AOI21xp33_ASAP7_75t_SL g1332 ( .A1(n_1325), .A2(n_1311), .B(n_1318), .Y(n_1332) );
NOR4xp25_ASAP7_75t_L g1333 ( .A(n_1326), .B(n_1315), .C(n_1314), .D(n_1319), .Y(n_1333) );
NAND4xp25_ASAP7_75t_L g1334 ( .A(n_1331), .B(n_1320), .C(n_1329), .D(n_1321), .Y(n_1334) );
NOR3xp33_ASAP7_75t_SL g1335 ( .A(n_1323), .B(n_1317), .C(n_1021), .Y(n_1335) );
INVxp67_ASAP7_75t_L g1336 ( .A(n_1330), .Y(n_1336) );
AOI211xp5_ASAP7_75t_L g1337 ( .A1(n_1324), .A2(n_1129), .B(n_1040), .C(n_1145), .Y(n_1337) );
NOR2xp33_ASAP7_75t_SL g1338 ( .A(n_1328), .B(n_1082), .Y(n_1338) );
NAND3xp33_ASAP7_75t_SL g1339 ( .A(n_1322), .B(n_1024), .C(n_961), .Y(n_1339) );
NAND3xp33_ASAP7_75t_SL g1340 ( .A(n_1333), .B(n_1327), .C(n_1024), .Y(n_1340) );
NOR3x1_ASAP7_75t_L g1341 ( .A(n_1334), .B(n_1128), .C(n_1139), .Y(n_1341) );
NOR2x1_ASAP7_75t_L g1342 ( .A(n_1339), .B(n_1032), .Y(n_1342) );
NOR2x1_ASAP7_75t_L g1343 ( .A(n_1335), .B(n_986), .Y(n_1343) );
OAI211xp5_ASAP7_75t_SL g1344 ( .A1(n_1336), .A2(n_936), .B(n_1015), .C(n_1044), .Y(n_1344) );
NAND3xp33_ASAP7_75t_SL g1345 ( .A(n_1332), .B(n_1132), .C(n_1096), .Y(n_1345) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1342), .Y(n_1346) );
NAND4xp75_ASAP7_75t_L g1347 ( .A(n_1341), .B(n_1338), .C(n_1337), .D(n_1099), .Y(n_1347) );
NOR2xp33_ASAP7_75t_L g1348 ( .A(n_1345), .B(n_1140), .Y(n_1348) );
AOI22xp5_ASAP7_75t_L g1349 ( .A1(n_1340), .A2(n_978), .B1(n_960), .B2(n_1117), .Y(n_1349) );
NOR3xp33_ASAP7_75t_L g1350 ( .A(n_1343), .B(n_936), .C(n_1002), .Y(n_1350) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1346), .Y(n_1351) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1348), .Y(n_1352) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1349), .Y(n_1353) );
INVx2_ASAP7_75t_L g1354 ( .A(n_1347), .Y(n_1354) );
INVx3_ASAP7_75t_L g1355 ( .A(n_1354), .Y(n_1355) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1351), .Y(n_1356) );
NAND2x1_ASAP7_75t_L g1357 ( .A(n_1352), .B(n_1350), .Y(n_1357) );
NAND2xp5_ASAP7_75t_L g1358 ( .A(n_1353), .B(n_1122), .Y(n_1358) );
AOI21xp5_ASAP7_75t_L g1359 ( .A1(n_1355), .A2(n_1344), .B(n_1015), .Y(n_1359) );
AOI21xp5_ASAP7_75t_L g1360 ( .A1(n_1356), .A2(n_1119), .B(n_1028), .Y(n_1360) );
NOR2xp67_ASAP7_75t_SL g1361 ( .A(n_1358), .B(n_1033), .Y(n_1361) );
INVx2_ASAP7_75t_L g1362 ( .A(n_1361), .Y(n_1362) );
NAND2xp5_ASAP7_75t_L g1363 ( .A(n_1359), .B(n_1357), .Y(n_1363) );
XNOR2xp5_ASAP7_75t_L g1364 ( .A(n_1360), .B(n_320), .Y(n_1364) );
AOI21xp5_ASAP7_75t_L g1365 ( .A1(n_1363), .A2(n_1044), .B(n_1034), .Y(n_1365) );
NAND3xp33_ASAP7_75t_L g1366 ( .A(n_1364), .B(n_1034), .C(n_322), .Y(n_1366) );
AOI222xp33_ASAP7_75t_L g1367 ( .A1(n_1362), .A2(n_1034), .B1(n_328), .B2(n_329), .C1(n_331), .C2(n_333), .Y(n_1367) );
NAND2x1_ASAP7_75t_L g1368 ( .A(n_1366), .B(n_321), .Y(n_1368) );
AOI22xp33_ASAP7_75t_SL g1369 ( .A1(n_1365), .A2(n_335), .B1(n_336), .B2(n_337), .Y(n_1369) );
AOI21xp33_ASAP7_75t_L g1370 ( .A1(n_1367), .A2(n_339), .B(n_340), .Y(n_1370) );
NOR2x1_ASAP7_75t_L g1371 ( .A(n_1368), .B(n_341), .Y(n_1371) );
NAND2xp5_ASAP7_75t_L g1372 ( .A(n_1369), .B(n_342), .Y(n_1372) );
OR2x6_ASAP7_75t_L g1373 ( .A(n_1370), .B(n_343), .Y(n_1373) );
AOI22xp33_ASAP7_75t_L g1374 ( .A1(n_1373), .A2(n_1372), .B1(n_1371), .B2(n_347), .Y(n_1374) );
endmodule