module fake_jpeg_17839_n_40 (n_3, n_2, n_1, n_0, n_4, n_5, n_40);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_3),
.B(n_1),
.Y(n_8)
);

BUFx5_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

AOI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_13),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_14),
.A2(n_5),
.B1(n_12),
.B2(n_7),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_16),
.Y(n_27)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_17),
.B(n_18),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_2),
.Y(n_18)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_10),
.Y(n_19)
);

NAND2x1_ASAP7_75t_SL g24 ( 
.A(n_19),
.B(n_20),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_2),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_5),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_17),
.A2(n_15),
.B1(n_18),
.B2(n_16),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_26),
.C(n_11),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_28),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_9),
.C(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_26),
.C(n_22),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_25),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_34),
.C(n_35),
.Y(n_36)
);

AND2x6_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

AOI222xp33_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_36),
.B1(n_31),
.B2(n_32),
.C1(n_24),
.C2(n_19),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_18),
.B(n_20),
.Y(n_40)
);


endmodule