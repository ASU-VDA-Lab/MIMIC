module fake_jpeg_29715_n_424 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_424);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_424;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_20),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_51),
.B(n_52),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_28),
.B(n_50),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_33),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_57),
.B(n_68),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_28),
.B(n_20),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_31),
.B(n_9),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_89),
.Y(n_107)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_86),
.Y(n_126)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_62),
.A2(n_49),
.B1(n_50),
.B2(n_47),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_94),
.A2(n_99),
.B1(n_106),
.B2(n_131),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_63),
.A2(n_49),
.B1(n_47),
.B2(n_31),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_67),
.A2(n_49),
.B1(n_38),
.B2(n_48),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_58),
.A2(n_38),
.B1(n_25),
.B2(n_27),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_122),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_23),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_23),
.Y(n_152)
);

NOR2x1_ASAP7_75t_R g122 ( 
.A(n_84),
.B(n_29),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_70),
.A2(n_48),
.B1(n_40),
.B2(n_41),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_53),
.A2(n_43),
.B(n_27),
.C(n_41),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_110),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_64),
.A2(n_45),
.B1(n_40),
.B2(n_48),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_134),
.A2(n_45),
.B1(n_69),
.B2(n_56),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_107),
.A2(n_134),
.B1(n_89),
.B2(n_83),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_135),
.A2(n_136),
.B1(n_161),
.B2(n_45),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_90),
.A2(n_80),
.B1(n_79),
.B2(n_71),
.Y(n_136)
);

AO22x1_ASAP7_75t_L g137 ( 
.A1(n_95),
.A2(n_56),
.B1(n_54),
.B2(n_72),
.Y(n_137)
);

OR2x4_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_158),
.Y(n_176)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_139),
.B(n_141),
.Y(n_188)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_140),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_124),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_142),
.Y(n_196)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_144),
.B(n_152),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_146),
.A2(n_117),
.B1(n_109),
.B2(n_34),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_101),
.Y(n_149)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_151),
.Y(n_180)
);

INVx11_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_154),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_93),
.B(n_44),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_160),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_157),
.Y(n_192)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_111),
.A2(n_43),
.B1(n_75),
.B2(n_73),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_159),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_128),
.B(n_126),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_117),
.A2(n_61),
.B1(n_65),
.B2(n_82),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_113),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_133),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_166),
.B(n_119),
.Y(n_182)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_167),
.A2(n_168),
.B1(n_108),
.B2(n_147),
.Y(n_178)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_120),
.Y(n_177)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

BUFx2_ASAP7_75t_SL g206 ( 
.A(n_178),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_181),
.A2(n_187),
.B1(n_161),
.B2(n_149),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_182),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_110),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_185),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_137),
.A2(n_118),
.B1(n_92),
.B2(n_108),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_184),
.A2(n_191),
.B1(n_195),
.B2(n_148),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_160),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_137),
.A2(n_127),
.B1(n_55),
.B2(n_113),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_150),
.A2(n_44),
.B1(n_34),
.B2(n_46),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_150),
.A2(n_29),
.B(n_36),
.C(n_46),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_197),
.B(n_150),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_160),
.C(n_135),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_198),
.B(n_216),
.C(n_179),
.Y(n_236)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_199),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_200),
.A2(n_203),
.B1(n_180),
.B2(n_173),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_176),
.A2(n_143),
.B1(n_164),
.B2(n_159),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_205),
.Y(n_232)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_171),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_211),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_165),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_214),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_176),
.A2(n_140),
.B1(n_142),
.B2(n_136),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_209),
.A2(n_210),
.B1(n_213),
.B2(n_218),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_176),
.A2(n_91),
.B1(n_130),
.B2(n_101),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_172),
.Y(n_212)
);

INVxp33_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_181),
.A2(n_158),
.B1(n_103),
.B2(n_125),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_138),
.Y(n_214)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_172),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_186),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_169),
.C(n_156),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_190),
.A2(n_125),
.B1(n_130),
.B2(n_129),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_219),
.A2(n_187),
.B1(n_190),
.B2(n_182),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_171),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_220),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_222),
.A2(n_226),
.B1(n_231),
.B2(n_233),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_219),
.A2(n_192),
.B1(n_189),
.B2(n_197),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_192),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_229),
.Y(n_245)
);

MAJx2_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_188),
.C(n_197),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_228),
.B(n_236),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_208),
.A2(n_195),
.B1(n_188),
.B2(n_175),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_201),
.A2(n_189),
.B1(n_186),
.B2(n_91),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_209),
.A2(n_103),
.B1(n_129),
.B2(n_157),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_235),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_201),
.B(n_180),
.Y(n_237)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_237),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_205),
.A2(n_193),
.B(n_179),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_238),
.A2(n_220),
.B(n_196),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_217),
.B(n_20),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_239),
.B(n_9),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_204),
.A2(n_153),
.B1(n_170),
.B2(n_173),
.Y(n_241)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_241),
.Y(n_248)
);

AND2x2_ASAP7_75t_SL g242 ( 
.A(n_214),
.B(n_196),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_242),
.Y(n_253)
);

BUFx24_ASAP7_75t_SL g244 ( 
.A(n_239),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_246),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_217),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_198),
.C(n_216),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_251),
.C(n_252),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_193),
.C(n_206),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_210),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_263),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_218),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_259),
.Y(n_273)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_206),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_260),
.A2(n_211),
.B(n_207),
.Y(n_293)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_261),
.Y(n_286)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_262),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_225),
.B(n_194),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_194),
.C(n_199),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_266),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_224),
.C(n_242),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_194),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_243),
.Y(n_281)
);

OAI22x1_ASAP7_75t_SL g268 ( 
.A1(n_226),
.A2(n_212),
.B1(n_215),
.B2(n_173),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_268),
.A2(n_212),
.B1(n_170),
.B2(n_234),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_222),
.B(n_215),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_269),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_247),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_272),
.B(n_262),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_249),
.A2(n_230),
.B1(n_221),
.B2(n_229),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_274),
.A2(n_275),
.B1(n_282),
.B2(n_248),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_249),
.A2(n_221),
.B1(n_224),
.B2(n_242),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_260),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_279),
.B(n_259),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_281),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_255),
.A2(n_233),
.B1(n_226),
.B2(n_241),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_247),
.B(n_222),
.Y(n_283)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

OAI21xp33_ASAP7_75t_L g284 ( 
.A1(n_245),
.A2(n_243),
.B(n_240),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_284),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_231),
.Y(n_285)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_285),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_231),
.Y(n_287)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_287),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_268),
.A2(n_235),
.B(n_223),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_289),
.A2(n_154),
.B(n_151),
.Y(n_312)
);

XOR2x1_ASAP7_75t_L g290 ( 
.A(n_252),
.B(n_235),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_290),
.B(n_29),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_253),
.B(n_245),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_291),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_248),
.A2(n_223),
.B1(n_235),
.B2(n_240),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_292),
.A2(n_294),
.B1(n_257),
.B2(n_272),
.Y(n_300)
);

A2O1A1Ixp33_ASAP7_75t_SL g316 ( 
.A1(n_293),
.A2(n_168),
.B(n_54),
.C(n_66),
.Y(n_316)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_261),
.Y(n_295)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_295),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_250),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_296),
.B(n_301),
.C(n_304),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_299),
.A2(n_294),
.B1(n_286),
.B2(n_288),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_300),
.A2(n_282),
.B1(n_275),
.B2(n_274),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_251),
.C(n_264),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_302),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_271),
.B(n_264),
.C(n_256),
.Y(n_304)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_265),
.Y(n_306)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_306),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_270),
.B(n_267),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_308),
.Y(n_329)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_277),
.Y(n_309)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_309),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_273),
.B(n_255),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_310),
.B(n_311),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_277),
.B(n_163),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_312),
.A2(n_316),
.B(n_319),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_314),
.B(n_320),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_280),
.B(n_48),
.C(n_40),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_318),
.B(n_59),
.C(n_35),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_279),
.A2(n_283),
.B(n_278),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_280),
.B(n_40),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_297),
.A2(n_278),
.B1(n_290),
.B2(n_292),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_321),
.A2(n_325),
.B1(n_340),
.B2(n_316),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_323),
.B(n_324),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_300),
.A2(n_285),
.B1(n_287),
.B2(n_295),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_298),
.A2(n_288),
.B1(n_286),
.B2(n_281),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_326),
.B(n_331),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_319),
.A2(n_289),
.B1(n_293),
.B2(n_276),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_332),
.B(n_320),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_307),
.A2(n_10),
.B1(n_19),
.B2(n_17),
.Y(n_333)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_333),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_315),
.A2(n_303),
.B1(n_305),
.B2(n_299),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_334),
.B(n_339),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_309),
.A2(n_8),
.B1(n_16),
.B2(n_14),
.Y(n_337)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_337),
.Y(n_347)
);

INVx11_ASAP7_75t_L g338 ( 
.A(n_316),
.Y(n_338)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_338),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_313),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_310),
.A2(n_12),
.B1(n_11),
.B2(n_9),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_301),
.B(n_296),
.C(n_304),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_343),
.B(n_318),
.C(n_314),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_344),
.B(n_356),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_329),
.B(n_317),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_348),
.B(n_352),
.Y(n_367)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_341),
.Y(n_351)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_351),
.Y(n_372)
);

O2A1O1Ixp33_ASAP7_75t_L g352 ( 
.A1(n_330),
.A2(n_312),
.B(n_313),
.C(n_306),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_326),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_354),
.B(n_321),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_355),
.B(n_342),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_336),
.B(n_311),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_356),
.B(n_359),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_327),
.B(n_316),
.C(n_35),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_357),
.B(n_360),
.C(n_361),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_358),
.A2(n_330),
.B1(n_323),
.B2(n_331),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_336),
.B(n_12),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_327),
.B(n_35),
.C(n_11),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_343),
.B(n_35),
.C(n_11),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_362),
.B(n_364),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_347),
.A2(n_338),
.B1(n_335),
.B2(n_325),
.Y(n_363)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_363),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_346),
.B(n_328),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_365),
.A2(n_353),
.B1(n_358),
.B2(n_340),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_355),
.B(n_328),
.C(n_334),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_368),
.B(n_357),
.C(n_359),
.Y(n_378)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_369),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_370),
.B(n_344),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_360),
.B(n_339),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_371),
.B(n_375),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_349),
.A2(n_322),
.B(n_341),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_373),
.A2(n_367),
.B(n_372),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_350),
.B(n_322),
.Y(n_375)
);

FAx1_ASAP7_75t_L g377 ( 
.A(n_365),
.B(n_350),
.CI(n_345),
.CON(n_377),
.SN(n_377)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_377),
.B(n_378),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_370),
.B(n_361),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_379),
.B(n_380),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_380),
.B(n_384),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_368),
.B(n_345),
.C(n_324),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_381),
.B(n_383),
.Y(n_390)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_382),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_366),
.B(n_353),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_385),
.A2(n_366),
.B1(n_352),
.B2(n_374),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_388),
.B(n_377),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_386),
.B(n_374),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_391),
.B(n_396),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_392),
.B(n_35),
.C(n_36),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_376),
.A2(n_332),
.B(n_342),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_393),
.A2(n_398),
.B(n_378),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_381),
.B(n_7),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_394),
.Y(n_406)
);

BUFx24_ASAP7_75t_SL g396 ( 
.A(n_377),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_387),
.A2(n_7),
.B(n_1),
.Y(n_398)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_400),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_397),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_401),
.B(n_402),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_395),
.A2(n_0),
.B(n_1),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_403),
.B(n_404),
.Y(n_412)
);

NOR3xp33_ASAP7_75t_SL g404 ( 
.A(n_390),
.B(n_0),
.C(n_1),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_389),
.A2(n_0),
.B(n_2),
.Y(n_405)
);

A2O1A1O1Ixp25_ASAP7_75t_L g413 ( 
.A1(n_405),
.A2(n_3),
.B(n_4),
.C(n_5),
.D(n_6),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_407),
.B(n_394),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_410),
.A2(n_411),
.B(n_413),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_401),
.A2(n_389),
.B1(n_4),
.B2(n_5),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_408),
.A2(n_399),
.B(n_406),
.Y(n_415)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_415),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_409),
.A2(n_3),
.B(n_4),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_416),
.A2(n_417),
.B(n_6),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_412),
.A2(n_5),
.B(n_6),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_418),
.B(n_414),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_420),
.B(n_419),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_421),
.A2(n_36),
.B(n_35),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_422),
.B(n_36),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_423),
.A2(n_36),
.B(n_6),
.Y(n_424)
);


endmodule