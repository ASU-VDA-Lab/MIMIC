module real_jpeg_30427_n_13 (n_8, n_116, n_0, n_2, n_114, n_10, n_9, n_12, n_6, n_121, n_11, n_112, n_120, n_7, n_117, n_3, n_119, n_5, n_4, n_115, n_122, n_1, n_118, n_113, n_13);

input n_8;
input n_116;
input n_0;
input n_2;
input n_114;
input n_10;
input n_9;
input n_12;
input n_6;
input n_121;
input n_11;
input n_112;
input n_120;
input n_7;
input n_117;
input n_3;
input n_119;
input n_5;
input n_4;
input n_115;
input n_122;
input n_1;
input n_118;
input n_113;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

AOI322xp5_ASAP7_75t_L g105 ( 
.A1(n_0),
.A2(n_36),
.A3(n_38),
.B1(n_44),
.B2(n_106),
.C1(n_108),
.C2(n_122),
.Y(n_105)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_1),
.B(n_46),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_2),
.B(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_2),
.Y(n_109)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_4),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g14 ( 
.A1(n_5),
.A2(n_15),
.B1(n_16),
.B2(n_21),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_6),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_7),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_7),
.B(n_96),
.Y(n_107)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_8),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_17),
.Y(n_16)
);

AOI221xp5_ASAP7_75t_L g67 ( 
.A1(n_10),
.A2(n_12),
.B1(n_68),
.B2(n_73),
.C(n_77),
.Y(n_67)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_10),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_11),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_11),
.B(n_54),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_12),
.B(n_68),
.C(n_73),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_22),
.Y(n_13)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI31xp67_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_59),
.A3(n_94),
.B(n_101),
.Y(n_24)
);

NOR3xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_43),
.C(n_53),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_26),
.A2(n_102),
.B(n_105),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_36),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR3xp33_ASAP7_75t_L g106 ( 
.A(n_28),
.B(n_53),
.C(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_29),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_42),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_113),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OA21x2_ASAP7_75t_SL g102 ( 
.A1(n_43),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_52),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2x1_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_88),
.C(n_89),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_81),
.B(n_87),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_67),
.B1(n_79),
.B2(n_80),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_118),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_86),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_86),
.Y(n_87)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_100),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_112),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_114),
.Y(n_47)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_115),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_116),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_117),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_119),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_120),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_121),
.Y(n_97)
);


endmodule