module fake_jpeg_30952_n_497 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_497);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_497;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_4),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_52),
.B(n_55),
.Y(n_126)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_53),
.Y(n_130)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_45),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_58),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_59),
.B(n_62),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_60),
.Y(n_154)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx2_ASAP7_75t_R g153 ( 
.A(n_64),
.Y(n_153)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_67),
.B(n_69),
.Y(n_141)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_8),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_71),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_35),
.B(n_8),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_72),
.B(n_75),
.Y(n_144)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx11_ASAP7_75t_SL g76 ( 
.A(n_19),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_78),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_21),
.B(n_9),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_79),
.B(n_82),
.Y(n_115)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_81),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_18),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g83 ( 
.A(n_17),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_17),
.Y(n_85)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_87),
.Y(n_151)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

AOI21xp33_ASAP7_75t_L g91 ( 
.A1(n_30),
.A2(n_9),
.B(n_1),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_36),
.C(n_31),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_21),
.B(n_10),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_95),
.Y(n_102)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_50),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_96),
.B(n_18),
.Y(n_120)
);

BUFx10_ASAP7_75t_L g97 ( 
.A(n_18),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_98),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_23),
.B(n_10),
.Y(n_98)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_33),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_20),
.B1(n_49),
.B2(n_38),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_101),
.A2(n_105),
.B1(n_113),
.B2(n_57),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_91),
.A2(n_63),
.B1(n_89),
.B2(n_85),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_104),
.A2(n_107),
.B1(n_117),
.B2(n_123),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_99),
.A2(n_20),
.B1(n_49),
.B2(n_38),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_51),
.A2(n_47),
.B1(n_40),
.B2(n_34),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_64),
.A2(n_35),
.B(n_23),
.C(n_34),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_108),
.B(n_112),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_71),
.A2(n_30),
.B1(n_36),
.B2(n_41),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_81),
.A2(n_47),
.B1(n_40),
.B2(n_33),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_116),
.B(n_7),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_L g117 ( 
.A1(n_84),
.A2(n_47),
.B1(n_40),
.B2(n_31),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_93),
.A2(n_41),
.B1(n_32),
.B2(n_33),
.Y(n_123)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_124),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_32),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_136),
.B(n_140),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_97),
.B(n_33),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_56),
.B(n_7),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_142),
.B(n_149),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_53),
.B(n_7),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_66),
.B(n_7),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_155),
.B(n_3),
.Y(n_202)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_156),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_131),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_157),
.B(n_158),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_108),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_159),
.A2(n_145),
.B1(n_137),
.B2(n_132),
.Y(n_210)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_160),
.Y(n_231)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_161),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_139),
.A2(n_60),
.B1(n_80),
.B2(n_73),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_163),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_117),
.A2(n_65),
.B1(n_95),
.B2(n_70),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_164),
.A2(n_204),
.B1(n_205),
.B2(n_154),
.Y(n_214)
);

OR2x2_ASAP7_75t_SL g165 ( 
.A(n_116),
.B(n_76),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_165),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_95),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_166),
.B(n_176),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_139),
.A2(n_58),
.B1(n_2),
.B2(n_3),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_167),
.Y(n_213)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_168),
.Y(n_224)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_169),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_125),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_170),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_115),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_173),
.B(n_181),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_141),
.B(n_11),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_174),
.B(n_190),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_110),
.Y(n_175)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_175),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_126),
.B(n_11),
.Y(n_176)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_177),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_178),
.B(n_183),
.Y(n_248)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_138),
.Y(n_179)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_179),
.Y(n_225)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_106),
.Y(n_180)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_180),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_153),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_102),
.B(n_12),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_153),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_184),
.B(n_186),
.Y(n_249)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_185),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_100),
.B(n_12),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_109),
.B(n_6),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_187),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_112),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_188),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_110),
.Y(n_189)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_189),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_119),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_191),
.Y(n_250)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_192),
.Y(n_251)
);

OA21x2_ASAP7_75t_L g193 ( 
.A1(n_145),
.A2(n_111),
.B(n_122),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_193),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_143),
.Y(n_195)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_195),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_135),
.Y(n_196)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_196),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_129),
.B(n_6),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_199),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_137),
.B(n_13),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_198),
.B(n_202),
.Y(n_235)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_147),
.B(n_13),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_203),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_135),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_111),
.A2(n_122),
.B1(n_114),
.B2(n_151),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_114),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_205)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_138),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_206),
.B(n_154),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_152),
.B(n_4),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_207),
.B(n_208),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_133),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_210),
.B(n_214),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_188),
.A2(n_148),
.B1(n_118),
.B2(n_152),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_217),
.A2(n_223),
.B1(n_189),
.B2(n_15),
.Y(n_295)
);

A2O1A1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_178),
.A2(n_133),
.B(n_127),
.C(n_143),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_219),
.A2(n_238),
.B(n_243),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_127),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_220),
.B(n_228),
.C(n_219),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_158),
.A2(n_190),
.B1(n_182),
.B2(n_162),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_118),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_227),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_125),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_132),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_237),
.B(n_242),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_182),
.B(n_0),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_171),
.B(n_0),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_243),
.B(n_244),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_171),
.B(n_121),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_172),
.B(n_121),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_246),
.B(n_196),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_247),
.Y(n_284)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_250),
.Y(n_255)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_255),
.Y(n_301)
);

AO22x1_ASAP7_75t_SL g256 ( 
.A1(n_223),
.A2(n_162),
.B1(n_172),
.B2(n_165),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_256),
.B(n_265),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_239),
.A2(n_205),
.B1(n_185),
.B2(n_180),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_258),
.A2(n_280),
.B1(n_252),
.B2(n_231),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_259),
.B(n_266),
.Y(n_317)
);

NAND2xp33_ASAP7_75t_SL g260 ( 
.A(n_244),
.B(n_193),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_260),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_212),
.B(n_181),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_261),
.B(n_262),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_212),
.Y(n_262)
);

AO21x2_ASAP7_75t_L g263 ( 
.A1(n_239),
.A2(n_193),
.B(n_170),
.Y(n_263)
);

OA22x2_ASAP7_75t_L g311 ( 
.A1(n_263),
.A2(n_286),
.B1(n_290),
.B2(n_253),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_264),
.B(n_287),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_173),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_232),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_174),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_267),
.B(n_272),
.Y(n_322)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_268),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_222),
.A2(n_198),
.B1(n_157),
.B2(n_195),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_269),
.A2(n_275),
.B(n_216),
.Y(n_320)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_218),
.Y(n_270)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_270),
.Y(n_310)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_271),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_248),
.B(n_208),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_220),
.B(n_191),
.C(n_192),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_273),
.B(n_277),
.C(n_281),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_245),
.A2(n_206),
.B(n_179),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_274),
.A2(n_278),
.B(n_279),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_245),
.A2(n_161),
.B(n_199),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_237),
.B(n_156),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_213),
.A2(n_170),
.B1(n_177),
.B2(n_160),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_222),
.A2(n_213),
.B1(n_214),
.B2(n_227),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_211),
.B(n_169),
.C(n_168),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_238),
.A2(n_234),
.B1(n_210),
.B2(n_240),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_282),
.A2(n_289),
.B1(n_295),
.B2(n_231),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_211),
.B(n_203),
.C(n_196),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_283),
.B(n_225),
.C(n_224),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_217),
.B(n_5),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_209),
.B(n_203),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_291),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_226),
.A2(n_215),
.B1(n_242),
.B2(n_209),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_249),
.B(n_14),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_233),
.B(n_175),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_247),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_293),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_235),
.B(n_175),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_294),
.B(n_16),
.Y(n_331)
);

OAI22x1_ASAP7_75t_L g296 ( 
.A1(n_263),
.A2(n_215),
.B1(n_235),
.B2(n_252),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_296),
.A2(n_306),
.B1(n_276),
.B2(n_281),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_270),
.Y(n_300)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_300),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_264),
.B(n_251),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_303),
.B(n_289),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_305),
.A2(n_312),
.B1(n_313),
.B2(n_323),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_261),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_307),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_261),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_309),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_311),
.B(n_320),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_293),
.A2(n_253),
.B1(n_241),
.B2(n_229),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_284),
.A2(n_241),
.B1(n_229),
.B2(n_236),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_315),
.B(n_299),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_287),
.A2(n_225),
.B(n_224),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_316),
.A2(n_325),
.B(n_263),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_273),
.B(n_254),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_318),
.B(n_328),
.C(n_285),
.Y(n_357)
);

OA21x2_ASAP7_75t_L g321 ( 
.A1(n_263),
.A2(n_254),
.B(n_230),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_321),
.B(n_331),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_280),
.A2(n_230),
.B1(n_236),
.B2(n_218),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_276),
.A2(n_216),
.B1(n_221),
.B2(n_14),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_324),
.A2(n_258),
.B1(n_286),
.B2(n_284),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_265),
.A2(n_274),
.B(n_276),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_291),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_326),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_277),
.B(n_221),
.C(n_14),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_255),
.Y(n_330)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_330),
.Y(n_338)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_268),
.Y(n_332)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_332),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_320),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_334),
.B(n_340),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_335),
.B(n_361),
.C(n_365),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_322),
.B(n_272),
.Y(n_336)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_336),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_337),
.B(n_256),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_312),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_327),
.A2(n_262),
.B(n_269),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_341),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_322),
.B(n_288),
.Y(n_342)
);

CKINVDCx14_ASAP7_75t_R g379 ( 
.A(n_342),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_343),
.A2(n_355),
.B1(n_363),
.B2(n_364),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_314),
.B(n_294),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_345),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_318),
.B(n_257),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_346),
.B(n_357),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_307),
.B(n_267),
.Y(n_347)
);

NAND3xp33_ASAP7_75t_L g390 ( 
.A(n_347),
.B(n_353),
.C(n_317),
.Y(n_390)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_301),
.Y(n_349)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_349),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_309),
.B(n_279),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_327),
.A2(n_274),
.B(n_276),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_354),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_306),
.A2(n_257),
.B1(n_256),
.B2(n_283),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_301),
.Y(n_356)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_356),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_314),
.B(n_290),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_359),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_290),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_362),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_299),
.B(n_292),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_304),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_319),
.B(n_303),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_365),
.B(n_285),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_366),
.B(n_368),
.C(n_370),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_335),
.B(n_361),
.C(n_357),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_340),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_369),
.A2(n_382),
.B1(n_343),
.B2(n_344),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_346),
.B(n_319),
.C(n_315),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_333),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_373),
.B(n_380),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_337),
.B(n_297),
.C(n_292),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_376),
.B(n_328),
.C(n_353),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_377),
.B(n_381),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_352),
.Y(n_378)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_378),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_333),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_351),
.A2(n_298),
.B1(n_324),
.B2(n_321),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_358),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_384),
.B(n_386),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_355),
.A2(n_305),
.B1(n_323),
.B2(n_321),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_385),
.A2(n_394),
.B1(n_367),
.B2(n_351),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_358),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_341),
.B(n_325),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_387),
.B(n_302),
.Y(n_412)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_390),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_363),
.A2(n_308),
.B1(n_295),
.B2(n_313),
.Y(n_394)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_395),
.Y(n_426)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_374),
.Y(n_397)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_397),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_366),
.B(n_350),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_399),
.B(n_408),
.Y(n_422)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_374),
.Y(n_400)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_400),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_401),
.A2(n_406),
.B1(n_409),
.B2(n_410),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_372),
.B(n_344),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_404),
.B(n_407),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_383),
.A2(n_334),
.B(n_350),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_405),
.A2(n_387),
.B(n_311),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_367),
.A2(n_352),
.B1(n_354),
.B2(n_350),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_389),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_394),
.A2(n_385),
.B1(n_389),
.B2(n_371),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_371),
.A2(n_311),
.B1(n_302),
.B2(n_256),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_412),
.B(n_370),
.Y(n_429)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_388),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_413),
.B(n_416),
.Y(n_421)
);

NAND2x1_ASAP7_75t_SL g415 ( 
.A(n_383),
.B(n_311),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_415),
.A2(n_263),
.B(n_275),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_393),
.A2(n_362),
.B1(n_356),
.B2(n_349),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_388),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_417),
.B(n_403),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_368),
.B(n_316),
.C(n_348),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_418),
.B(n_375),
.C(n_377),
.Y(n_431)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_423),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_401),
.A2(n_391),
.B1(n_379),
.B2(n_382),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_424),
.B(n_425),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_403),
.B(n_392),
.Y(n_425)
);

INVx13_ASAP7_75t_L g428 ( 
.A(n_414),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_428),
.B(n_402),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_432),
.Y(n_443)
);

NOR2x1_ASAP7_75t_L g430 ( 
.A(n_406),
.B(n_369),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_430),
.A2(n_435),
.B(n_436),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_431),
.B(n_434),
.Y(n_452)
);

XNOR2x1_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_376),
.Y(n_434)
);

XOR2x2_ASAP7_75t_L g436 ( 
.A(n_415),
.B(n_399),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_398),
.B(n_375),
.C(n_381),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_437),
.B(n_398),
.C(n_408),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_419),
.B(n_411),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_438),
.B(n_441),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_439),
.B(n_434),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_419),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_431),
.A2(n_404),
.B(n_405),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_444),
.A2(n_450),
.B(n_451),
.Y(n_463)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_445),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_424),
.B(n_409),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_446),
.B(n_453),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_437),
.B(n_396),
.C(n_412),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_447),
.B(n_448),
.C(n_429),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_422),
.B(n_396),
.C(n_395),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_435),
.A2(n_407),
.B(n_410),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_426),
.A2(n_417),
.B(n_400),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_422),
.B(n_397),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_442),
.B(n_428),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_454),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_457),
.B(n_462),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_458),
.A2(n_443),
.B(n_339),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_440),
.B(n_420),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_460),
.B(n_466),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_439),
.B(n_420),
.C(n_436),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_461),
.B(n_465),
.C(n_467),
.Y(n_472)
);

AOI21x1_ASAP7_75t_L g462 ( 
.A1(n_449),
.A2(n_432),
.B(n_436),
.Y(n_462)
);

OAI21xp33_ASAP7_75t_L g464 ( 
.A1(n_449),
.A2(n_426),
.B(n_430),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_464),
.A2(n_450),
.B1(n_427),
.B2(n_433),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_448),
.B(n_452),
.C(n_447),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_451),
.B(n_428),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_452),
.B(n_421),
.C(n_430),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_455),
.B(n_433),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_470),
.B(n_475),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_473),
.B(n_474),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_465),
.B(n_443),
.C(n_427),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_463),
.B(n_467),
.Y(n_475)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_476),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_459),
.A2(n_348),
.B1(n_338),
.B2(n_329),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_477),
.B(n_332),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_461),
.B(n_339),
.C(n_338),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_478),
.A2(n_456),
.B(n_464),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_479),
.B(n_481),
.Y(n_489)
);

AOI22xp33_ASAP7_75t_SL g482 ( 
.A1(n_473),
.A2(n_263),
.B1(n_260),
.B2(n_310),
.Y(n_482)
);

CKINVDCx14_ASAP7_75t_R g486 ( 
.A(n_482),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_472),
.A2(n_474),
.B(n_468),
.Y(n_484)
);

AO221x1_ASAP7_75t_L g487 ( 
.A1(n_484),
.A2(n_472),
.B1(n_471),
.B2(n_478),
.C(n_457),
.Y(n_487)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_487),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_483),
.B(n_471),
.C(n_469),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_488),
.B(n_310),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_488),
.B(n_485),
.C(n_480),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_490),
.B(n_492),
.C(n_330),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_491),
.A2(n_489),
.B1(n_486),
.B2(n_482),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_493),
.A2(n_494),
.B(n_304),
.Y(n_495)
);

AOI21xp33_ASAP7_75t_L g496 ( 
.A1(n_495),
.A2(n_329),
.B(n_271),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_496),
.B(n_286),
.Y(n_497)
);


endmodule