module fake_jpeg_4612_n_186 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_186);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_0),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_29),
.A2(n_12),
.B1(n_22),
.B2(n_19),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_32),
.A2(n_23),
.B1(n_15),
.B2(n_14),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_34),
.A2(n_36),
.B(n_37),
.Y(n_57)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_32),
.A2(n_12),
.B1(n_22),
.B2(n_19),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_30),
.A2(n_22),
.B1(n_19),
.B2(n_13),
.Y(n_37)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_45),
.Y(n_64)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_52),
.B1(n_17),
.B2(n_20),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_48),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_29),
.C(n_27),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_24),
.B(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_31),
.B1(n_17),
.B2(n_14),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_13),
.B1(n_23),
.B2(n_15),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_15),
.B1(n_23),
.B2(n_13),
.Y(n_62)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_56),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_33),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_58),
.B(n_40),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_43),
.B1(n_42),
.B2(n_40),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_59),
.A2(n_54),
.B1(n_45),
.B2(n_44),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_46),
.Y(n_83)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_63),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_62),
.Y(n_77)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_67),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_55),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_68),
.A2(n_54),
.B1(n_50),
.B2(n_48),
.Y(n_85)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_60),
.C(n_57),
.Y(n_76)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_74),
.B(n_68),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_83),
.C(n_72),
.Y(n_98)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_81),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_79),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_71),
.B(n_50),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_82),
.Y(n_90)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_57),
.B(n_24),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_78),
.B(n_72),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_74),
.B(n_66),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_96),
.B(n_102),
.Y(n_109)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_93),
.B(n_99),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_66),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_69),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_75),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_95),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_63),
.B(n_51),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_96),
.C(n_97),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_80),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_70),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_103),
.Y(n_112)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_108),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_67),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_118),
.B(n_97),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_95),
.B(n_82),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_107),
.Y(n_123)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

NAND5xp2_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_85),
.C(n_77),
.D(n_61),
.E(n_64),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_92),
.B(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_115),
.Y(n_128)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_117),
.Y(n_129)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_98),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_112),
.B(n_105),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_121),
.A2(n_116),
.B(n_104),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_132),
.C(n_20),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_117),
.A2(n_118),
.B1(n_101),
.B2(n_119),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_125),
.A2(n_127),
.B1(n_108),
.B2(n_105),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_106),
.B(n_93),
.Y(n_126)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_100),
.B1(n_92),
.B2(n_65),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_61),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_20),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_115),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_131),
.B(n_128),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_39),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_27),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_25),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_142),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_137),
.A2(n_140),
.B1(n_145),
.B2(n_122),
.Y(n_153)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_139),
.A2(n_144),
.B(n_128),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_123),
.A2(n_113),
.B1(n_25),
.B2(n_2),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_134),
.B(n_88),
.Y(n_141)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_88),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_146),
.C(n_132),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_88),
.B1(n_21),
.B2(n_16),
.Y(n_145)
);

AO22x1_ASAP7_75t_L g158 ( 
.A1(n_148),
.A2(n_151),
.B1(n_146),
.B2(n_143),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_130),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_121),
.B1(n_139),
.B2(n_129),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_154),
.B1(n_21),
.B2(n_20),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_153),
.B(n_7),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_129),
.B1(n_122),
.B2(n_133),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_7),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_21),
.C(n_31),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_147),
.B(n_120),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_157),
.B(n_160),
.Y(n_169)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_20),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_161),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_163),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_156),
.B(n_20),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_150),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_148),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_5),
.C(n_1),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_151),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_171),
.A2(n_5),
.B(n_1),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_174),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_173),
.B(n_175),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_168),
.A2(n_4),
.B(n_1),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_9),
.C(n_2),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_21),
.Y(n_176)
);

XOR2x2_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_170),
.Y(n_178)
);

AOI322xp5_ASAP7_75t_L g182 ( 
.A1(n_178),
.A2(n_181),
.A3(n_3),
.B1(n_4),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_182)
);

AOI322xp5_ASAP7_75t_L g181 ( 
.A1(n_177),
.A2(n_169),
.A3(n_3),
.B1(n_4),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_182),
.B(n_183),
.Y(n_184)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_179),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_180),
.B1(n_11),
.B2(n_0),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_0),
.Y(n_186)
);


endmodule