module fake_jpeg_22635_n_281 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_281);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_281;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_18),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_7),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_44),
.B(n_19),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_51),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_35),
.B1(n_21),
.B2(n_28),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_60),
.B1(n_62),
.B2(n_72),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_35),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_44),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_27),
.Y(n_57)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_35),
.B1(n_28),
.B2(n_26),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_58),
.A2(n_33),
.B1(n_20),
.B2(n_23),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_31),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_68),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_21),
.B1(n_28),
.B2(n_26),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_24),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_28),
.B1(n_34),
.B2(n_26),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_45),
.A2(n_21),
.B1(n_34),
.B2(n_26),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_34),
.B1(n_31),
.B2(n_32),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_27),
.Y(n_66)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_32),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_27),
.Y(n_71)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_39),
.A2(n_34),
.B1(n_29),
.B2(n_17),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_75),
.B(n_79),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_20),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_88),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_25),
.B1(n_31),
.B2(n_32),
.Y(n_79)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_91),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_69),
.A2(n_25),
.B1(n_30),
.B2(n_17),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_85),
.A2(n_87),
.B1(n_50),
.B2(n_24),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_25),
.B(n_20),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_86),
.A2(n_56),
.B(n_61),
.Y(n_115)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_55),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_42),
.C(n_41),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_45),
.B1(n_42),
.B2(n_41),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_89),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_20),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_99),
.Y(n_109)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_45),
.B1(n_42),
.B2(n_41),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_30),
.B1(n_22),
.B2(n_17),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_48),
.A2(n_30),
.B1(n_22),
.B2(n_33),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_54),
.A2(n_22),
.B1(n_33),
.B2(n_20),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_97),
.B1(n_100),
.B2(n_66),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_20),
.C(n_24),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_0),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_20),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_57),
.A2(n_24),
.B1(n_23),
.B2(n_8),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_103),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_51),
.Y(n_103)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_70),
.Y(n_119)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_24),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_24),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_124),
.B1(n_129),
.B2(n_108),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_115),
.A2(n_132),
.B(n_23),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_13),
.B(n_16),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g153 ( 
.A1(n_118),
.A2(n_133),
.B(n_135),
.Y(n_153)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_65),
.Y(n_120)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_51),
.Y(n_122)
);

NOR2xp67_ASAP7_75t_R g141 ( 
.A(n_122),
.B(n_103),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_123),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_83),
.A2(n_97),
.B1(n_88),
.B2(n_73),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_81),
.B(n_83),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_126),
.B(n_134),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_77),
.B(n_65),
.Y(n_128)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_104),
.A2(n_70),
.B1(n_65),
.B2(n_54),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_78),
.B(n_50),
.Y(n_130)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_80),
.B(n_92),
.Y(n_131)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_81),
.B(n_9),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_63),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_93),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_122),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_162),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_124),
.A2(n_89),
.B1(n_98),
.B2(n_76),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_138),
.A2(n_145),
.B1(n_160),
.B2(n_109),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_148),
.B(n_125),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_112),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_142),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_143),
.A2(n_155),
.B1(n_158),
.B2(n_163),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_89),
.B1(n_102),
.B2(n_91),
.Y(n_145)
);

OAI32xp33_ASAP7_75t_L g146 ( 
.A1(n_109),
.A2(n_99),
.A3(n_90),
.B1(n_89),
.B2(n_93),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_147),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_R g148 ( 
.A(n_122),
.B(n_93),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_84),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_152),
.B(n_119),
.Y(n_184)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_154),
.B(n_159),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_113),
.A2(n_63),
.B1(n_55),
.B2(n_23),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_156),
.A2(n_135),
.B1(n_132),
.B2(n_161),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_111),
.A2(n_63),
.B1(n_55),
.B2(n_23),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_23),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_136),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_110),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_161),
.Y(n_169)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_117),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_111),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_175),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_121),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_167),
.A2(n_149),
.B(n_154),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_168),
.A2(n_170),
.B1(n_173),
.B2(n_181),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_145),
.A2(n_147),
.B1(n_138),
.B2(n_137),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_156),
.A2(n_125),
.B1(n_126),
.B2(n_121),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_174),
.A2(n_157),
.B(n_144),
.Y(n_191)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_183),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_143),
.B(n_135),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_188),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_130),
.Y(n_179)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_163),
.Y(n_180)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_158),
.A2(n_116),
.B1(n_114),
.B2(n_135),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_182),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_157),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_187),
.Y(n_210)
);

OAI21xp33_ASAP7_75t_L g185 ( 
.A1(n_153),
.A2(n_133),
.B(n_134),
.Y(n_185)
);

AOI221xp5_ASAP7_75t_L g211 ( 
.A1(n_185),
.A2(n_10),
.B1(n_13),
.B2(n_6),
.C(n_7),
.Y(n_211)
);

OAI22x1_ASAP7_75t_SL g186 ( 
.A1(n_141),
.A2(n_123),
.B1(n_114),
.B2(n_127),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_186),
.A2(n_139),
.B1(n_151),
.B2(n_4),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_150),
.B(n_127),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_114),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_123),
.C(n_3),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_189),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_198),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_186),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_192),
.Y(n_222)
);

AND5x1_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_150),
.C(n_149),
.D(n_151),
.E(n_140),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_194),
.A2(n_211),
.B1(n_204),
.B2(n_200),
.Y(n_228)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_165),
.Y(n_196)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_173),
.B(n_164),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_169),
.C(n_190),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_205),
.A2(n_175),
.B1(n_182),
.B2(n_166),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_174),
.A2(n_139),
.B(n_3),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_207),
.A2(n_189),
.B1(n_184),
.B2(n_171),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_178),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_208),
.A2(n_209),
.B1(n_176),
.B2(n_180),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_178),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_199),
.B(n_183),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_212),
.B(n_229),
.Y(n_230)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_217),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_219),
.Y(n_241)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_203),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_221),
.C(n_226),
.Y(n_240)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_210),
.Y(n_220)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_177),
.C(n_168),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_223),
.A2(n_225),
.B1(n_227),
.B2(n_228),
.Y(n_234)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_224),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_171),
.C(n_170),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_200),
.A2(n_188),
.B1(n_169),
.B2(n_165),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_196),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_198),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_233),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_193),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_222),
.A2(n_195),
.B1(n_192),
.B2(n_207),
.Y(n_235)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_201),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_237),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_191),
.Y(n_237)
);

AOI31xp67_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_206),
.A3(n_205),
.B(n_195),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_242),
.B(n_235),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_167),
.C(n_209),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_240),
.C(n_218),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_252),
.C(n_253),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_214),
.Y(n_245)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_246),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_248),
.Y(n_256)
);

INVx11_ASAP7_75t_L g248 ( 
.A(n_241),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_213),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_255),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_219),
.C(n_227),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_213),
.C(n_224),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_234),
.C(n_220),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_251),
.A2(n_215),
.B1(n_236),
.B2(n_233),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_262),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_255),
.A2(n_237),
.B1(n_231),
.B2(n_167),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_253),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_262)
);

FAx1_ASAP7_75t_SL g263 ( 
.A(n_252),
.B(n_5),
.CI(n_6),
.CON(n_263),
.SN(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_244),
.C(n_254),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_269),
.C(n_262),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_264),
.B(n_254),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_266),
.B(n_263),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_258),
.B(n_248),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_258),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_257),
.A2(n_250),
.B(n_12),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_268),
.A2(n_256),
.B(n_16),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_250),
.C(n_10),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_270),
.A2(n_261),
.B(n_263),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_271),
.A2(n_272),
.B(n_273),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_275),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_265),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_260),
.C(n_276),
.Y(n_279)
);

BUFx24_ASAP7_75t_SL g280 ( 
.A(n_279),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_277),
.Y(n_281)
);


endmodule