module fake_aes_3565_n_25 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_25);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_25;
wire n_20;
wire n_23;
wire n_22;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
AND2x2_ASAP7_75t_L g12 ( .A(n_4), .B(n_11), .Y(n_12) );
INVx3_ASAP7_75t_L g13 ( .A(n_0), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_9), .B(n_8), .Y(n_14) );
AND2x4_ASAP7_75t_L g15 ( .A(n_6), .B(n_5), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_13), .Y(n_16) );
OA21x2_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_15), .B(n_14), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_18), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_19), .B(n_17), .Y(n_20) );
OAI21xp5_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_15), .B(n_12), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
OAI22x1_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_23) );
OAI22xp5_ASAP7_75t_SL g24 ( .A1(n_23), .A2(n_3), .B1(n_7), .B2(n_10), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
endmodule