module real_jpeg_7736_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

HAxp5_ASAP7_75t_SL g12 ( 
.A(n_1),
.B(n_8),
.CON(n_12),
.SN(n_12)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

OR2x2_ASAP7_75t_SL g27 ( 
.A(n_1),
.B(n_3),
.Y(n_27)
);

OA21x2_ASAP7_75t_L g8 ( 
.A1(n_2),
.A2(n_9),
.B(n_10),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_2),
.B(n_9),
.Y(n_10)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_25),
.Y(n_31)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

AOI211xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_13),
.B(n_26),
.C(n_28),
.Y(n_6)
);

OAI21xp5_ASAP7_75t_SL g7 ( 
.A1(n_8),
.A2(n_11),
.B(n_12),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_8),
.B(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g15 ( 
.A1(n_9),
.A2(n_16),
.B(n_24),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_9),
.B(n_16),
.Y(n_24)
);

BUFx24_ASAP7_75t_SL g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_25),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

OA21x2_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B(n_23),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_22),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);


endmodule