module real_aes_2455_n_382 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_382);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_382;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_577;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_852;
wire n_766;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_571;
wire n_1034;
wire n_549;
wire n_491;
wire n_694;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_989;
wire n_773;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_856;
wire n_594;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_678;
wire n_427;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_994;
wire n_744;
wire n_384;
wire n_938;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_1049;
wire n_466;
wire n_636;
wire n_559;
wire n_872;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_904;
wire n_683;
wire n_570;
wire n_675;
wire n_840;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_1025;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_671;
wire n_973;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_867;
wire n_745;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_417;
wire n_754;
wire n_607;
wire n_449;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_947;
wire n_970;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_617;
wire n_402;
wire n_733;
wire n_552;
wire n_602;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1037;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_999;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_985;
wire n_777;
wire n_488;
wire n_501;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_898;
wire n_734;
wire n_604;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_1003;
wire n_1028;
wire n_1000;
wire n_533;
wire n_727;
wire n_1014;
wire n_397;
wire n_749;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_915;
wire n_470;
wire n_851;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_845;
wire n_850;
wire n_1043;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_928;
wire n_637;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_623;
wire n_1032;
wire n_721;
wire n_446;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_639;
wire n_587;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1036;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1024;
wire n_842;
wire n_849;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_0), .A2(n_333), .B1(n_529), .B2(n_530), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_1), .A2(n_218), .B1(n_536), .B2(n_571), .Y(n_570) );
AOI22xp33_ASAP7_75t_SL g799 ( .A1(n_2), .A2(n_276), .B1(n_553), .B2(n_592), .Y(n_799) );
AOI22xp33_ASAP7_75t_SL g812 ( .A1(n_3), .A2(n_170), .B1(n_680), .B2(n_681), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_4), .A2(n_122), .B1(n_548), .B2(n_584), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g1039 ( .A1(n_5), .A2(n_317), .B1(n_546), .B2(n_548), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_6), .A2(n_129), .B1(n_606), .B2(n_793), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g874 ( .A(n_7), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_8), .B(n_515), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g1038 ( .A(n_9), .Y(n_1038) );
AOI22xp33_ASAP7_75t_SL g923 ( .A1(n_10), .A2(n_255), .B1(n_529), .B2(n_530), .Y(n_923) );
AOI22xp5_ASAP7_75t_L g974 ( .A1(n_11), .A2(n_50), .B1(n_548), .B2(n_584), .Y(n_974) );
AOI22xp5_ASAP7_75t_L g891 ( .A1(n_12), .A2(n_98), .B1(n_447), .B2(n_521), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_13), .A2(n_283), .B1(n_610), .B2(n_623), .Y(n_1024) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_14), .A2(n_364), .B1(n_667), .B2(n_765), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_15), .A2(n_200), .B1(n_538), .B2(n_539), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_16), .A2(n_237), .B1(n_896), .B2(n_898), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_17), .A2(n_82), .B1(n_482), .B2(n_980), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_18), .A2(n_103), .B1(n_621), .B2(n_696), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_19), .A2(n_145), .B1(n_554), .B2(n_670), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_20), .A2(n_329), .B1(n_603), .B2(n_900), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_21), .A2(n_192), .B1(n_428), .B2(n_584), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_22), .A2(n_84), .B1(n_630), .B2(n_744), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_23), .A2(n_182), .B1(n_492), .B2(n_600), .Y(n_1027) );
AOI22xp33_ASAP7_75t_SL g926 ( .A1(n_24), .A2(n_180), .B1(n_536), .B2(n_868), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_25), .A2(n_352), .B1(n_662), .B2(n_749), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_26), .A2(n_156), .B1(n_557), .B2(n_668), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_27), .A2(n_65), .B1(n_553), .B2(n_554), .Y(n_987) );
XOR2x2_ASAP7_75t_L g930 ( .A(n_28), .B(n_931), .Y(n_930) );
AO222x2_ASAP7_75t_L g877 ( .A1(n_29), .A2(n_151), .B1(n_239), .B2(n_517), .C1(n_850), .C2(n_852), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_30), .A2(n_339), .B1(n_855), .B2(n_856), .Y(n_880) );
INVx1_ASAP7_75t_SL g414 ( .A(n_31), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g1012 ( .A(n_31), .B(n_43), .Y(n_1012) );
OA22x2_ASAP7_75t_L g652 ( .A1(n_32), .A2(n_653), .B1(n_654), .B2(n_655), .Y(n_652) );
CKINVDCx20_ASAP7_75t_R g653 ( .A(n_32), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g960 ( .A1(n_33), .A2(n_178), .B1(n_611), .B2(n_842), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_34), .A2(n_378), .B1(n_606), .B2(n_607), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_35), .B(n_586), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_36), .A2(n_291), .B1(n_538), .B2(n_539), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_37), .A2(n_123), .B1(n_855), .B2(n_856), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_38), .A2(n_216), .B1(n_630), .B2(n_632), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_39), .A2(n_232), .B1(n_569), .B2(n_742), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_40), .A2(n_188), .B1(n_524), .B2(n_989), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_41), .A2(n_369), .B1(n_667), .B2(n_668), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_42), .A2(n_332), .B1(n_621), .B2(n_692), .Y(n_757) );
AO22x2_ASAP7_75t_L g416 ( .A1(n_43), .A2(n_358), .B1(n_413), .B2(n_417), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_44), .A2(n_209), .B1(n_623), .B2(n_710), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_45), .A2(n_118), .B1(n_606), .B2(n_662), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_46), .A2(n_56), .B1(n_553), .B2(n_592), .Y(n_954) );
AOI22xp5_ASAP7_75t_L g823 ( .A1(n_47), .A2(n_331), .B1(n_623), .B2(n_710), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_48), .A2(n_371), .B1(n_607), .B2(n_621), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_49), .A2(n_284), .B1(n_621), .B2(n_712), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_51), .A2(n_343), .B1(n_603), .B2(n_690), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_52), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g415 ( .A(n_53), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_54), .A2(n_243), .B1(n_611), .B2(n_621), .Y(n_840) );
AOI22xp5_ASAP7_75t_L g927 ( .A1(n_55), .A2(n_312), .B1(n_535), .B2(n_539), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_57), .A2(n_297), .B1(n_557), .B2(n_893), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_58), .A2(n_295), .B1(n_603), .B2(n_632), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_59), .A2(n_308), .B1(n_538), .B2(n_867), .Y(n_924) );
AOI22xp33_ASAP7_75t_SL g820 ( .A1(n_60), .A2(n_318), .B1(n_621), .B2(n_658), .Y(n_820) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_61), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_62), .A2(n_136), .B1(n_760), .B2(n_900), .Y(n_941) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_63), .A2(n_355), .B1(n_562), .B2(n_563), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_64), .A2(n_303), .B1(n_568), .B2(n_569), .Y(n_996) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_66), .A2(n_249), .B1(n_584), .B2(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_67), .A2(n_351), .B1(n_662), .B2(n_695), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_68), .A2(n_211), .B1(n_695), .B2(n_696), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_69), .A2(n_345), .B1(n_505), .B2(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_70), .B(n_586), .Y(n_972) );
AO22x2_ASAP7_75t_L g423 ( .A1(n_71), .A2(n_194), .B1(n_413), .B2(n_424), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_72), .A2(n_197), .B1(n_481), .B2(n_600), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_73), .A2(n_88), .B1(n_481), .B2(n_904), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_74), .A2(n_313), .B1(n_600), .B2(n_623), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_75), .A2(n_236), .B1(n_603), .B2(n_632), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_76), .A2(n_353), .B1(n_592), .B2(n_670), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_77), .A2(n_167), .B1(n_524), .B2(n_525), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_78), .A2(n_169), .B1(n_603), .B2(n_1047), .Y(n_1046) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_79), .A2(n_199), .B1(n_621), .B2(n_692), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_80), .A2(n_161), .B1(n_469), .B2(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_SL g883 ( .A1(n_81), .A2(n_119), .B1(n_529), .B2(n_530), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_83), .A2(n_288), .B1(n_867), .B2(n_868), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_85), .A2(n_256), .B1(n_453), .B2(n_458), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_86), .A2(n_252), .B1(n_517), .B2(n_518), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g1052 ( .A1(n_87), .A2(n_114), .B1(n_482), .B2(n_980), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_89), .A2(n_198), .B1(n_557), .B2(n_1043), .Y(n_1042) );
AOI22xp33_ASAP7_75t_SL g736 ( .A1(n_90), .A2(n_195), .B1(n_554), .B2(n_737), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_91), .A2(n_235), .B1(n_569), .B2(n_710), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_92), .A2(n_372), .B1(n_548), .B2(n_584), .Y(n_1021) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_93), .A2(n_305), .B1(n_458), .B2(n_667), .Y(n_719) );
AOI22xp5_ASAP7_75t_L g1014 ( .A1(n_94), .A2(n_1015), .B1(n_1016), .B2(n_1028), .Y(n_1014) );
CKINVDCx20_ASAP7_75t_R g1028 ( .A(n_94), .Y(n_1028) );
AOI22xp5_ASAP7_75t_L g958 ( .A1(n_95), .A2(n_280), .B1(n_690), .B2(n_959), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_96), .A2(n_142), .B1(n_487), .B2(n_698), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_97), .A2(n_327), .B1(n_454), .B2(n_668), .Y(n_738) );
AO222x2_ASAP7_75t_L g917 ( .A1(n_99), .A2(n_208), .B1(n_362), .B2(n_522), .C1(n_525), .C2(n_850), .Y(n_917) );
AOI22xp33_ASAP7_75t_SL g785 ( .A1(n_100), .A2(n_133), .B1(n_786), .B2(n_788), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g520 ( .A1(n_101), .A2(n_230), .B1(n_521), .B2(n_522), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g1048 ( .A1(n_102), .A2(n_298), .B1(n_476), .B2(n_1049), .Y(n_1048) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_104), .A2(n_254), .B1(n_569), .B2(n_980), .Y(n_979) );
AOI22xp33_ASAP7_75t_SL g920 ( .A1(n_105), .A2(n_258), .B1(n_517), .B2(n_518), .Y(n_920) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_106), .Y(n_495) );
AOI222xp33_ASAP7_75t_L g720 ( .A1(n_107), .A2(n_179), .B1(n_344), .B2(n_548), .C1(n_672), .C2(n_721), .Y(n_720) );
OA22x2_ASAP7_75t_L g399 ( .A1(n_108), .A2(n_400), .B1(n_401), .B2(n_402), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_108), .Y(n_400) );
AOI222xp33_ASAP7_75t_L g836 ( .A1(n_109), .A2(n_147), .B1(n_275), .B2(n_557), .C1(n_672), .C2(n_686), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_110), .A2(n_163), .B1(n_525), .B2(n_858), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_111), .A2(n_271), .B1(n_639), .B2(n_893), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_112), .A2(n_234), .B1(n_760), .B2(n_900), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_113), .A2(n_130), .B1(n_626), .B2(n_749), .Y(n_940) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_115), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_116), .A2(n_238), .B1(n_505), .B2(n_603), .Y(n_660) );
AO22x2_ASAP7_75t_L g420 ( .A1(n_117), .A2(n_287), .B1(n_413), .B2(n_421), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g1020 ( .A1(n_120), .A2(n_302), .B1(n_668), .B2(n_801), .Y(n_1020) );
OAI22x1_ASAP7_75t_L g984 ( .A1(n_121), .A2(n_985), .B1(n_999), .B2(n_1000), .Y(n_984) );
CKINVDCx16_ASAP7_75t_R g1000 ( .A(n_121), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_124), .A2(n_159), .B1(n_686), .B2(n_801), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_125), .A2(n_377), .B1(n_562), .B2(n_611), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_126), .A2(n_265), .B1(n_606), .B2(n_793), .Y(n_1026) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_127), .A2(n_150), .B1(n_610), .B2(n_611), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_128), .A2(n_244), .B1(n_680), .B2(n_681), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_131), .A2(n_247), .B1(n_692), .B2(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g722 ( .A(n_132), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_134), .A2(n_350), .B1(n_530), .B2(n_862), .Y(n_861) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_135), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_137), .A2(n_202), .B1(n_536), .B2(n_571), .Y(n_865) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_138), .A2(n_337), .B1(n_427), .B2(n_433), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_139), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_140), .B(n_586), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g838 ( .A1(n_141), .A2(n_229), .B1(n_592), .B2(n_670), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_143), .A2(n_233), .B1(n_482), .B2(n_749), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_144), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_146), .A2(n_270), .B1(n_548), .B2(n_584), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g938 ( .A1(n_148), .A2(n_328), .B1(n_611), .B2(n_710), .Y(n_938) );
XOR2x2_ASAP7_75t_L g1033 ( .A(n_149), .B(n_1034), .Y(n_1033) );
INVxp67_ASAP7_75t_L g1059 ( .A(n_149), .Y(n_1059) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_152), .A2(n_173), .B1(n_557), .B2(n_686), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_153), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g884 ( .A1(n_154), .A2(n_160), .B1(n_867), .B2(n_868), .Y(n_884) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_155), .A2(n_336), .B1(n_680), .B2(n_681), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g977 ( .A1(n_157), .A2(n_223), .B1(n_710), .B2(n_712), .Y(n_977) );
AOI22xp5_ASAP7_75t_L g766 ( .A1(n_158), .A2(n_242), .B1(n_584), .B2(n_665), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_162), .A2(n_220), .B1(n_712), .B2(n_993), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_164), .B(n_550), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_165), .A2(n_240), .B1(n_610), .B2(n_658), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_166), .A2(n_289), .B1(n_505), .B2(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_168), .B(n_406), .Y(n_1019) );
AOI22xp33_ASAP7_75t_SL g821 ( .A1(n_171), .A2(n_304), .B1(n_603), .B2(n_632), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_172), .A2(n_346), .B1(n_557), .B2(n_765), .Y(n_934) );
OA22x2_ASAP7_75t_L g831 ( .A1(n_174), .A2(n_832), .B1(n_833), .B2(n_834), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_174), .Y(n_832) );
INVx1_ASAP7_75t_L g806 ( .A(n_175), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_176), .A2(n_354), .B1(n_532), .B2(n_747), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_177), .Y(n_731) );
AOI22xp33_ASAP7_75t_SL g669 ( .A1(n_181), .A2(n_227), .B1(n_592), .B2(n_670), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_183), .A2(n_379), .B1(n_433), .B2(n_642), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g906 ( .A(n_184), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_185), .A2(n_205), .B1(n_553), .B2(n_680), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_186), .A2(n_299), .B1(n_441), .B2(n_447), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_187), .A2(n_259), .B1(n_553), .B2(n_592), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_189), .A2(n_367), .B1(n_548), .B2(n_584), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_190), .A2(n_381), .B1(n_492), .B2(n_842), .Y(n_902) );
AOI22xp33_ASAP7_75t_SL g790 ( .A1(n_191), .A2(n_314), .B1(n_600), .B2(n_791), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_193), .A2(n_253), .B1(n_558), .B2(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g1011 ( .A(n_194), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_196), .A2(n_228), .B1(n_538), .B2(n_539), .Y(n_863) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_201), .A2(n_359), .B1(n_553), .B2(n_554), .Y(n_552) );
INVx1_ASAP7_75t_L g796 ( .A(n_203), .Y(n_796) );
AOI22xp33_ASAP7_75t_SL g919 ( .A1(n_204), .A2(n_324), .B1(n_855), .B2(n_858), .Y(n_919) );
OAI22xp5_ASAP7_75t_L g968 ( .A1(n_206), .A2(n_969), .B1(n_970), .B2(n_982), .Y(n_968) );
INVxp67_ASAP7_75t_L g982 ( .A(n_206), .Y(n_982) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_207), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_210), .A2(n_267), .B1(n_584), .B2(n_665), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_212), .A2(n_279), .B1(n_620), .B2(n_622), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_213), .A2(n_316), .B1(n_625), .B2(n_626), .Y(n_624) );
OA22x2_ASAP7_75t_L g752 ( .A1(n_214), .A2(n_753), .B1(n_754), .B2(n_768), .Y(n_752) );
INVxp67_ASAP7_75t_L g768 ( .A(n_214), .Y(n_768) );
OA22x2_ASAP7_75t_L g770 ( .A1(n_214), .A2(n_753), .B1(n_754), .B2(n_768), .Y(n_770) );
XNOR2x1_ASAP7_75t_L g579 ( .A(n_215), .B(n_580), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g837 ( .A1(n_217), .A2(n_374), .B1(n_584), .B2(n_665), .Y(n_837) );
INVx2_ASAP7_75t_L g389 ( .A(n_219), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_221), .A2(n_370), .B1(n_535), .B2(n_536), .Y(n_886) );
OA22x2_ASAP7_75t_L g673 ( .A1(n_222), .A2(n_674), .B1(n_700), .B2(n_701), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_222), .Y(n_700) );
AOI22xp33_ASAP7_75t_SL g962 ( .A1(n_224), .A2(n_272), .B1(n_481), .B2(n_606), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_225), .A2(n_245), .B1(n_695), .B2(n_716), .Y(n_715) );
AOI22xp33_ASAP7_75t_SL g1041 ( .A1(n_226), .A2(n_347), .B1(n_448), .B2(n_670), .Y(n_1041) );
AOI22xp5_ASAP7_75t_L g841 ( .A1(n_231), .A2(n_322), .B1(n_623), .B2(n_842), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_241), .A2(n_282), .B1(n_565), .B2(n_690), .Y(n_689) );
CKINVDCx16_ASAP7_75t_R g869 ( .A(n_246), .Y(n_869) );
AOI22xp5_ASAP7_75t_L g779 ( .A1(n_248), .A2(n_780), .B1(n_781), .B2(n_802), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_248), .Y(n_780) );
OAI22xp5_ASAP7_75t_L g913 ( .A1(n_250), .A2(n_914), .B1(n_915), .B2(n_928), .Y(n_913) );
INVx1_ASAP7_75t_L g928 ( .A(n_250), .Y(n_928) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_251), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g851 ( .A1(n_257), .A2(n_340), .B1(n_517), .B2(n_852), .Y(n_851) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_260), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g952 ( .A1(n_261), .A2(n_268), .B1(n_548), .B2(n_584), .Y(n_952) );
AOI22xp33_ASAP7_75t_SL g879 ( .A1(n_262), .A2(n_285), .B1(n_525), .B2(n_858), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_263), .A2(n_349), .B1(n_569), .B2(n_621), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_264), .A2(n_300), .B1(n_546), .B2(n_548), .Y(n_545) );
AOI211xp5_ASAP7_75t_L g382 ( .A1(n_266), .A2(n_383), .B(n_392), .C(n_1013), .Y(n_382) );
XNOR2x1_ASAP7_75t_L g946 ( .A(n_269), .B(n_947), .Y(n_946) );
CKINVDCx20_ASAP7_75t_R g588 ( .A(n_273), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_274), .A2(n_357), .B1(n_568), .B2(n_569), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_277), .B(n_586), .Y(n_933) );
OA22x2_ASAP7_75t_L g614 ( .A1(n_278), .A2(n_615), .B1(n_616), .B2(n_617), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_278), .Y(n_615) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_281), .Y(n_479) );
AOI22xp33_ASAP7_75t_SL g784 ( .A1(n_286), .A2(n_335), .B1(n_610), .B2(n_611), .Y(n_784) );
NOR2xp33_ASAP7_75t_L g1009 ( .A(n_287), .B(n_1010), .Y(n_1009) );
AOI222xp33_ASAP7_75t_L g997 ( .A1(n_290), .A2(n_301), .B1(n_341), .B2(n_850), .C1(n_852), .C2(n_998), .Y(n_997) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_292), .B(n_586), .Y(n_683) );
CKINVDCx20_ASAP7_75t_R g596 ( .A(n_293), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_294), .A2(n_380), .B1(n_603), .B2(n_759), .Y(n_1025) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_296), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g951 ( .A(n_306), .Y(n_951) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_307), .A2(n_325), .B1(n_759), .B2(n_760), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_309), .A2(n_334), .B1(n_606), .B2(n_662), .Y(n_844) );
INVx1_ASAP7_75t_L g750 ( .A(n_310), .Y(n_750) );
INVx3_ASAP7_75t_L g413 ( .A(n_311), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_315), .A2(n_326), .B1(n_535), .B2(n_536), .Y(n_534) );
AOI222xp33_ASAP7_75t_L g905 ( .A1(n_319), .A2(n_356), .B1(n_365), .B2(n_427), .C1(n_433), .C2(n_586), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_320), .A2(n_366), .B1(n_454), .B2(n_765), .Y(n_813) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_321), .Y(n_425) );
CKINVDCx20_ASAP7_75t_R g594 ( .A(n_323), .Y(n_594) );
CKINVDCx20_ASAP7_75t_R g572 ( .A(n_330), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_338), .A2(n_361), .B1(n_441), .B2(n_554), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_342), .B(n_672), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_348), .A2(n_376), .B1(n_557), .B2(n_558), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_360), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g1007 ( .A(n_360), .Y(n_1007) );
INVx1_ASAP7_75t_L g386 ( .A(n_363), .Y(n_386) );
AND2x2_ASAP7_75t_R g1030 ( .A(n_363), .B(n_1007), .Y(n_1030) );
INVxp67_ASAP7_75t_L g391 ( .A(n_368), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_373), .B(n_850), .Y(n_849) );
CKINVDCx20_ASAP7_75t_R g590 ( .A(n_375), .Y(n_590) );
BUFx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NOR2x1_ASAP7_75t_R g384 ( .A(n_385), .B(n_387), .Y(n_384) );
OR2x2_ASAP7_75t_L g1058 ( .A(n_385), .B(n_388), .Y(n_1058) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g1006 ( .A(n_386), .B(n_1007), .Y(n_1006) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_772), .B1(n_1002), .B2(n_1003), .C(n_1004), .Y(n_392) );
INVx1_ASAP7_75t_L g1002 ( .A(n_393), .Y(n_1002) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_395), .B1(n_647), .B2(n_771), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_576), .B1(n_645), .B2(n_646), .Y(n_395) );
INVx2_ASAP7_75t_L g645 ( .A(n_396), .Y(n_645) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OAI22x1_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_508), .B1(n_509), .B2(n_575), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g575 ( .A(n_399), .Y(n_575) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND3x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_462), .C(n_483), .Y(n_402) );
NOR2xp67_ASAP7_75t_SL g403 ( .A(n_404), .B(n_439), .Y(n_403) );
OAI21xp5_ASAP7_75t_SL g404 ( .A1(n_405), .A2(n_425), .B(n_426), .Y(n_404) );
OAI222xp33_ASAP7_75t_L g728 ( .A1(n_405), .A2(n_729), .B1(n_731), .B2(n_732), .C1(n_733), .C2(n_734), .Y(n_728) );
OAI21xp33_ASAP7_75t_L g795 ( .A1(n_405), .A2(n_796), .B(n_797), .Y(n_795) );
INVx3_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g637 ( .A(n_407), .Y(n_637) );
INVx3_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVx4_ASAP7_75t_SL g515 ( .A(n_408), .Y(n_515) );
INVx3_ASAP7_75t_L g550 ( .A(n_408), .Y(n_550) );
INVx3_ASAP7_75t_L g586 ( .A(n_408), .Y(n_586) );
INVx4_ASAP7_75t_SL g672 ( .A(n_408), .Y(n_672) );
BUFx2_ASAP7_75t_L g1037 ( .A(n_408), .Y(n_1037) );
INVx6_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_418), .Y(n_409) );
AND2x4_ASAP7_75t_L g449 ( .A(n_410), .B(n_450), .Y(n_449) );
AND2x4_ASAP7_75t_L g460 ( .A(n_410), .B(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g522 ( .A(n_410), .B(n_450), .Y(n_522) );
AND2x2_ASAP7_75t_L g525 ( .A(n_410), .B(n_461), .Y(n_525) );
AND2x4_ASAP7_75t_L g850 ( .A(n_410), .B(n_418), .Y(n_850) );
AND2x2_ASAP7_75t_L g856 ( .A(n_410), .B(n_450), .Y(n_856) );
AND2x2_ASAP7_75t_L g989 ( .A(n_410), .B(n_461), .Y(n_989) );
AND2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_416), .Y(n_410) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_411), .Y(n_432) );
AND2x2_ASAP7_75t_L g437 ( .A(n_411), .B(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g457 ( .A(n_411), .Y(n_457) );
OAI22x1_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_413), .B1(n_414), .B2(n_415), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g417 ( .A(n_413), .Y(n_417) );
INVx2_ASAP7_75t_L g421 ( .A(n_413), .Y(n_421) );
INVx1_ASAP7_75t_L g424 ( .A(n_413), .Y(n_424) );
INVx2_ASAP7_75t_L g438 ( .A(n_416), .Y(n_438) );
AND2x2_ASAP7_75t_L g456 ( .A(n_416), .B(n_457), .Y(n_456) );
BUFx2_ASAP7_75t_L g506 ( .A(n_416), .Y(n_506) );
AND2x4_ASAP7_75t_L g466 ( .A(n_418), .B(n_437), .Y(n_466) );
AND2x4_ASAP7_75t_L g478 ( .A(n_418), .B(n_471), .Y(n_478) );
AND2x2_ASAP7_75t_L g489 ( .A(n_418), .B(n_456), .Y(n_489) );
AND2x2_ASAP7_75t_L g535 ( .A(n_418), .B(n_437), .Y(n_535) );
AND2x6_ASAP7_75t_L g538 ( .A(n_418), .B(n_456), .Y(n_538) );
AND2x2_ASAP7_75t_L g571 ( .A(n_418), .B(n_437), .Y(n_571) );
AND2x2_ASAP7_75t_L g867 ( .A(n_418), .B(n_471), .Y(n_867) );
AND2x4_ASAP7_75t_L g418 ( .A(n_419), .B(n_422), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g431 ( .A(n_420), .B(n_423), .Y(n_431) );
AND2x4_ASAP7_75t_L g436 ( .A(n_420), .B(n_422), .Y(n_436) );
INVx1_ASAP7_75t_L g446 ( .A(n_420), .Y(n_446) );
INVxp67_ASAP7_75t_L g461 ( .A(n_422), .Y(n_461) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g445 ( .A(n_423), .B(n_446), .Y(n_445) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx3_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g665 ( .A(n_429), .Y(n_665) );
INVx2_ASAP7_75t_L g678 ( .A(n_429), .Y(n_678) );
INVx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx12f_ASAP7_75t_L g548 ( .A(n_430), .Y(n_548) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
AND2x4_ASAP7_75t_L g482 ( .A(n_431), .B(n_471), .Y(n_482) );
AND2x4_ASAP7_75t_L g505 ( .A(n_431), .B(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_SL g518 ( .A(n_431), .B(n_432), .Y(n_518) );
AND2x4_ASAP7_75t_L g530 ( .A(n_431), .B(n_506), .Y(n_530) );
AND2x4_ASAP7_75t_L g536 ( .A(n_431), .B(n_471), .Y(n_536) );
AND2x2_ASAP7_75t_SL g852 ( .A(n_431), .B(n_432), .Y(n_852) );
BUFx6f_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
BUFx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g547 ( .A(n_435), .Y(n_547) );
BUFx5_ASAP7_75t_L g584 ( .A(n_435), .Y(n_584) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
AND2x4_ASAP7_75t_L g455 ( .A(n_436), .B(n_456), .Y(n_455) );
AND2x4_ASAP7_75t_L g470 ( .A(n_436), .B(n_471), .Y(n_470) );
AND2x4_ASAP7_75t_L g517 ( .A(n_436), .B(n_437), .Y(n_517) );
AND2x2_ASAP7_75t_L g524 ( .A(n_436), .B(n_456), .Y(n_524) );
AND2x2_ASAP7_75t_L g858 ( .A(n_436), .B(n_456), .Y(n_858) );
AND2x2_ASAP7_75t_L g868 ( .A(n_436), .B(n_471), .Y(n_868) );
AND2x2_ASAP7_75t_L g444 ( .A(n_437), .B(n_445), .Y(n_444) );
AND2x4_ASAP7_75t_L g855 ( .A(n_437), .B(n_445), .Y(n_855) );
AND2x4_ASAP7_75t_L g471 ( .A(n_438), .B(n_457), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g439 ( .A(n_440), .B(n_452), .Y(n_439) );
BUFx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx4_ASAP7_75t_L g521 ( .A(n_443), .Y(n_521) );
INVx2_ASAP7_75t_L g681 ( .A(n_443), .Y(n_681) );
INVx3_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_444), .Y(n_553) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_444), .Y(n_670) );
AND2x4_ASAP7_75t_L g494 ( .A(n_445), .B(n_471), .Y(n_494) );
AND2x2_ASAP7_75t_L g502 ( .A(n_445), .B(n_456), .Y(n_502) );
AND2x2_ASAP7_75t_SL g529 ( .A(n_445), .B(n_456), .Y(n_529) );
AND2x6_ASAP7_75t_L g539 ( .A(n_445), .B(n_471), .Y(n_539) );
AND2x2_ASAP7_75t_L g862 ( .A(n_445), .B(n_456), .Y(n_862) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_446), .Y(n_451) );
BUFx6f_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
BUFx3_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g555 ( .A(n_449), .Y(n_555) );
BUFx4f_ASAP7_75t_L g592 ( .A(n_449), .Y(n_592) );
BUFx6f_ASAP7_75t_SL g680 ( .A(n_449), .Y(n_680) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g595 ( .A(n_454), .Y(n_595) );
BUFx2_ASAP7_75t_L g639 ( .A(n_454), .Y(n_639) );
BUFx4f_ASAP7_75t_SL g801 ( .A(n_454), .Y(n_801) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx3_ASAP7_75t_L g557 ( .A(n_455), .Y(n_557) );
BUFx2_ASAP7_75t_L g667 ( .A(n_455), .Y(n_667) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g558 ( .A(n_459), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_459), .A2(n_594), .B1(n_595), .B2(n_596), .Y(n_593) );
INVx2_ASAP7_75t_SL g668 ( .A(n_459), .Y(n_668) );
INVx2_ASAP7_75t_SL g686 ( .A(n_459), .Y(n_686) );
INVx1_ASAP7_75t_L g765 ( .A(n_459), .Y(n_765) );
INVx2_ASAP7_75t_L g893 ( .A(n_459), .Y(n_893) );
INVx2_ASAP7_75t_L g1043 ( .A(n_459), .Y(n_1043) );
INVx6_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_463), .B(n_472), .Y(n_462) );
OAI22xp33_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B1(n_467), .B2(n_468), .Y(n_463) );
INVx2_ASAP7_75t_L g606 ( .A(n_465), .Y(n_606) );
INVx2_ASAP7_75t_L g695 ( .A(n_465), .Y(n_695) );
INVx3_ASAP7_75t_L g749 ( .A(n_465), .Y(n_749) );
INVx2_ASAP7_75t_L g904 ( .A(n_465), .Y(n_904) );
INVx6_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx3_ASAP7_75t_L g625 ( .A(n_466), .Y(n_625) );
BUFx3_ASAP7_75t_L g980 ( .A(n_466), .Y(n_980) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx6f_ASAP7_75t_L g898 ( .A(n_469), .Y(n_898) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_470), .Y(n_569) );
BUFx3_ASAP7_75t_L g623 ( .A(n_470), .Y(n_623) );
INVx2_ASAP7_75t_L g699 ( .A(n_470), .Y(n_699) );
OAI22xp33_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_474), .B1(n_479), .B2(n_480), .Y(n_472) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
INVx3_ASAP7_75t_SL g532 ( .A(n_477), .Y(n_532) );
INVx2_ASAP7_75t_L g568 ( .A(n_477), .Y(n_568) );
INVx4_ASAP7_75t_L g601 ( .A(n_477), .Y(n_601) );
INVx2_ASAP7_75t_SL g621 ( .A(n_477), .Y(n_621) );
INVx8_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
BUFx2_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g627 ( .A(n_482), .Y(n_627) );
BUFx3_ASAP7_75t_L g696 ( .A(n_482), .Y(n_696) );
BUFx3_ASAP7_75t_L g716 ( .A(n_482), .Y(n_716) );
BUFx2_ASAP7_75t_SL g793 ( .A(n_482), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_484), .B(n_496), .Y(n_483) );
OAI22xp33_ASAP7_75t_SL g484 ( .A1(n_485), .A2(n_490), .B1(n_491), .B2(n_495), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx3_ASAP7_75t_L g562 ( .A(n_488), .Y(n_562) );
INVx2_ASAP7_75t_SL g610 ( .A(n_488), .Y(n_610) );
INVx2_ASAP7_75t_L g710 ( .A(n_488), .Y(n_710) );
INVx2_ASAP7_75t_SL g842 ( .A(n_488), .Y(n_842) );
INVx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx2_ASAP7_75t_L g742 ( .A(n_489), .Y(n_742) );
BUFx2_ASAP7_75t_L g993 ( .A(n_489), .Y(n_993) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_SL g563 ( .A(n_493), .Y(n_563) );
INVx2_ASAP7_75t_SL g611 ( .A(n_493), .Y(n_611) );
INVx1_ASAP7_75t_SL g658 ( .A(n_493), .Y(n_658) );
INVx2_ASAP7_75t_L g692 ( .A(n_493), .Y(n_692) );
INVx2_ASAP7_75t_L g712 ( .A(n_493), .Y(n_712) );
INVx2_ASAP7_75t_L g1049 ( .A(n_493), .Y(n_1049) );
INVx8_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
OAI22xp33_ASAP7_75t_SL g496 ( .A1(n_497), .A2(n_503), .B1(n_504), .B2(n_507), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g959 ( .A(n_499), .Y(n_959) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx6f_ASAP7_75t_L g760 ( .A(n_500), .Y(n_760) );
INVx1_ASAP7_75t_L g787 ( .A(n_500), .Y(n_787) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g631 ( .A(n_501), .Y(n_631) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx3_ASAP7_75t_L g565 ( .A(n_502), .Y(n_565) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_502), .Y(n_603) );
INVx2_ASAP7_75t_L g632 ( .A(n_504), .Y(n_632) );
INVx3_ASAP7_75t_L g690 ( .A(n_504), .Y(n_690) );
INVx2_ASAP7_75t_L g788 ( .A(n_504), .Y(n_788) );
INVx2_ASAP7_75t_L g1047 ( .A(n_504), .Y(n_1047) );
INVx5_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
BUFx3_ASAP7_75t_L g744 ( .A(n_505), .Y(n_744) );
BUFx2_ASAP7_75t_L g759 ( .A(n_505), .Y(n_759) );
BUFx2_ASAP7_75t_L g900 ( .A(n_505), .Y(n_900) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AO22x2_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_541), .B1(n_573), .B2(n_574), .Y(n_509) );
INVx1_ASAP7_75t_SL g574 ( .A(n_510), .Y(n_574) );
XOR2x2_ASAP7_75t_L g578 ( .A(n_510), .B(n_579), .Y(n_578) );
XOR2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_540), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_512), .B(n_526), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_519), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_516), .Y(n_513) );
INVx1_ASAP7_75t_SL g815 ( .A(n_515), .Y(n_815) );
HB1xp67_ASAP7_75t_L g998 ( .A(n_517), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_523), .Y(n_519) );
INVx2_ASAP7_75t_SL g589 ( .A(n_521), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_527), .B(n_533), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_531), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_537), .Y(n_533) );
INVx2_ASAP7_75t_L g573 ( .A(n_541), .Y(n_573) );
XOR2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_572), .Y(n_541) );
NAND2x1p5_ASAP7_75t_L g542 ( .A(n_543), .B(n_559), .Y(n_542) );
NOR2x1_ASAP7_75t_L g543 ( .A(n_544), .B(n_551), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_549), .Y(n_544) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_546), .Y(n_730) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g721 ( .A(n_547), .Y(n_721) );
BUFx3_ASAP7_75t_L g642 ( .A(n_548), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_556), .Y(n_551) );
BUFx6f_ASAP7_75t_SL g737 ( .A(n_553), .Y(n_737) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NOR2x1_ASAP7_75t_L g559 ( .A(n_560), .B(n_566), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_564), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_570), .Y(n_566) );
INVx1_ASAP7_75t_L g608 ( .A(n_569), .Y(n_608) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_569), .Y(n_747) );
INVx1_ASAP7_75t_L g646 ( .A(n_576), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_612), .B1(n_613), .B2(n_643), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g644 ( .A(n_578), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_597), .Y(n_580) );
NOR3xp33_ASAP7_75t_L g581 ( .A(n_582), .B(n_587), .C(n_593), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_583), .B(n_585), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B1(n_590), .B2(n_591), .Y(n_587) );
INVxp67_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_598), .B(n_604), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_602), .Y(n_598) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g897 ( .A(n_601), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_609), .Y(n_604) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
BUFx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NOR3x1_ASAP7_75t_SL g617 ( .A(n_618), .B(n_628), .C(n_634), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_624), .Y(n_618) );
BUFx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
BUFx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_SL g662 ( .A(n_627), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_633), .Y(n_628) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NAND4xp25_ASAP7_75t_SL g634 ( .A(n_635), .B(n_638), .C(n_640), .D(n_641), .Y(n_634) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g733 ( .A(n_642), .Y(n_733) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g771 ( .A(n_647), .Y(n_771) );
OA22x2_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_649), .B1(n_723), .B2(n_724), .Y(n_647) );
INVx2_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
OA22x2_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_651), .B1(n_705), .B2(n_706), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_673), .B1(n_703), .B2(n_704), .Y(n_651) );
INVx1_ASAP7_75t_L g703 ( .A(n_652), .Y(n_703) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NOR2x1_ASAP7_75t_L g655 ( .A(n_656), .B(n_663), .Y(n_655) );
NAND4xp25_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .C(n_660), .D(n_661), .Y(n_656) );
NAND4xp25_ASAP7_75t_L g663 ( .A(n_664), .B(n_666), .C(n_669), .D(n_671), .Y(n_663) );
INVx1_ASAP7_75t_L g950 ( .A(n_672), .Y(n_950) );
INVx2_ASAP7_75t_L g704 ( .A(n_673), .Y(n_704) );
AO22x2_ASAP7_75t_SL g804 ( .A1(n_673), .A2(n_704), .B1(n_805), .B2(n_826), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_687), .Y(n_674) );
NOR3xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_682), .C(n_684), .Y(n_675) );
NOR4xp25_ASAP7_75t_L g701 ( .A(n_676), .B(n_688), .C(n_693), .D(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_679), .Y(n_676) );
INVxp67_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_683), .B(n_685), .Y(n_702) );
INVxp67_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_688), .B(n_693), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_691), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_697), .Y(n_693) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g791 ( .A(n_699), .Y(n_791) );
INVx3_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
XOR2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_722), .Y(n_706) );
NAND4xp75_ASAP7_75t_L g707 ( .A(n_708), .B(n_713), .C(n_717), .D(n_720), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_709), .B(n_711), .Y(n_708) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
AND2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_751), .B1(n_769), .B2(n_770), .Y(n_724) );
INVx3_ASAP7_75t_L g769 ( .A(n_725), .Y(n_769) );
XOR2x2_ASAP7_75t_L g725 ( .A(n_726), .B(n_750), .Y(n_725) );
NAND2xp5_ASAP7_75t_SL g726 ( .A(n_727), .B(n_739), .Y(n_726) );
NOR2x1_ASAP7_75t_L g727 ( .A(n_728), .B(n_735), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_736), .B(n_738), .Y(n_735) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_740), .B(n_745), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_741), .B(n_743), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_748), .Y(n_745) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx2_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
NOR2x1_ASAP7_75t_L g754 ( .A(n_755), .B(n_762), .Y(n_754) );
NAND4xp25_ASAP7_75t_SL g755 ( .A(n_756), .B(n_757), .C(n_758), .D(n_761), .Y(n_755) );
NAND4xp25_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .C(n_766), .D(n_767), .Y(n_762) );
INVx1_ASAP7_75t_L g1003 ( .A(n_772), .Y(n_1003) );
XNOR2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_908), .Y(n_772) );
AOI22xp5_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_775), .B1(n_827), .B2(n_828), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_777), .B1(n_803), .B2(n_804), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
BUFx3_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVxp33_ASAP7_75t_SL g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_SL g802 ( .A(n_781), .Y(n_802) );
AND2x2_ASAP7_75t_L g781 ( .A(n_782), .B(n_794), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_789), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_784), .B(n_785), .Y(n_783) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_790), .B(n_792), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g794 ( .A(n_795), .B(n_798), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx2_ASAP7_75t_L g826 ( .A(n_805), .Y(n_826) );
OAI21x1_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_807), .B(n_825), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_806), .B(n_809), .Y(n_825) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_810), .B(n_818), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g810 ( .A(n_811), .B(n_814), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .Y(n_811) );
OAI21xp33_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_816), .B(n_817), .Y(n_814) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_819), .B(n_822), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .Y(n_822) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
XNOR2xp5_ASAP7_75t_SL g828 ( .A(n_829), .B(n_870), .Y(n_828) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
XNOR2x1_ASAP7_75t_L g830 ( .A(n_831), .B(n_845), .Y(n_830) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
NOR2x1_ASAP7_75t_L g834 ( .A(n_835), .B(n_839), .Y(n_834) );
NAND3xp33_ASAP7_75t_L g835 ( .A(n_836), .B(n_837), .C(n_838), .Y(n_835) );
NAND4xp25_ASAP7_75t_L g839 ( .A(n_840), .B(n_841), .C(n_843), .D(n_844), .Y(n_839) );
XOR2x2_ASAP7_75t_L g845 ( .A(n_846), .B(n_869), .Y(n_845) );
NAND2x1p5_ASAP7_75t_L g846 ( .A(n_847), .B(n_859), .Y(n_846) );
NOR2x1_ASAP7_75t_L g847 ( .A(n_848), .B(n_853), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_849), .B(n_851), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_854), .B(n_857), .Y(n_853) );
NOR2x1_ASAP7_75t_L g859 ( .A(n_860), .B(n_864), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_861), .B(n_863), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_865), .B(n_866), .Y(n_864) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_872), .B1(n_888), .B2(n_907), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx2_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
XNOR2x1_ASAP7_75t_L g873 ( .A(n_874), .B(n_875), .Y(n_873) );
AND2x2_ASAP7_75t_L g875 ( .A(n_876), .B(n_881), .Y(n_875) );
NOR2xp33_ASAP7_75t_L g876 ( .A(n_877), .B(n_878), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_879), .B(n_880), .Y(n_878) );
NOR2xp33_ASAP7_75t_L g881 ( .A(n_882), .B(n_885), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_883), .B(n_884), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_886), .B(n_887), .Y(n_885) );
INVx2_ASAP7_75t_SL g907 ( .A(n_888), .Y(n_907) );
XNOR2x1_ASAP7_75t_L g888 ( .A(n_889), .B(n_906), .Y(n_888) );
NAND4xp75_ASAP7_75t_L g889 ( .A(n_890), .B(n_894), .C(n_901), .D(n_905), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_891), .B(n_892), .Y(n_890) );
AND2x2_ASAP7_75t_L g894 ( .A(n_895), .B(n_899), .Y(n_894) );
INVx1_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
AND2x2_ASAP7_75t_L g901 ( .A(n_902), .B(n_903), .Y(n_901) );
OAI22xp5_ASAP7_75t_SL g908 ( .A1(n_909), .A2(n_965), .B1(n_966), .B2(n_1001), .Y(n_908) );
INVx1_ASAP7_75t_L g1001 ( .A(n_909), .Y(n_1001) );
OAI22xp5_ASAP7_75t_SL g909 ( .A1(n_910), .A2(n_911), .B1(n_943), .B2(n_964), .Y(n_909) );
INVx2_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
AO22x2_ASAP7_75t_L g911 ( .A1(n_912), .A2(n_929), .B1(n_930), .B2(n_942), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
BUFx2_ASAP7_75t_L g942 ( .A(n_913), .Y(n_942) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
NAND2xp5_ASAP7_75t_SL g915 ( .A(n_916), .B(n_921), .Y(n_915) );
NOR2xp33_ASAP7_75t_L g916 ( .A(n_917), .B(n_918), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_919), .B(n_920), .Y(n_918) );
NOR2xp33_ASAP7_75t_L g921 ( .A(n_922), .B(n_925), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_923), .B(n_924), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_926), .B(n_927), .Y(n_925) );
INVx1_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
NOR2xp67_ASAP7_75t_L g931 ( .A(n_932), .B(n_937), .Y(n_931) );
NAND4xp25_ASAP7_75t_SL g932 ( .A(n_933), .B(n_934), .C(n_935), .D(n_936), .Y(n_932) );
NAND4xp25_ASAP7_75t_L g937 ( .A(n_938), .B(n_939), .C(n_940), .D(n_941), .Y(n_937) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
INVx2_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g964 ( .A(n_945), .Y(n_964) );
INVx1_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
AND2x4_ASAP7_75t_L g947 ( .A(n_948), .B(n_956), .Y(n_947) );
NOR2xp67_ASAP7_75t_L g948 ( .A(n_949), .B(n_953), .Y(n_948) );
OAI21xp5_ASAP7_75t_SL g949 ( .A1(n_950), .A2(n_951), .B(n_952), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_954), .B(n_955), .Y(n_953) );
NOR2x1_ASAP7_75t_L g956 ( .A(n_957), .B(n_961), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_958), .B(n_960), .Y(n_957) );
NAND2xp5_ASAP7_75t_L g961 ( .A(n_962), .B(n_963), .Y(n_961) );
INVx2_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
OA22x2_ASAP7_75t_L g966 ( .A1(n_967), .A2(n_968), .B1(n_983), .B2(n_984), .Y(n_966) );
INVx2_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
NOR2xp67_ASAP7_75t_L g970 ( .A(n_971), .B(n_976), .Y(n_970) );
NAND4xp25_ASAP7_75t_L g971 ( .A(n_972), .B(n_973), .C(n_974), .D(n_975), .Y(n_971) );
NAND4xp25_ASAP7_75t_L g976 ( .A(n_977), .B(n_978), .C(n_979), .D(n_981), .Y(n_976) );
INVx2_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
NAND4xp25_ASAP7_75t_SL g985 ( .A(n_986), .B(n_990), .C(n_994), .D(n_997), .Y(n_985) );
AND4x1_ASAP7_75t_L g999 ( .A(n_986), .B(n_990), .C(n_994), .D(n_997), .Y(n_999) );
AND2x2_ASAP7_75t_L g986 ( .A(n_987), .B(n_988), .Y(n_986) );
AND2x2_ASAP7_75t_L g990 ( .A(n_991), .B(n_992), .Y(n_990) );
AND2x2_ASAP7_75t_L g994 ( .A(n_995), .B(n_996), .Y(n_994) );
INVx1_ASAP7_75t_SL g1004 ( .A(n_1005), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_1006), .B(n_1008), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g1055 ( .A(n_1006), .B(n_1009), .Y(n_1055) );
INVx1_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1012), .Y(n_1010) );
OAI222xp33_ASAP7_75t_R g1013 ( .A1(n_1014), .A2(n_1029), .B1(n_1031), .B2(n_1053), .C1(n_1056), .C2(n_1059), .Y(n_1013) );
CKINVDCx20_ASAP7_75t_R g1015 ( .A(n_1016), .Y(n_1015) );
HB1xp67_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
OR2x2_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1023), .Y(n_1017) );
NAND4xp25_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1020), .C(n_1021), .D(n_1022), .Y(n_1018) );
NAND4xp25_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1025), .C(n_1026), .D(n_1027), .Y(n_1023) );
INVx1_ASAP7_75t_SL g1029 ( .A(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
HB1xp67_ASAP7_75t_L g1032 ( .A(n_1033), .Y(n_1032) );
NAND2x1_ASAP7_75t_SL g1034 ( .A(n_1035), .B(n_1044), .Y(n_1034) );
NOR2x1_ASAP7_75t_L g1035 ( .A(n_1036), .B(n_1040), .Y(n_1035) );
OAI21xp5_ASAP7_75t_SL g1036 ( .A1(n_1037), .A2(n_1038), .B(n_1039), .Y(n_1036) );
NAND2xp5_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1042), .Y(n_1040) );
NOR2x1_ASAP7_75t_L g1044 ( .A(n_1045), .B(n_1050), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1048), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1050 ( .A(n_1051), .B(n_1052), .Y(n_1050) );
INVx1_ASAP7_75t_SL g1053 ( .A(n_1054), .Y(n_1053) );
CKINVDCx6p67_ASAP7_75t_R g1054 ( .A(n_1055), .Y(n_1054) );
CKINVDCx20_ASAP7_75t_R g1056 ( .A(n_1057), .Y(n_1056) );
CKINVDCx20_ASAP7_75t_R g1057 ( .A(n_1058), .Y(n_1057) );
endmodule