module real_jpeg_21374_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_342, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_342;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_0),
.A2(n_22),
.B1(n_24),
.B2(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_0),
.A2(n_26),
.B1(n_28),
.B2(n_31),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_0),
.A2(n_31),
.B1(n_46),
.B2(n_47),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_0),
.A2(n_31),
.B1(n_40),
.B2(n_41),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_1),
.A2(n_22),
.B1(n_24),
.B2(n_57),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_57),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_1),
.A2(n_40),
.B1(n_41),
.B2(n_57),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_1),
.A2(n_26),
.B1(n_28),
.B2(n_57),
.Y(n_296)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_3),
.A2(n_22),
.B1(n_24),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_3),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_3),
.A2(n_26),
.B1(n_28),
.B2(n_125),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_3),
.A2(n_40),
.B1(n_41),
.B2(n_125),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_125),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_4),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_4),
.B(n_25),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_L g175 ( 
.A1(n_4),
.A2(n_14),
.B(n_47),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_4),
.A2(n_40),
.B1(n_41),
.B2(n_123),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_4),
.A2(n_96),
.B1(n_151),
.B2(n_184),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_4),
.B(n_76),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_4),
.B(n_28),
.Y(n_210)
);

AOI21xp33_ASAP7_75t_L g214 ( 
.A1(n_4),
.A2(n_28),
.B(n_210),
.Y(n_214)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_5),
.Y(n_99)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_5),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_6),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_6),
.A2(n_23),
.B1(n_40),
.B2(n_41),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_6),
.A2(n_23),
.B1(n_26),
.B2(n_28),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_6),
.A2(n_23),
.B1(n_46),
.B2(n_47),
.Y(n_202)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_8),
.A2(n_26),
.B1(n_28),
.B2(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_8),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_8),
.A2(n_22),
.B1(n_24),
.B2(n_118),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_8),
.A2(n_46),
.B1(n_47),
.B2(n_118),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_8),
.A2(n_40),
.B1(n_41),
.B2(n_118),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_9),
.A2(n_26),
.B1(n_28),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_9),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_120),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_9),
.A2(n_40),
.B1(n_41),
.B2(n_120),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_9),
.A2(n_22),
.B1(n_24),
.B2(n_120),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_11),
.A2(n_22),
.B1(n_24),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_11),
.A2(n_40),
.B1(n_41),
.B2(n_55),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_55),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_11),
.A2(n_26),
.B1(n_28),
.B2(n_55),
.Y(n_275)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_25)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_14),
.A2(n_40),
.B(n_44),
.C(n_45),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_14),
.B(n_40),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_15),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_84),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_82),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_34),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_19),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_29),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_20),
.A2(n_53),
.B(n_258),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_25),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_21),
.Y(n_304)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

O2A1O1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_25),
.B(n_27),
.C(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_27),
.Y(n_33)
);

HAxp5_ASAP7_75t_SL g122 ( 
.A(n_22),
.B(n_123),
.CON(n_122),
.SN(n_122)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_25),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_25),
.B(n_30),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_25),
.A2(n_32),
.B1(n_122),
.B2(n_124),
.Y(n_121)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_26),
.A2(n_33),
.B1(n_122),
.B2(n_129),
.Y(n_128)
);

AOI32xp33_ASAP7_75t_L g209 ( 
.A1(n_26),
.A2(n_40),
.A3(n_66),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_27),
.B(n_28),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_28),
.A2(n_63),
.B(n_64),
.C(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_28),
.B(n_64),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_29),
.A2(n_54),
.B(n_58),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_32),
.A2(n_79),
.B(n_80),
.Y(n_78)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_35),
.B(n_83),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_74),
.C(n_78),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_36),
.A2(n_37),
.B1(n_336),
.B2(n_338),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_51),
.C(n_59),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_38),
.A2(n_316),
.B1(n_317),
.B2(n_318),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_38),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_38),
.A2(n_59),
.B1(n_60),
.B2(n_316),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_45),
.B(n_49),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_39),
.A2(n_49),
.B(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_39),
.A2(n_45),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_39),
.A2(n_45),
.B1(n_179),
.B2(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_39),
.A2(n_45),
.B1(n_199),
.B2(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_39),
.A2(n_217),
.B(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_39),
.A2(n_45),
.B1(n_105),
.B2(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_39),
.A2(n_113),
.B(n_250),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_41),
.B1(n_64),
.B2(n_66),
.Y(n_63)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_41),
.A2(n_48),
.B(n_123),
.C(n_175),
.Y(n_174)
);

NAND2xp33_ASAP7_75t_SL g211 ( 
.A(n_41),
.B(n_64),
.Y(n_211)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_45),
.A2(n_105),
.B(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_45),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_45),
.B(n_123),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_46),
.B(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_46),
.B(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_50),
.B(n_114),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_51),
.A2(n_52),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_58),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_53),
.A2(n_58),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_53),
.A2(n_58),
.B1(n_137),
.B2(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_53),
.A2(n_81),
.B(n_304),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_56),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_68),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_62),
.A2(n_69),
.B(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_67),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_63),
.A2(n_70),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_63),
.A2(n_70),
.B1(n_157),
.B2(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_63),
.B(n_73),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_63),
.A2(n_68),
.B(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_63),
.A2(n_70),
.B1(n_275),
.B2(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_67),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_69),
.A2(n_76),
.B(n_77),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_69),
.A2(n_76),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_69),
.A2(n_77),
.B(n_261),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_69),
.A2(n_261),
.B(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_337),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_78),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_333),
.B(n_339),
.Y(n_84)
);

OAI321xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_309),
.A3(n_328),
.B1(n_331),
.B2(n_332),
.C(n_342),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_288),
.B(n_308),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_266),
.B(n_287),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_159),
.B(n_241),
.C(n_265),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_142),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_90),
.B(n_142),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_126),
.B2(n_141),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_110),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_93),
.B(n_110),
.C(n_141),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_104),
.B2(n_109),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_94),
.B(n_109),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_100),
.B(n_101),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_96),
.A2(n_100),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_96),
.A2(n_99),
.B1(n_168),
.B2(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_96),
.A2(n_171),
.B(n_201),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_96),
.A2(n_151),
.B(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_97),
.B(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_97),
.A2(n_167),
.B1(n_169),
.B2(n_170),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_97),
.A2(n_102),
.B(n_202),
.Y(n_208)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_98),
.B(n_202),
.Y(n_201)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_103),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_104),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_106),
.B(n_233),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_107),
.B(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.C(n_121),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_116),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_117),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_119),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_121),
.B(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_123),
.B(n_151),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_124),
.Y(n_136)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_133),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_127),
.B(n_134),
.C(n_139),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_130),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_138),
.B2(n_139),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.C(n_147),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_143),
.B(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_154),
.C(n_155),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_149),
.A2(n_150),
.B1(n_154),
.B2(n_228),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_152),
.B(n_201),
.Y(n_248)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_154),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_155),
.B(n_227),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_240),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_235),
.B(n_239),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_222),
.B(n_234),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_204),
.B(n_221),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_191),
.B(n_203),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_180),
.B(n_190),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_172),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_172),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_174),
.B(n_176),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_185),
.B(n_189),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_183),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_192),
.B(n_193),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_200),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_198),
.C(n_200),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_202),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_206),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_212),
.B1(n_219),
.B2(n_220),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_207),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_209),
.Y(n_231)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_212),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_215),
.B1(n_216),
.B2(n_218),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_213),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_218),
.C(n_219),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_223),
.B(n_224),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_229),
.B2(n_230),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_231),
.C(n_232),
.Y(n_236)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_236),
.B(n_237),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_242),
.B(n_243),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_263),
.B2(n_264),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_251),
.B2(n_252),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_252),
.C(n_264),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_249),
.Y(n_272)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_255),
.B2(n_262),
.Y(n_252)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_259),
.B2(n_260),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_260),
.C(n_262),
.Y(n_286)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_263),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_267),
.B(n_268),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_286),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_279),
.B2(n_280),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_280),
.C(n_286),
.Y(n_289)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_272),
.B(n_276),
.C(n_278),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_274),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_284),
.B2(n_285),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_281),
.A2(n_282),
.B1(n_303),
.B2(n_305),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_281),
.A2(n_299),
.B(n_303),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_284),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_284),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_289),
.B(n_290),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_306),
.B2(n_307),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_298),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_293),
.B(n_298),
.C(n_307),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_295),
.B(n_297),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_295),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_296),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_311),
.C(n_320),
.Y(n_310)
);

FAx1_ASAP7_75t_SL g330 ( 
.A(n_297),
.B(n_311),
.CI(n_320),
.CON(n_330),
.SN(n_330)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_301),
.B2(n_302),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_303),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_306),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_321),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_321),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_312),
.A2(n_313),
.B1(n_323),
.B2(n_326),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_313),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_316),
.C(n_318),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_313),
.B(n_326),
.C(n_327),
.Y(n_334)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_318),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_327),
.Y(n_321)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_323),
.Y(n_326)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_329),
.B(n_330),
.Y(n_331)
);

BUFx24_ASAP7_75t_SL g340 ( 
.A(n_330),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_335),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_336),
.Y(n_338)
);


endmodule