module fake_jpeg_1361_n_242 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_242);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_242;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_33),
.B(n_32),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_42),
.B(n_44),
.Y(n_85)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_25),
.B(n_0),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_47),
.B(n_62),
.Y(n_90)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_28),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_51),
.B(n_60),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_23),
.Y(n_79)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_28),
.B(n_14),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_22),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_21),
.B(n_1),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_65),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_34),
.Y(n_64)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_34),
.B1(n_31),
.B2(n_37),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_66),
.A2(n_73),
.B1(n_24),
.B2(n_17),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_37),
.C(n_36),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_67),
.B(n_64),
.Y(n_115)
);

OR2x2_ASAP7_75t_SL g70 ( 
.A(n_63),
.B(n_36),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_70),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_21),
.B1(n_31),
.B2(n_40),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_45),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_83),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_79),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_47),
.A2(n_64),
.B1(n_35),
.B2(n_46),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_41),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_32),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_20),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_89),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_43),
.A2(n_21),
.B1(n_38),
.B2(n_40),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_88),
.A2(n_41),
.B1(n_61),
.B2(n_53),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_29),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_49),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_94),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_29),
.Y(n_94)
);

NOR2x1_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_35),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_101),
.A2(n_117),
.B1(n_124),
.B2(n_127),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_86),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_102),
.B(n_103),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_27),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_129),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_115),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_66),
.B1(n_50),
.B2(n_87),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_68),
.B1(n_76),
.B2(n_98),
.Y(n_132)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

NOR2x1_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_65),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_116),
.Y(n_130)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_27),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_81),
.A2(n_24),
.B1(n_17),
.B2(n_58),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_118),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_59),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_121),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_90),
.A2(n_52),
.B1(n_19),
.B2(n_4),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_13),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_13),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_81),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_124)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_67),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_78),
.B(n_5),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_132),
.A2(n_96),
.B1(n_82),
.B2(n_93),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_117),
.B1(n_105),
.B2(n_115),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_134),
.A2(n_129),
.B1(n_114),
.B2(n_112),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_137),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_72),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_104),
.B(n_70),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_143),
.B(n_99),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_110),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_145),
.B(n_123),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_98),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_105),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_74),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_119),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_R g149 ( 
.A1(n_106),
.A2(n_81),
.B1(n_74),
.B2(n_76),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_121),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_155),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_131),
.A2(n_102),
.B1(n_103),
.B2(n_119),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_156),
.A2(n_173),
.B1(n_174),
.B2(n_150),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_162),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_106),
.C(n_120),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_165),
.C(n_154),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_142),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_160),
.B(n_161),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_120),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_163),
.Y(n_181)
);

AOI322xp5_ASAP7_75t_SL g191 ( 
.A1(n_164),
.A2(n_7),
.A3(n_8),
.B1(n_10),
.B2(n_153),
.C1(n_141),
.C2(n_152),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_111),
.C(n_109),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_169),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_128),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g188 ( 
.A1(n_167),
.A2(n_172),
.B(n_169),
.Y(n_188)
);

NOR2x1_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_99),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_170),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_129),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_93),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_171),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_133),
.B(n_125),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_134),
.A2(n_82),
.B1(n_96),
.B2(n_113),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_153),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_136),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_154),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_165),
.C(n_168),
.Y(n_201)
);

AOI322xp5_ASAP7_75t_L g177 ( 
.A1(n_170),
.A2(n_148),
.A3(n_154),
.B1(n_131),
.B2(n_138),
.C1(n_151),
.C2(n_132),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_177),
.B(n_188),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_175),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_186),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_168),
.Y(n_204)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_136),
.Y(n_187)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_187),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_140),
.Y(n_189)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_189),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_191),
.B(n_171),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_193),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_159),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_197),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_152),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_164),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_207),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_204),
.C(n_206),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_192),
.A2(n_166),
.B1(n_157),
.B2(n_174),
.Y(n_202)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_141),
.C(n_166),
.Y(n_206)
);

AOI322xp5_ASAP7_75t_L g208 ( 
.A1(n_203),
.A2(n_180),
.A3(n_185),
.B1(n_192),
.B2(n_189),
.C1(n_187),
.C2(n_186),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_212),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_176),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_217),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_205),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_205),
.A2(n_196),
.B(n_192),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_214),
.A2(n_179),
.B(n_181),
.Y(n_225)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_185),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_213),
.A2(n_194),
.B1(n_200),
.B2(n_180),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_219),
.A2(n_221),
.B1(n_150),
.B2(n_151),
.Y(n_231)
);

AOI211xp5_ASAP7_75t_L g220 ( 
.A1(n_213),
.A2(n_202),
.B(n_194),
.C(n_182),
.Y(n_220)
);

OAI21xp33_ASAP7_75t_L g230 ( 
.A1(n_220),
.A2(n_201),
.B(n_173),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_214),
.A2(n_179),
.B1(n_171),
.B2(n_177),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_184),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_223),
.B(n_216),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_225),
.A2(n_215),
.B(n_181),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_211),
.C(n_217),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_226),
.B(n_228),
.Y(n_232)
);

AOI31xp67_ASAP7_75t_SL g234 ( 
.A1(n_227),
.A2(n_230),
.A3(n_220),
.B(n_221),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_211),
.C(n_210),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_231),
.C(n_218),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_230),
.A2(n_222),
.B(n_225),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_233),
.A2(n_139),
.B(n_8),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_234),
.A2(n_226),
.B1(n_228),
.B2(n_139),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_219),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_236),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_237),
.A2(n_238),
.B(n_232),
.Y(n_239)
);

AO21x1_ASAP7_75t_L g241 ( 
.A1(n_239),
.A2(n_7),
.B(n_10),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_240),
.Y(n_242)
);


endmodule