module fake_ariane_2220_n_1637 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1637);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1637;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_888;
wire n_845;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_91),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_15),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_16),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_76),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_113),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_134),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_71),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_96),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_149),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_30),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_36),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_43),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_103),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_3),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_24),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_86),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_129),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_84),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_67),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_58),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_81),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_118),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_16),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_11),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_15),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_31),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_43),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_12),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_139),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_0),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_89),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_88),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_51),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_53),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_19),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_137),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_19),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_98),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_57),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_99),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_23),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_107),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_17),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_110),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_17),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_12),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_66),
.Y(n_212)
);

BUFx8_ASAP7_75t_SL g213 ( 
.A(n_125),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_36),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_144),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_117),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_5),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_119),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_158),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_93),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_69),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_60),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_130),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_8),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_73),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_147),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_62),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_145),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_2),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_61),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_123),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_153),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_102),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_78),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_95),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_51),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_9),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_114),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_74),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_77),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_11),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_142),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_59),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_25),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_23),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_33),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_79),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_34),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_82),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_148),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_68),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_49),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_50),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_75),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_39),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_1),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_150),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_108),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_18),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_135),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_133),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_41),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_138),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_54),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_49),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_140),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_159),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_124),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_22),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_105),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_64),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_1),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_115),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_162),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_3),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_52),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_21),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_120),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_32),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_127),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_63),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_72),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_65),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_122),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_30),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_13),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_0),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_141),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_41),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_29),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_83),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_128),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_143),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_87),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_40),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_131),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_116),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_31),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_56),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_26),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_161),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_97),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_6),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_42),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_121),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_32),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_27),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_25),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_26),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_109),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_126),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_48),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_33),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_7),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_100),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_160),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_29),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_152),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_90),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_4),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_111),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_80),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_24),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_21),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_276),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_165),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_245),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_264),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_197),
.B(n_2),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_165),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_213),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_312),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_273),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_284),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_206),
.Y(n_335)
);

NOR2xp67_ASAP7_75t_L g336 ( 
.A(n_255),
.B(n_4),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_210),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_211),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_165),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_173),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_246),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_214),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_165),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_255),
.B(n_5),
.Y(n_344)
);

NOR2xp67_ASAP7_75t_L g345 ( 
.A(n_289),
.B(n_6),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_165),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_292),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_166),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_196),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_166),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_173),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_312),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_224),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_166),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_166),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_166),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_289),
.B(n_7),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_237),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_241),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_200),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_200),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_196),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_200),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_223),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_200),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_248),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_200),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_244),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_252),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_253),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_223),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_262),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_244),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_315),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_265),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_269),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_272),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_315),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_259),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_174),
.Y(n_380)
);

INVxp67_ASAP7_75t_SL g381 ( 
.A(n_323),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_174),
.Y(n_382)
);

INVxp33_ASAP7_75t_SL g383 ( 
.A(n_177),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_177),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_187),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_191),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_191),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_256),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_259),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_307),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_307),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_256),
.Y(n_392)
);

NOR2xp67_ASAP7_75t_L g393 ( 
.A(n_187),
.B(n_8),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_256),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_222),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_222),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_167),
.B(n_9),
.Y(n_397)
);

OR2x2_ASAP7_75t_L g398 ( 
.A(n_323),
.B(n_10),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_189),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_230),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_230),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_180),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_319),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_189),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_192),
.Y(n_405)
);

INVx4_ASAP7_75t_L g406 ( 
.A(n_402),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_333),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_347),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_341),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_R g410 ( 
.A(n_331),
.B(n_204),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_328),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_334),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_326),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_352),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_332),
.B(n_181),
.Y(n_415)
);

OA21x2_ASAP7_75t_L g416 ( 
.A1(n_397),
.A2(n_183),
.B(n_182),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_381),
.B(n_194),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_349),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_335),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_175),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_326),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_362),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_371),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_337),
.Y(n_424)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_371),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_338),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_395),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_395),
.Y(n_428)
);

INVx4_ASAP7_75t_L g429 ( 
.A(n_398),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_368),
.B(n_373),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_330),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_R g432 ( 
.A(n_342),
.B(n_205),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_330),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_353),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_336),
.B(n_178),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_339),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_358),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_339),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_R g439 ( 
.A(n_359),
.B(n_209),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_396),
.Y(n_440)
);

INVx6_ASAP7_75t_L g441 ( 
.A(n_398),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_404),
.A2(n_300),
.B1(n_202),
.B2(n_286),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_364),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_366),
.Y(n_444)
);

BUFx8_ASAP7_75t_L g445 ( 
.A(n_396),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_343),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_400),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_343),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_380),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_369),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_346),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_374),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_370),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_383),
.B(n_203),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_400),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_401),
.B(n_207),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_372),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_375),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_345),
.B(n_401),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_386),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_403),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_346),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_403),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_348),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_373),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_379),
.Y(n_466)
);

CKINVDCx8_ASAP7_75t_R g467 ( 
.A(n_405),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_378),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_379),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_348),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_376),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_350),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_377),
.B(n_212),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_350),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_354),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_387),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_354),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_454),
.A2(n_329),
.B1(n_384),
.B2(n_382),
.Y(n_478)
);

INVx5_ASAP7_75t_L g479 ( 
.A(n_413),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_448),
.Y(n_480)
);

OAI22xp33_ASAP7_75t_L g481 ( 
.A1(n_441),
.A2(n_325),
.B1(n_394),
.B2(n_385),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_423),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_406),
.B(n_344),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_448),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_409),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_414),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_406),
.B(n_357),
.Y(n_487)
);

INVx5_ASAP7_75t_L g488 ( 
.A(n_413),
.Y(n_488)
);

BUFx10_ASAP7_75t_L g489 ( 
.A(n_419),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_413),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_406),
.B(n_399),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_429),
.B(n_340),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_430),
.Y(n_493)
);

OR2x6_ASAP7_75t_L g494 ( 
.A(n_459),
.B(n_393),
.Y(n_494)
);

AND2x2_ASAP7_75t_SL g495 ( 
.A(n_429),
.B(n_319),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_473),
.B(n_351),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_430),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_413),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_407),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_427),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_448),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_428),
.Y(n_502)
);

OAI22xp33_ASAP7_75t_SL g503 ( 
.A1(n_441),
.A2(n_327),
.B1(n_195),
.B2(n_295),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_425),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_418),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_440),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_432),
.B(n_221),
.Y(n_507)
);

INVxp33_ASAP7_75t_L g508 ( 
.A(n_449),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_447),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_425),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_455),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_425),
.B(n_355),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_429),
.B(n_388),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_459),
.B(n_355),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_439),
.B(n_226),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_461),
.Y(n_516)
);

BUFx10_ASAP7_75t_L g517 ( 
.A(n_419),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_463),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_465),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_420),
.B(n_389),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_441),
.B(n_415),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_466),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_469),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_459),
.B(n_356),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_435),
.A2(n_285),
.B1(n_290),
.B2(n_303),
.Y(n_525)
);

BUFx4f_ASAP7_75t_L g526 ( 
.A(n_416),
.Y(n_526)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_460),
.B(n_202),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_451),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_420),
.B(n_389),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_441),
.A2(n_300),
.B1(n_286),
.B2(n_287),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_413),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_421),
.Y(n_532)
);

OR2x6_ASAP7_75t_L g533 ( 
.A(n_442),
.B(n_390),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_424),
.B(n_227),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_417),
.B(n_356),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g536 ( 
.A(n_467),
.B(n_392),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_435),
.A2(n_198),
.B1(n_188),
.B2(n_236),
.Y(n_537)
);

NOR2x1p5_ASAP7_75t_L g538 ( 
.A(n_424),
.B(n_287),
.Y(n_538)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_426),
.B(n_295),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_426),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_434),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_451),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_451),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_435),
.B(n_360),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_431),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_434),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_456),
.B(n_390),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_437),
.B(n_228),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_416),
.A2(n_324),
.B1(n_229),
.B2(n_298),
.Y(n_549)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_416),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_421),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_436),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_433),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_431),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_416),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_436),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_437),
.B(n_391),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_444),
.B(n_391),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_444),
.B(n_190),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_450),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_450),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_433),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_436),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_436),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_453),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_464),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_438),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_446),
.B(n_361),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_464),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_438),
.Y(n_570)
);

OR2x6_ASAP7_75t_L g571 ( 
.A(n_468),
.B(n_445),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_438),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_445),
.A2(n_217),
.B1(n_277),
.B2(n_208),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_477),
.B(n_361),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_477),
.B(n_472),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_453),
.B(n_235),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_472),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_445),
.A2(n_275),
.B1(n_279),
.B2(n_170),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_475),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_475),
.B(n_363),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_462),
.B(n_363),
.Y(n_581)
);

BUFx4f_ASAP7_75t_L g582 ( 
.A(n_462),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_462),
.B(n_365),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g584 ( 
.A(n_457),
.B(n_304),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_462),
.A2(n_271),
.B1(n_311),
.B2(n_306),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_462),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_457),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_470),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_470),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_470),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_470),
.Y(n_591)
);

AND2x2_ASAP7_75t_SL g592 ( 
.A(n_476),
.B(n_239),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_470),
.Y(n_593)
);

INVxp67_ASAP7_75t_SL g594 ( 
.A(n_474),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_474),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_458),
.A2(n_304),
.B1(n_306),
.B2(n_308),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_474),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_SL g598 ( 
.A1(n_407),
.A2(n_308),
.B1(n_309),
.B2(n_313),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_458),
.B(n_309),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_471),
.B(n_467),
.Y(n_600)
);

BUFx4f_ASAP7_75t_L g601 ( 
.A(n_474),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_471),
.B(n_365),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_408),
.B(n_240),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_410),
.B(n_249),
.Y(n_604)
);

NAND2xp33_ASAP7_75t_L g605 ( 
.A(n_408),
.B(n_280),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_468),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_411),
.B(n_250),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_411),
.B(n_258),
.Y(n_608)
);

INVx5_ASAP7_75t_L g609 ( 
.A(n_422),
.Y(n_609)
);

BUFx8_ASAP7_75t_SL g610 ( 
.A(n_412),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_412),
.B(n_260),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_443),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_452),
.B(n_261),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_454),
.B(n_268),
.Y(n_614)
);

OR2x2_ASAP7_75t_L g615 ( 
.A(n_460),
.B(n_313),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_425),
.Y(n_616)
);

BUFx10_ASAP7_75t_L g617 ( 
.A(n_419),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_480),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_521),
.B(n_164),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_495),
.B(n_164),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_480),
.Y(n_621)
);

O2A1O1Ixp5_ASAP7_75t_L g622 ( 
.A1(n_614),
.A2(n_293),
.B(n_305),
.C(n_297),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_484),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_496),
.B(n_314),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_495),
.B(n_314),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_526),
.B(n_168),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_484),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_540),
.B(n_317),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_501),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_547),
.B(n_168),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_534),
.B(n_548),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_606),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_526),
.B(n_169),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_547),
.B(n_169),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_526),
.B(n_171),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_501),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_528),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_485),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_534),
.B(n_317),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_528),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_542),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_542),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_576),
.B(n_171),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_549),
.A2(n_320),
.B1(n_288),
.B2(n_296),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_490),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_543),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_550),
.A2(n_320),
.B1(n_283),
.B2(n_294),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_548),
.B(n_172),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_614),
.A2(n_557),
.B1(n_558),
.B2(n_478),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_557),
.A2(n_186),
.B1(n_322),
.B2(n_321),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_558),
.B(n_172),
.Y(n_651)
);

INVx8_ASAP7_75t_L g652 ( 
.A(n_571),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_602),
.A2(n_186),
.B1(n_322),
.B2(n_321),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_543),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_545),
.Y(n_655)
);

NOR2x1p5_ASAP7_75t_L g656 ( 
.A(n_541),
.B(n_176),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_545),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_616),
.B(n_179),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_616),
.B(n_481),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_602),
.A2(n_193),
.B1(n_318),
.B2(n_316),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_539),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_539),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_532),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_482),
.B(n_493),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_551),
.Y(n_665)
);

OAI221xp5_ASAP7_75t_L g666 ( 
.A1(n_525),
.A2(n_282),
.B1(n_281),
.B2(n_291),
.C(n_310),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_553),
.Y(n_667)
);

NAND3xp33_ASAP7_75t_SL g668 ( 
.A(n_598),
.B(n_184),
.C(n_318),
.Y(n_668)
);

INVxp67_ASAP7_75t_R g669 ( 
.A(n_499),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_562),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_491),
.B(n_184),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_483),
.B(n_487),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_497),
.B(n_492),
.Y(n_673)
);

INVxp33_ASAP7_75t_L g674 ( 
.A(n_610),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_486),
.B(n_185),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_606),
.B(n_367),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_616),
.B(n_193),
.Y(n_677)
);

BUFx5_ASAP7_75t_L g678 ( 
.A(n_504),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_554),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_500),
.B(n_199),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_606),
.B(n_199),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_502),
.B(n_201),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_541),
.B(n_201),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_512),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_504),
.B(n_278),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_510),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_490),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_506),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_609),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_509),
.B(n_278),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_546),
.B(n_299),
.Y(n_691)
);

OAI221xp5_ASAP7_75t_L g692 ( 
.A1(n_537),
.A2(n_302),
.B1(n_301),
.B2(n_299),
.C(n_243),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_511),
.B(n_302),
.Y(n_693)
);

NAND2x1_ASAP7_75t_L g694 ( 
.A(n_556),
.B(n_280),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_516),
.B(n_301),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_609),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_594),
.A2(n_238),
.B(n_274),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_575),
.A2(n_234),
.B(n_270),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_546),
.B(n_280),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_584),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_518),
.B(n_215),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_609),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_510),
.B(n_10),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_554),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_519),
.B(n_216),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_531),
.A2(n_242),
.B(n_267),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_522),
.B(n_523),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_520),
.B(n_218),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_520),
.B(n_219),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_529),
.B(n_220),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_566),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_556),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_494),
.B(n_13),
.Y(n_713)
);

NOR2xp67_ASAP7_75t_SL g714 ( 
.A(n_560),
.B(n_251),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_494),
.B(n_14),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_514),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_529),
.B(n_225),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_524),
.B(n_231),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_584),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_566),
.Y(n_720)
);

NAND2xp33_ASAP7_75t_L g721 ( 
.A(n_490),
.B(n_254),
.Y(n_721)
);

HB1xp67_ASAP7_75t_L g722 ( 
.A(n_609),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_560),
.B(n_280),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_568),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_569),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_569),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_550),
.A2(n_280),
.B1(n_266),
.B2(n_263),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_494),
.B(n_14),
.Y(n_728)
);

NOR3xp33_ASAP7_75t_L g729 ( 
.A(n_587),
.B(n_513),
.C(n_596),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_550),
.A2(n_257),
.B1(n_247),
.B2(n_233),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_571),
.B(n_18),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_535),
.B(n_232),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_544),
.B(n_20),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_561),
.B(n_20),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_610),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_507),
.B(n_22),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_507),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_515),
.B(n_28),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_561),
.B(n_35),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_490),
.Y(n_740)
);

INVx2_ASAP7_75t_SL g741 ( 
.A(n_599),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_587),
.B(n_37),
.Y(n_742)
);

A2O1A1Ixp33_ASAP7_75t_L g743 ( 
.A1(n_603),
.A2(n_37),
.B(n_38),
.C(n_39),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_599),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_609),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_515),
.B(n_38),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_531),
.A2(n_92),
.B(n_155),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_494),
.B(n_40),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_574),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_577),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_579),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_580),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_556),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_600),
.B(n_42),
.Y(n_754)
);

INVx4_ASAP7_75t_L g755 ( 
.A(n_571),
.Y(n_755)
);

O2A1O1Ixp5_ASAP7_75t_L g756 ( 
.A1(n_564),
.A2(n_572),
.B(n_593),
.C(n_597),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_527),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_564),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_607),
.B(n_530),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_581),
.Y(n_760)
);

OAI221xp5_ASAP7_75t_L g761 ( 
.A1(n_585),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.C(n_47),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_583),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_565),
.B(n_44),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_555),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_527),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_565),
.B(n_48),
.Y(n_766)
);

INVxp67_ASAP7_75t_L g767 ( 
.A(n_608),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_498),
.B(n_50),
.Y(n_768)
);

OR2x6_ASAP7_75t_L g769 ( 
.A(n_571),
.B(n_52),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_586),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_607),
.B(n_55),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_555),
.A2(n_70),
.B1(n_85),
.B2(n_94),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_586),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_498),
.B(n_101),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_611),
.B(n_156),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_604),
.B(n_104),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_589),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_485),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_555),
.B(n_106),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_L g780 ( 
.A1(n_649),
.A2(n_533),
.B1(n_559),
.B2(n_573),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_654),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_672),
.A2(n_559),
.B(n_582),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_767),
.B(n_604),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_664),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_672),
.B(n_617),
.Y(n_785)
);

OAI22xp5_ASAP7_75t_L g786 ( 
.A1(n_764),
.A2(n_533),
.B1(n_578),
.B2(n_508),
.Y(n_786)
);

O2A1O1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_624),
.A2(n_533),
.B(n_605),
.C(n_508),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_628),
.B(n_617),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_624),
.B(n_617),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_688),
.Y(n_790)
);

O2A1O1Ixp33_ASAP7_75t_L g791 ( 
.A1(n_743),
.A2(n_533),
.B(n_605),
.C(n_615),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_631),
.B(n_489),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_764),
.A2(n_538),
.B1(n_592),
.B2(n_615),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_633),
.A2(n_601),
.B(n_563),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_661),
.B(n_517),
.Y(n_795)
);

AOI21x1_ASAP7_75t_L g796 ( 
.A1(n_633),
.A2(n_591),
.B(n_589),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_663),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_631),
.B(n_517),
.Y(n_798)
);

OR2x2_ASAP7_75t_L g799 ( 
.A(n_638),
.B(n_778),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_671),
.B(n_517),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_635),
.A2(n_601),
.B(n_552),
.Y(n_801)
);

O2A1O1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_743),
.A2(n_503),
.B(n_613),
.C(n_552),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_632),
.Y(n_803)
);

INVxp67_ASAP7_75t_SL g804 ( 
.A(n_645),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_671),
.B(n_489),
.Y(n_805)
);

BUFx4f_ASAP7_75t_L g806 ( 
.A(n_652),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_635),
.A2(n_552),
.B(n_567),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_759),
.B(n_489),
.Y(n_808)
);

NAND3xp33_ASAP7_75t_L g809 ( 
.A(n_625),
.B(n_612),
.C(n_536),
.Y(n_809)
);

CKINVDCx8_ASAP7_75t_R g810 ( 
.A(n_735),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_759),
.A2(n_592),
.B1(n_531),
.B2(n_563),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_662),
.B(n_613),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_618),
.A2(n_563),
.B(n_570),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_L g814 ( 
.A1(n_647),
.A2(n_567),
.B1(n_570),
.B2(n_593),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_629),
.A2(n_567),
.B(n_570),
.Y(n_815)
);

BUFx2_ASAP7_75t_SL g816 ( 
.A(n_689),
.Y(n_816)
);

INVx4_ASAP7_75t_L g817 ( 
.A(n_652),
.Y(n_817)
);

A2O1A1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_625),
.A2(n_771),
.B(n_639),
.C(n_648),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_643),
.B(n_716),
.Y(n_819)
);

NOR2xp67_ASAP7_75t_L g820 ( 
.A(n_700),
.B(n_597),
.Y(n_820)
);

CKINVDCx6p67_ASAP7_75t_R g821 ( 
.A(n_769),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_637),
.A2(n_597),
.B(n_593),
.Y(n_822)
);

BUFx4f_ASAP7_75t_L g823 ( 
.A(n_652),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_640),
.A2(n_572),
.B(n_564),
.Y(n_824)
);

NOR3xp33_ASAP7_75t_L g825 ( 
.A(n_668),
.B(n_572),
.C(n_505),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_641),
.A2(n_595),
.B(n_590),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_719),
.B(n_741),
.Y(n_827)
);

NAND3xp33_ASAP7_75t_L g828 ( 
.A(n_648),
.B(n_505),
.C(n_595),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_646),
.A2(n_590),
.B(n_588),
.Y(n_829)
);

AOI21x1_ASAP7_75t_L g830 ( 
.A1(n_776),
.A2(n_590),
.B(n_588),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_621),
.A2(n_590),
.B(n_588),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_754),
.B(n_590),
.Y(n_832)
);

NAND2x1p5_ASAP7_75t_L g833 ( 
.A(n_696),
.B(n_702),
.Y(n_833)
);

O2A1O1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_673),
.A2(n_488),
.B(n_479),
.C(n_588),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_647),
.A2(n_588),
.B1(n_498),
.B2(n_488),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_665),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_623),
.A2(n_498),
.B(n_488),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_630),
.B(n_498),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_627),
.A2(n_488),
.B(n_479),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_756),
.A2(n_488),
.B(n_479),
.Y(n_840)
);

AOI21x1_ASAP7_75t_L g841 ( 
.A1(n_657),
.A2(n_479),
.B(n_132),
.Y(n_841)
);

NAND3xp33_ASAP7_75t_L g842 ( 
.A(n_639),
.B(n_479),
.C(n_136),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_644),
.A2(n_112),
.B1(n_146),
.B2(n_151),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_644),
.A2(n_154),
.B1(n_620),
.B2(n_775),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_634),
.B(n_724),
.Y(n_845)
);

OR2x2_ASAP7_75t_L g846 ( 
.A(n_744),
.B(n_757),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_632),
.B(n_681),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_712),
.Y(n_848)
);

OAI21xp5_ASAP7_75t_L g849 ( 
.A1(n_684),
.A2(n_733),
.B(n_636),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_669),
.B(n_765),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_620),
.A2(n_729),
.B1(n_659),
.B2(n_771),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_642),
.A2(n_707),
.B(n_677),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_749),
.B(n_619),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_683),
.B(n_691),
.Y(n_854)
);

OAI21x1_ASAP7_75t_L g855 ( 
.A1(n_679),
.A2(n_711),
.B(n_704),
.Y(n_855)
);

NOR3xp33_ASAP7_75t_L g856 ( 
.A(n_734),
.B(n_739),
.C(n_763),
.Y(n_856)
);

NOR3xp33_ASAP7_75t_L g857 ( 
.A(n_734),
.B(n_739),
.C(n_763),
.Y(n_857)
);

A2O1A1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_703),
.A2(n_748),
.B(n_713),
.C(n_715),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_685),
.B(n_651),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_683),
.B(n_691),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_659),
.B(n_681),
.Y(n_861)
);

O2A1O1Ixp33_ASAP7_75t_SL g862 ( 
.A1(n_658),
.A2(n_677),
.B(n_768),
.C(n_774),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_766),
.B(n_685),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_645),
.Y(n_864)
);

O2A1O1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_708),
.A2(n_717),
.B(n_710),
.C(n_709),
.Y(n_865)
);

NOR2xp67_ASAP7_75t_SL g866 ( 
.A(n_742),
.B(n_761),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_703),
.A2(n_667),
.B(n_670),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_658),
.A2(n_712),
.B(n_758),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_753),
.A2(n_758),
.B(n_686),
.Y(n_869)
);

AOI33xp33_ASAP7_75t_L g870 ( 
.A1(n_650),
.A2(n_737),
.A3(n_660),
.B1(n_653),
.B2(n_730),
.B3(n_727),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_753),
.A2(n_686),
.B(n_718),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_751),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_745),
.B(n_715),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_732),
.A2(n_701),
.B(n_705),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_645),
.Y(n_875)
);

NAND3xp33_ASAP7_75t_L g876 ( 
.A(n_730),
.B(n_727),
.C(n_692),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_752),
.B(n_762),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_713),
.B(n_728),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_731),
.B(n_728),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_760),
.B(n_676),
.Y(n_880)
);

NAND3xp33_ASAP7_75t_L g881 ( 
.A(n_748),
.B(n_736),
.C(n_738),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_676),
.B(n_680),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_682),
.B(n_695),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_690),
.B(n_693),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_720),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_622),
.A2(n_746),
.B(n_772),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_725),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_698),
.A2(n_777),
.B(n_773),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_770),
.A2(n_675),
.B(n_645),
.Y(n_889)
);

NOR2x1_ASAP7_75t_L g890 ( 
.A(n_656),
.B(n_755),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_687),
.A2(n_740),
.B(n_726),
.Y(n_891)
);

NOR2x1_ASAP7_75t_L g892 ( 
.A(n_755),
.B(n_769),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_687),
.A2(n_740),
.B(n_697),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_687),
.A2(n_740),
.B(n_706),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_687),
.A2(n_740),
.B(n_750),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_722),
.Y(n_896)
);

INVx4_ASAP7_75t_L g897 ( 
.A(n_769),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_774),
.A2(n_694),
.B(n_723),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_699),
.A2(n_723),
.B(n_721),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_678),
.B(n_714),
.Y(n_900)
);

INVx5_ASAP7_75t_L g901 ( 
.A(n_731),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_722),
.B(n_747),
.Y(n_902)
);

A2O1A1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_666),
.A2(n_759),
.B(n_631),
.C(n_625),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_678),
.A2(n_672),
.B(n_633),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_678),
.B(n_674),
.Y(n_905)
);

O2A1O1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_678),
.A2(n_767),
.B(n_624),
.C(n_614),
.Y(n_906)
);

AO22x1_ASAP7_75t_L g907 ( 
.A1(n_678),
.A2(n_407),
.B1(n_600),
.B2(n_333),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_672),
.A2(n_633),
.B(n_626),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_672),
.A2(n_633),
.B(n_626),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_767),
.B(n_521),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_672),
.A2(n_779),
.B(n_526),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_672),
.A2(n_633),
.B(n_626),
.Y(n_912)
);

NOR2xp67_ASAP7_75t_L g913 ( 
.A(n_767),
.B(n_609),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_SL g914 ( 
.A(n_735),
.B(n_407),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_672),
.A2(n_633),
.B(n_626),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_759),
.A2(n_631),
.B1(n_625),
.B2(n_767),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_672),
.A2(n_779),
.B(n_526),
.Y(n_917)
);

NAND3xp33_ASAP7_75t_L g918 ( 
.A(n_624),
.B(n_767),
.C(n_424),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_759),
.A2(n_631),
.B(n_625),
.C(n_624),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_767),
.B(n_521),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_672),
.A2(n_633),
.B(n_626),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_645),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_778),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_767),
.A2(n_624),
.B(n_614),
.C(n_743),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_778),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_767),
.B(n_521),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_759),
.A2(n_631),
.B1(n_625),
.B2(n_767),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_767),
.B(n_333),
.Y(n_928)
);

AOI22x1_ASAP7_75t_L g929 ( 
.A1(n_663),
.A2(n_665),
.B1(n_670),
.B2(n_667),
.Y(n_929)
);

OAI21x1_ASAP7_75t_L g930 ( 
.A1(n_756),
.A2(n_657),
.B(n_655),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_672),
.A2(n_779),
.B(n_526),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_672),
.A2(n_633),
.B(n_626),
.Y(n_932)
);

CKINVDCx10_ASAP7_75t_R g933 ( 
.A(n_735),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_767),
.B(n_521),
.Y(n_934)
);

OAI221xp5_ASAP7_75t_L g935 ( 
.A1(n_759),
.A2(n_649),
.B1(n_624),
.B2(n_639),
.C(n_631),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_672),
.A2(n_633),
.B(n_626),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_649),
.B(n_495),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_767),
.B(n_521),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_767),
.B(n_333),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_767),
.B(n_521),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_767),
.B(n_521),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_649),
.B(n_495),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_628),
.B(n_540),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_767),
.B(n_521),
.Y(n_944)
);

INVx5_ASAP7_75t_L g945 ( 
.A(n_645),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_645),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_632),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_672),
.A2(n_633),
.B(n_626),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_632),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_767),
.B(n_333),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_632),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_664),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_664),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_672),
.B(n_724),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_911),
.A2(n_931),
.B(n_917),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_935),
.B(n_785),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_818),
.B(n_851),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_943),
.B(n_879),
.Y(n_958)
);

CKINVDCx20_ASAP7_75t_R g959 ( 
.A(n_810),
.Y(n_959)
);

OAI21x1_ASAP7_75t_L g960 ( 
.A1(n_904),
.A2(n_841),
.B(n_893),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_954),
.B(n_920),
.Y(n_961)
);

NOR2xp67_ASAP7_75t_L g962 ( 
.A(n_918),
.B(n_901),
.Y(n_962)
);

INVxp67_ASAP7_75t_L g963 ( 
.A(n_846),
.Y(n_963)
);

A2O1A1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_919),
.A2(n_903),
.B(n_927),
.C(n_916),
.Y(n_964)
);

NAND3xp33_ASAP7_75t_SL g965 ( 
.A(n_808),
.B(n_787),
.C(n_928),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_908),
.A2(n_912),
.B(n_909),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_926),
.B(n_934),
.Y(n_967)
);

OAI21x1_ASAP7_75t_L g968 ( 
.A1(n_894),
.A2(n_921),
.B(n_915),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_827),
.B(n_812),
.Y(n_969)
);

OAI21x1_ASAP7_75t_L g970 ( 
.A1(n_932),
.A2(n_948),
.B(n_936),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_911),
.A2(n_931),
.B(n_917),
.Y(n_971)
);

OAI21xp33_ASAP7_75t_L g972 ( 
.A1(n_939),
.A2(n_950),
.B(n_870),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_938),
.B(n_940),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_874),
.A2(n_853),
.B(n_782),
.Y(n_974)
);

BUFx3_ASAP7_75t_L g975 ( 
.A(n_806),
.Y(n_975)
);

OAI21x1_ASAP7_75t_L g976 ( 
.A1(n_829),
.A2(n_898),
.B(n_855),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_817),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_941),
.B(n_944),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_876),
.A2(n_852),
.B(n_865),
.Y(n_979)
);

AO31x2_ASAP7_75t_L g980 ( 
.A1(n_844),
.A2(n_861),
.A3(n_811),
.B(n_835),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_819),
.A2(n_871),
.B(n_832),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_878),
.B(n_792),
.Y(n_982)
);

OAI21x1_ASAP7_75t_L g983 ( 
.A1(n_889),
.A2(n_888),
.B(n_899),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_883),
.A2(n_884),
.B(n_906),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_806),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_845),
.B(n_859),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_789),
.B(n_798),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_780),
.A2(n_786),
.B1(n_793),
.B2(n_937),
.Y(n_988)
);

BUFx2_ASAP7_75t_L g989 ( 
.A(n_925),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_924),
.A2(n_791),
.B(n_858),
.C(n_854),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_862),
.A2(n_900),
.B(n_838),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_780),
.B(n_786),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_877),
.A2(n_849),
.B(n_844),
.Y(n_993)
);

OAI21x1_ASAP7_75t_L g994 ( 
.A1(n_849),
.A2(n_801),
.B(n_794),
.Y(n_994)
);

BUFx2_ASAP7_75t_L g995 ( 
.A(n_850),
.Y(n_995)
);

OAI21x1_ASAP7_75t_L g996 ( 
.A1(n_840),
.A2(n_807),
.B(n_895),
.Y(n_996)
);

OAI21x1_ASAP7_75t_SL g997 ( 
.A1(n_929),
.A2(n_886),
.B(n_868),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_799),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_783),
.B(n_907),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_784),
.B(n_952),
.Y(n_1000)
);

OAI21x1_ASAP7_75t_L g1001 ( 
.A1(n_840),
.A2(n_891),
.B(n_826),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_817),
.Y(n_1002)
);

OAI22x1_ASAP7_75t_L g1003 ( 
.A1(n_901),
.A2(n_942),
.B1(n_897),
.B2(n_860),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_793),
.B(n_863),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_788),
.B(n_795),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_L g1006 ( 
.A1(n_831),
.A2(n_837),
.B(n_813),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_856),
.A2(n_857),
.B(n_886),
.C(n_866),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_815),
.A2(n_834),
.B(n_839),
.Y(n_1008)
);

OAI21x1_ASAP7_75t_L g1009 ( 
.A1(n_869),
.A2(n_824),
.B(n_822),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_953),
.B(n_880),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_902),
.A2(n_847),
.B(n_882),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_790),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_902),
.A2(n_951),
.B(n_949),
.Y(n_1013)
);

OAI21x1_ASAP7_75t_L g1014 ( 
.A1(n_835),
.A2(n_842),
.B(n_814),
.Y(n_1014)
);

INVx3_ASAP7_75t_L g1015 ( 
.A(n_945),
.Y(n_1015)
);

AO21x1_ASAP7_75t_L g1016 ( 
.A1(n_843),
.A2(n_811),
.B(n_873),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_945),
.B(n_946),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_814),
.A2(n_781),
.B(n_833),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_901),
.B(n_797),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_881),
.A2(n_802),
.B(n_843),
.C(n_836),
.Y(n_1020)
);

OAI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_872),
.A2(n_848),
.B(n_896),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_892),
.B(n_897),
.Y(n_1022)
);

OR2x2_ASAP7_75t_L g1023 ( 
.A(n_809),
.B(n_828),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_L g1024 ( 
.A1(n_875),
.A2(n_803),
.B(n_949),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_803),
.A2(n_951),
.B(n_947),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_848),
.A2(n_947),
.B(n_804),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_945),
.B(n_946),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_885),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_905),
.A2(n_887),
.B(n_890),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_913),
.A2(n_820),
.B(n_922),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_864),
.A2(n_922),
.B(n_823),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_825),
.B(n_823),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_816),
.B(n_864),
.Y(n_1033)
);

OA21x2_ASAP7_75t_L g1034 ( 
.A1(n_821),
.A2(n_914),
.B(n_933),
.Y(n_1034)
);

OAI21x1_ASAP7_75t_L g1035 ( 
.A1(n_830),
.A2(n_930),
.B(n_796),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_830),
.A2(n_930),
.B(n_796),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_911),
.A2(n_931),
.B(n_917),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_830),
.A2(n_930),
.B(n_796),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_830),
.A2(n_930),
.B(n_796),
.Y(n_1039)
);

INVxp67_ASAP7_75t_L g1040 ( 
.A(n_846),
.Y(n_1040)
);

BUFx10_ASAP7_75t_L g1041 ( 
.A(n_928),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_830),
.A2(n_930),
.B(n_796),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_911),
.A2(n_931),
.B(n_917),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_817),
.B(n_901),
.Y(n_1044)
);

BUFx12f_ASAP7_75t_L g1045 ( 
.A(n_923),
.Y(n_1045)
);

OAI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_935),
.A2(n_927),
.B1(n_916),
.B2(n_780),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_919),
.A2(n_954),
.B(n_818),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_954),
.B(n_910),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_954),
.B(n_910),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_919),
.A2(n_954),
.B(n_818),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_943),
.B(n_879),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_923),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_L g1053 ( 
.A1(n_830),
.A2(n_930),
.B(n_796),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_830),
.A2(n_930),
.B(n_796),
.Y(n_1054)
);

AOI211x1_ASAP7_75t_L g1055 ( 
.A1(n_935),
.A2(n_954),
.B(n_866),
.C(n_867),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_830),
.A2(n_930),
.B(n_796),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_790),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_817),
.Y(n_1058)
);

INVx3_ASAP7_75t_SL g1059 ( 
.A(n_799),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_923),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_954),
.B(n_910),
.Y(n_1061)
);

NAND2x1p5_ASAP7_75t_L g1062 ( 
.A(n_901),
.B(n_817),
.Y(n_1062)
);

INVx2_ASAP7_75t_SL g1063 ( 
.A(n_925),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_935),
.B(n_785),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_830),
.A2(n_930),
.B(n_796),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_954),
.B(n_910),
.Y(n_1066)
);

AOI211x1_ASAP7_75t_L g1067 ( 
.A1(n_935),
.A2(n_954),
.B(n_866),
.C(n_867),
.Y(n_1067)
);

AO31x2_ASAP7_75t_L g1068 ( 
.A1(n_818),
.A2(n_844),
.A3(n_909),
.B(n_908),
.Y(n_1068)
);

O2A1O1Ixp5_ASAP7_75t_L g1069 ( 
.A1(n_818),
.A2(n_800),
.B(n_805),
.C(n_911),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_919),
.A2(n_954),
.B(n_818),
.Y(n_1070)
);

OR2x2_ASAP7_75t_L g1071 ( 
.A(n_799),
.B(n_411),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_790),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_817),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_945),
.Y(n_1074)
);

INVx4_ASAP7_75t_L g1075 ( 
.A(n_901),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_830),
.A2(n_930),
.B(n_796),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_954),
.B(n_910),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_945),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_830),
.A2(n_930),
.B(n_796),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_SL g1080 ( 
.A1(n_966),
.A2(n_956),
.B(n_1064),
.C(n_1070),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_1045),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_956),
.B(n_1064),
.Y(n_1082)
);

INVx3_ASAP7_75t_SL g1083 ( 
.A(n_959),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_959),
.Y(n_1084)
);

INVx1_ASAP7_75t_SL g1085 ( 
.A(n_995),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_989),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_1045),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1012),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_957),
.A2(n_1050),
.B(n_971),
.Y(n_1089)
);

OR2x6_ASAP7_75t_L g1090 ( 
.A(n_1044),
.B(n_992),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1057),
.Y(n_1091)
);

INVx1_ASAP7_75t_SL g1092 ( 
.A(n_998),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1072),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_1074),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1004),
.A2(n_972),
.B1(n_992),
.B2(n_1046),
.Y(n_1095)
);

OA21x2_ASAP7_75t_L g1096 ( 
.A1(n_968),
.A2(n_983),
.B(n_970),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_975),
.B(n_985),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_1044),
.B(n_1022),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_955),
.A2(n_1043),
.B(n_1037),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_988),
.A2(n_1004),
.B1(n_1046),
.B2(n_1016),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_961),
.B(n_1048),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_993),
.A2(n_964),
.B(n_1020),
.C(n_990),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_1071),
.A2(n_969),
.B1(n_1023),
.B2(n_965),
.Y(n_1103)
);

OR2x6_ASAP7_75t_L g1104 ( 
.A(n_1022),
.B(n_1075),
.Y(n_1104)
);

INVxp67_ASAP7_75t_SL g1105 ( 
.A(n_963),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_1041),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1049),
.B(n_1061),
.Y(n_1107)
);

CKINVDCx16_ASAP7_75t_R g1108 ( 
.A(n_1041),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_986),
.A2(n_1028),
.B1(n_1066),
.B2(n_1077),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_967),
.B(n_973),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_964),
.A2(n_990),
.B1(n_1007),
.B2(n_1067),
.Y(n_1111)
);

AOI221xp5_ASAP7_75t_L g1112 ( 
.A1(n_1055),
.A2(n_978),
.B1(n_1020),
.B2(n_1007),
.C(n_982),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_982),
.B(n_987),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1005),
.B(n_1040),
.Y(n_1114)
);

NOR2x1_ASAP7_75t_SL g1115 ( 
.A(n_1074),
.B(n_1078),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_1041),
.Y(n_1116)
);

CKINVDCx16_ASAP7_75t_R g1117 ( 
.A(n_1052),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1000),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_984),
.B(n_1010),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_1060),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1011),
.B(n_974),
.Y(n_1121)
);

NAND2xp33_ASAP7_75t_SL g1122 ( 
.A(n_1059),
.B(n_977),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_1074),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_999),
.B(n_980),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1019),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_981),
.A2(n_1013),
.B(n_1069),
.Y(n_1126)
);

OR2x2_ASAP7_75t_L g1127 ( 
.A(n_1034),
.B(n_1032),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_980),
.B(n_1021),
.Y(n_1128)
);

INVx1_ASAP7_75t_SL g1129 ( 
.A(n_1033),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_977),
.B(n_1058),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_962),
.A2(n_979),
.B1(n_1002),
.B2(n_1073),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_1062),
.B(n_1015),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_980),
.A2(n_1026),
.B1(n_1025),
.B2(n_991),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1015),
.B(n_1078),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_1074),
.B(n_1078),
.Y(n_1135)
);

INVx5_ASAP7_75t_L g1136 ( 
.A(n_1078),
.Y(n_1136)
);

OAI22xp33_ASAP7_75t_L g1137 ( 
.A1(n_1003),
.A2(n_1031),
.B1(n_1027),
.B2(n_1017),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_997),
.A2(n_968),
.B(n_970),
.Y(n_1138)
);

AOI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1014),
.A2(n_1018),
.B1(n_1029),
.B2(n_1030),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1068),
.B(n_1018),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1068),
.B(n_1024),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_1024),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_1068),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_994),
.Y(n_1144)
);

CKINVDCx11_ASAP7_75t_R g1145 ( 
.A(n_994),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_996),
.B(n_1001),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_SL g1147 ( 
.A(n_1008),
.B(n_1006),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_960),
.A2(n_1009),
.B(n_1079),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_976),
.A2(n_960),
.B1(n_1035),
.B2(n_1036),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_976),
.Y(n_1150)
);

AND2x6_ASAP7_75t_L g1151 ( 
.A(n_1035),
.B(n_1036),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_1038),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_1039),
.B(n_1042),
.Y(n_1153)
);

BUFx12f_ASAP7_75t_L g1154 ( 
.A(n_1039),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_1053),
.Y(n_1155)
);

BUFx12f_ASAP7_75t_L g1156 ( 
.A(n_1053),
.Y(n_1156)
);

AND2x6_ASAP7_75t_L g1157 ( 
.A(n_1054),
.B(n_1056),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_1054),
.B(n_1056),
.Y(n_1158)
);

NAND3xp33_ASAP7_75t_L g1159 ( 
.A(n_1065),
.B(n_1079),
.C(n_1076),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_975),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_992),
.A2(n_935),
.B1(n_916),
.B2(n_927),
.Y(n_1161)
);

OR2x6_ASAP7_75t_SL g1162 ( 
.A(n_1071),
.B(n_778),
.Y(n_1162)
);

A2O1A1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_956),
.A2(n_818),
.B(n_935),
.C(n_919),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_1074),
.Y(n_1164)
);

INVx6_ASAP7_75t_L g1165 ( 
.A(n_1045),
.Y(n_1165)
);

INVx2_ASAP7_75t_SL g1166 ( 
.A(n_1045),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_958),
.B(n_1051),
.Y(n_1167)
);

OR2x2_ASAP7_75t_L g1168 ( 
.A(n_958),
.B(n_1051),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1012),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_959),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_972),
.A2(n_919),
.B(n_818),
.C(n_935),
.Y(n_1171)
);

AOI221xp5_ASAP7_75t_L g1172 ( 
.A1(n_1046),
.A2(n_935),
.B1(n_780),
.B2(n_972),
.C(n_919),
.Y(n_1172)
);

O2A1O1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_972),
.A2(n_919),
.B(n_818),
.C(n_935),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_956),
.B(n_1064),
.Y(n_1174)
);

NOR2x1_ASAP7_75t_SL g1175 ( 
.A(n_1074),
.B(n_1078),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_956),
.B(n_1064),
.Y(n_1176)
);

INVxp67_ASAP7_75t_SL g1177 ( 
.A(n_963),
.Y(n_1177)
);

BUFx10_ASAP7_75t_L g1178 ( 
.A(n_1063),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1012),
.Y(n_1179)
);

NAND3xp33_ASAP7_75t_L g1180 ( 
.A(n_956),
.B(n_935),
.C(n_818),
.Y(n_1180)
);

INVx2_ASAP7_75t_SL g1181 ( 
.A(n_1045),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_958),
.B(n_1051),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_SL g1183 ( 
.A1(n_1016),
.A2(n_1050),
.B(n_1047),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_956),
.A2(n_818),
.B(n_935),
.C(n_919),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_956),
.B(n_1064),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_956),
.B(n_1064),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_972),
.A2(n_919),
.B(n_818),
.C(n_935),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_956),
.A2(n_818),
.B(n_935),
.C(n_919),
.Y(n_1188)
);

BUFx2_ASAP7_75t_SL g1189 ( 
.A(n_1084),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_1170),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1088),
.Y(n_1191)
);

CKINVDCx6p67_ASAP7_75t_R g1192 ( 
.A(n_1083),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_1136),
.Y(n_1193)
);

BUFx12f_ASAP7_75t_L g1194 ( 
.A(n_1106),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1091),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1093),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_1086),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1161),
.A2(n_1172),
.B1(n_1095),
.B2(n_1100),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1148),
.A2(n_1138),
.B(n_1126),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1161),
.A2(n_1172),
.B1(n_1180),
.B2(n_1186),
.Y(n_1200)
);

INVx11_ASAP7_75t_L g1201 ( 
.A(n_1154),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1082),
.A2(n_1176),
.B1(n_1185),
.B2(n_1174),
.Y(n_1202)
);

CKINVDCx11_ASAP7_75t_R g1203 ( 
.A(n_1162),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1169),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1174),
.A2(n_1185),
.B1(n_1176),
.B2(n_1186),
.Y(n_1205)
);

INVx4_ASAP7_75t_L g1206 ( 
.A(n_1090),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_1092),
.Y(n_1207)
);

BUFx2_ASAP7_75t_L g1208 ( 
.A(n_1156),
.Y(n_1208)
);

CKINVDCx11_ASAP7_75t_R g1209 ( 
.A(n_1117),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1179),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1118),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1125),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_1116),
.Y(n_1213)
);

AO21x1_ASAP7_75t_L g1214 ( 
.A1(n_1171),
.A2(n_1187),
.B(n_1173),
.Y(n_1214)
);

AOI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1110),
.A2(n_1103),
.B1(n_1112),
.B2(n_1182),
.Y(n_1215)
);

BUFx12f_ASAP7_75t_L g1216 ( 
.A(n_1120),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_1108),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1112),
.A2(n_1127),
.B1(n_1111),
.B2(n_1167),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_1092),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_1150),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1143),
.Y(n_1221)
);

OR2x2_ASAP7_75t_L g1222 ( 
.A(n_1124),
.B(n_1128),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1141),
.Y(n_1223)
);

INVx8_ASAP7_75t_L g1224 ( 
.A(n_1104),
.Y(n_1224)
);

BUFx12f_ASAP7_75t_L g1225 ( 
.A(n_1178),
.Y(n_1225)
);

INVx4_ASAP7_75t_L g1226 ( 
.A(n_1094),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1163),
.A2(n_1188),
.B(n_1184),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1129),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1183),
.A2(n_1107),
.B1(n_1101),
.B2(n_1124),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1129),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1119),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_1145),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1101),
.A2(n_1107),
.B1(n_1114),
.B2(n_1109),
.Y(n_1233)
);

BUFx8_ASAP7_75t_L g1234 ( 
.A(n_1081),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1119),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_1168),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1113),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1142),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1099),
.A2(n_1121),
.B(n_1089),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1158),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1080),
.B(n_1105),
.Y(n_1241)
);

OAI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1085),
.A2(n_1177),
.B1(n_1165),
.B2(n_1087),
.Y(n_1242)
);

INVx3_ASAP7_75t_L g1243 ( 
.A(n_1094),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1165),
.A2(n_1089),
.B1(n_1181),
.B2(n_1166),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1131),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1131),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1102),
.Y(n_1247)
);

BUFx2_ASAP7_75t_R g1248 ( 
.A(n_1135),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_SL g1249 ( 
.A1(n_1133),
.A2(n_1160),
.B1(n_1115),
.B2(n_1175),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1121),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1134),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1155),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1123),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1123),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_1160),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1164),
.B(n_1140),
.Y(n_1256)
);

AO21x2_ASAP7_75t_L g1257 ( 
.A1(n_1149),
.A2(n_1159),
.B(n_1139),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1146),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1146),
.Y(n_1259)
);

CKINVDCx6p67_ASAP7_75t_R g1260 ( 
.A(n_1178),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_1151),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1160),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1132),
.B(n_1130),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1137),
.Y(n_1264)
);

INVxp67_ASAP7_75t_L g1265 ( 
.A(n_1097),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1122),
.Y(n_1266)
);

INVx1_ASAP7_75t_SL g1267 ( 
.A(n_1151),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1144),
.A2(n_1152),
.B1(n_1153),
.B2(n_1096),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1151),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1147),
.B(n_1151),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_SL g1271 ( 
.A1(n_1147),
.A2(n_992),
.B1(n_780),
.B2(n_935),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1157),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1157),
.B(n_992),
.Y(n_1273)
);

AOI22xp5_ASAP7_75t_SL g1274 ( 
.A1(n_1082),
.A2(n_780),
.B1(n_992),
.B2(n_786),
.Y(n_1274)
);

CKINVDCx6p67_ASAP7_75t_R g1275 ( 
.A(n_1083),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1092),
.Y(n_1276)
);

AND2x4_ASAP7_75t_L g1277 ( 
.A(n_1090),
.B(n_1098),
.Y(n_1277)
);

CKINVDCx10_ASAP7_75t_R g1278 ( 
.A(n_1117),
.Y(n_1278)
);

CKINVDCx11_ASAP7_75t_R g1279 ( 
.A(n_1083),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1223),
.B(n_1273),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1238),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1223),
.B(n_1273),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_1207),
.Y(n_1283)
);

OAI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1227),
.A2(n_1200),
.B(n_1198),
.Y(n_1284)
);

INVx3_ASAP7_75t_L g1285 ( 
.A(n_1258),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1250),
.Y(n_1286)
);

OR2x6_ASAP7_75t_L g1287 ( 
.A(n_1224),
.B(n_1206),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1231),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1219),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1237),
.B(n_1202),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1276),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1235),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1256),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1238),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1222),
.Y(n_1295)
);

INVx4_ASAP7_75t_L g1296 ( 
.A(n_1201),
.Y(n_1296)
);

AOI21xp33_ASAP7_75t_L g1297 ( 
.A1(n_1214),
.A2(n_1274),
.B(n_1241),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_1209),
.Y(n_1298)
);

BUFx12f_ASAP7_75t_L g1299 ( 
.A(n_1209),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1222),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1193),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1190),
.B(n_1197),
.Y(n_1302)
);

AOI21xp33_ASAP7_75t_L g1303 ( 
.A1(n_1214),
.A2(n_1264),
.B(n_1228),
.Y(n_1303)
);

NAND2x1_ASAP7_75t_L g1304 ( 
.A(n_1245),
.B(n_1246),
.Y(n_1304)
);

CKINVDCx20_ASAP7_75t_R g1305 ( 
.A(n_1279),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1191),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1220),
.B(n_1240),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1269),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1195),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1272),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_1201),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1221),
.B(n_1259),
.Y(n_1312)
);

AOI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1199),
.A2(n_1239),
.B(n_1268),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1271),
.B(n_1196),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1236),
.B(n_1232),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1204),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1210),
.Y(n_1317)
);

INVx1_ASAP7_75t_SL g1318 ( 
.A(n_1255),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1261),
.B(n_1229),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1212),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1211),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1252),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1252),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1205),
.B(n_1233),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1251),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1267),
.B(n_1218),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1232),
.B(n_1230),
.Y(n_1327)
);

AOI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1208),
.A2(n_1266),
.B(n_1270),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1232),
.B(n_1206),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1270),
.B(n_1247),
.Y(n_1330)
);

INVx5_ASAP7_75t_L g1331 ( 
.A(n_1224),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1253),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1254),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1257),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1277),
.B(n_1257),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_1293),
.B(n_1208),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1295),
.B(n_1197),
.Y(n_1337)
);

BUFx8_ASAP7_75t_L g1338 ( 
.A(n_1299),
.Y(n_1338)
);

OR2x2_ASAP7_75t_L g1339 ( 
.A(n_1295),
.B(n_1215),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1325),
.B(n_1242),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1283),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1289),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1280),
.B(n_1243),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1281),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1291),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1280),
.B(n_1243),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1282),
.B(n_1243),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1281),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1284),
.A2(n_1244),
.B1(n_1217),
.B2(n_1192),
.Y(n_1349)
);

INVx3_ASAP7_75t_L g1350 ( 
.A(n_1304),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1282),
.B(n_1263),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1294),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_SL g1353 ( 
.A1(n_1314),
.A2(n_1324),
.B1(n_1326),
.B2(n_1319),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1306),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1300),
.B(n_1189),
.Y(n_1355)
);

BUFx2_ASAP7_75t_L g1356 ( 
.A(n_1294),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1306),
.Y(n_1357)
);

INVx1_ASAP7_75t_SL g1358 ( 
.A(n_1318),
.Y(n_1358)
);

OR2x6_ASAP7_75t_L g1359 ( 
.A(n_1287),
.B(n_1224),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1309),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1297),
.A2(n_1217),
.B1(n_1192),
.B2(n_1275),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1290),
.B(n_1262),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1309),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1335),
.B(n_1226),
.Y(n_1364)
);

BUFx6f_ASAP7_75t_L g1365 ( 
.A(n_1301),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1304),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1312),
.B(n_1275),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1332),
.Y(n_1368)
);

INVx2_ASAP7_75t_SL g1369 ( 
.A(n_1329),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1333),
.Y(n_1370)
);

AOI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1361),
.A2(n_1328),
.B(n_1313),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1368),
.B(n_1288),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1370),
.B(n_1292),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1342),
.B(n_1345),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1341),
.B(n_1286),
.Y(n_1375)
);

OAI22x1_ASAP7_75t_L g1376 ( 
.A1(n_1340),
.A2(n_1328),
.B1(n_1315),
.B2(n_1316),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1364),
.B(n_1307),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1364),
.B(n_1307),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1343),
.B(n_1346),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1344),
.B(n_1320),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1356),
.B(n_1321),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1343),
.B(n_1308),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1349),
.A2(n_1298),
.B1(n_1299),
.B2(n_1302),
.Y(n_1383)
);

OAI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1362),
.A2(n_1303),
.B(n_1327),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_SL g1385 ( 
.A1(n_1353),
.A2(n_1311),
.B(n_1203),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_SL g1386 ( 
.A1(n_1359),
.A2(n_1287),
.B(n_1367),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1348),
.B(n_1316),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_L g1388 ( 
.A(n_1337),
.B(n_1279),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1367),
.A2(n_1249),
.B1(n_1305),
.B2(n_1296),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1348),
.B(n_1317),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1336),
.A2(n_1296),
.B1(n_1248),
.B2(n_1311),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1352),
.B(n_1317),
.Y(n_1392)
);

OA211x2_ASAP7_75t_L g1393 ( 
.A1(n_1338),
.A2(n_1296),
.B(n_1265),
.C(n_1278),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1346),
.B(n_1308),
.Y(n_1394)
);

NOR3xp33_ASAP7_75t_SL g1395 ( 
.A(n_1338),
.B(n_1213),
.C(n_1190),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1354),
.Y(n_1396)
);

NAND3xp33_ASAP7_75t_L g1397 ( 
.A(n_1339),
.B(n_1334),
.C(n_1310),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_SL g1398 ( 
.A(n_1338),
.B(n_1194),
.Y(n_1398)
);

NAND3xp33_ASAP7_75t_L g1399 ( 
.A(n_1355),
.B(n_1334),
.C(n_1310),
.Y(n_1399)
);

NAND3xp33_ASAP7_75t_L g1400 ( 
.A(n_1355),
.B(n_1334),
.C(n_1330),
.Y(n_1400)
);

NAND2xp33_ASAP7_75t_L g1401 ( 
.A(n_1365),
.B(n_1350),
.Y(n_1401)
);

NAND3xp33_ASAP7_75t_L g1402 ( 
.A(n_1336),
.B(n_1322),
.C(n_1323),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1347),
.B(n_1285),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_L g1404 ( 
.A(n_1338),
.B(n_1194),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1396),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1396),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_SL g1407 ( 
.A(n_1384),
.B(n_1369),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1372),
.B(n_1354),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1373),
.Y(n_1409)
);

OR2x6_ASAP7_75t_L g1410 ( 
.A(n_1386),
.B(n_1359),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1380),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1379),
.B(n_1347),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1381),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1402),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1377),
.B(n_1351),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1377),
.B(n_1378),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1387),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1376),
.Y(n_1418)
);

INVx5_ASAP7_75t_L g1419 ( 
.A(n_1403),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1375),
.Y(n_1420)
);

BUFx2_ASAP7_75t_L g1421 ( 
.A(n_1382),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1390),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1392),
.B(n_1357),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1374),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1399),
.B(n_1366),
.Y(n_1425)
);

INVxp67_ASAP7_75t_SL g1426 ( 
.A(n_1376),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1382),
.B(n_1360),
.Y(n_1427)
);

BUFx2_ASAP7_75t_L g1428 ( 
.A(n_1394),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1399),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1371),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1403),
.B(n_1366),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1405),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1405),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1425),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1406),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1419),
.B(n_1371),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1425),
.Y(n_1437)
);

NAND2x1p5_ASAP7_75t_L g1438 ( 
.A(n_1425),
.B(n_1331),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1406),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1414),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1425),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1423),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1419),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1408),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1414),
.B(n_1400),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1429),
.B(n_1420),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1408),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1420),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1427),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1425),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1419),
.B(n_1401),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1430),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1419),
.B(n_1401),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1429),
.B(n_1360),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1430),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1419),
.B(n_1388),
.Y(n_1456)
);

INVx3_ASAP7_75t_SL g1457 ( 
.A(n_1410),
.Y(n_1457)
);

INVx3_ASAP7_75t_L g1458 ( 
.A(n_1419),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1411),
.B(n_1363),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1416),
.B(n_1421),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1427),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1411),
.B(n_1397),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1428),
.B(n_1363),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1409),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1460),
.B(n_1428),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1460),
.B(n_1415),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1432),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1440),
.B(n_1424),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1432),
.Y(n_1469)
);

NAND2x1_ASAP7_75t_L g1470 ( 
.A(n_1443),
.B(n_1431),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1440),
.B(n_1398),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1446),
.B(n_1445),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_1456),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1433),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1460),
.B(n_1415),
.Y(n_1475)
);

INVx2_ASAP7_75t_SL g1476 ( 
.A(n_1456),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1456),
.B(n_1415),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1446),
.B(n_1424),
.Y(n_1478)
);

INVx4_ASAP7_75t_L g1479 ( 
.A(n_1443),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_R g1480 ( 
.A(n_1436),
.B(n_1404),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1444),
.B(n_1417),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1444),
.B(n_1417),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1451),
.B(n_1412),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1452),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1451),
.B(n_1412),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1452),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1447),
.B(n_1422),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1447),
.B(n_1422),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1445),
.B(n_1413),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1433),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1435),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1435),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1439),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1445),
.B(n_1413),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1439),
.Y(n_1495)
);

INVxp67_ASAP7_75t_L g1496 ( 
.A(n_1454),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1452),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1452),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1459),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1453),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1459),
.Y(n_1501)
);

AOI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1457),
.A2(n_1426),
.B1(n_1385),
.B2(n_1418),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1466),
.B(n_1443),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1467),
.Y(n_1504)
);

INVx4_ASAP7_75t_L g1505 ( 
.A(n_1479),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1472),
.B(n_1463),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1502),
.A2(n_1438),
.B1(n_1462),
.B2(n_1407),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1471),
.A2(n_1438),
.B1(n_1462),
.B2(n_1426),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1465),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1472),
.B(n_1463),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1496),
.B(n_1463),
.Y(n_1511)
);

INVx2_ASAP7_75t_SL g1512 ( 
.A(n_1473),
.Y(n_1512)
);

BUFx3_ASAP7_75t_L g1513 ( 
.A(n_1465),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1468),
.B(n_1449),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1466),
.B(n_1443),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1467),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1484),
.A2(n_1418),
.B1(n_1430),
.B2(n_1457),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1469),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1484),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1486),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1489),
.B(n_1461),
.Y(n_1521)
);

INVx2_ASAP7_75t_SL g1522 ( 
.A(n_1473),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1475),
.B(n_1458),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1489),
.B(n_1461),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1469),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1494),
.B(n_1448),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1490),
.Y(n_1527)
);

INVx1_ASAP7_75t_SL g1528 ( 
.A(n_1494),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1490),
.Y(n_1529)
);

INVx1_ASAP7_75t_SL g1530 ( 
.A(n_1476),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1474),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1478),
.B(n_1454),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1475),
.B(n_1448),
.Y(n_1533)
);

AOI222xp33_ASAP7_75t_L g1534 ( 
.A1(n_1486),
.A2(n_1418),
.B1(n_1455),
.B2(n_1383),
.C1(n_1457),
.C2(n_1442),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1477),
.B(n_1458),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1491),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1477),
.B(n_1458),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1476),
.Y(n_1538)
);

AOI222xp33_ASAP7_75t_L g1539 ( 
.A1(n_1528),
.A2(n_1498),
.B1(n_1497),
.B2(n_1455),
.C1(n_1457),
.C2(n_1501),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1509),
.Y(n_1540)
);

INVx1_ASAP7_75t_SL g1541 ( 
.A(n_1509),
.Y(n_1541)
);

AOI221xp5_ASAP7_75t_SL g1542 ( 
.A1(n_1507),
.A2(n_1437),
.B1(n_1434),
.B2(n_1450),
.C(n_1441),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1513),
.B(n_1483),
.Y(n_1543)
);

INVxp67_ASAP7_75t_L g1544 ( 
.A(n_1513),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1530),
.B(n_1531),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1506),
.B(n_1481),
.Y(n_1546)
);

XOR2xp5_ASAP7_75t_L g1547 ( 
.A(n_1508),
.B(n_1393),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1510),
.A2(n_1438),
.B1(n_1462),
.B2(n_1500),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1537),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1512),
.A2(n_1438),
.B1(n_1500),
.B2(n_1434),
.Y(n_1550)
);

AOI222xp33_ASAP7_75t_L g1551 ( 
.A1(n_1517),
.A2(n_1498),
.B1(n_1497),
.B2(n_1455),
.C1(n_1499),
.C2(n_1501),
.Y(n_1551)
);

OAI21xp5_ASAP7_75t_SL g1552 ( 
.A1(n_1534),
.A2(n_1436),
.B(n_1458),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1504),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_L g1554 ( 
.A(n_1505),
.B(n_1479),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1512),
.B(n_1499),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1504),
.Y(n_1556)
);

OAI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1526),
.A2(n_1389),
.B1(n_1391),
.B2(n_1441),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1522),
.B(n_1464),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1505),
.B(n_1213),
.Y(n_1559)
);

NAND3xp33_ASAP7_75t_L g1560 ( 
.A(n_1522),
.B(n_1487),
.C(n_1482),
.Y(n_1560)
);

O2A1O1Ixp33_ASAP7_75t_L g1561 ( 
.A1(n_1538),
.A2(n_1455),
.B(n_1488),
.C(n_1493),
.Y(n_1561)
);

OAI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1521),
.A2(n_1437),
.B1(n_1434),
.B2(n_1441),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1516),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1538),
.B(n_1464),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1541),
.B(n_1524),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1544),
.B(n_1532),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1553),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1543),
.B(n_1503),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1544),
.B(n_1503),
.Y(n_1569)
);

AOI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1557),
.A2(n_1519),
.B1(n_1520),
.B2(n_1514),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1540),
.B(n_1515),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1549),
.B(n_1515),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1545),
.B(n_1532),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1556),
.Y(n_1574)
);

NOR2x1_ASAP7_75t_L g1575 ( 
.A(n_1559),
.B(n_1505),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1546),
.B(n_1533),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1555),
.B(n_1511),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1554),
.B(n_1523),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1554),
.B(n_1523),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1560),
.B(n_1516),
.Y(n_1580)
);

INVx1_ASAP7_75t_SL g1581 ( 
.A(n_1547),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1551),
.B(n_1518),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1563),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1558),
.Y(n_1584)
);

AOI21xp33_ASAP7_75t_L g1585 ( 
.A1(n_1582),
.A2(n_1539),
.B(n_1561),
.Y(n_1585)
);

XOR2x2_ASAP7_75t_L g1586 ( 
.A(n_1570),
.B(n_1542),
.Y(n_1586)
);

AOI211xp5_ASAP7_75t_L g1587 ( 
.A1(n_1580),
.A2(n_1557),
.B(n_1552),
.C(n_1562),
.Y(n_1587)
);

NOR3xp33_ASAP7_75t_L g1588 ( 
.A(n_1581),
.B(n_1566),
.C(n_1573),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1577),
.A2(n_1564),
.B(n_1562),
.Y(n_1589)
);

INVx1_ASAP7_75t_SL g1590 ( 
.A(n_1569),
.Y(n_1590)
);

NAND4xp75_ASAP7_75t_L g1591 ( 
.A(n_1575),
.B(n_1393),
.C(n_1520),
.D(n_1519),
.Y(n_1591)
);

AOI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1584),
.A2(n_1548),
.B1(n_1529),
.B2(n_1518),
.C(n_1536),
.Y(n_1592)
);

AOI211xp5_ASAP7_75t_L g1593 ( 
.A1(n_1565),
.A2(n_1571),
.B(n_1569),
.C(n_1572),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1568),
.B(n_1535),
.Y(n_1594)
);

NAND4xp25_ASAP7_75t_SL g1595 ( 
.A(n_1568),
.B(n_1436),
.C(n_1437),
.D(n_1434),
.Y(n_1595)
);

OAI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1565),
.A2(n_1450),
.B1(n_1441),
.B2(n_1437),
.Y(n_1596)
);

NAND2xp33_ASAP7_75t_SL g1597 ( 
.A(n_1594),
.B(n_1571),
.Y(n_1597)
);

NAND3xp33_ASAP7_75t_SL g1598 ( 
.A(n_1587),
.B(n_1579),
.C(n_1578),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1590),
.Y(n_1599)
);

NOR3xp33_ASAP7_75t_L g1600 ( 
.A(n_1588),
.B(n_1574),
.C(n_1567),
.Y(n_1600)
);

NAND4xp75_ASAP7_75t_L g1601 ( 
.A(n_1585),
.B(n_1572),
.C(n_1579),
.D(n_1578),
.Y(n_1601)
);

INVxp67_ASAP7_75t_L g1602 ( 
.A(n_1591),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1593),
.Y(n_1603)
);

OA22x2_ASAP7_75t_L g1604 ( 
.A1(n_1586),
.A2(n_1576),
.B1(n_1583),
.B2(n_1550),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1589),
.B(n_1525),
.Y(n_1605)
);

NOR3xp33_ASAP7_75t_L g1606 ( 
.A(n_1592),
.B(n_1527),
.C(n_1525),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1599),
.B(n_1596),
.Y(n_1607)
);

O2A1O1Ixp33_ASAP7_75t_L g1608 ( 
.A1(n_1598),
.A2(n_1527),
.B(n_1536),
.C(n_1529),
.Y(n_1608)
);

NOR3xp33_ASAP7_75t_SL g1609 ( 
.A(n_1601),
.B(n_1595),
.C(n_1480),
.Y(n_1609)
);

AOI221xp5_ASAP7_75t_L g1610 ( 
.A1(n_1605),
.A2(n_1495),
.B1(n_1491),
.B2(n_1493),
.C(n_1492),
.Y(n_1610)
);

NAND5xp2_ASAP7_75t_L g1611 ( 
.A(n_1603),
.B(n_1395),
.C(n_1480),
.D(n_1483),
.E(n_1485),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1607),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1608),
.B(n_1600),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1610),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1609),
.A2(n_1604),
.B1(n_1597),
.B2(n_1602),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1611),
.Y(n_1616)
);

AOI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1607),
.A2(n_1606),
.B1(n_1537),
.B2(n_1535),
.Y(n_1617)
);

BUFx2_ASAP7_75t_L g1618 ( 
.A(n_1617),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1612),
.B(n_1537),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1616),
.Y(n_1620)
);

NAND3x1_ASAP7_75t_L g1621 ( 
.A(n_1615),
.B(n_1458),
.C(n_1216),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1613),
.B(n_1535),
.Y(n_1622)
);

XOR2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1620),
.B(n_1614),
.Y(n_1623)
);

XOR2xp5_ASAP7_75t_L g1624 ( 
.A(n_1618),
.B(n_1216),
.Y(n_1624)
);

NOR2x1_ASAP7_75t_L g1625 ( 
.A(n_1619),
.B(n_1479),
.Y(n_1625)
);

INVxp67_ASAP7_75t_L g1626 ( 
.A(n_1624),
.Y(n_1626)
);

XOR2xp5_ASAP7_75t_L g1627 ( 
.A(n_1626),
.B(n_1622),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1627),
.B(n_1625),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1627),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1629),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1628),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1630),
.B(n_1628),
.Y(n_1632)
);

INVxp33_ASAP7_75t_SL g1633 ( 
.A(n_1631),
.Y(n_1633)
);

OAI222xp33_ASAP7_75t_L g1634 ( 
.A1(n_1632),
.A2(n_1623),
.B1(n_1621),
.B2(n_1537),
.C1(n_1495),
.C2(n_1492),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1634),
.A2(n_1633),
.B1(n_1225),
.B2(n_1234),
.Y(n_1635)
);

OAI221xp5_ASAP7_75t_R g1636 ( 
.A1(n_1635),
.A2(n_1260),
.B1(n_1225),
.B2(n_1470),
.C(n_1234),
.Y(n_1636)
);

AOI211xp5_ASAP7_75t_L g1637 ( 
.A1(n_1636),
.A2(n_1234),
.B(n_1260),
.C(n_1358),
.Y(n_1637)
);


endmodule