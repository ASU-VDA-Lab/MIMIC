module real_jpeg_6961_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_11;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_9;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_1),
.B(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_31),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_1),
.B(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_1),
.A2(n_27),
.B1(n_62),
.B2(n_66),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_1),
.B(n_74),
.C(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_1),
.B(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_1),
.B(n_106),
.C(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_1),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_139)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_1),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_3),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_5),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_6),
.A2(n_17),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_6),
.A2(n_36),
.B1(n_81),
.B2(n_84),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_6),
.A2(n_36),
.B1(n_153),
.B2(n_158),
.Y(n_152)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_7),
.Y(n_74)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_120),
.Y(n_8)
);

AOI21xp5_ASAP7_75t_L g9 ( 
.A1(n_10),
.A2(n_91),
.B(n_119),
.Y(n_9)
);

OAI21xp5_ASAP7_75t_L g10 ( 
.A1(n_11),
.A2(n_55),
.B(n_90),
.Y(n_10)
);

AOI21xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_40),
.B(n_54),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_23),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_21),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_16),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_22),
.A2(n_24),
.B1(n_26),
.B2(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_26),
.B1(n_32),
.B2(n_35),
.Y(n_23)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_24),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_26),
.B(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_33),
.B(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_42),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_41),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_41),
.B(n_96),
.C(n_112),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_43),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2x1_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_48),
.B2(n_52),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_57),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_85),
.B2(n_89),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_58),
.B(n_89),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_58),
.A2(n_59),
.B1(n_138),
.B2(n_161),
.Y(n_137)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_79),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_70),
.Y(n_60)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVx5_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_75),
.B2(n_77),
.Y(n_71)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_85),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_118),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_118),
.Y(n_119)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_111),
.B1(n_112),
.B2(n_117),
.Y(n_95)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g138 ( 
.A1(n_98),
.A2(n_139),
.B1(n_144),
.B2(n_152),
.Y(n_138)
);

NAND2x1_ASAP7_75t_L g144 ( 
.A(n_98),
.B(n_145),
.Y(n_144)
);

AOI22x1_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_102),
.B1(n_106),
.B2(n_108),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_105),
.Y(n_150)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_162),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_123),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_137),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_133),
.B2(n_136),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_133),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_138),
.Y(n_161)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_148),
.B1(n_149),
.B2(n_151),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);


endmodule