module fake_jpeg_16503_n_206 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_0),
.B(n_14),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_33),
.Y(n_42)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_30),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_1),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_37),
.B(n_25),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_27),
.Y(n_77)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_50),
.B(n_32),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_65),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_38),
.B(n_22),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_57),
.A2(n_64),
.B(n_29),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_55),
.A2(n_17),
.B1(n_19),
.B2(n_36),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_31),
.B1(n_54),
.B2(n_48),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_19),
.B1(n_23),
.B2(n_20),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_59),
.A2(n_75),
.B1(n_16),
.B2(n_20),
.Y(n_80)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_38),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_63),
.B(n_33),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_39),
.B(n_38),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_52),
.B(n_34),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_25),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_72),
.Y(n_83)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_40),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_33),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_41),
.A2(n_40),
.B1(n_32),
.B2(n_36),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_41),
.A2(n_18),
.B1(n_29),
.B2(n_27),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_21),
.B1(n_24),
.B2(n_15),
.Y(n_90)
);

NAND2xp33_ASAP7_75t_SL g81 ( 
.A(n_77),
.B(n_15),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_43),
.A2(n_36),
.B1(n_33),
.B2(n_35),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_51),
.B1(n_47),
.B2(n_33),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_79),
.A2(n_87),
.B1(n_78),
.B2(n_73),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_80),
.A2(n_90),
.B1(n_62),
.B2(n_10),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_88),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_96),
.Y(n_110)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_59),
.A2(n_31),
.B1(n_23),
.B2(n_16),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_64),
.A2(n_35),
.B(n_18),
.C(n_24),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_95),
.B1(n_100),
.B2(n_99),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_99),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_51),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_21),
.Y(n_98)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_61),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_61),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_101),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_51),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_57),
.C(n_47),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_114),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_106),
.B1(n_111),
.B2(n_115),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_109),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_96),
.A2(n_77),
.B1(n_70),
.B2(n_67),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_86),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_108),
.B(n_118),
.Y(n_140)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_78),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_77),
.B1(n_60),
.B2(n_73),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_47),
.C(n_78),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_83),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_SL g127 ( 
.A1(n_116),
.A2(n_95),
.B(n_90),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_62),
.Y(n_119)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_9),
.Y(n_120)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_4),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_121),
.A2(n_4),
.B(n_6),
.Y(n_128)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_122),
.A2(n_80),
.B1(n_82),
.B2(n_87),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_124),
.A2(n_138),
.B1(n_11),
.B2(n_12),
.Y(n_159)
);

OA21x2_ASAP7_75t_L g125 ( 
.A1(n_116),
.A2(n_89),
.B(n_95),
.Y(n_125)
);

OA21x2_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_127),
.B(n_116),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_116),
.C(n_8),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_117),
.A2(n_95),
.B(n_93),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_141),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_122),
.A2(n_93),
.B(n_91),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_91),
.B(n_7),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_9),
.Y(n_139)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_113),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_142),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_109),
.A2(n_8),
.B(n_11),
.Y(n_143)
);

INVxp33_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_110),
.C(n_102),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_149),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_106),
.C(n_121),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_111),
.C(n_115),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_150),
.B(n_149),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_137),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_153),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_154),
.A2(n_155),
.B(n_131),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_105),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_156),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_159),
.B(n_140),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_162),
.A2(n_168),
.B(n_144),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_164),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_148),
.B(n_130),
.Y(n_165)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_165),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_129),
.Y(n_166)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_158),
.B(n_138),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_167),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_155),
.A2(n_125),
.B(n_136),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_169),
.B(n_154),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_126),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_170),
.Y(n_177)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_144),
.B1(n_157),
.B2(n_154),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_145),
.C(n_132),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_176),
.C(n_160),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_174),
.A2(n_168),
.B1(n_157),
.B2(n_161),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_125),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_143),
.Y(n_189)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_181),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_186),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_188),
.C(n_176),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_178),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_173),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_169),
.B1(n_163),
.B2(n_151),
.Y(n_185)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_185),
.Y(n_195)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_175),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_189),
.B(n_174),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_192),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_172),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_193),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_194),
.A2(n_185),
.B(n_187),
.Y(n_196)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_196),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_193),
.A2(n_151),
.B(n_182),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_195),
.C(n_191),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_201),
.C(n_198),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_199),
.B(n_188),
.C(n_128),
.Y(n_201)
);

AOI21xp33_ASAP7_75t_SL g205 ( 
.A1(n_203),
.A2(n_204),
.B(n_13),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_180),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_13),
.Y(n_206)
);


endmodule