module real_aes_6144_n_104 (n_17, n_28, n_994, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_995, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_994;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_995;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_357;
wire n_635;
wire n_287;
wire n_503;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_987;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_974;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_260;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_983;
wire n_767;
wire n_138;
wire n_696;
wire n_955;
wire n_889;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_958;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_961;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_743;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_795;
wire n_116;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_106;
wire n_791;
wire n_981;
wire n_976;
wire n_559;
wire n_636;
wire n_466;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_984;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_962;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_960;
wire n_164;
wire n_671;
wire n_973;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_142;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_985;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_957;
wire n_296;
wire n_702;
wire n_954;
wire n_969;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_965;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_972;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_498;
wire n_691;
wire n_481;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_922;
wire n_926;
wire n_149;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_134;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_982;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_967;
wire n_473;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_968;
wire n_646;
wire n_650;
wire n_105;
wire n_710;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
wire n_862;
INVx1_ASAP7_75t_L g697 ( .A(n_0), .Y(n_697) );
INVx1_ASAP7_75t_L g252 ( .A(n_1), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g144 ( .A1(n_2), .A2(n_18), .B1(n_145), .B2(n_148), .Y(n_144) );
INVx2_ASAP7_75t_L g212 ( .A(n_3), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_4), .B(n_590), .Y(n_675) );
INVx1_ASAP7_75t_SL g277 ( .A(n_5), .Y(n_277) );
INVxp67_ASAP7_75t_L g125 ( .A(n_6), .Y(n_125) );
BUFx2_ASAP7_75t_L g578 ( .A(n_6), .Y(n_578) );
INVx1_ASAP7_75t_L g976 ( .A(n_6), .Y(n_976) );
NAND2xp5_ASAP7_75t_SL g676 ( .A(n_7), .B(n_259), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_8), .A2(n_42), .B1(n_589), .B2(n_665), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_9), .A2(n_48), .B1(n_187), .B2(n_606), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g724 ( .A1(n_10), .A2(n_68), .B1(n_632), .B2(n_719), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_11), .B(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_12), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g692 ( .A(n_13), .Y(n_692) );
OAI22xp5_ASAP7_75t_SL g116 ( .A1(n_14), .A2(n_69), .B1(n_117), .B2(n_118), .Y(n_116) );
INVxp33_ASAP7_75t_SL g118 ( .A(n_14), .Y(n_118) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_15), .A2(n_56), .B1(n_258), .B2(n_259), .Y(n_257) );
INVx1_ASAP7_75t_L g695 ( .A(n_16), .Y(n_695) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_17), .A2(n_72), .B(n_161), .Y(n_160) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_17), .A2(n_72), .B(n_161), .Y(n_167) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_19), .A2(n_70), .B1(n_632), .B2(n_719), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_20), .B(n_146), .Y(n_223) );
AOI22xp5_ASAP7_75t_L g202 ( .A1(n_21), .A2(n_83), .B1(n_203), .B2(n_205), .Y(n_202) );
INVx2_ASAP7_75t_L g194 ( .A(n_22), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g961 ( .A1(n_23), .A2(n_962), .B1(n_965), .B2(n_966), .Y(n_961) );
CKINVDCx5p33_ASAP7_75t_R g965 ( .A(n_23), .Y(n_965) );
INVx1_ASAP7_75t_L g689 ( .A(n_24), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g151 ( .A1(n_25), .A2(n_29), .B1(n_152), .B2(n_154), .Y(n_151) );
BUFx3_ASAP7_75t_L g113 ( .A(n_26), .Y(n_113) );
BUFx8_ASAP7_75t_SL g989 ( .A(n_26), .Y(n_989) );
O2A1O1Ixp5_ASAP7_75t_L g186 ( .A1(n_27), .A2(n_149), .B(n_187), .C(n_191), .Y(n_186) );
AOI22xp33_ASAP7_75t_L g207 ( .A1(n_28), .A2(n_64), .B1(n_188), .B2(n_208), .Y(n_207) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_30), .Y(n_300) );
AO22x1_ASAP7_75t_L g672 ( .A1(n_31), .A2(n_81), .B1(n_281), .B2(n_673), .Y(n_672) );
CKINVDCx5p33_ASAP7_75t_R g593 ( .A(n_32), .Y(n_593) );
AND2x2_ASAP7_75t_L g605 ( .A(n_33), .B(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_34), .B(n_281), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g972 ( .A(n_35), .Y(n_972) );
AOI22xp5_ASAP7_75t_L g265 ( .A1(n_36), .A2(n_84), .B1(n_266), .B2(n_269), .Y(n_265) );
INVx1_ASAP7_75t_L g130 ( .A(n_37), .Y(n_130) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_38), .A2(n_87), .B1(n_554), .B2(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g555 ( .A(n_38), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_38), .B(n_135), .Y(n_957) );
INVx1_ASAP7_75t_L g180 ( .A(n_39), .Y(n_180) );
AOI22x1_ASAP7_75t_L g630 ( .A1(n_40), .A2(n_101), .B1(n_631), .B2(n_632), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_41), .B(n_634), .Y(n_666) );
AND2x2_ASAP7_75t_L g109 ( .A(n_43), .B(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_44), .B(n_176), .Y(n_247) );
INVx2_ASAP7_75t_L g192 ( .A(n_45), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_46), .Y(n_301) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_47), .B(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g222 ( .A(n_49), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_50), .B(n_245), .Y(n_244) );
INVx1_ASAP7_75t_SL g280 ( .A(n_51), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_52), .B(n_154), .Y(n_649) );
INVx1_ASAP7_75t_L g295 ( .A(n_53), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_54), .B(n_182), .Y(n_596) );
INVx1_ASAP7_75t_L g161 ( .A(n_55), .Y(n_161) );
AND2x4_ASAP7_75t_L g163 ( .A(n_57), .B(n_164), .Y(n_163) );
AND2x4_ASAP7_75t_L g184 ( .A(n_57), .B(n_164), .Y(n_184) );
INVx1_ASAP7_75t_L g284 ( .A(n_58), .Y(n_284) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_59), .Y(n_150) );
INVx2_ASAP7_75t_L g721 ( .A(n_60), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_61), .A2(n_76), .B1(n_589), .B2(n_631), .Y(n_661) );
CKINVDCx14_ASAP7_75t_R g678 ( .A(n_62), .Y(n_678) );
AND2x2_ASAP7_75t_L g612 ( .A(n_63), .B(n_281), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_65), .B(n_228), .Y(n_227) );
AO22x1_ASAP7_75t_SL g960 ( .A1(n_66), .A2(n_961), .B1(n_967), .B2(n_968), .Y(n_960) );
INVx1_ASAP7_75t_L g967 ( .A(n_66), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_67), .B(n_245), .Y(n_650) );
INVx1_ASAP7_75t_L g117 ( .A(n_69), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_69), .B(n_239), .Y(n_643) );
NAND2x1p5_ASAP7_75t_L g616 ( .A(n_71), .B(n_602), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g962 ( .A1(n_73), .A2(n_88), .B1(n_963), .B2(n_964), .Y(n_962) );
INVx1_ASAP7_75t_L g963 ( .A(n_73), .Y(n_963) );
CKINVDCx14_ASAP7_75t_R g636 ( .A(n_74), .Y(n_636) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_75), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_77), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_78), .B(n_590), .Y(n_647) );
OR2x6_ASAP7_75t_L g127 ( .A(n_79), .B(n_128), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_80), .B(n_155), .Y(n_282) );
INVx1_ASAP7_75t_L g129 ( .A(n_82), .Y(n_129) );
INVx1_ASAP7_75t_L g110 ( .A(n_85), .Y(n_110) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_86), .Y(n_147) );
BUFx5_ASAP7_75t_L g153 ( .A(n_86), .Y(n_153) );
INVx1_ASAP7_75t_L g190 ( .A(n_86), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_87), .Y(n_554) );
INVx1_ASAP7_75t_L g964 ( .A(n_88), .Y(n_964) );
INVx2_ASAP7_75t_L g699 ( .A(n_89), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_90), .B(n_228), .Y(n_278) );
INVx2_ASAP7_75t_L g225 ( .A(n_91), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g552 ( .A(n_92), .Y(n_552) );
INVx1_ASAP7_75t_L g232 ( .A(n_93), .Y(n_232) );
NAND2xp33_ASAP7_75t_L g608 ( .A(n_94), .B(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g303 ( .A(n_95), .Y(n_303) );
INVx2_ASAP7_75t_SL g164 ( .A(n_96), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_97), .B(n_293), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_98), .B(n_615), .Y(n_646) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_99), .B(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_100), .B(n_239), .Y(n_238) );
AO32x2_ASAP7_75t_L g142 ( .A1(n_102), .A2(n_143), .A3(n_158), .B1(n_162), .B2(n_165), .Y(n_142) );
AO22x2_ASAP7_75t_L g308 ( .A1(n_102), .A2(n_143), .B1(n_309), .B2(n_311), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_103), .B(n_600), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_114), .B1(n_563), .B2(n_570), .C(n_984), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
BUFx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
OR2x2_ASAP7_75t_SL g107 ( .A(n_108), .B(n_111), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_108), .B(n_569), .Y(n_568) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
OA21x2_ASAP7_75t_L g987 ( .A1(n_109), .A2(n_988), .B(n_990), .Y(n_987) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
CKINVDCx6p67_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_113), .Y(n_569) );
OAI21xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_131), .B(n_557), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_119), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_116), .B(n_120), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g984 ( .A(n_117), .B(n_985), .Y(n_984) );
INVxp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_R g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx10_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
BUFx8_ASAP7_75t_SL g562 ( .A(n_123), .Y(n_562) );
INVx2_ASAP7_75t_SL g566 ( .A(n_123), .Y(n_566) );
BUFx6f_ASAP7_75t_L g992 ( .A(n_123), .Y(n_992) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
INVx8_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OR2x6_ASAP7_75t_L g975 ( .A(n_127), .B(n_976), .Y(n_975) );
OAI32xp33_ASAP7_75t_L g977 ( .A1(n_127), .A2(n_959), .A3(n_971), .B1(n_978), .B2(n_995), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AOI21xp5_ASAP7_75t_SL g557 ( .A1(n_133), .A2(n_558), .B(n_559), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_135), .B1(n_549), .B2(n_550), .Y(n_133) );
INVxp67_ASAP7_75t_SL g134 ( .A(n_135), .Y(n_134) );
OR2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_454), .Y(n_135) );
INVxp33_ASAP7_75t_L g956 ( .A(n_136), .Y(n_956) );
NAND4xp25_ASAP7_75t_L g136 ( .A(n_137), .B(n_350), .C(n_397), .D(n_429), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g137 ( .A(n_138), .B(n_334), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_304), .Y(n_138) );
OAI21xp33_ASAP7_75t_SL g139 ( .A1(n_140), .A2(n_213), .B(n_235), .Y(n_139) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_168), .Y(n_140) );
INVx1_ASAP7_75t_L g349 ( .A(n_141), .Y(n_349) );
AND2x2_ASAP7_75t_SL g354 ( .A(n_141), .B(n_217), .Y(n_354) );
AND2x2_ASAP7_75t_L g433 ( .A(n_141), .B(n_327), .Y(n_433) );
OR2x2_ASAP7_75t_L g457 ( .A(n_141), .B(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g475 ( .A(n_141), .B(n_357), .Y(n_475) );
AND2x2_ASAP7_75t_L g497 ( .A(n_141), .B(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g513 ( .A(n_141), .Y(n_513) );
BUFx8_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g381 ( .A(n_142), .Y(n_381) );
AND2x2_ASAP7_75t_L g529 ( .A(n_142), .B(n_380), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_149), .B1(n_151), .B2(n_156), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_145), .B(n_192), .Y(n_191) );
INVx2_ASAP7_75t_SL g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g174 ( .A(n_146), .Y(n_174) );
INVx1_ASAP7_75t_L g208 ( .A(n_146), .Y(n_208) );
INVx2_ASAP7_75t_L g253 ( .A(n_146), .Y(n_253) );
INVx1_ASAP7_75t_L g609 ( .A(n_146), .Y(n_609) );
INVx1_ASAP7_75t_L g615 ( .A(n_146), .Y(n_615) );
INVx6_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g148 ( .A(n_147), .Y(n_148) );
INVx3_ASAP7_75t_L g155 ( .A(n_147), .Y(n_155) );
INVx2_ASAP7_75t_L g268 ( .A(n_147), .Y(n_268) );
INVx2_ASAP7_75t_L g182 ( .A(n_148), .Y(n_182) );
INVxp67_ASAP7_75t_SL g269 ( .A(n_148), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_149), .A2(n_242), .B(n_244), .Y(n_241) );
INVx4_ASAP7_75t_L g298 ( .A(n_149), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_149), .A2(n_589), .B1(n_591), .B2(n_594), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_149), .A2(n_646), .B(n_647), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_149), .B(n_660), .Y(n_659) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_150), .Y(n_157) );
INVx4_ASAP7_75t_L g177 ( .A(n_150), .Y(n_177) );
INVx3_ASAP7_75t_L g210 ( .A(n_150), .Y(n_210) );
INVx1_ASAP7_75t_L g271 ( .A(n_150), .Y(n_271) );
INVxp67_ASAP7_75t_L g610 ( .A(n_150), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_150), .B(n_689), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_150), .B(n_692), .Y(n_691) );
OAI22xp33_ASAP7_75t_L g299 ( .A1(n_152), .A2(n_253), .B1(n_300), .B2(n_301), .Y(n_299) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g245 ( .A(n_153), .Y(n_245) );
INVx1_ASAP7_75t_L g249 ( .A(n_153), .Y(n_249) );
INVx2_ASAP7_75t_L g258 ( .A(n_153), .Y(n_258) );
INVx2_ASAP7_75t_L g281 ( .A(n_153), .Y(n_281) );
INVx2_ASAP7_75t_L g590 ( .A(n_153), .Y(n_590) );
INVx1_ASAP7_75t_L g276 ( .A(n_154), .Y(n_276) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g205 ( .A(n_155), .Y(n_205) );
INVx1_ASAP7_75t_L g243 ( .A(n_155), .Y(n_243) );
INVx1_ASAP7_75t_L g259 ( .A(n_155), .Y(n_259) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g206 ( .A(n_157), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_157), .A2(n_225), .B(n_226), .C(n_227), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_157), .B(n_261), .Y(n_260) );
A2O1A1Ixp33_ASAP7_75t_L g275 ( .A1(n_157), .A2(n_276), .B(n_277), .C(n_278), .Y(n_275) );
INVxp67_ASAP7_75t_L g598 ( .A(n_157), .Y(n_598) );
INVx2_ASAP7_75t_SL g618 ( .A(n_157), .Y(n_618) );
INVx1_ASAP7_75t_L g651 ( .A(n_157), .Y(n_651) );
AO31x2_ASAP7_75t_L g170 ( .A1(n_158), .A2(n_171), .A3(n_185), .B(n_193), .Y(n_170) );
INVx2_ASAP7_75t_L g311 ( .A(n_158), .Y(n_311) );
BUFx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_159), .B(n_194), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_159), .B(n_212), .Y(n_211) );
INVx3_ASAP7_75t_L g239 ( .A(n_159), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_159), .B(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx4_ASAP7_75t_L g200 ( .A(n_160), .Y(n_200) );
BUFx3_ASAP7_75t_L g322 ( .A(n_160), .Y(n_322) );
OAI21x1_ASAP7_75t_L g587 ( .A1(n_162), .A2(n_588), .B(n_595), .Y(n_587) );
AO31x2_ASAP7_75t_L g626 ( .A1(n_162), .A2(n_627), .A3(n_633), .B(n_635), .Y(n_626) );
AO31x2_ASAP7_75t_L g712 ( .A1(n_162), .A2(n_627), .A3(n_633), .B(n_635), .Y(n_712) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g197 ( .A(n_163), .B(n_198), .Y(n_197) );
INVx3_ASAP7_75t_L g230 ( .A(n_163), .Y(n_230) );
AND2x2_ASAP7_75t_L g309 ( .A(n_163), .B(n_310), .Y(n_309) );
INVx3_ASAP7_75t_L g621 ( .A(n_163), .Y(n_621) );
INVx1_ASAP7_75t_L g670 ( .A(n_163), .Y(n_670) );
INVxp67_ASAP7_75t_L g286 ( .A(n_165), .Y(n_286) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_166), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_167), .B(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g233 ( .A(n_167), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_167), .B(n_230), .Y(n_254) );
NOR2xp67_ASAP7_75t_L g261 ( .A(n_167), .B(n_230), .Y(n_261) );
BUFx3_ASAP7_75t_L g263 ( .A(n_167), .Y(n_263) );
INVx1_ASAP7_75t_L g310 ( .A(n_167), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_167), .B(n_230), .Y(n_660) );
INVx2_ASAP7_75t_L g685 ( .A(n_167), .Y(n_685) );
AND2x2_ASAP7_75t_L g437 ( .A(n_168), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g518 ( .A(n_168), .B(n_374), .Y(n_518) );
INVxp67_ASAP7_75t_SL g534 ( .A(n_168), .Y(n_534) );
AND2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_195), .Y(n_168) );
INVx1_ASAP7_75t_L g394 ( .A(n_169), .Y(n_394) );
INVx2_ASAP7_75t_SL g491 ( .A(n_169), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_169), .B(n_381), .Y(n_504) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g234 ( .A(n_170), .Y(n_234) );
OR2x2_ASAP7_75t_L g314 ( .A(n_170), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g327 ( .A(n_170), .B(n_218), .Y(n_327) );
AND2x2_ASAP7_75t_L g357 ( .A(n_170), .B(n_312), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_170), .B(n_315), .Y(n_410) );
AOI221x1_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_175), .B1(n_179), .B2(n_181), .C(n_183), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_178), .Y(n_175) );
AND2x2_ASAP7_75t_L g179 ( .A(n_176), .B(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_177), .B(n_252), .Y(n_251) );
NOR2xp33_ASAP7_75t_SL g694 ( .A(n_177), .B(n_695), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_177), .B(n_697), .Y(n_696) );
NAND3xp33_ASAP7_75t_SL g717 ( .A(n_177), .B(n_620), .C(n_685), .Y(n_717) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_182), .B(n_691), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_182), .A2(n_281), .B1(n_694), .B2(n_696), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_183), .B(n_209), .Y(n_291) );
NOR3xp33_ASAP7_75t_L g294 ( .A(n_183), .B(n_209), .C(n_295), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_183), .B(n_298), .Y(n_297) );
INVx4_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g228 ( .A(n_189), .Y(n_228) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g204 ( .A(n_190), .Y(n_204) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_195), .Y(n_340) );
INVx2_ASAP7_75t_L g373 ( .A(n_195), .Y(n_373) );
AND2x2_ASAP7_75t_L g540 ( .A(n_195), .B(n_312), .Y(n_540) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g216 ( .A(n_196), .Y(n_216) );
INVx1_ASAP7_75t_L g315 ( .A(n_196), .Y(n_315) );
AOI21x1_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_201), .B(n_211), .Y(n_196) );
AOI21xp33_ASAP7_75t_SL g619 ( .A1(n_198), .A2(n_620), .B(n_622), .Y(n_619) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_199), .B(n_230), .Y(n_274) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx3_ASAP7_75t_L g602 ( .A(n_200), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_206), .B1(n_207), .B2(n_209), .Y(n_201) );
INVx2_ASAP7_75t_L g673 ( .A(n_203), .Y(n_673) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx2_ASAP7_75t_L g226 ( .A(n_204), .Y(n_226) );
INVx1_ASAP7_75t_L g665 ( .A(n_205), .Y(n_665) );
INVx1_ASAP7_75t_L g719 ( .A(n_205), .Y(n_719) );
AOI21x1_ASAP7_75t_L g671 ( .A1(n_206), .A2(n_672), .B(n_674), .Y(n_671) );
INVx1_ASAP7_75t_L g221 ( .A(n_208), .Y(n_221) );
NAND3xp33_ASAP7_75t_L g723 ( .A(n_209), .B(n_620), .C(n_685), .Y(n_723) );
INVx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_210), .A2(n_221), .B(n_222), .C(n_223), .Y(n_220) );
A2O1A1Ixp33_ASAP7_75t_L g279 ( .A1(n_210), .A2(n_280), .B(n_281), .C(n_282), .Y(n_279) );
INVx2_ASAP7_75t_L g462 ( .A(n_213), .Y(n_462) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_217), .Y(n_213) );
NAND2x1p5_ASAP7_75t_L g326 ( .A(n_214), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_214), .B(n_307), .Y(n_412) );
INVx4_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
HB1xp67_ASAP7_75t_SL g352 ( .A(n_215), .Y(n_352) );
AND2x2_ASAP7_75t_L g471 ( .A(n_215), .B(n_357), .Y(n_471) );
AND2x2_ASAP7_75t_L g484 ( .A(n_215), .B(n_217), .Y(n_484) );
INVx2_ASAP7_75t_L g487 ( .A(n_215), .Y(n_487) );
BUFx3_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g380 ( .A(n_216), .Y(n_380) );
INVx2_ASAP7_75t_L g458 ( .A(n_217), .Y(n_458) );
AND2x4_ASAP7_75t_L g217 ( .A(n_218), .B(n_234), .Y(n_217) );
INVx2_ASAP7_75t_L g312 ( .A(n_218), .Y(n_312) );
INVx1_ASAP7_75t_L g375 ( .A(n_218), .Y(n_375) );
BUFx3_ASAP7_75t_L g393 ( .A(n_218), .Y(n_393) );
AND2x4_ASAP7_75t_L g438 ( .A(n_218), .B(n_381), .Y(n_438) );
INVx3_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AO31x2_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_224), .A3(n_229), .B(n_231), .Y(n_219) );
NOR2xp67_ASAP7_75t_L g289 ( .A(n_226), .B(n_290), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_232), .B(n_233), .Y(n_231) );
NOR2xp33_ASAP7_75t_SL g283 ( .A(n_233), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g634 ( .A(n_233), .Y(n_634) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_272), .Y(n_235) );
AND2x2_ASAP7_75t_L g500 ( .A(n_236), .B(n_332), .Y(n_500) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_255), .Y(n_236) );
INVx2_ASAP7_75t_L g324 ( .A(n_237), .Y(n_324) );
INVx1_ASAP7_75t_L g347 ( .A(n_237), .Y(n_347) );
AND2x2_ASAP7_75t_L g363 ( .A(n_237), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g426 ( .A(n_237), .Y(n_426) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_237), .Y(n_537) );
AND2x4_ASAP7_75t_L g237 ( .A(n_238), .B(n_240), .Y(n_237) );
NOR2x1_ASAP7_75t_L g652 ( .A(n_239), .B(n_621), .Y(n_652) );
OAI21xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_246), .B(n_254), .Y(n_240) );
OAI21xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_248), .B(n_250), .Y(n_246) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_253), .Y(n_250) );
INVx2_ASAP7_75t_L g606 ( .A(n_253), .Y(n_606) );
AND2x2_ASAP7_75t_L g323 ( .A(n_255), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g343 ( .A(n_255), .Y(n_343) );
INVx2_ASAP7_75t_L g361 ( .A(n_255), .Y(n_361) );
INVx1_ASAP7_75t_L g385 ( .A(n_255), .Y(n_385) );
NAND2x1p5_ASAP7_75t_L g255 ( .A(n_256), .B(n_264), .Y(n_255) );
AND2x2_ASAP7_75t_SL g331 ( .A(n_256), .B(n_264), .Y(n_331) );
OA21x2_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_260), .B(n_262), .Y(n_256) );
INVx2_ASAP7_75t_L g632 ( .A(n_258), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_261), .B(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_270), .Y(n_264) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g293 ( .A(n_268), .Y(n_293) );
INVx1_ASAP7_75t_L g629 ( .A(n_271), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_271), .B(n_660), .Y(n_663) );
INVx1_ASAP7_75t_L g411 ( .A(n_272), .Y(n_411) );
AND2x2_ASAP7_75t_L g460 ( .A(n_272), .B(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g548 ( .A(n_272), .B(n_323), .Y(n_548) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_285), .Y(n_272) );
OR2x2_ASAP7_75t_L g319 ( .A(n_273), .B(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g333 ( .A(n_273), .Y(n_333) );
INVx2_ASAP7_75t_L g364 ( .A(n_273), .Y(n_364) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_273), .Y(n_390) );
INVx1_ASAP7_75t_L g424 ( .A(n_273), .Y(n_424) );
INVx1_ASAP7_75t_L g470 ( .A(n_273), .Y(n_470) );
AO31x2_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_275), .A3(n_279), .B(n_283), .Y(n_273) );
OR2x2_ASAP7_75t_L g369 ( .A(n_285), .B(n_324), .Y(n_369) );
AND2x2_ASAP7_75t_L g425 ( .A(n_285), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g493 ( .A(n_285), .B(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g516 ( .A(n_285), .B(n_361), .Y(n_516) );
AO21x2_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_287), .B(n_302), .Y(n_285) );
AO21x2_ASAP7_75t_L g320 ( .A1(n_287), .A2(n_302), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_296), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_291), .B1(n_292), .B2(n_294), .Y(n_288) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_298), .B(n_592), .Y(n_591) );
OAI22x1_ASAP7_75t_L g627 ( .A1(n_298), .A2(n_628), .B1(n_629), .B2(n_630), .Y(n_627) );
AOI22xp33_ASAP7_75t_SL g304 ( .A1(n_305), .A2(n_316), .B1(n_325), .B2(n_328), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_306), .B(n_313), .Y(n_305) );
OAI221xp5_ASAP7_75t_L g510 ( .A1(n_306), .A2(n_446), .B1(n_511), .B2(n_514), .C(n_517), .Y(n_510) );
INVx4_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x4_ASAP7_75t_L g452 ( .A(n_307), .B(n_453), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_307), .B(n_534), .Y(n_533) );
AND2x4_ASAP7_75t_L g307 ( .A(n_308), .B(n_312), .Y(n_307) );
INVx1_ASAP7_75t_L g337 ( .A(n_308), .Y(n_337) );
INVx1_ASAP7_75t_L g376 ( .A(n_308), .Y(n_376) );
AND2x4_ASAP7_75t_L g404 ( .A(n_308), .B(n_393), .Y(n_404) );
AND2x2_ASAP7_75t_L g428 ( .A(n_313), .B(n_392), .Y(n_428) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g453 ( .A(n_314), .Y(n_453) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_315), .Y(n_405) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp67_ASAP7_75t_L g317 ( .A(n_318), .B(n_323), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g419 ( .A(n_319), .B(n_384), .Y(n_419) );
AND2x2_ASAP7_75t_L g332 ( .A(n_320), .B(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g362 ( .A(n_320), .Y(n_362) );
BUFx2_ASAP7_75t_L g396 ( .A(n_320), .Y(n_396) );
NOR2xp67_ASAP7_75t_SL g635 ( .A(n_321), .B(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g677 ( .A(n_321), .B(n_678), .Y(n_677) );
INVx3_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OA21x2_ASAP7_75t_L g586 ( .A1(n_322), .A2(n_587), .B(n_599), .Y(n_586) );
OA21x2_ASAP7_75t_L g710 ( .A1(n_322), .A2(n_587), .B(n_599), .Y(n_710) );
AND2x2_ASAP7_75t_L g440 ( .A(n_323), .B(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_323), .B(n_396), .Y(n_450) );
AND2x2_ASAP7_75t_L g501 ( .A(n_323), .B(n_395), .Y(n_501) );
AND2x2_ASAP7_75t_L g524 ( .A(n_323), .B(n_414), .Y(n_524) );
INVx3_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g336 ( .A(n_327), .B(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g378 ( .A(n_327), .Y(n_378) );
INVx2_ASAP7_75t_L g444 ( .A(n_327), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_328), .A2(n_518), .B1(n_519), .B2(n_520), .Y(n_517) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2x1p5_ASAP7_75t_L g329 ( .A(n_330), .B(n_332), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_330), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g469 ( .A(n_331), .B(n_347), .Y(n_469) );
INVx2_ASAP7_75t_L g494 ( .A(n_331), .Y(n_494) );
AND2x2_ASAP7_75t_L g527 ( .A(n_331), .B(n_347), .Y(n_527) );
AND2x4_ASAP7_75t_L g339 ( .A(n_332), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g466 ( .A(n_332), .Y(n_466) );
INVxp67_ASAP7_75t_SL g368 ( .A(n_333), .Y(n_368) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_333), .Y(n_473) );
OAI32xp33_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_338), .A3(n_341), .B1(n_344), .B2(n_348), .Y(n_334) );
OAI22xp33_ASAP7_75t_L g543 ( .A1(n_335), .A2(n_544), .B1(n_545), .B2(n_547), .Y(n_543) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_339), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g443 ( .A(n_340), .Y(n_443) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI311xp33_ASAP7_75t_L g429 ( .A1(n_342), .A2(n_430), .A3(n_431), .B(n_434), .C(n_445), .Y(n_429) );
BUFx3_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g422 ( .A(n_343), .B(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND5xp2_ASAP7_75t_L g388 ( .A(n_346), .B(n_389), .C(n_391), .D(n_394), .E(n_395), .Y(n_388) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NOR3xp33_ASAP7_75t_L g350 ( .A(n_351), .B(n_365), .C(n_387), .Y(n_350) );
AOI31xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_353), .A3(n_355), .B(n_358), .Y(n_351) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g512 ( .A(n_357), .B(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g528 ( .A(n_357), .B(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g546 ( .A(n_357), .B(n_373), .Y(n_546) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_363), .Y(n_359) );
AND2x4_ASAP7_75t_L g535 ( .A(n_360), .B(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_361), .Y(n_448) );
BUFx2_ASAP7_75t_L g461 ( .A(n_361), .Y(n_461) );
AND2x4_ASAP7_75t_L g414 ( .A(n_362), .B(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g474 ( .A(n_362), .B(n_426), .Y(n_474) );
AND2x2_ASAP7_75t_L g515 ( .A(n_363), .B(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g521 ( .A(n_363), .B(n_385), .Y(n_521) );
INVx1_ASAP7_75t_L g415 ( .A(n_364), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_370), .B1(n_377), .B2(n_382), .Y(n_365) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g401 ( .A(n_367), .Y(n_401) );
OAI322xp33_ASAP7_75t_L g406 ( .A1(n_367), .A2(n_407), .A3(n_408), .B1(n_411), .B2(n_412), .C1(n_413), .C2(n_416), .Y(n_406) );
OR2x6_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVxp67_ASAP7_75t_L g386 ( .A(n_369), .Y(n_386) );
INVxp67_ASAP7_75t_SL g449 ( .A(n_369), .Y(n_449) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx3_ASAP7_75t_L g432 ( .A(n_373), .Y(n_432) );
AND2x2_ASAP7_75t_L g519 ( .A(n_373), .B(n_392), .Y(n_519) );
INVx1_ASAP7_75t_L g407 ( .A(n_374), .Y(n_407) );
AND2x4_ASAP7_75t_SL g374 ( .A(n_375), .B(n_376), .Y(n_374) );
OR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx1_ASAP7_75t_L g417 ( .A(n_379), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
AND2x2_ASAP7_75t_L g490 ( .A(n_381), .B(n_491), .Y(n_490) );
INVx3_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_384), .B(n_386), .Y(n_383) );
AND2x2_ASAP7_75t_L g389 ( .A(n_384), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g400 ( .A(n_384), .Y(n_400) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVxp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_392), .B(n_487), .Y(n_486) );
INVx2_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AOI211xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_402), .B(n_406), .C(n_418), .Y(n_397) );
AND2x4_ASAP7_75t_L g398 ( .A(n_399), .B(n_401), .Y(n_398) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
OR2x2_ASAP7_75t_L g531 ( .A(n_405), .B(n_504), .Y(n_531) );
OAI211xp5_ASAP7_75t_L g522 ( .A1(n_407), .A2(n_523), .B(n_525), .C(n_532), .Y(n_522) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g498 ( .A(n_410), .Y(n_498) );
INVx1_ASAP7_75t_L g430 ( .A(n_414), .Y(n_430) );
AND2x2_ASAP7_75t_L g480 ( .A(n_414), .B(n_461), .Y(n_480) );
AND2x4_ASAP7_75t_L g507 ( .A(n_414), .B(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g526 ( .A(n_414), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AOI21xp33_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_420), .B(n_427), .Y(n_418) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g421 ( .A(n_422), .B(n_425), .Y(n_421) );
INVxp67_ASAP7_75t_L g441 ( .A(n_423), .Y(n_441) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_423), .Y(n_483) );
AND2x2_ASAP7_75t_L g542 ( .A(n_423), .B(n_537), .Y(n_542) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g435 ( .A(n_425), .Y(n_435) );
AND2x2_ASAP7_75t_L g478 ( .A(n_426), .B(n_470), .Y(n_478) );
INVx1_ASAP7_75t_L g508 ( .A(n_426), .Y(n_508) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_436), .B1(n_439), .B2(n_442), .Y(n_434) );
INVx2_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OR2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_450), .B(n_451), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AND2x4_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
INVx1_ASAP7_75t_L g506 ( .A(n_448), .Y(n_506) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVxp33_ASAP7_75t_L g955 ( .A(n_454), .Y(n_955) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_509), .Y(n_454) );
NOR3xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_476), .C(n_495), .Y(n_455) );
OAI221xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_459), .B1(n_462), .B2(n_463), .C(n_467), .Y(n_456) );
OAI211xp5_ASAP7_75t_L g476 ( .A1(n_457), .A2(n_477), .B(n_479), .C(n_485), .Y(n_476) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g465 ( .A(n_461), .Y(n_465) );
INVxp67_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
NOR2x1p5_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_471), .B1(n_472), .B2(n_475), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_469), .B(n_483), .Y(n_482) );
NOR2xp67_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x4_ASAP7_75t_L g492 ( .A(n_478), .B(n_493), .Y(n_492) );
OAI21xp33_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B(n_484), .Y(n_479) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OAI21xp33_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_488), .B(n_492), .Y(n_485) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_489), .B(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
OAI22xp33_ASAP7_75t_SL g495 ( .A1(n_496), .A2(n_499), .B1(n_502), .B2(n_505), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_501), .A2(n_526), .B1(n_528), .B2(n_530), .Y(n_525) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVxp67_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
NOR3xp33_ASAP7_75t_L g509 ( .A(n_510), .B(n_522), .C(n_543), .Y(n_509) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x4_ASAP7_75t_L g541 ( .A(n_516), .B(n_542), .Y(n_541) );
BUFx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g544 ( .A(n_526), .Y(n_544) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_535), .B1(n_538), .B2(n_541), .Y(n_532) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_552), .B1(n_553), .B2(n_556), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g556 ( .A(n_553), .Y(n_556) );
AOI31xp33_ASAP7_75t_L g954 ( .A1(n_555), .A2(n_578), .A3(n_955), .B(n_956), .Y(n_954) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
CKINVDCx5p33_ASAP7_75t_R g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
BUFx3_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_980), .Y(n_571) );
AOI21xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_958), .B(n_977), .Y(n_572) );
INVx1_ASAP7_75t_L g983 ( .A(n_573), .Y(n_983) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x4_ASAP7_75t_L g574 ( .A(n_575), .B(n_953), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_579), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
BUFx8_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_848), .Y(n_579) );
NAND4xp25_ASAP7_75t_SL g580 ( .A(n_581), .B(n_739), .C(n_785), .D(n_817), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_680), .B(n_700), .Y(n_581) );
OAI21xp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_637), .B(n_653), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_583), .A2(n_797), .B1(n_801), .B2(n_803), .Y(n_796) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_623), .Y(n_584) );
INVx2_ASAP7_75t_L g729 ( .A(n_585), .Y(n_729) );
AND2x2_ASAP7_75t_L g846 ( .A(n_585), .B(n_847), .Y(n_846) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_603), .Y(n_585) );
AND2x2_ASAP7_75t_L g763 ( .A(n_586), .B(n_657), .Y(n_763) );
AND2x2_ASAP7_75t_L g813 ( .A(n_586), .B(n_783), .Y(n_813) );
NAND2x1_ASAP7_75t_L g840 ( .A(n_586), .B(n_625), .Y(n_840) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AOI21xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_597), .B(n_598), .Y(n_595) );
OR2x2_ASAP7_75t_L g669 ( .A(n_600), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g720 ( .A(n_601), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g765 ( .A(n_603), .B(n_712), .Y(n_765) );
AND2x2_ASAP7_75t_L g788 ( .A(n_603), .B(n_712), .Y(n_788) );
AND2x4_ASAP7_75t_L g834 ( .A(n_603), .B(n_709), .Y(n_834) );
AO21x2_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_611), .B(n_619), .Y(n_603) );
AO21x2_ASAP7_75t_L g706 ( .A1(n_604), .A2(n_611), .B(n_619), .Y(n_706) );
OAI21x1_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_607), .B(n_610), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_606), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g631 ( .A(n_609), .Y(n_631) );
OAI21x1_ASAP7_75t_SL g611 ( .A1(n_612), .A2(n_613), .B(n_617), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_616), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g622 ( .A(n_616), .Y(n_622) );
AOI21x1_ASAP7_75t_L g674 ( .A1(n_618), .A2(n_675), .B(n_676), .Y(n_674) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g727 ( .A(n_623), .Y(n_727) );
AND2x2_ASAP7_75t_L g908 ( .A(n_623), .B(n_834), .Y(n_908) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g679 ( .A(n_624), .Y(n_679) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g835 ( .A(n_625), .B(n_824), .Y(n_835) );
INVx1_ASAP7_75t_L g903 ( .A(n_625), .Y(n_903) );
AND2x2_ASAP7_75t_L g950 ( .A(n_625), .B(n_706), .Y(n_950) );
INVx3_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g889 ( .A(n_626), .B(n_756), .Y(n_889) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g859 ( .A(n_640), .B(n_747), .Y(n_859) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g777 ( .A(n_641), .B(n_668), .Y(n_777) );
AND2x2_ASAP7_75t_L g809 ( .A(n_641), .B(n_715), .Y(n_809) );
INVx3_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g667 ( .A(n_642), .B(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g737 ( .A(n_642), .B(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g792 ( .A(n_642), .Y(n_792) );
AND2x4_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
OAI21x1_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_648), .B(n_652), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_650), .B(n_651), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_654), .B(n_679), .Y(n_653) );
INVx1_ASAP7_75t_L g906 ( .A(n_654), .Y(n_906) );
AND2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_667), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g787 ( .A(n_656), .Y(n_787) );
INVx1_ASAP7_75t_L g830 ( .A(n_656), .Y(n_830) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g731 ( .A(n_657), .Y(n_731) );
AND2x2_ASAP7_75t_L g755 ( .A(n_657), .B(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_657), .B(n_705), .Y(n_802) );
INVx2_ASAP7_75t_L g824 ( .A(n_657), .Y(n_824) );
NAND2x1p5_ASAP7_75t_L g657 ( .A(n_658), .B(n_662), .Y(n_657) );
AND2x2_ASAP7_75t_L g783 ( .A(n_658), .B(n_662), .Y(n_783) );
OR2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_661), .Y(n_658) );
OA21x2_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_664), .B(n_666), .Y(n_662) );
AND2x2_ASAP7_75t_L g713 ( .A(n_667), .B(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g749 ( .A(n_667), .Y(n_749) );
AND2x2_ASAP7_75t_L g759 ( .A(n_667), .B(n_760), .Y(n_759) );
INVx2_ASAP7_75t_SL g738 ( .A(n_668), .Y(n_738) );
OAI21x1_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_671), .B(n_677), .Y(n_668) );
OAI21xp5_ASAP7_75t_L g770 ( .A1(n_669), .A2(n_671), .B(n_677), .Y(n_770) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_670), .B(n_684), .Y(n_683) );
OR2x2_ASAP7_75t_L g753 ( .A(n_679), .B(n_754), .Y(n_753) );
NAND3xp33_ASAP7_75t_L g947 ( .A(n_680), .B(n_948), .C(n_951), .Y(n_947) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g893 ( .A(n_681), .B(n_894), .Y(n_893) );
AND2x2_ASAP7_75t_L g897 ( .A(n_681), .B(n_798), .Y(n_897) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g714 ( .A(n_682), .B(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g735 ( .A(n_682), .Y(n_735) );
OR2x2_ASAP7_75t_L g769 ( .A(n_682), .B(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g776 ( .A(n_682), .Y(n_776) );
AND2x2_ASAP7_75t_L g808 ( .A(n_682), .B(n_738), .Y(n_808) );
AO21x2_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_686), .B(n_698), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND3xp33_ASAP7_75t_SL g686 ( .A(n_687), .B(n_690), .C(n_693), .Y(n_686) );
AOI31xp33_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_725), .A3(n_730), .B(n_732), .Y(n_700) );
INVx1_ASAP7_75t_L g740 ( .A(n_701), .Y(n_740) );
OAI21xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_707), .B(n_713), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
OR2x2_ASAP7_75t_L g934 ( .A(n_704), .B(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVxp67_ASAP7_75t_L g784 ( .A(n_706), .Y(n_784) );
INVx2_ASAP7_75t_L g816 ( .A(n_706), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_707), .B(n_730), .Y(n_742) );
OAI21xp33_ASAP7_75t_L g922 ( .A1(n_707), .A2(n_923), .B(n_924), .Y(n_922) );
INVx2_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_711), .Y(n_708) );
INVxp67_ASAP7_75t_SL g822 ( .A(n_709), .Y(n_822) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g756 ( .A(n_710), .Y(n_756) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AND2x4_ASAP7_75t_L g815 ( .A(n_712), .B(n_816), .Y(n_815) );
AND2x2_ASAP7_75t_L g745 ( .A(n_714), .B(n_746), .Y(n_745) );
NAND2x1_ASAP7_75t_SL g810 ( .A(n_714), .B(n_737), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_714), .B(n_798), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_714), .B(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g938 ( .A(n_714), .Y(n_938) );
INVx2_ASAP7_75t_L g736 ( .A(n_715), .Y(n_736) );
AND2x2_ASAP7_75t_L g751 ( .A(n_715), .B(n_735), .Y(n_751) );
INVx1_ASAP7_75t_L g761 ( .A(n_715), .Y(n_761) );
NOR2x1_ASAP7_75t_L g775 ( .A(n_715), .B(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g779 ( .A(n_715), .Y(n_779) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_715), .Y(n_795) );
INVx1_ASAP7_75t_L g858 ( .A(n_715), .Y(n_858) );
OR2x6_ASAP7_75t_L g715 ( .A(n_716), .B(n_722), .Y(n_715) );
OAI21x1_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B(n_720), .Y(n_716) );
NOR2xp67_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
OR2x2_ASAP7_75t_L g940 ( .A(n_729), .B(n_847), .Y(n_940) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_732), .A2(n_821), .B1(n_823), .B2(n_825), .Y(n_820) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_734), .B(n_737), .Y(n_733) );
AND2x2_ASAP7_75t_L g826 ( .A(n_734), .B(n_798), .Y(n_826) );
AND2x2_ASAP7_75t_L g924 ( .A(n_734), .B(n_777), .Y(n_924) );
AND2x2_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
AND2x2_ASAP7_75t_L g778 ( .A(n_737), .B(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g747 ( .A(n_738), .Y(n_747) );
INVx1_ASAP7_75t_L g894 ( .A(n_738), .Y(n_894) );
AOI221x1_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_741), .B1(n_743), .B2(n_752), .C(n_757), .Y(n_739) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_748), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AOI22xp5_ASAP7_75t_L g836 ( .A1(n_745), .A2(n_759), .B1(n_837), .B2(n_838), .Y(n_836) );
INVxp67_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
OR2x2_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
OR2x2_ASAP7_75t_L g844 ( .A(n_749), .B(n_760), .Y(n_844) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
AND2x2_ASAP7_75t_L g843 ( .A(n_751), .B(n_777), .Y(n_843) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g866 ( .A(n_755), .Y(n_866) );
INVx1_ASAP7_75t_L g772 ( .A(n_756), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_756), .B(n_824), .Y(n_935) );
OAI221xp5_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_762), .B1(n_766), .B2(n_771), .C(n_773), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
OR2x2_ASAP7_75t_SL g803 ( .A(n_760), .B(n_804), .Y(n_803) );
HB1xp67_ASAP7_75t_L g905 ( .A(n_760), .Y(n_905) );
OR2x2_ASAP7_75t_L g943 ( .A(n_760), .B(n_859), .Y(n_943) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g767 ( .A(n_761), .B(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_763), .B(n_814), .Y(n_880) );
AND2x2_ASAP7_75t_L g902 ( .A(n_763), .B(n_903), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_763), .B(n_950), .Y(n_949) );
AND2x2_ASAP7_75t_L g829 ( .A(n_764), .B(n_830), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_764), .B(n_865), .Y(n_864) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
OR2x2_ASAP7_75t_L g771 ( .A(n_765), .B(n_772), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_765), .A2(n_806), .B1(n_810), .B2(n_811), .Y(n_805) );
INVxp67_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
OAI21xp33_ASAP7_75t_L g871 ( .A1(n_767), .A2(n_872), .B(n_877), .Y(n_871) );
AND2x2_ASAP7_75t_L g832 ( .A(n_768), .B(n_795), .Y(n_832) );
INVx1_ASAP7_75t_L g931 ( .A(n_768), .Y(n_931) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
OR2x2_ASAP7_75t_L g791 ( .A(n_769), .B(n_792), .Y(n_791) );
BUFx2_ASAP7_75t_L g876 ( .A(n_770), .Y(n_876) );
AND3x2_ASAP7_75t_L g780 ( .A(n_772), .B(n_781), .C(n_784), .Y(n_780) );
OR2x2_ASAP7_75t_L g801 ( .A(n_772), .B(n_802), .Y(n_801) );
OAI21xp5_ASAP7_75t_SL g773 ( .A1(n_774), .A2(n_778), .B(n_780), .Y(n_773) );
AND2x4_ASAP7_75t_L g774 ( .A(n_775), .B(n_777), .Y(n_774) );
INVx2_ASAP7_75t_L g800 ( .A(n_775), .Y(n_800) );
INVx2_ASAP7_75t_L g804 ( .A(n_777), .Y(n_804) );
INVx1_ASAP7_75t_L g862 ( .A(n_777), .Y(n_862) );
AND2x2_ASAP7_75t_L g910 ( .A(n_779), .B(n_792), .Y(n_910) );
AND2x2_ASAP7_75t_L g852 ( .A(n_781), .B(n_815), .Y(n_852) );
INVx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
OR2x2_ASAP7_75t_L g839 ( .A(n_782), .B(n_840), .Y(n_839) );
INVx2_ASAP7_75t_L g847 ( .A(n_782), .Y(n_847) );
INVx2_ASAP7_75t_SL g782 ( .A(n_783), .Y(n_782) );
HB1xp67_ASAP7_75t_L g819 ( .A(n_784), .Y(n_819) );
AOI211xp5_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_789), .B(n_796), .C(n_805), .Y(n_785) );
AND2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
OR2x2_ASAP7_75t_L g790 ( .A(n_791), .B(n_793), .Y(n_790) );
OAI221xp5_ASAP7_75t_SL g827 ( .A1(n_791), .A2(n_828), .B1(n_831), .B2(n_833), .C(n_836), .Y(n_827) );
INVxp67_ASAP7_75t_L g853 ( .A(n_791), .Y(n_853) );
INVx2_ASAP7_75t_L g798 ( .A(n_792), .Y(n_798) );
HB1xp67_ASAP7_75t_L g892 ( .A(n_792), .Y(n_892) );
HB1xp67_ASAP7_75t_L g918 ( .A(n_793), .Y(n_918) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
HB1xp67_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_798), .B(n_799), .Y(n_797) );
OR2x2_ASAP7_75t_L g942 ( .A(n_798), .B(n_800), .Y(n_942) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g923 ( .A(n_802), .Y(n_923) );
OR2x2_ASAP7_75t_L g937 ( .A(n_804), .B(n_938), .Y(n_937) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
AND2x4_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_808), .B(n_858), .Y(n_882) );
BUFx3_ASAP7_75t_L g911 ( .A(n_808), .Y(n_911) );
INVx2_ASAP7_75t_L g930 ( .A(n_809), .Y(n_930) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
NOR2xp67_ASAP7_75t_SL g812 ( .A(n_813), .B(n_814), .Y(n_812) );
AND2x4_ASAP7_75t_L g877 ( .A(n_813), .B(n_815), .Y(n_877) );
INVx3_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
BUFx3_ASAP7_75t_L g900 ( .A(n_815), .Y(n_900) );
INVx1_ASAP7_75t_L g888 ( .A(n_816), .Y(n_888) );
NOR3xp33_ASAP7_75t_L g817 ( .A(n_818), .B(n_827), .C(n_841), .Y(n_817) );
AND2x2_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
HB1xp67_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
AND2x2_ASAP7_75t_L g837 ( .A(n_824), .B(n_834), .Y(n_837) );
INVx2_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_830), .B(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g916 ( .A(n_830), .Y(n_916) );
INVx2_ASAP7_75t_SL g831 ( .A(n_832), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_834), .B(n_835), .Y(n_833) );
BUFx3_ASAP7_75t_L g870 ( .A(n_834), .Y(n_870) );
AND2x4_ASAP7_75t_SL g917 ( .A(n_834), .B(n_903), .Y(n_917) );
INVx2_ASAP7_75t_L g855 ( .A(n_835), .Y(n_855) );
INVx2_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
HB1xp67_ASAP7_75t_L g945 ( .A(n_840), .Y(n_945) );
AOI21xp33_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_844), .B(n_845), .Y(n_841) );
OAI222xp33_ASAP7_75t_L g883 ( .A1(n_842), .A2(n_884), .B1(n_890), .B2(n_895), .C1(n_899), .C2(n_901), .Y(n_883) );
INVx2_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_849), .B(n_912), .Y(n_848) );
NOR4xp25_ASAP7_75t_L g849 ( .A(n_850), .B(n_867), .C(n_883), .D(n_904), .Y(n_849) );
NAND2xp5_ASAP7_75t_SL g850 ( .A(n_851), .B(n_860), .Y(n_850) );
AOI21xp5_ASAP7_75t_L g851 ( .A1(n_852), .A2(n_853), .B(n_854), .Y(n_851) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_855), .B(n_856), .Y(n_854) );
OR2x2_ASAP7_75t_L g856 ( .A(n_857), .B(n_859), .Y(n_856) );
HB1xp67_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
AND2x2_ASAP7_75t_L g898 ( .A(n_858), .B(n_876), .Y(n_898) );
HB1xp67_ASAP7_75t_L g920 ( .A(n_859), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_861), .B(n_863), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx2_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
OAI211xp5_ASAP7_75t_L g867 ( .A1(n_868), .A2(n_869), .B(n_871), .C(n_878), .Y(n_867) );
INVx2_ASAP7_75t_L g927 ( .A(n_870), .Y(n_927) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVxp67_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_879), .B(n_881), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_885), .B(n_916), .Y(n_946) );
INVx2_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
NAND2x1p5_ASAP7_75t_L g886 ( .A(n_887), .B(n_889), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
AND2x2_ASAP7_75t_L g891 ( .A(n_892), .B(n_893), .Y(n_891) );
INVx1_ASAP7_75t_L g952 ( .A(n_894), .Y(n_952) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
AND2x2_ASAP7_75t_L g896 ( .A(n_897), .B(n_898), .Y(n_896) );
INVx1_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
OAI32xp33_ASAP7_75t_L g904 ( .A1(n_905), .A2(n_906), .A3(n_907), .B1(n_909), .B2(n_994), .Y(n_904) );
INVx2_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
OAI221xp5_ASAP7_75t_L g944 ( .A1(n_909), .A2(n_929), .B1(n_945), .B2(n_946), .C(n_947), .Y(n_944) );
NAND2x2_ASAP7_75t_L g909 ( .A(n_910), .B(n_911), .Y(n_909) );
AOI211x1_ASAP7_75t_L g912 ( .A1(n_913), .A2(n_919), .B(n_921), .C(n_944), .Y(n_912) );
AND2x2_ASAP7_75t_L g913 ( .A(n_914), .B(n_918), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
NAND2xp67_ASAP7_75t_L g915 ( .A(n_916), .B(n_917), .Y(n_915) );
HB1xp67_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
NAND3xp33_ASAP7_75t_L g921 ( .A(n_922), .B(n_925), .C(n_932), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_926), .B(n_928), .Y(n_925) );
INVxp67_ASAP7_75t_SL g926 ( .A(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
OR2x2_ASAP7_75t_L g929 ( .A(n_930), .B(n_931), .Y(n_929) );
AOI22xp5_ASAP7_75t_L g932 ( .A1(n_933), .A2(n_936), .B1(n_939), .B2(n_941), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
INVx2_ASAP7_75t_SL g936 ( .A(n_937), .Y(n_936) );
INVx2_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_942), .B(n_943), .Y(n_941) );
INVxp67_ASAP7_75t_SL g948 ( .A(n_949), .Y(n_948) );
INVx1_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
NAND2x1_ASAP7_75t_L g953 ( .A(n_954), .B(n_957), .Y(n_953) );
NOR2xp33_ASAP7_75t_L g958 ( .A(n_959), .B(n_969), .Y(n_958) );
CKINVDCx20_ASAP7_75t_R g959 ( .A(n_960), .Y(n_959) );
INVx1_ASAP7_75t_L g979 ( .A(n_960), .Y(n_979) );
INVx1_ASAP7_75t_L g968 ( .A(n_961), .Y(n_968) );
INVx1_ASAP7_75t_L g966 ( .A(n_962), .Y(n_966) );
NOR2xp33_ASAP7_75t_L g981 ( .A(n_969), .B(n_982), .Y(n_981) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
NOR2xp33_ASAP7_75t_L g971 ( .A(n_972), .B(n_973), .Y(n_971) );
BUFx3_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
BUFx2_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
CKINVDCx5p33_ASAP7_75t_R g978 ( .A(n_979), .Y(n_978) );
INVx1_ASAP7_75t_L g982 ( .A(n_979), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g980 ( .A(n_981), .B(n_983), .Y(n_980) );
INVx1_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
CKINVDCx20_ASAP7_75t_R g988 ( .A(n_989), .Y(n_988) );
INVx2_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
INVx5_ASAP7_75t_SL g991 ( .A(n_992), .Y(n_991) );
endmodule