module fake_jpeg_29894_n_534 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_534);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_534;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_14),
.B(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_18),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_51),
.B(n_53),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx11_ASAP7_75t_L g157 ( 
.A(n_55),
.Y(n_157)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_59),
.B(n_72),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_67),
.Y(n_132)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_70),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_71),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_18),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_73),
.Y(n_152)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

BUFx4f_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_46),
.Y(n_76)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_76),
.Y(n_143)
);

NAND2x1_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_0),
.Y(n_77)
);

INVx5_ASAP7_75t_SL g123 ( 
.A(n_77),
.Y(n_123)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_81),
.Y(n_147)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_82),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_83),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_29),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_84),
.Y(n_109)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_37),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_86),
.B(n_90),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_31),
.B(n_17),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_91),
.Y(n_151)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_93),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_94),
.Y(n_162)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

BUFx4f_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_96),
.Y(n_128)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

BUFx4f_ASAP7_75t_SL g199 ( 
.A(n_104),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_79),
.B(n_40),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_115),
.B(n_141),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_67),
.A2(n_45),
.B1(n_24),
.B2(n_19),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_116),
.A2(n_137),
.B1(n_85),
.B2(n_87),
.Y(n_188)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

INVx11_ASAP7_75t_L g217 ( 
.A(n_131),
.Y(n_217)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_66),
.A2(n_45),
.B1(n_30),
.B2(n_28),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_138),
.Y(n_179)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_93),
.B(n_40),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_52),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_145),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_61),
.Y(n_153)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_63),
.B(n_31),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_160),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_75),
.Y(n_160)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_118),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_165),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_123),
.A2(n_99),
.B1(n_64),
.B2(n_91),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_166),
.A2(n_171),
.B1(n_202),
.B2(n_213),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_134),
.Y(n_167)
);

INVx5_ASAP7_75t_SL g248 ( 
.A(n_167),
.Y(n_248)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_169),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

INVx11_ASAP7_75t_L g264 ( 
.A(n_170),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_123),
.A2(n_62),
.B1(n_73),
.B2(n_70),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_172),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_173),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_107),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_174),
.B(n_177),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_144),
.A2(n_58),
.B1(n_69),
.B2(n_71),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_175),
.A2(n_206),
.B1(n_220),
.B2(n_223),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_117),
.B(n_19),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_104),
.Y(n_178)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_178),
.Y(n_275)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_124),
.Y(n_182)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_182),
.Y(n_236)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_108),
.Y(n_183)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_125),
.Y(n_184)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_184),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g185 ( 
.A(n_121),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_185),
.Y(n_231)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_125),
.Y(n_186)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

BUFx16f_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_187),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_188),
.B(n_205),
.Y(n_235)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_120),
.Y(n_189)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_189),
.Y(n_254)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_122),
.Y(n_190)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_190),
.Y(n_257)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_135),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_192),
.Y(n_250)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_124),
.Y(n_193)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_193),
.Y(n_252)
);

NOR2x1_ASAP7_75t_L g194 ( 
.A(n_105),
.B(n_96),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_194),
.B(n_195),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_117),
.B(n_154),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_113),
.Y(n_196)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_196),
.Y(n_265)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_136),
.Y(n_198)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_198),
.Y(n_269)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_114),
.Y(n_200)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_200),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_154),
.B(n_45),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_201),
.B(n_203),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_151),
.A2(n_83),
.B1(n_45),
.B2(n_55),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_109),
.B(n_45),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_109),
.B(n_77),
.C(n_65),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_204),
.B(n_219),
.C(n_21),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_142),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_137),
.A2(n_156),
.B1(n_21),
.B2(n_27),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_127),
.Y(n_207)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_207),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_110),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_212),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_162),
.B(n_19),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_168),
.Y(n_241)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_107),
.Y(n_210)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_210),
.Y(n_263)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_132),
.Y(n_211)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_211),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_116),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_132),
.A2(n_56),
.B1(n_30),
.B2(n_28),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_163),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_214),
.B(n_216),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_119),
.B(n_24),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_215),
.B(n_218),
.Y(n_266)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_126),
.B(n_24),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_149),
.B(n_32),
.C(n_30),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_111),
.A2(n_106),
.B1(n_112),
.B2(n_148),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_161),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_221),
.B(n_222),
.Y(n_262)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_102),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_103),
.A2(n_23),
.B1(n_48),
.B2(n_41),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_157),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_224),
.B(n_128),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_159),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_227),
.B(n_237),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_187),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_229),
.B(n_241),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_212),
.A2(n_159),
.B1(n_152),
.B2(n_150),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_230),
.A2(n_273),
.B1(n_175),
.B2(n_220),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_103),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_129),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_238),
.B(n_246),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_187),
.A2(n_111),
.B1(n_130),
.B2(n_158),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_242),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_176),
.B(n_150),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_197),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_247),
.B(n_271),
.Y(n_288)
);

O2A1O1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_171),
.A2(n_22),
.B(n_23),
.C(n_25),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_249),
.B(n_216),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_SL g255 ( 
.A(n_219),
.B(n_33),
.C(n_35),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_256),
.C(n_261),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_166),
.B(n_82),
.Y(n_261)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_267),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_202),
.A2(n_152),
.B1(n_129),
.B2(n_22),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_268),
.A2(n_225),
.B1(n_235),
.B2(n_260),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_205),
.B(n_48),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_192),
.B(n_41),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_170),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_213),
.A2(n_27),
.B1(n_25),
.B2(n_35),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_276),
.B(n_280),
.Y(n_331)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_277),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_262),
.Y(n_280)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_228),
.Y(n_283)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_283),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_235),
.A2(n_232),
.B(n_238),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_284),
.A2(n_231),
.B(n_274),
.Y(n_353)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_236),
.Y(n_285)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_285),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_240),
.A2(n_182),
.B1(n_193),
.B2(n_191),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_286),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_226),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_289),
.B(n_291),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_227),
.B(n_180),
.C(n_164),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_290),
.B(n_307),
.C(n_278),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_253),
.B(n_198),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_292),
.A2(n_302),
.B1(n_321),
.B2(n_248),
.Y(n_351)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_251),
.Y(n_293)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_293),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_269),
.Y(n_294)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_294),
.Y(n_337)
);

AND2x6_ASAP7_75t_L g295 ( 
.A(n_255),
.B(n_35),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_295),
.B(n_297),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_236),
.Y(n_296)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_296),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_246),
.B(n_167),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_250),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_298),
.Y(n_333)
);

INVx8_ASAP7_75t_L g299 ( 
.A(n_275),
.Y(n_299)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_299),
.Y(n_343)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_228),
.Y(n_300)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_300),
.Y(n_348)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_233),
.Y(n_301)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_301),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_235),
.A2(n_181),
.B1(n_173),
.B2(n_179),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_243),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_303),
.B(n_314),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_305),
.B(n_254),
.Y(n_326)
);

BUFx12_ASAP7_75t_L g306 ( 
.A(n_270),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_306),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_256),
.B(n_197),
.C(n_128),
.Y(n_307)
);

OA22x2_ASAP7_75t_L g325 ( 
.A1(n_308),
.A2(n_311),
.B1(n_292),
.B2(n_287),
.Y(n_325)
);

INVx6_ASAP7_75t_L g309 ( 
.A(n_252),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_309),
.A2(n_316),
.B1(n_319),
.B2(n_320),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_259),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_310),
.B(n_312),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_225),
.A2(n_217),
.B1(n_191),
.B2(n_178),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_311),
.A2(n_248),
.B1(n_250),
.B2(n_234),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_237),
.B(n_37),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_244),
.B(n_37),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_313),
.B(n_315),
.Y(n_330)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_243),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_261),
.B(n_241),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_233),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_260),
.B(n_217),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_317),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_241),
.B(n_0),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_318),
.B(n_0),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_264),
.Y(n_319)
);

INVx5_ASAP7_75t_L g320 ( 
.A(n_270),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_249),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_279),
.B(n_245),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_324),
.B(n_327),
.C(n_334),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_325),
.B(n_339),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_326),
.B(n_351),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_279),
.B(n_245),
.Y(n_327)
);

OAI32xp33_ASAP7_75t_L g329 ( 
.A1(n_304),
.A2(n_252),
.A3(n_254),
.B1(n_257),
.B2(n_263),
.Y(n_329)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_329),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_332),
.B(n_349),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_308),
.B(n_257),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_336),
.A2(n_314),
.B(n_303),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_304),
.B(n_263),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_340),
.A2(n_281),
.B1(n_299),
.B2(n_293),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_284),
.A2(n_269),
.B(n_231),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_341),
.A2(n_353),
.B(n_199),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_278),
.B(n_258),
.C(n_274),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_345),
.B(n_358),
.C(n_359),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_315),
.B(n_258),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_347),
.B(n_354),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_296),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_290),
.B(n_265),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_307),
.B(n_265),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_312),
.B(n_239),
.C(n_275),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_313),
.B(n_239),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_360),
.B(n_302),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_310),
.B(n_234),
.Y(n_361)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_361),
.Y(n_382)
);

O2A1O1Ixp33_ASAP7_75t_L g363 ( 
.A1(n_352),
.A2(n_305),
.B(n_281),
.C(n_295),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_363),
.A2(n_371),
.B(n_379),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_364),
.B(n_185),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_334),
.B(n_318),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_365),
.B(n_358),
.C(n_324),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_335),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_366),
.B(n_375),
.Y(n_420)
);

CKINVDCx12_ASAP7_75t_R g367 ( 
.A(n_342),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_367),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_368),
.A2(n_391),
.B1(n_396),
.B2(n_338),
.Y(n_421)
);

BUFx12f_ASAP7_75t_L g373 ( 
.A(n_355),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_SL g424 ( 
.A1(n_373),
.A2(n_392),
.B1(n_393),
.B2(n_185),
.Y(n_424)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_346),
.Y(n_375)
);

AND2x6_ASAP7_75t_L g376 ( 
.A(n_344),
.B(n_288),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_SL g404 ( 
.A(n_376),
.B(n_353),
.C(n_329),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_335),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_378),
.B(n_380),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_352),
.A2(n_320),
.B(n_282),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_350),
.B(n_309),
.Y(n_380)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_335),
.Y(n_383)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_383),
.Y(n_399)
);

A2O1A1O1Ixp25_ASAP7_75t_L g411 ( 
.A1(n_384),
.A2(n_341),
.B(n_339),
.C(n_326),
.D(n_325),
.Y(n_411)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_346),
.Y(n_385)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_385),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_331),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_386),
.B(n_389),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_333),
.B(n_306),
.Y(n_387)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_387),
.Y(n_402)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_322),
.Y(n_388)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_388),
.Y(n_413)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_348),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_336),
.A2(n_285),
.B1(n_277),
.B2(n_319),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_390),
.A2(n_351),
.B1(n_356),
.B2(n_362),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_336),
.A2(n_306),
.B1(n_199),
.B2(n_264),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_357),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_361),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_328),
.B(n_17),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_394),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_328),
.B(n_17),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_395),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_332),
.B(n_16),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_398),
.B(n_403),
.C(n_406),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_369),
.B(n_327),
.C(n_354),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_404),
.B(n_418),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_369),
.B(n_374),
.C(n_365),
.Y(n_406)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_409),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_374),
.B(n_345),
.C(n_347),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_410),
.B(n_427),
.C(n_377),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_411),
.A2(n_368),
.B(n_376),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_372),
.A2(n_325),
.B1(n_330),
.B2(n_359),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_412),
.A2(n_419),
.B1(n_422),
.B2(n_426),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_330),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_415),
.B(n_417),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_397),
.B(n_360),
.Y(n_417)
);

A2O1A1Ixp33_ASAP7_75t_L g418 ( 
.A1(n_381),
.A2(n_325),
.B(n_355),
.C(n_337),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_372),
.A2(n_340),
.B1(n_362),
.B2(n_343),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_421),
.B(n_363),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_370),
.A2(n_323),
.B1(n_16),
.B2(n_15),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_364),
.B(n_199),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_423),
.B(n_425),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_424),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_381),
.A2(n_170),
.B1(n_16),
.B2(n_34),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_383),
.B(n_34),
.C(n_1),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_370),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_428),
.A2(n_422),
.B1(n_388),
.B2(n_416),
.Y(n_453)
);

MAJx2_ASAP7_75t_L g431 ( 
.A(n_406),
.B(n_393),
.C(n_382),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_431),
.B(n_445),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_407),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_432),
.B(n_450),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_435),
.A2(n_452),
.B1(n_414),
.B2(n_428),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_408),
.B(n_373),
.Y(n_436)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_436),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_398),
.B(n_384),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_437),
.B(n_441),
.C(n_442),
.Y(n_459)
);

INVx11_ASAP7_75t_L g440 ( 
.A(n_420),
.Y(n_440)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_440),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_410),
.B(n_382),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_423),
.B(n_403),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_401),
.B(n_391),
.Y(n_443)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_443),
.Y(n_470)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_413),
.Y(n_444)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_444),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_425),
.B(n_417),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_446),
.B(n_448),
.C(n_449),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_412),
.B(n_371),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_399),
.B(n_379),
.C(n_390),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_402),
.B(n_392),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_415),
.B(n_389),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_451),
.B(n_34),
.C(n_6),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_453),
.B(n_4),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_405),
.B(n_373),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_454),
.B(n_373),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_434),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_455),
.B(n_456),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_429),
.A2(n_419),
.B1(n_409),
.B2(n_418),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_448),
.A2(n_426),
.B1(n_411),
.B2(n_414),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_463),
.B(n_464),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_466),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_452),
.A2(n_435),
.B1(n_447),
.B2(n_438),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_467),
.B(n_472),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_443),
.A2(n_427),
.B1(n_400),
.B2(n_375),
.Y(n_468)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_468),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_451),
.A2(n_385),
.B1(n_3),
.B2(n_4),
.Y(n_469)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_469),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_437),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_471),
.B(n_441),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_449),
.B(n_5),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_473),
.B(n_7),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_474),
.B(n_442),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_430),
.B(n_5),
.C(n_6),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_475),
.B(n_446),
.C(n_431),
.Y(n_478)
);

BUFx12_ASAP7_75t_L g476 ( 
.A(n_475),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_476),
.B(n_489),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_478),
.B(n_488),
.Y(n_504)
);

AOI21xp33_ASAP7_75t_L g479 ( 
.A1(n_470),
.A2(n_430),
.B(n_440),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_479),
.A2(n_488),
.B(n_478),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_482),
.B(n_459),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_R g483 ( 
.A(n_463),
.B(n_439),
.C(n_445),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_483),
.A2(n_462),
.B(n_456),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_486),
.B(n_487),
.Y(n_499)
);

NAND3xp33_ASAP7_75t_L g487 ( 
.A(n_460),
.B(n_439),
.C(n_433),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_459),
.B(n_433),
.C(n_7),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_458),
.B(n_5),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_461),
.B(n_7),
.Y(n_491)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_491),
.Y(n_498)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_492),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_493),
.B(n_494),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_477),
.A2(n_457),
.B1(n_472),
.B2(n_473),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_495),
.A2(n_480),
.B1(n_482),
.B2(n_471),
.Y(n_510)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_497),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_483),
.B(n_465),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_506),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_477),
.A2(n_468),
.B1(n_457),
.B2(n_465),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_501),
.B(n_502),
.Y(n_511)
);

BUFx24_ASAP7_75t_SL g502 ( 
.A(n_484),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_490),
.A2(n_461),
.B1(n_462),
.B2(n_469),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_505),
.B(n_476),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_485),
.B(n_474),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_501),
.A2(n_485),
.B(n_481),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_507),
.B(n_508),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_499),
.A2(n_481),
.B(n_480),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_510),
.B(n_514),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_496),
.B(n_504),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_513),
.B(n_515),
.Y(n_518)
);

NAND2x1_ASAP7_75t_SL g515 ( 
.A(n_494),
.B(n_476),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_516),
.B(n_498),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_517),
.B(n_519),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_509),
.B(n_503),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_509),
.B(n_493),
.C(n_506),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_522),
.B(n_500),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_520),
.B(n_507),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_523),
.B(n_518),
.C(n_515),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_521),
.B(n_511),
.C(n_512),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_525),
.B(n_526),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_528),
.A2(n_518),
.B(n_523),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_529),
.B(n_527),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_530),
.A2(n_524),
.B1(n_8),
.B2(n_10),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_531),
.B(n_8),
.C(n_10),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_10),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_533),
.B(n_10),
.Y(n_534)
);


endmodule