module fake_jpeg_21946_n_101 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_101);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_101;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_10),
.B(n_4),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_6),
.B(n_0),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_19),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_25),
.A2(n_33),
.B1(n_19),
.B2(n_16),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_23),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_27),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_30),
.Y(n_41)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_2),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_32),
.B(n_23),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_22),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_16),
.Y(n_43)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_43),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_42),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_26),
.B(n_18),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_49),
.Y(n_56)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_24),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_21),
.C(n_13),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_8),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_33),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_29),
.A2(n_21),
.B1(n_24),
.B2(n_12),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_11),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_27),
.B(n_20),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_46),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_63),
.C(n_40),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_54),
.B1(n_57),
.B2(n_61),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_34),
.B1(n_30),
.B2(n_21),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_32),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_55),
.B(n_58),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_25),
.B1(n_12),
.B2(n_20),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_15),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_8),
.Y(n_60)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_37),
.A2(n_31),
.B1(n_4),
.B2(n_3),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_10),
.Y(n_64)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_65),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_62),
.A2(n_39),
.B(n_48),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_72),
.C(n_74),
.Y(n_81)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_59),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_41),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_75),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_41),
.B(n_44),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_37),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_77),
.B(n_78),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_83),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_63),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_84),
.C(n_66),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_72),
.A2(n_53),
.B1(n_57),
.B2(n_50),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_70),
.A2(n_61),
.B1(n_40),
.B2(n_35),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_79),
.B(n_68),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_88),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_83),
.B(n_68),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_81),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_93),
.C(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_92),
.B(n_69),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_80),
.B1(n_81),
.B2(n_84),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

NOR2x1_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_96),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_76),
.C(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_97),
.B(n_90),
.Y(n_99)
);

OAI321xp33_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_97),
.A3(n_91),
.B1(n_98),
.B2(n_69),
.C(n_73),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_35),
.Y(n_101)
);


endmodule