module real_aes_17407_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_815;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
CKINVDCx5p33_ASAP7_75t_R g548 ( .A(n_0), .Y(n_548) );
AND2x4_ASAP7_75t_L g105 ( .A(n_1), .B(n_106), .Y(n_105) );
AOI22xp5_ASAP7_75t_L g267 ( .A1(n_2), .A2(n_4), .B1(n_268), .B2(n_269), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_3), .A2(n_23), .B1(n_217), .B2(n_251), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g153 ( .A1(n_5), .A2(n_53), .B1(n_154), .B2(n_155), .Y(n_153) );
BUFx3_ASAP7_75t_L g601 ( .A(n_6), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_7), .A2(n_13), .B1(n_169), .B2(n_170), .Y(n_168) );
INVx1_ASAP7_75t_L g106 ( .A(n_8), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_9), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_10), .B(n_194), .Y(n_579) );
OR2x2_ASAP7_75t_L g112 ( .A(n_11), .B(n_32), .Y(n_112) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_12), .Y(n_146) );
INVx1_ASAP7_75t_L g838 ( .A(n_14), .Y(n_838) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_15), .B(n_145), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_16), .B(n_185), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_17), .A2(n_86), .B1(n_145), .B2(n_251), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g832 ( .A1(n_18), .A2(n_19), .B1(n_833), .B2(n_834), .Y(n_832) );
INVx1_ASAP7_75t_L g834 ( .A(n_18), .Y(n_834) );
INVx1_ASAP7_75t_L g833 ( .A(n_19), .Y(n_833) );
OAI21x1_ASAP7_75t_L g159 ( .A1(n_20), .A2(n_49), .B(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_21), .B(n_496), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_22), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_24), .B(n_217), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_25), .B(n_142), .Y(n_209) );
INVx4_ASAP7_75t_R g193 ( .A(n_26), .Y(n_193) );
AO32x1_ASAP7_75t_L g517 ( .A1(n_27), .A2(n_205), .A3(n_206), .B1(n_518), .B2(n_521), .Y(n_517) );
AO32x2_ASAP7_75t_L g609 ( .A1(n_27), .A2(n_205), .A3(n_206), .B1(n_518), .B2(n_521), .Y(n_609) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_28), .B(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g273 ( .A(n_29), .Y(n_273) );
A2O1A1Ixp33_ASAP7_75t_SL g248 ( .A1(n_30), .A2(n_141), .B(n_169), .C(n_249), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_31), .A2(n_46), .B1(n_169), .B2(n_173), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_33), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_34), .A2(n_52), .B1(n_195), .B2(n_217), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_35), .A2(n_91), .B1(n_173), .B2(n_251), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_36), .B(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_37), .B(n_529), .Y(n_533) );
INVx1_ASAP7_75t_L g213 ( .A(n_38), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_39), .B(n_169), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_40), .A2(n_68), .B1(n_173), .B2(n_557), .Y(n_556) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_41), .Y(n_227) );
INVx2_ASAP7_75t_L g117 ( .A(n_42), .Y(n_117) );
BUFx3_ASAP7_75t_L g111 ( .A(n_43), .Y(n_111) );
INVx1_ASAP7_75t_L g125 ( .A(n_43), .Y(n_125) );
INVx1_ASAP7_75t_L g489 ( .A(n_44), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_45), .B(n_535), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_47), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g172 ( .A1(n_48), .A2(n_85), .B1(n_169), .B2(n_173), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_50), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g593 ( .A(n_51), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_54), .A2(n_79), .B1(n_148), .B2(n_529), .Y(n_589) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_55), .Y(n_179) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_56), .A2(n_83), .B1(n_145), .B2(n_251), .Y(n_597) );
INVx1_ASAP7_75t_L g160 ( .A(n_57), .Y(n_160) );
AND2x4_ASAP7_75t_L g163 ( .A(n_58), .B(n_164), .Y(n_163) );
AOI22xp5_ASAP7_75t_L g129 ( .A1(n_59), .A2(n_78), .B1(n_130), .B2(n_131), .Y(n_129) );
INVx1_ASAP7_75t_L g131 ( .A(n_59), .Y(n_131) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_60), .A2(n_90), .B1(n_173), .B2(n_266), .Y(n_265) );
AO22x1_ASAP7_75t_L g143 ( .A1(n_61), .A2(n_73), .B1(n_144), .B2(n_147), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_62), .B(n_251), .Y(n_578) );
INVx1_ASAP7_75t_L g164 ( .A(n_63), .Y(n_164) );
AND2x2_ASAP7_75t_L g252 ( .A(n_64), .B(n_205), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_65), .B(n_205), .Y(n_584) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_66), .A2(n_151), .B(n_154), .C(n_547), .Y(n_546) );
NAND3xp33_ASAP7_75t_L g583 ( .A(n_67), .B(n_251), .C(n_582), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_69), .B(n_154), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_70), .Y(n_243) );
AND2x2_ASAP7_75t_L g549 ( .A(n_71), .B(n_199), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_72), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_74), .B(n_217), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_75), .A2(n_96), .B1(n_145), .B2(n_148), .Y(n_591) );
INVx2_ASAP7_75t_L g142 ( .A(n_76), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_77), .B(n_229), .Y(n_570) );
INVx1_ASAP7_75t_L g130 ( .A(n_78), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_80), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_81), .B(n_205), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_82), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_84), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_87), .B(n_582), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_88), .A2(n_100), .B1(n_173), .B2(n_195), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_89), .B(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_92), .B(n_205), .Y(n_224) );
INVx1_ASAP7_75t_L g109 ( .A(n_93), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_93), .B(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_94), .B(n_185), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_L g188 ( .A1(n_95), .A2(n_154), .B(n_175), .C(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g198 ( .A(n_97), .B(n_199), .Y(n_198) );
NAND2xp33_ASAP7_75t_L g232 ( .A(n_98), .B(n_194), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g567 ( .A(n_99), .Y(n_567) );
AOI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_113), .B(n_837), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx5_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
BUFx3_ASAP7_75t_L g839 ( .A(n_104), .Y(n_839) );
AND2x6_ASAP7_75t_L g104 ( .A(n_105), .B(n_107), .Y(n_104) );
INVx1_ASAP7_75t_L g498 ( .A(n_107), .Y(n_498) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g829 ( .A(n_108), .Y(n_829) );
HB1xp67_ASAP7_75t_L g831 ( .A(n_108), .Y(n_831) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NOR2x1_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
INVx1_ASAP7_75t_L g505 ( .A(n_111), .Y(n_505) );
INVx1_ASAP7_75t_L g126 ( .A(n_112), .Y(n_126) );
OR2x6_ASAP7_75t_L g113 ( .A(n_114), .B(n_499), .Y(n_113) );
OAI21xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_118), .B(n_493), .Y(n_114) );
BUFx3_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x6_ASAP7_75t_SL g503 ( .A(n_116), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_117), .B(n_498), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_127), .B(n_488), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx3_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
CKINVDCx8_ASAP7_75t_R g492 ( .A(n_122), .Y(n_492) );
AND2x6_ASAP7_75t_SL g122 ( .A(n_123), .B(n_126), .Y(n_122) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_126), .B(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
XNOR2x1_ASAP7_75t_L g128 ( .A(n_129), .B(n_132), .Y(n_128) );
AO22x2_ASAP7_75t_L g507 ( .A1(n_132), .A2(n_508), .B1(n_828), .B2(n_830), .Y(n_507) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_398), .Y(n_132) );
NOR3xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_327), .C(n_369), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_301), .Y(n_134) );
AOI22xp33_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_200), .B1(n_276), .B2(n_287), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OR2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_181), .Y(n_137) );
AOI21xp33_ASAP7_75t_L g320 ( .A1(n_138), .A2(n_321), .B(n_323), .Y(n_320) );
AOI21xp33_ASAP7_75t_L g393 ( .A1(n_138), .A2(n_394), .B(n_395), .Y(n_393) );
OR2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_165), .Y(n_138) );
INVx2_ASAP7_75t_L g313 ( .A(n_139), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_139), .B(n_166), .Y(n_343) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_143), .B(n_149), .C(n_161), .Y(n_140) );
INVx6_ASAP7_75t_L g171 ( .A(n_141), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_141), .A2(n_232), .B(n_233), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_141), .B(n_143), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_141), .A2(n_247), .B1(n_519), .B2(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_141), .A2(n_578), .B(n_579), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_141), .A2(n_171), .B1(n_597), .B2(n_598), .Y(n_596) );
BUFx8_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g152 ( .A(n_142), .Y(n_152) );
INVx1_ASAP7_75t_L g175 ( .A(n_142), .Y(n_175) );
INVx1_ASAP7_75t_L g212 ( .A(n_142), .Y(n_212) );
INVxp67_ASAP7_75t_SL g144 ( .A(n_145), .Y(n_144) );
INVx3_ASAP7_75t_L g535 ( .A(n_145), .Y(n_535) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g148 ( .A(n_146), .Y(n_148) );
INVx1_ASAP7_75t_L g154 ( .A(n_146), .Y(n_154) );
INVx1_ASAP7_75t_L g156 ( .A(n_146), .Y(n_156) );
INVx3_ASAP7_75t_L g169 ( .A(n_146), .Y(n_169) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_146), .Y(n_173) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_146), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_146), .Y(n_195) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_146), .Y(n_217) );
INVx1_ASAP7_75t_L g245 ( .A(n_146), .Y(n_245) );
INVx2_ASAP7_75t_L g251 ( .A(n_146), .Y(n_251) );
OAI21xp33_ASAP7_75t_SL g208 ( .A1(n_147), .A2(n_209), .B(n_210), .Y(n_208) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_148), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g284 ( .A(n_149), .Y(n_284) );
OAI21x1_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_153), .B(n_157), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_150), .A2(n_215), .B(n_216), .Y(n_214) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_150), .A2(n_171), .B1(n_256), .B2(n_257), .Y(n_255) );
AOI21x1_ASAP7_75t_L g527 ( .A1(n_150), .A2(n_528), .B(n_530), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_150), .A2(n_171), .B1(n_556), .B2(n_558), .Y(n_555) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g230 ( .A(n_152), .Y(n_230) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_156), .B(n_190), .Y(n_189) );
OAI21xp33_ASAP7_75t_L g161 ( .A1(n_157), .A2(n_158), .B(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g176 ( .A(n_158), .Y(n_176) );
INVx2_ASAP7_75t_L g180 ( .A(n_158), .Y(n_180) );
INVx2_ASAP7_75t_L g186 ( .A(n_158), .Y(n_186) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_159), .Y(n_206) );
INVx1_ASAP7_75t_L g286 ( .A(n_161), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_162), .A2(n_241), .B(n_248), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_162), .A2(n_541), .B(n_546), .Y(n_540) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
BUFx10_ASAP7_75t_L g177 ( .A(n_163), .Y(n_177) );
BUFx10_ASAP7_75t_L g219 ( .A(n_163), .Y(n_219) );
INVx1_ASAP7_75t_L g271 ( .A(n_163), .Y(n_271) );
AO31x2_ASAP7_75t_L g553 ( .A1(n_163), .A2(n_554), .A3(n_555), .B(n_559), .Y(n_553) );
AND2x2_ASAP7_75t_L g383 ( .A(n_165), .B(n_222), .Y(n_383) );
INVx1_ASAP7_75t_L g416 ( .A(n_165), .Y(n_416) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_L g278 ( .A(n_166), .B(n_223), .Y(n_278) );
AND2x2_ASAP7_75t_L g309 ( .A(n_166), .B(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g318 ( .A(n_166), .Y(n_318) );
OR2x2_ASAP7_75t_L g337 ( .A(n_166), .B(n_183), .Y(n_337) );
AND2x2_ASAP7_75t_L g352 ( .A(n_166), .B(n_183), .Y(n_352) );
AO31x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_176), .A3(n_177), .B(n_178), .Y(n_166) );
OAI22x1_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_171), .B1(n_172), .B2(n_174), .Y(n_167) );
INVx4_ASAP7_75t_L g170 ( .A(n_169), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_170), .A2(n_227), .B(n_228), .C(n_229), .Y(n_226) );
OAI22xp5_ASAP7_75t_L g264 ( .A1(n_171), .A2(n_174), .B1(n_265), .B2(n_267), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_171), .A2(n_533), .B(n_534), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_171), .A2(n_589), .B1(n_590), .B2(n_591), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_173), .B(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g268 ( .A(n_173), .Y(n_268) );
INVx2_ASAP7_75t_L g531 ( .A(n_173), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_174), .B(n_192), .Y(n_191) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g545 ( .A(n_175), .Y(n_545) );
INVx1_ASAP7_75t_SL g590 ( .A(n_175), .Y(n_590) );
INVx2_ASAP7_75t_L g575 ( .A(n_176), .Y(n_575) );
INVx2_ASAP7_75t_L g197 ( .A(n_177), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
INVx2_ASAP7_75t_L g199 ( .A(n_180), .Y(n_199) );
BUFx2_ASAP7_75t_L g239 ( .A(n_180), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_180), .B(n_260), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_180), .B(n_273), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_180), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_182), .B(n_351), .Y(n_394) );
OR2x2_ASAP7_75t_L g482 ( .A(n_182), .B(n_343), .Y(n_482) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g310 ( .A(n_183), .Y(n_310) );
AND2x2_ASAP7_75t_L g319 ( .A(n_183), .B(n_282), .Y(n_319) );
AND2x2_ASAP7_75t_L g322 ( .A(n_183), .B(n_223), .Y(n_322) );
AND2x2_ASAP7_75t_L g341 ( .A(n_183), .B(n_222), .Y(n_341) );
AND2x4_ASAP7_75t_L g360 ( .A(n_183), .B(n_283), .Y(n_360) );
AO21x2_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_187), .B(n_198), .Y(n_183) );
AOI21x1_ASAP7_75t_L g539 ( .A1(n_184), .A2(n_540), .B(n_549), .Y(n_539) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_191), .B(n_197), .Y(n_187) );
OAI22xp33_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B1(n_195), .B2(n_196), .Y(n_192) );
INVx2_ASAP7_75t_L g266 ( .A(n_194), .Y(n_266) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_195), .A2(n_217), .B1(n_543), .B2(n_544), .Y(n_542) );
INVx1_ASAP7_75t_L g571 ( .A(n_195), .Y(n_571) );
OAI21xp33_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_220), .B(n_261), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_201), .B(n_355), .Y(n_458) );
CKINVDCx14_ASAP7_75t_R g201 ( .A(n_202), .Y(n_201) );
BUFx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_203), .B(n_275), .Y(n_274) );
INVx3_ASAP7_75t_L g291 ( .A(n_203), .Y(n_291) );
OR2x2_ASAP7_75t_L g299 ( .A(n_203), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_203), .B(n_292), .Y(n_324) );
AND2x2_ASAP7_75t_L g349 ( .A(n_203), .B(n_263), .Y(n_349) );
AND2x2_ASAP7_75t_L g367 ( .A(n_203), .B(n_297), .Y(n_367) );
INVx1_ASAP7_75t_L g406 ( .A(n_203), .Y(n_406) );
AND2x2_ASAP7_75t_L g408 ( .A(n_203), .B(n_409), .Y(n_408) );
NAND2x1p5_ASAP7_75t_SL g427 ( .A(n_203), .B(n_348), .Y(n_427) );
AND2x4_ASAP7_75t_L g203 ( .A(n_204), .B(n_207), .Y(n_203) );
NOR2x1_ASAP7_75t_L g234 ( .A(n_205), .B(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g258 ( .A(n_205), .Y(n_258) );
INVx4_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g218 ( .A(n_206), .B(n_219), .Y(n_218) );
INVx2_ASAP7_75t_SL g525 ( .A(n_206), .Y(n_525) );
BUFx3_ASAP7_75t_L g554 ( .A(n_206), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_206), .B(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g564 ( .A(n_206), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_206), .B(n_600), .Y(n_599) );
OAI21xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_214), .B(n_218), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
BUFx4f_ASAP7_75t_L g247 ( .A(n_212), .Y(n_247) );
INVx1_ASAP7_75t_L g582 ( .A(n_212), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_217), .B(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g557 ( .A(n_217), .Y(n_557) );
INVx1_ASAP7_75t_L g235 ( .A(n_219), .Y(n_235) );
AO31x2_ASAP7_75t_L g254 ( .A1(n_219), .A2(n_255), .A3(n_258), .B(n_259), .Y(n_254) );
OAI21x1_ASAP7_75t_L g565 ( .A1(n_219), .A2(n_566), .B(n_569), .Y(n_565) );
OAI21x1_ASAP7_75t_L g576 ( .A1(n_219), .A2(n_577), .B(n_580), .Y(n_576) );
AOI31xp67_ASAP7_75t_L g595 ( .A1(n_219), .A2(n_258), .A3(n_596), .B(n_599), .Y(n_595) );
OAI32xp33_ASAP7_75t_L g311 ( .A1(n_220), .A2(n_303), .A3(n_312), .B1(n_314), .B2(n_316), .Y(n_311) );
OR2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_236), .Y(n_220) );
INVx1_ASAP7_75t_L g351 ( .A(n_221), .Y(n_351) );
AND2x2_ASAP7_75t_L g359 ( .A(n_221), .B(n_360), .Y(n_359) );
BUFx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g358 ( .A(n_222), .B(n_282), .Y(n_358) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
BUFx3_ASAP7_75t_L g308 ( .A(n_223), .Y(n_308) );
AND2x2_ASAP7_75t_L g317 ( .A(n_223), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g423 ( .A(n_223), .Y(n_423) );
NAND2x1p5_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
OAI21x1_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_231), .B(n_234), .Y(n_225) );
INVx2_ASAP7_75t_SL g229 ( .A(n_230), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_230), .A2(n_570), .B1(n_571), .B2(n_572), .Y(n_569) );
INVx2_ASAP7_75t_L g293 ( .A(n_236), .Y(n_293) );
OR2x2_ASAP7_75t_L g303 ( .A(n_236), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g425 ( .A(n_236), .Y(n_425) );
OR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_253), .Y(n_236) );
AND2x2_ASAP7_75t_L g326 ( .A(n_237), .B(n_254), .Y(n_326) );
INVx2_ASAP7_75t_L g348 ( .A(n_237), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_237), .B(n_263), .Y(n_368) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g275 ( .A(n_238), .Y(n_275) );
AOI21x1_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_252), .Y(n_238) );
AO31x2_ASAP7_75t_L g263 ( .A1(n_239), .A2(n_264), .A3(n_270), .B(n_272), .Y(n_263) );
OAI21xp5_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_244), .B(n_247), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
INVx2_ASAP7_75t_L g269 ( .A(n_245), .Y(n_269) );
O2A1O1Ixp5_ASAP7_75t_L g566 ( .A1(n_247), .A2(n_269), .B(n_567), .C(n_568), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
INVx2_ASAP7_75t_SL g529 ( .A(n_251), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_253), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g357 ( .A(n_253), .Y(n_357) );
INVx2_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
BUFx2_ASAP7_75t_L g297 ( .A(n_254), .Y(n_297) );
OR2x2_ASAP7_75t_L g363 ( .A(n_254), .B(n_263), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_254), .B(n_263), .Y(n_396) );
INVx2_ASAP7_75t_L g344 ( .A(n_261), .Y(n_344) );
OR2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_274), .Y(n_261) );
OR2x2_ASAP7_75t_L g331 ( .A(n_262), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g409 ( .A(n_262), .Y(n_409) );
INVx1_ASAP7_75t_L g292 ( .A(n_263), .Y(n_292) );
INVx1_ASAP7_75t_L g300 ( .A(n_263), .Y(n_300) );
INVx1_ASAP7_75t_L g315 ( .A(n_263), .Y(n_315) );
AO31x2_ASAP7_75t_L g587 ( .A1(n_270), .A2(n_554), .A3(n_588), .B(n_592), .Y(n_587) );
INVx2_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
INVx2_ASAP7_75t_SL g521 ( .A(n_271), .Y(n_521) );
OR2x2_ASAP7_75t_L g419 ( .A(n_274), .B(n_396), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_275), .B(n_291), .Y(n_332) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_275), .Y(n_334) );
OR2x2_ASAP7_75t_L g433 ( .A(n_275), .B(n_357), .Y(n_433) );
INVxp67_ASAP7_75t_L g457 ( .A(n_275), .Y(n_457) );
INVx2_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
NAND2x1_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_278), .B(n_319), .Y(n_386) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g335 ( .A(n_280), .B(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g448 ( .A(n_281), .Y(n_448) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g477 ( .A(n_282), .B(n_310), .Y(n_477) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g403 ( .A(n_283), .B(n_310), .Y(n_403) );
AOI21x1_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_285), .B(n_286), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_294), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_293), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_290), .B(n_326), .Y(n_440) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVx2_ASAP7_75t_L g304 ( .A(n_291), .Y(n_304) );
AND2x2_ASAP7_75t_L g354 ( .A(n_291), .B(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_291), .B(n_348), .Y(n_397) );
OR2x2_ASAP7_75t_L g469 ( .A(n_291), .B(n_356), .Y(n_469) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g389 ( .A(n_295), .B(n_390), .Y(n_389) );
AND2x4_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx2_ASAP7_75t_L g380 ( .A(n_296), .Y(n_380) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g370 ( .A(n_299), .B(n_371), .Y(n_370) );
INVxp67_ASAP7_75t_SL g381 ( .A(n_299), .Y(n_381) );
OR2x2_ASAP7_75t_L g432 ( .A(n_299), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g487 ( .A(n_299), .Y(n_487) );
AOI211xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_305), .B(n_311), .C(n_320), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g376 ( .A(n_304), .B(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_304), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g449 ( .A(n_304), .B(n_326), .Y(n_449) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_307), .B(n_352), .Y(n_374) );
NAND2x1p5_ASAP7_75t_L g391 ( .A(n_307), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g459 ( .A(n_307), .B(n_460), .Y(n_459) );
INVx3_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx2_ASAP7_75t_L g402 ( .A(n_308), .Y(n_402) );
AND2x2_ASAP7_75t_L g430 ( .A(n_309), .B(n_358), .Y(n_430) );
INVx2_ASAP7_75t_L g453 ( .A(n_309), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_309), .B(n_351), .Y(n_485) );
AND2x4_ASAP7_75t_SL g439 ( .A(n_312), .B(n_317), .Y(n_439) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g392 ( .A(n_313), .B(n_318), .Y(n_392) );
OR2x2_ASAP7_75t_L g444 ( .A(n_313), .B(n_337), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_314), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_314), .B(n_326), .Y(n_480) );
BUFx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g428 ( .A(n_315), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
INVx1_ASAP7_75t_L g411 ( .A(n_317), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_317), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g461 ( .A(n_318), .Y(n_461) );
BUFx2_ASAP7_75t_L g329 ( .A(n_319), .Y(n_329) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g447 ( .A(n_322), .B(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g371 ( .A(n_326), .Y(n_371) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_326), .Y(n_388) );
NAND3xp33_ASAP7_75t_SL g327 ( .A(n_328), .B(n_338), .C(n_353), .Y(n_327) );
AOI22xp33_ASAP7_75t_SL g328 ( .A1(n_329), .A2(n_330), .B1(n_333), .B2(n_335), .Y(n_328) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AOI222xp33_ASAP7_75t_L g441 ( .A1(n_335), .A2(n_361), .B1(n_442), .B2(n_445), .C1(n_447), .C2(n_449), .Y(n_441) );
AND2x2_ASAP7_75t_L g473 ( .A(n_336), .B(n_422), .Y(n_473) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g421 ( .A(n_337), .B(n_422), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_344), .B1(n_345), .B2(n_350), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx2_ASAP7_75t_SL g417 ( .A(n_341), .Y(n_417) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_349), .Y(n_345) );
AND2x2_ASAP7_75t_L g404 ( .A(n_346), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g362 ( .A(n_347), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g356 ( .A(n_348), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g471 ( .A(n_349), .Y(n_471) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_352), .B(n_448), .Y(n_467) );
INVx1_ASAP7_75t_L g484 ( .A(n_352), .Y(n_484) );
AOI222xp33_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_358), .B1(n_359), .B2(n_361), .C1(n_364), .C2(n_365), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_360), .Y(n_364) );
AND2x2_ASAP7_75t_L g382 ( .A(n_360), .B(n_383), .Y(n_382) );
INVx3_ASAP7_75t_L g413 ( .A(n_360), .Y(n_413) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g377 ( .A(n_363), .Y(n_377) );
OR2x2_ASAP7_75t_L g446 ( .A(n_363), .B(n_427), .Y(n_446) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
OAI211xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_372), .B(n_375), .C(n_384), .Y(n_369) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OAI21xp33_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_378), .B(n_382), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g462 ( .A1(n_376), .A2(n_414), .B1(n_463), .B2(n_466), .C(n_468), .Y(n_462) );
AND2x4_ASAP7_75t_L g405 ( .A(n_377), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
INVx1_ASAP7_75t_L g436 ( .A(n_383), .Y(n_436) );
AOI211x1_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_387), .B(n_389), .C(n_393), .Y(n_384) );
INVxp67_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g454 ( .A(n_392), .Y(n_454) );
NAND3xp33_ASAP7_75t_L g442 ( .A(n_395), .B(n_443), .C(n_444), .Y(n_442) );
OR2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
INVx1_ASAP7_75t_L g478 ( .A(n_396), .Y(n_478) );
NOR2x1_ASAP7_75t_L g398 ( .A(n_399), .B(n_450), .Y(n_398) );
NAND4xp25_ASAP7_75t_L g399 ( .A(n_400), .B(n_407), .C(n_429), .D(n_441), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_404), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
AND2x2_ASAP7_75t_L g460 ( .A(n_403), .B(n_461), .Y(n_460) );
AOI221x1_ASAP7_75t_L g429 ( .A1(n_405), .A2(n_430), .B1(n_431), .B2(n_434), .C(n_437), .Y(n_429) );
AND2x2_ASAP7_75t_L g455 ( .A(n_405), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g465 ( .A(n_406), .Y(n_465) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_410), .B1(n_414), .B2(n_418), .C(n_420), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_412), .B(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_417), .A2(n_421), .B1(n_424), .B2(n_426), .Y(n_420) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AOI21xp5_ASAP7_75t_L g437 ( .A1(n_421), .A2(n_438), .B(n_440), .Y(n_437) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g443 ( .A(n_423), .Y(n_443) );
OR2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVxp67_ASAP7_75t_L g464 ( .A(n_433), .Y(n_464) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OAI22xp33_ASAP7_75t_L g483 ( .A1(n_446), .A2(n_484), .B1(n_485), .B2(n_486), .Y(n_483) );
NAND3xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_462), .C(n_474), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_455), .B1(n_458), .B2(n_459), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
INVxp67_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g470 ( .A(n_457), .B(n_471), .Y(n_470) );
NAND2x1_ASAP7_75t_L g486 ( .A(n_457), .B(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
INVx2_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_470), .B(n_472), .Y(n_468) );
INVx1_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
AOI221xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_478), .B1(n_479), .B2(n_481), .C(n_483), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx3_ASAP7_75t_R g481 ( .A(n_482), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_488), .B(n_494), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
INVx4_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx3_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_495), .Y(n_494) );
BUFx10_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_506), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx5_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OAI22xp33_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_832), .B1(n_835), .B2(n_836), .Y(n_506) );
INVx1_ASAP7_75t_L g835 ( .A(n_507), .Y(n_835) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_715), .Y(n_508) );
AND4x1_ASAP7_75t_L g509 ( .A(n_510), .B(n_624), .C(n_662), .D(n_700), .Y(n_509) );
NOR2x1_ASAP7_75t_L g510 ( .A(n_511), .B(n_602), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_550), .B(n_561), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x4_ASAP7_75t_L g513 ( .A(n_514), .B(n_522), .Y(n_513) );
NAND2xp5_ASAP7_75t_R g673 ( .A(n_514), .B(n_621), .Y(n_673) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g774 ( .A(n_516), .B(n_652), .Y(n_774) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
OR2x2_ASAP7_75t_L g552 ( .A(n_517), .B(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g635 ( .A(n_517), .Y(n_635) );
AND2x2_ASAP7_75t_L g649 ( .A(n_517), .B(n_553), .Y(n_649) );
OAI21x1_ASAP7_75t_L g526 ( .A1(n_521), .A2(n_527), .B(n_532), .Y(n_526) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_537), .Y(n_522) );
BUFx2_ASAP7_75t_L g551 ( .A(n_523), .Y(n_551) );
AND2x2_ASAP7_75t_L g607 ( .A(n_523), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g622 ( .A(n_523), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_523), .B(n_553), .Y(n_639) );
INVx3_ASAP7_75t_L g652 ( .A(n_523), .Y(n_652) );
AND2x2_ASAP7_75t_L g687 ( .A(n_523), .B(n_609), .Y(n_687) );
INVx2_ASAP7_75t_L g699 ( .A(n_523), .Y(n_699) );
INVx1_ASAP7_75t_L g703 ( .A(n_523), .Y(n_703) );
INVxp67_ASAP7_75t_L g740 ( .A(n_523), .Y(n_740) );
OR2x2_ASAP7_75t_L g753 ( .A(n_523), .B(n_636), .Y(n_753) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
OAI21x1_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_526), .B(n_536), .Y(n_524) );
OAI21xp5_ASAP7_75t_L g580 ( .A1(n_531), .A2(n_581), .B(n_583), .Y(n_580) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g605 ( .A(n_538), .Y(n_605) );
INVx1_ASAP7_75t_L g692 ( .A(n_538), .Y(n_692) );
AND2x2_ASAP7_75t_L g707 ( .A(n_538), .B(n_553), .Y(n_707) );
INVx1_ASAP7_75t_L g722 ( .A(n_538), .Y(n_722) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g636 ( .A(n_539), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_542), .B(n_545), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_550), .A2(n_811), .B1(n_813), .B2(n_815), .Y(n_810) );
OR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_551), .B(n_691), .Y(n_768) );
BUFx2_ASAP7_75t_L g782 ( .A(n_551), .Y(n_782) );
AND2x2_ASAP7_75t_L g800 ( .A(n_551), .B(n_656), .Y(n_800) );
INVx2_ASAP7_75t_L g682 ( .A(n_552), .Y(n_682) );
OR2x2_ASAP7_75t_L g698 ( .A(n_552), .B(n_699), .Y(n_698) );
INVx3_ASAP7_75t_L g606 ( .A(n_553), .Y(n_606) );
AND2x2_ASAP7_75t_L g691 ( .A(n_553), .B(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_585), .Y(n_561) );
OR2x2_ASAP7_75t_L g747 ( .A(n_562), .B(n_704), .Y(n_747) );
OR2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_574), .Y(n_562) );
AND2x2_ASAP7_75t_L g618 ( .A(n_563), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g659 ( .A(n_563), .Y(n_659) );
INVx2_ASAP7_75t_SL g667 ( .A(n_563), .Y(n_667) );
BUFx2_ASAP7_75t_L g679 ( .A(n_563), .Y(n_679) );
OR2x2_ASAP7_75t_L g767 ( .A(n_563), .B(n_587), .Y(n_767) );
OA21x2_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_565), .B(n_573), .Y(n_563) );
OA21x2_ASAP7_75t_L g632 ( .A1(n_564), .A2(n_565), .B(n_573), .Y(n_632) );
AND2x2_ASAP7_75t_L g611 ( .A(n_574), .B(n_594), .Y(n_611) );
AND2x2_ASAP7_75t_L g647 ( .A(n_574), .B(n_632), .Y(n_647) );
OAI21xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .B(n_584), .Y(n_574) );
OAI21x1_ASAP7_75t_L g617 ( .A1(n_575), .A2(n_576), .B(n_584), .Y(n_617) );
INVx1_ASAP7_75t_L g685 ( .A(n_585), .Y(n_685) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_586), .B(n_679), .Y(n_678) );
AND2x4_ASAP7_75t_L g791 ( .A(n_586), .B(n_771), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_586), .B(n_614), .Y(n_815) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_594), .Y(n_586) );
INVx1_ASAP7_75t_L g619 ( .A(n_587), .Y(n_619) );
INVx2_ASAP7_75t_L g629 ( .A(n_587), .Y(n_629) );
AND2x2_ASAP7_75t_L g643 ( .A(n_587), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g658 ( .A(n_587), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g672 ( .A(n_587), .B(n_632), .Y(n_672) );
OR2x2_ASAP7_75t_L g704 ( .A(n_587), .B(n_644), .Y(n_704) );
INVx1_ASAP7_75t_L g788 ( .A(n_587), .Y(n_788) );
AND2x2_ASAP7_75t_L g631 ( .A(n_594), .B(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g669 ( .A(n_594), .Y(n_669) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g645 ( .A(n_595), .Y(n_645) );
CKINVDCx5p33_ASAP7_75t_R g600 ( .A(n_601), .Y(n_600) );
OAI22xp33_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_610), .B1(n_612), .B2(n_620), .Y(n_602) );
NAND2x1p5_ASAP7_75t_L g603 ( .A(n_604), .B(n_607), .Y(n_603) );
AND2x4_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx1_ASAP7_75t_L g749 ( .A(n_605), .Y(n_749) );
INVx1_ASAP7_75t_L g623 ( .A(n_606), .Y(n_623) );
AND2x4_ASAP7_75t_L g656 ( .A(n_606), .B(n_609), .Y(n_656) );
AND2x2_ASAP7_75t_L g765 ( .A(n_606), .B(n_636), .Y(n_765) );
AND2x2_ASAP7_75t_L g817 ( .A(n_607), .B(n_691), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_607), .B(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVxp67_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g671 ( .A(n_611), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g804 ( .A(n_611), .B(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_618), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_614), .B(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g723 ( .A(n_614), .Y(n_723) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g789 ( .A(n_615), .Y(n_789) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g676 ( .A(n_616), .Y(n_676) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g661 ( .A(n_617), .B(n_645), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_618), .B(n_660), .Y(n_776) );
AND2x2_ASAP7_75t_L g668 ( .A(n_619), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx1_ASAP7_75t_L g808 ( .A(n_623), .Y(n_808) );
AOI221xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_633), .B1(n_640), .B2(n_648), .C(n_653), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_630), .Y(n_626) );
AND2x2_ASAP7_75t_L g726 ( .A(n_627), .B(n_647), .Y(n_726) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_628), .B(n_647), .Y(n_695) );
OR2x2_ASAP7_75t_L g710 ( .A(n_628), .B(n_661), .Y(n_710) );
INVx2_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g675 ( .A(n_629), .B(n_676), .Y(n_675) );
INVxp67_ASAP7_75t_L g786 ( .A(n_631), .Y(n_786) );
INVx1_ASAP7_75t_L g746 ( .A(n_632), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_637), .Y(n_633) );
AND2x2_ASAP7_75t_L g806 ( .A(n_634), .B(n_807), .Y(n_806) );
OR2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
AND2x2_ASAP7_75t_L g760 ( .A(n_635), .B(n_722), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_636), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g681 ( .A(n_636), .Y(n_681) );
INVx1_ASAP7_75t_L g733 ( .A(n_636), .Y(n_733) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OAI21xp33_ASAP7_75t_L g701 ( .A1(n_641), .A2(n_667), .B(n_702), .Y(n_701) );
OR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_646), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g696 ( .A(n_643), .B(n_679), .Y(n_696) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_643), .Y(n_736) );
AND2x2_ASAP7_75t_L g820 ( .A(n_643), .B(n_757), .Y(n_820) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g827 ( .A(n_646), .B(n_744), .Y(n_827) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
INVx2_ASAP7_75t_SL g728 ( .A(n_649), .Y(n_728) );
AND2x2_ASAP7_75t_L g732 ( .A(n_649), .B(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g792 ( .A(n_649), .B(n_652), .Y(n_792) );
AND2x2_ASAP7_75t_L g814 ( .A(n_649), .B(n_739), .Y(n_814) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g711 ( .A(n_652), .B(n_656), .Y(n_711) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_655), .B(n_657), .Y(n_654) );
BUFx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AND2x4_ASAP7_75t_L g705 ( .A(n_656), .B(n_681), .Y(n_705) );
AND2x2_ASAP7_75t_L g738 ( .A(n_656), .B(n_739), .Y(n_738) );
INVx3_ASAP7_75t_L g755 ( .A(n_656), .Y(n_755) );
INVx1_ASAP7_75t_L g824 ( .A(n_657), .Y(n_824) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_660), .Y(n_657) );
AND2x4_ASAP7_75t_L g688 ( .A(n_658), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g730 ( .A(n_660), .B(n_679), .Y(n_730) );
AND2x2_ASAP7_75t_L g756 ( .A(n_660), .B(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OR2x2_ASAP7_75t_L g766 ( .A(n_661), .B(n_767), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_663), .B(n_683), .Y(n_662) );
A2O1A1Ixp33_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_670), .B(n_673), .C(n_674), .Y(n_663) );
INVx2_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_668), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_666), .B(n_812), .Y(n_811) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_667), .B(n_714), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_667), .B(n_736), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_668), .B(n_771), .Y(n_770) );
AND2x2_ASAP7_75t_L g689 ( .A(n_669), .B(n_676), .Y(n_689) );
INVx1_ASAP7_75t_L g744 ( .A(n_669), .Y(n_744) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OAI21xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_677), .B(n_680), .Y(n_674) );
NAND2x1p5_ASAP7_75t_L g745 ( .A(n_676), .B(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g757 ( .A(n_679), .Y(n_757) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
AND2x4_ASAP7_75t_L g781 ( .A(n_682), .B(n_749), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_693), .Y(n_683) );
A2O1A1Ixp33_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_686), .B(n_688), .C(n_690), .Y(n_684) );
BUFx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g748 ( .A(n_687), .B(n_749), .Y(n_748) );
BUFx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
OAI21xp5_ASAP7_75t_SL g693 ( .A1(n_694), .A2(n_696), .B(n_697), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_699), .Y(n_708) );
OR2x2_ASAP7_75t_L g727 ( .A(n_699), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g809 ( .A(n_699), .Y(n_809) );
AOI222xp33_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_705), .B1(n_706), .B2(n_709), .C1(n_711), .C2(n_712), .Y(n_700) );
NOR2x1_ASAP7_75t_L g718 ( .A(n_702), .B(n_719), .Y(n_718) );
OR2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
NAND2x1p5_ASAP7_75t_L g759 ( .A(n_703), .B(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g714 ( .A(n_704), .Y(n_714) );
INVx1_ASAP7_75t_L g812 ( .A(n_704), .Y(n_812) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_707), .B(n_773), .Y(n_772) );
BUFx2_ASAP7_75t_L g790 ( .A(n_707), .Y(n_790) );
AND2x4_ASAP7_75t_L g797 ( .A(n_707), .B(n_774), .Y(n_797) );
INVx2_ASAP7_75t_L g826 ( .A(n_707), .Y(n_826) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
OAI22xp33_ASAP7_75t_L g762 ( .A1(n_710), .A2(n_763), .B1(n_766), .B2(n_768), .Y(n_762) );
AOI211xp5_ASAP7_75t_L g816 ( .A1(n_712), .A2(n_817), .B(n_818), .C(n_822), .Y(n_816) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NOR2xp67_ASAP7_75t_SL g715 ( .A(n_716), .B(n_777), .Y(n_715) );
NAND4xp25_ASAP7_75t_L g716 ( .A(n_717), .B(n_734), .C(n_741), .D(n_761), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_723), .B(n_724), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_727), .B1(n_729), .B2(n_731), .Y(n_724) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_728), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_729), .B(n_795), .Y(n_794) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g739 ( .A(n_733), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_737), .Y(n_734) );
AND2x2_ASAP7_75t_L g737 ( .A(n_738), .B(n_740), .Y(n_737) );
INVx1_ASAP7_75t_L g764 ( .A(n_740), .Y(n_764) );
AOI221xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_748), .B1(n_750), .B2(n_756), .C(n_758), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_747), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_743), .B(n_759), .Y(n_758) );
OR2x2_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
AND2x2_ASAP7_75t_L g796 ( .A(n_744), .B(n_771), .Y(n_796) );
INVx2_ASAP7_75t_L g771 ( .A(n_745), .Y(n_771) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
NAND2x1_ASAP7_75t_SL g751 ( .A(n_752), .B(n_754), .Y(n_751) );
INVx1_ASAP7_75t_L g821 ( .A(n_752), .Y(n_821) );
INVx3_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g823 ( .A(n_760), .Y(n_823) );
NOR2xp33_ASAP7_75t_L g761 ( .A(n_762), .B(n_769), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
INVx1_ASAP7_75t_L g805 ( .A(n_767), .Y(n_805) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_772), .B1(n_775), .B2(n_776), .Y(n_769) );
AND2x2_ASAP7_75t_L g802 ( .A(n_771), .B(n_788), .Y(n_802) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g783 ( .A(n_776), .Y(n_783) );
NAND3xp33_ASAP7_75t_L g777 ( .A(n_778), .B(n_793), .C(n_816), .Y(n_777) );
AOI222xp33_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_783), .B1(n_784), .B2(n_790), .C1(n_791), .C2(n_792), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_780), .B(n_782), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
OR2x2_ASAP7_75t_L g785 ( .A(n_786), .B(n_787), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_789), .Y(n_787) );
AOI211xp5_ASAP7_75t_L g793 ( .A1(n_794), .A2(n_797), .B(n_798), .C(n_810), .Y(n_793) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_801), .B1(n_803), .B2(n_806), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .Y(n_807) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_819), .B(n_821), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_823), .A2(n_824), .B1(n_825), .B2(n_827), .Y(n_822) );
INVx4_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_SL g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g836 ( .A(n_832), .Y(n_836) );
NOR2xp33_ASAP7_75t_L g837 ( .A(n_838), .B(n_839), .Y(n_837) );
endmodule