module real_aes_12544_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_656;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_617;
wire n_139;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_686;
wire n_79;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
OA21x2_ASAP7_75t_L g110 ( .A1(n_0), .A2(n_43), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g187 ( .A(n_0), .Y(n_187) );
OAI222xp33_ASAP7_75t_L g600 ( .A1(n_1), .A2(n_65), .B1(n_71), .B2(n_601), .C1(n_607), .C2(n_608), .Y(n_600) );
INVx1_ASAP7_75t_L g618 ( .A(n_1), .Y(n_618) );
AND2x2_ASAP7_75t_L g141 ( .A(n_2), .B(n_142), .Y(n_141) );
AOI221xp5_ASAP7_75t_L g180 ( .A1(n_3), .A2(n_72), .B1(n_89), .B2(n_165), .C(n_181), .Y(n_180) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_3), .A2(n_705), .B1(n_706), .B2(n_707), .Y(n_704) );
INVx1_ASAP7_75t_L g707 ( .A(n_3), .Y(n_707) );
BUFx3_ASAP7_75t_L g522 ( .A(n_4), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_5), .A2(n_710), .B1(n_711), .B2(n_712), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_5), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_6), .B(n_148), .Y(n_268) );
INVx3_ASAP7_75t_L g519 ( .A(n_7), .Y(n_519) );
INVx2_ASAP7_75t_L g529 ( .A(n_8), .Y(n_529) );
INVx1_ASAP7_75t_L g547 ( .A(n_8), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_9), .A2(n_700), .B1(n_701), .B2(n_702), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_9), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_10), .B(n_115), .Y(n_168) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_10), .A2(n_512), .B1(n_738), .B2(n_741), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_11), .B(n_259), .Y(n_258) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_12), .Y(n_706) );
INVx1_ASAP7_75t_L g95 ( .A(n_13), .Y(n_95) );
BUFx3_ASAP7_75t_L g117 ( .A(n_13), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_14), .B(n_127), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_15), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_16), .A2(n_75), .B1(n_541), .B2(n_542), .Y(n_540) );
OAI321xp33_ASAP7_75t_L g616 ( .A1(n_16), .A2(n_617), .A3(n_626), .B1(n_638), .B2(n_642), .C(n_648), .Y(n_616) );
BUFx10_ASAP7_75t_L g725 ( .A(n_17), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_18), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_19), .B(n_133), .Y(n_213) );
OAI21xp33_ASAP7_75t_L g296 ( .A1(n_19), .A2(n_53), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g597 ( .A(n_20), .Y(n_597) );
OAI211xp5_ASAP7_75t_L g514 ( .A1(n_21), .A2(n_515), .B(n_537), .C(n_615), .Y(n_514) );
O2A1O1Ixp5_ASAP7_75t_L g182 ( .A1(n_22), .A2(n_170), .B(n_172), .C(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g564 ( .A(n_23), .Y(n_564) );
OAI322xp33_ASAP7_75t_L g651 ( .A1(n_23), .A2(n_71), .A3(n_652), .B1(n_656), .B2(n_664), .C1(n_670), .C2(n_675), .Y(n_651) );
AND2x2_ASAP7_75t_L g536 ( .A(n_24), .B(n_30), .Y(n_536) );
INVx1_ASAP7_75t_L g641 ( .A(n_24), .Y(n_641) );
AND2x2_ASAP7_75t_L g645 ( .A(n_24), .B(n_646), .Y(n_645) );
INVxp33_ASAP7_75t_L g669 ( .A(n_24), .Y(n_669) );
INVx1_ASAP7_75t_L g86 ( .A(n_25), .Y(n_86) );
INVx2_ASAP7_75t_L g534 ( .A(n_26), .Y(n_534) );
INVx1_ASAP7_75t_L g586 ( .A(n_27), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_28), .B(n_120), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_29), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_30), .B(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g646 ( .A(n_30), .Y(n_646) );
INVx1_ASAP7_75t_L g571 ( .A(n_31), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_32), .B(n_127), .Y(n_126) );
AND2x4_ASAP7_75t_L g85 ( .A(n_33), .B(n_86), .Y(n_85) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_33), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g548 ( .A1(n_34), .A2(n_47), .B1(n_549), .B2(n_553), .C(n_559), .Y(n_548) );
INVx1_ASAP7_75t_L g661 ( .A(n_34), .Y(n_661) );
NAND2x1_ASAP7_75t_L g267 ( .A(n_35), .B(n_142), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_36), .Y(n_223) );
INVx1_ASAP7_75t_L g264 ( .A(n_37), .Y(n_264) );
INVx1_ASAP7_75t_L g527 ( .A(n_38), .Y(n_527) );
INVx1_ASAP7_75t_L g552 ( .A(n_38), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_39), .Y(n_237) );
AOI221xp5_ASAP7_75t_L g587 ( .A1(n_40), .A2(n_70), .B1(n_588), .B2(n_589), .C(n_590), .Y(n_587) );
OAI222xp33_ASAP7_75t_L g682 ( .A1(n_40), .A2(n_47), .B1(n_70), .B2(n_683), .C1(n_686), .C2(n_688), .Y(n_682) );
AND2x2_ASAP7_75t_L g140 ( .A(n_41), .B(n_125), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_42), .B(n_119), .Y(n_198) );
INVx1_ASAP7_75t_L g186 ( .A(n_43), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_44), .B(n_148), .Y(n_247) );
INVx1_ASAP7_75t_L g111 ( .A(n_45), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_46), .B(n_125), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_48), .B(n_133), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_49), .B(n_201), .Y(n_266) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_49), .Y(n_701) );
NAND2xp5_ASAP7_75t_SL g118 ( .A(n_50), .B(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_51), .B(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g147 ( .A(n_52), .B(n_148), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_53), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_54), .B(n_170), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_54), .A2(n_697), .B1(n_715), .B2(n_731), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_54), .A2(n_697), .B1(n_739), .B2(n_740), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_55), .B(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_56), .B(n_119), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_57), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_58), .B(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_59), .B(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_60), .B(n_134), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g124 ( .A(n_61), .B(n_125), .Y(n_124) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_62), .A2(n_69), .B1(n_713), .B2(n_714), .Y(n_712) );
CKINVDCx5p33_ASAP7_75t_R g714 ( .A(n_62), .Y(n_714) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_63), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_64), .B(n_164), .Y(n_206) );
INVx1_ASAP7_75t_L g627 ( .A(n_65), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_66), .B(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g90 ( .A(n_67), .Y(n_90) );
BUFx3_ASAP7_75t_L g130 ( .A(n_67), .Y(n_130) );
INVx1_ASAP7_75t_L g145 ( .A(n_67), .Y(n_145) );
INVx2_ASAP7_75t_L g533 ( .A(n_68), .Y(n_533) );
AND2x2_ASAP7_75t_L g632 ( .A(n_68), .B(n_534), .Y(n_632) );
INVxp67_ASAP7_75t_SL g680 ( .A(n_68), .Y(n_680) );
INVx1_ASAP7_75t_L g713 ( .A(n_69), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_73), .B(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g521 ( .A(n_74), .Y(n_521) );
INVx1_ASAP7_75t_L g655 ( .A(n_75), .Y(n_655) );
INVx1_ASAP7_75t_L g583 ( .A(n_76), .Y(n_583) );
XNOR2xp5_ASAP7_75t_L g511 ( .A(n_77), .B(n_512), .Y(n_511) );
AOI21xp33_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_96), .B(n_510), .Y(n_78) );
BUFx6f_ASAP7_75t_L g79 ( .A(n_80), .Y(n_79) );
NOR2xp33_ASAP7_75t_L g80 ( .A(n_81), .B(n_87), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
BUFx2_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
BUFx6f_ASAP7_75t_SL g131 ( .A(n_85), .Y(n_131) );
INVx3_ASAP7_75t_L g156 ( .A(n_85), .Y(n_156) );
INVx2_ASAP7_75t_L g208 ( .A(n_85), .Y(n_208) );
INVx1_ASAP7_75t_L g228 ( .A(n_85), .Y(n_228) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_86), .Y(n_693) );
AO21x2_ASAP7_75t_L g743 ( .A1(n_87), .A2(n_692), .B(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g87 ( .A(n_88), .B(n_91), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g226 ( .A(n_89), .Y(n_226) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_89), .A2(n_233), .B1(n_235), .B2(n_239), .Y(n_232) );
INVx2_ASAP7_75t_SL g238 ( .A(n_89), .Y(n_238) );
BUFx3_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx1_ASAP7_75t_L g122 ( .A(n_90), .Y(n_122) );
HB1xp67_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_93), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx2_ASAP7_75t_L g125 ( .A(n_94), .Y(n_125) );
INVx2_ASAP7_75t_L g170 ( .A(n_94), .Y(n_170) );
INVx2_ASAP7_75t_L g222 ( .A(n_94), .Y(n_222) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx2_ASAP7_75t_L g166 ( .A(n_95), .Y(n_166) );
INVx4_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
AND2x4_ASAP7_75t_L g97 ( .A(n_98), .B(n_391), .Y(n_97) );
NOR4xp75_ASAP7_75t_L g98 ( .A(n_99), .B(n_313), .C(n_344), .D(n_372), .Y(n_98) );
OAI211xp5_ASAP7_75t_SL g99 ( .A1(n_100), .A2(n_175), .B(n_248), .C(n_277), .Y(n_99) );
INVxp67_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
AND2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_136), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_103), .B(n_450), .Y(n_468) );
NOR2xp67_ASAP7_75t_L g502 ( .A(n_103), .B(n_306), .Y(n_502) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_L g249 ( .A(n_104), .B(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g288 ( .A(n_104), .Y(n_288) );
INVx1_ASAP7_75t_L g309 ( .A(n_104), .Y(n_309) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_104), .Y(n_320) );
AND2x2_ASAP7_75t_L g416 ( .A(n_104), .B(n_417), .Y(n_416) );
INVx3_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AND2x2_ASAP7_75t_L g333 ( .A(n_105), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g389 ( .A(n_105), .B(n_307), .Y(n_389) );
AND2x2_ASAP7_75t_L g440 ( .A(n_105), .B(n_252), .Y(n_440) );
BUFx3_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g342 ( .A(n_106), .Y(n_342) );
OAI21x1_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_112), .B(n_132), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx3_ASAP7_75t_L g297 ( .A(n_109), .Y(n_297) );
BUFx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g135 ( .A(n_110), .Y(n_135) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_110), .Y(n_148) );
INVx1_ASAP7_75t_L g188 ( .A(n_111), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_123), .B(n_131), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_118), .B(n_121), .Y(n_113) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_116), .B(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g224 ( .A(n_116), .Y(n_224) );
INVx1_ASAP7_75t_L g234 ( .A(n_116), .Y(n_234) );
INVx2_ASAP7_75t_L g243 ( .A(n_116), .Y(n_243) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g120 ( .A(n_117), .Y(n_120) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_117), .Y(n_128) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g162 ( .A(n_120), .Y(n_162) );
INVx2_ASAP7_75t_L g201 ( .A(n_120), .Y(n_201) );
INVx2_ASAP7_75t_L g218 ( .A(n_120), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_121), .A2(n_161), .B(n_163), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_121), .A2(n_204), .B(n_206), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_121), .A2(n_241), .B(n_244), .Y(n_240) );
BUFx10_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_126), .B(n_129), .Y(n_123) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx3_ASAP7_75t_L g142 ( .A(n_128), .Y(n_142) );
INVx3_ASAP7_75t_L g261 ( .A(n_128), .Y(n_261) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g220 ( .A(n_130), .Y(n_220) );
INVx2_ASAP7_75t_L g259 ( .A(n_130), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_130), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g174 ( .A(n_131), .Y(n_174) );
OAI21x1_ASAP7_75t_L g256 ( .A1(n_131), .A2(n_257), .B(n_265), .Y(n_256) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_134), .B(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g406 ( .A(n_136), .B(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g335 ( .A(n_137), .Y(n_335) );
INVx2_ASAP7_75t_L g343 ( .A(n_137), .Y(n_343) );
AND2x2_ASAP7_75t_L g439 ( .A(n_137), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g493 ( .A(n_137), .Y(n_493) );
OR2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_157), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_138), .B(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_138), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g303 ( .A(n_138), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g307 ( .A(n_138), .Y(n_307) );
INVx2_ASAP7_75t_L g323 ( .A(n_138), .Y(n_323) );
AO21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_146), .B(n_153), .Y(n_138) );
OAI21xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_141), .B(n_143), .Y(n_139) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g152 ( .A(n_144), .Y(n_152) );
BUFx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g172 ( .A(n_145), .Y(n_172) );
NOR2xp67_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
AOI21xp33_ASAP7_75t_L g153 ( .A1(n_147), .A2(n_154), .B(n_155), .Y(n_153) );
INVxp33_ASAP7_75t_L g154 ( .A(n_148), .Y(n_154) );
INVx1_ASAP7_75t_L g191 ( .A(n_148), .Y(n_191) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_148), .Y(n_195) );
INVx1_ASAP7_75t_L g255 ( .A(n_148), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_152), .Y(n_149) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NOR3xp33_ASAP7_75t_L g179 ( .A(n_156), .B(n_180), .C(n_182), .Y(n_179) );
INVx3_ASAP7_75t_L g304 ( .A(n_157), .Y(n_304) );
INVx1_ASAP7_75t_L g318 ( .A(n_157), .Y(n_318) );
AND2x2_ASAP7_75t_L g322 ( .A(n_157), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g417 ( .A(n_157), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g444 ( .A(n_157), .Y(n_444) );
AND2x4_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
OAI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_167), .B(n_173), .Y(n_159) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx3_ASAP7_75t_L g181 ( .A(n_166), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_171), .Y(n_167) );
AOI21x1_ASAP7_75t_L g265 ( .A1(n_171), .A2(n_266), .B(n_267), .Y(n_265) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g202 ( .A(n_172), .Y(n_202) );
INVx2_ASAP7_75t_SL g175 ( .A(n_176), .Y(n_175) );
AOI32xp33_ASAP7_75t_L g365 ( .A1(n_176), .A2(n_366), .A3(n_368), .B1(n_369), .B2(n_371), .Y(n_365) );
AND2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_210), .Y(n_176) );
INVx1_ASAP7_75t_L g349 ( .A(n_177), .Y(n_349) );
AND2x2_ASAP7_75t_L g454 ( .A(n_177), .B(n_272), .Y(n_454) );
AND2x2_ASAP7_75t_L g507 ( .A(n_177), .B(n_281), .Y(n_507) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_192), .Y(n_177) );
INVx2_ASAP7_75t_L g276 ( .A(n_178), .Y(n_276) );
AND2x2_ASAP7_75t_L g279 ( .A(n_178), .B(n_280), .Y(n_279) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_178), .Y(n_476) );
AO21x2_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_185), .B(n_189), .Y(n_178) );
NAND2xp33_ASAP7_75t_L g298 ( .A(n_179), .B(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g205 ( .A(n_181), .Y(n_205) );
AO21x2_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_188), .Y(n_185) );
AOI21x1_ASAP7_75t_L g229 ( .A1(n_186), .A2(n_187), .B(n_188), .Y(n_229) );
NOR2xp33_ASAP7_75t_R g189 ( .A(n_190), .B(n_191), .Y(n_189) );
INVx2_ASAP7_75t_L g275 ( .A(n_192), .Y(n_275) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVxp67_ASAP7_75t_L g400 ( .A(n_193), .Y(n_400) );
OAI21x1_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_196), .B(n_209), .Y(n_193) );
OAI21x1_ASAP7_75t_L g230 ( .A1(n_194), .A2(n_231), .B(n_247), .Y(n_230) );
OAI21xp5_ASAP7_75t_L g280 ( .A1(n_194), .A2(n_196), .B(n_209), .Y(n_280) );
OAI21x1_ASAP7_75t_L g294 ( .A1(n_194), .A2(n_231), .B(n_247), .Y(n_294) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
OAI21x1_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_203), .B(n_207), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_202), .Y(n_197) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_SL g246 ( .A(n_208), .Y(n_246) );
AND2x2_ASAP7_75t_L g385 ( .A(n_210), .B(n_386), .Y(n_385) );
NAND2x1p5_ASAP7_75t_L g423 ( .A(n_210), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g445 ( .A(n_210), .B(n_279), .Y(n_445) );
AND2x4_ASAP7_75t_SL g461 ( .A(n_210), .B(n_274), .Y(n_461) );
AND2x2_ASAP7_75t_L g482 ( .A(n_210), .B(n_311), .Y(n_482) );
AND2x4_ASAP7_75t_L g210 ( .A(n_211), .B(n_230), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g273 ( .A(n_212), .Y(n_273) );
INVx2_ASAP7_75t_L g282 ( .A(n_212), .Y(n_282) );
AND2x2_ASAP7_75t_L g337 ( .A(n_212), .B(n_230), .Y(n_337) );
AND2x2_ASAP7_75t_L g364 ( .A(n_212), .B(n_329), .Y(n_364) );
AND2x4_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
NAND3xp33_ASAP7_75t_L g295 ( .A(n_214), .B(n_296), .C(n_298), .Y(n_295) );
NAND3xp33_ASAP7_75t_L g214 ( .A(n_215), .B(n_221), .C(n_227), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_219), .C(n_220), .Y(n_215) );
INVx2_ASAP7_75t_SL g217 ( .A(n_218), .Y(n_217) );
OAI221xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B1(n_224), .B2(n_225), .C(n_226), .Y(n_221) );
INVx2_ASAP7_75t_L g245 ( .A(n_222), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
INVx2_ASAP7_75t_L g300 ( .A(n_229), .Y(n_300) );
INVx1_ASAP7_75t_L g283 ( .A(n_230), .Y(n_283) );
OAI21x1_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_240), .B(n_246), .Y(n_231) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_238), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_269), .Y(n_248) );
INVxp67_ASAP7_75t_SL g441 ( .A(n_249), .Y(n_441) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g362 ( .A(n_251), .Y(n_362) );
INVx1_ASAP7_75t_L g287 ( .A(n_252), .Y(n_287) );
INVx2_ASAP7_75t_L g334 ( .A(n_252), .Y(n_334) );
INVx1_ASAP7_75t_L g359 ( .A(n_252), .Y(n_359) );
AND2x2_ASAP7_75t_L g371 ( .A(n_252), .B(n_342), .Y(n_371) );
AND2x4_ASAP7_75t_SL g377 ( .A(n_252), .B(n_323), .Y(n_377) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_252), .Y(n_381) );
INVxp67_ASAP7_75t_L g418 ( .A(n_252), .Y(n_418) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OAI21x1_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_256), .B(n_268), .Y(n_253) );
INVx1_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
OAI21xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_260), .B(n_262), .Y(n_257) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OAI22xp33_ASAP7_75t_L g465 ( .A1(n_270), .A2(n_466), .B1(n_468), .B2(n_469), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_274), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_272), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_272), .B(n_348), .Y(n_489) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g352 ( .A(n_274), .Y(n_352) );
AND2x2_ASAP7_75t_L g390 ( .A(n_274), .B(n_281), .Y(n_390) );
AND2x2_ASAP7_75t_L g509 ( .A(n_274), .B(n_293), .Y(n_509) );
AND2x4_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx2_ASAP7_75t_L g290 ( .A(n_275), .Y(n_290) );
AND2x2_ASAP7_75t_L g311 ( .A(n_276), .B(n_312), .Y(n_311) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_276), .Y(n_495) );
AOI222xp33_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_284), .B1(n_289), .B2(n_301), .C1(n_305), .C2(n_310), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
AND2x2_ASAP7_75t_L g336 ( .A(n_279), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g363 ( .A(n_279), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g368 ( .A(n_279), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_279), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g470 ( .A(n_279), .B(n_414), .Y(n_470) );
INVx1_ASAP7_75t_L g312 ( .A(n_280), .Y(n_312) );
AND2x2_ASAP7_75t_L g353 ( .A(n_281), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g437 ( .A(n_281), .B(n_339), .Y(n_437) );
AND2x2_ASAP7_75t_L g500 ( .A(n_281), .B(n_311), .Y(n_500) );
AND2x4_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx1_ASAP7_75t_L g414 ( .A(n_282), .Y(n_414) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g473 ( .A(n_285), .B(n_351), .Y(n_473) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_287), .Y(n_407) );
NOR2x1p5_ASAP7_75t_SL g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx1_ASAP7_75t_L g424 ( .A(n_290), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_290), .B(n_364), .Y(n_479) );
OAI221xp5_ASAP7_75t_L g436 ( .A1(n_291), .A2(n_437), .B1(n_438), .B2(n_441), .C(n_442), .Y(n_436) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_295), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_293), .B(n_309), .Y(n_308) );
INVxp67_ASAP7_75t_SL g411 ( .A(n_293), .Y(n_411) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_293), .Y(n_422) );
OR2x2_ASAP7_75t_L g490 ( .A(n_293), .B(n_295), .Y(n_490) );
BUFx3_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g329 ( .A(n_294), .Y(n_329) );
INVx1_ASAP7_75t_L g401 ( .A(n_295), .Y(n_401) );
INVx1_ASAP7_75t_L g431 ( .A(n_295), .Y(n_431) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NOR3xp33_ASAP7_75t_L g314 ( .A(n_301), .B(n_315), .C(n_321), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_301), .A2(n_347), .B1(n_350), .B2(n_352), .Y(n_346) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g379 ( .A(n_303), .B(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_303), .B(n_383), .Y(n_421) );
AND2x2_ASAP7_75t_L g434 ( .A(n_303), .B(n_354), .Y(n_434) );
OR2x2_ASAP7_75t_L g306 ( .A(n_304), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g351 ( .A(n_304), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
INVx3_ASAP7_75t_L g450 ( .A(n_306), .Y(n_450) );
INVx1_ASAP7_75t_L g383 ( .A(n_309), .Y(n_383) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x4_ASAP7_75t_L g327 ( .A(n_311), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_311), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g339 ( .A(n_312), .Y(n_339) );
OAI21xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_324), .B(n_330), .Y(n_313) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_319), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g375 ( .A(n_317), .B(n_376), .Y(n_375) );
AND2x4_ASAP7_75t_L g467 ( .A(n_317), .B(n_362), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_317), .B(n_376), .Y(n_503) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g358 ( .A(n_318), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g505 ( .A(n_321), .Y(n_505) );
BUFx3_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g366 ( .A(n_322), .B(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_322), .B(n_333), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_322), .B(n_341), .Y(n_425) );
BUFx2_ASAP7_75t_L g429 ( .A(n_323), .Y(n_429) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_327), .B(n_416), .Y(n_415) );
INVxp67_ASAP7_75t_L g432 ( .A(n_327), .Y(n_432) );
INVx1_ASAP7_75t_L g402 ( .A(n_328), .Y(n_402) );
AND2x2_ASAP7_75t_L g475 ( .A(n_328), .B(n_476), .Y(n_475) );
BUFx3_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AOI22xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_336), .B1(n_338), .B2(n_340), .Y(n_330) );
NOR2x1_ASAP7_75t_L g331 ( .A(n_332), .B(n_335), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g464 ( .A(n_333), .B(n_444), .Y(n_464) );
AND2x2_ASAP7_75t_L g341 ( .A(n_334), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g403 ( .A(n_335), .Y(n_403) );
AND2x2_ASAP7_75t_L g338 ( .A(n_337), .B(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g386 ( .A(n_339), .Y(n_386) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
AND2x2_ASAP7_75t_L g428 ( .A(n_341), .B(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_341), .B(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g491 ( .A(n_341), .Y(n_491) );
INVx2_ASAP7_75t_L g354 ( .A(n_342), .Y(n_354) );
NAND2x1_ASAP7_75t_SL g344 ( .A(n_345), .B(n_365), .Y(n_344) );
AOI22xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_353), .B1(n_355), .B2(n_363), .Y(n_345) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OAI32xp33_ASAP7_75t_L g420 ( .A1(n_352), .A2(n_421), .A3(n_422), .B1(n_423), .B2(n_425), .Y(n_420) );
NOR2x1_ASAP7_75t_L g357 ( .A(n_354), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g367 ( .A(n_354), .Y(n_367) );
AND2x2_ASAP7_75t_L g459 ( .A(n_354), .B(n_377), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g355 ( .A(n_356), .B(n_360), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g388 ( .A(n_359), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g396 ( .A(n_359), .Y(n_396) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx3_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g370 ( .A(n_364), .Y(n_370) );
OAI21xp5_ASAP7_75t_L g442 ( .A1(n_366), .A2(n_443), .B(n_445), .Y(n_442) );
AND2x2_ASAP7_75t_L g488 ( .A(n_367), .B(n_377), .Y(n_488) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OAI21xp33_ASAP7_75t_L g387 ( .A1(n_371), .A2(n_388), .B(n_390), .Y(n_387) );
A2O1A1Ixp33_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_378), .B(n_384), .C(n_387), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2x1_ASAP7_75t_L g378 ( .A(n_379), .B(n_382), .Y(n_378) );
INVx1_ASAP7_75t_L g481 ( .A(n_379), .Y(n_481) );
INVxp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_381), .Y(n_485) );
NAND2x1_ASAP7_75t_L g472 ( .A(n_382), .B(n_467), .Y(n_472) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g448 ( .A(n_388), .Y(n_448) );
NOR2x1_ASAP7_75t_L g391 ( .A(n_392), .B(n_455), .Y(n_391) );
NAND4xp25_ASAP7_75t_L g392 ( .A(n_393), .B(n_419), .C(n_435), .D(n_446), .Y(n_392) );
AOI21xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_403), .B(n_404), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_395), .B(n_397), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g451 ( .A(n_396), .B(n_444), .Y(n_451) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_402), .Y(n_398) );
INVx1_ASAP7_75t_L g462 ( .A(n_399), .Y(n_462) );
AND2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
NAND2x1p5_ASAP7_75t_L g453 ( .A(n_402), .B(n_454), .Y(n_453) );
OAI21xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_408), .B(n_415), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_412), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_411), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_420), .B(n_426), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_430), .B1(n_432), .B2(n_433), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g443 ( .A(n_440), .B(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g497 ( .A(n_440), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_451), .B(n_452), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
AND2x4_ASAP7_75t_L g483 ( .A(n_450), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AOI221xp5_ASAP7_75t_L g498 ( .A1(n_454), .A2(n_499), .B1(n_501), .B2(n_503), .C(n_504), .Y(n_498) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_477), .C(n_498), .Y(n_455) );
NOR3xp33_ASAP7_75t_SL g456 ( .A(n_457), .B(n_465), .C(n_471), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_460), .B1(n_462), .B2(n_463), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_463), .A2(n_505), .B1(n_506), .B2(n_508), .Y(n_504) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B(n_474), .Y(n_471) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_480), .B1(n_482), .B2(n_483), .C(n_486), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVxp67_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OAI221xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_489), .B1(n_490), .B2(n_491), .C(n_492), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND3xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .C(n_496), .Y(n_492) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx2_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
OAI221xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B1(n_689), .B2(n_696), .C(n_737), .Y(n_510) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
OA21x2_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_523), .B(n_530), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
NAND2x1p5_ASAP7_75t_L g535 ( .A(n_519), .B(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g614 ( .A(n_519), .Y(n_614) );
AND2x4_ASAP7_75t_L g644 ( .A(n_519), .B(n_645), .Y(n_644) );
AND3x1_ASAP7_75t_L g666 ( .A(n_519), .B(n_667), .C(n_669), .Y(n_666) );
AND2x4_ASAP7_75t_SL g681 ( .A(n_519), .B(n_536), .Y(n_681) );
INVx2_ASAP7_75t_L g603 ( .A(n_520), .Y(n_603) );
OR2x2_ASAP7_75t_L g607 ( .A(n_520), .B(n_581), .Y(n_607) );
OR2x6_ASAP7_75t_SL g609 ( .A(n_520), .B(n_556), .Y(n_609) );
OR2x6_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
BUFx2_ASAP7_75t_L g562 ( .A(n_521), .Y(n_562) );
INVx1_ASAP7_75t_L g570 ( .A(n_521), .Y(n_570) );
AND2x4_ASAP7_75t_L g561 ( .A(n_522), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g569 ( .A(n_522), .B(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g591 ( .A(n_522), .B(n_570), .Y(n_591) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx3_ASAP7_75t_L g541 ( .A(n_525), .Y(n_541) );
INVx4_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx12f_ASAP7_75t_L g588 ( .A(n_526), .Y(n_588) );
AND2x4_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
INVx1_ASAP7_75t_L g546 ( .A(n_527), .Y(n_546) );
AND2x4_ASAP7_75t_L g582 ( .A(n_527), .B(n_547), .Y(n_582) );
AND2x4_ASAP7_75t_L g557 ( .A(n_528), .B(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g551 ( .A(n_529), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g606 ( .A(n_529), .B(n_558), .Y(n_606) );
OR2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_535), .Y(n_530) );
INVx1_ASAP7_75t_L g620 ( .A(n_531), .Y(n_620) );
INVx3_ASAP7_75t_L g654 ( .A(n_531), .Y(n_654) );
OR2x6_ASAP7_75t_L g685 ( .A(n_531), .B(n_643), .Y(n_685) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
INVx2_ASAP7_75t_L g624 ( .A(n_533), .Y(n_624) );
AND2x4_ASAP7_75t_L g636 ( .A(n_533), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g625 ( .A(n_534), .Y(n_625) );
INVx2_ASAP7_75t_L g637 ( .A(n_534), .Y(n_637) );
OR2x6_ASAP7_75t_L g649 ( .A(n_535), .B(n_650), .Y(n_649) );
OR2x6_ASAP7_75t_L g672 ( .A(n_535), .B(n_673), .Y(n_672) );
OAI21xp5_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_600), .B(n_610), .Y(n_537) );
NAND4xp25_ASAP7_75t_SL g538 ( .A(n_539), .B(n_563), .C(n_578), .D(n_592), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_548), .Y(n_539) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx3_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g585 ( .A(n_545), .Y(n_585) );
AND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
INVx1_ASAP7_75t_L g566 ( .A(n_547), .Y(n_566) );
INVx5_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g595 ( .A(n_551), .Y(n_595) );
INVx2_ASAP7_75t_L g558 ( .A(n_552), .Y(n_558) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
BUFx2_ASAP7_75t_L g589 ( .A(n_555), .Y(n_589) );
INVx4_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_557), .Y(n_599) );
INVx1_ASAP7_75t_L g576 ( .A(n_558), .Y(n_576) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
BUFx6f_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_565), .B1(n_571), .B2(n_572), .Y(n_563) );
INVx2_ASAP7_75t_SL g730 ( .A(n_565), .Y(n_730) );
AND2x4_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
NAND3xp33_ASAP7_75t_L g723 ( .A(n_566), .B(n_590), .C(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g577 ( .A(n_568), .Y(n_577) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
BUFx3_ASAP7_75t_L g596 ( .A(n_569), .Y(n_596) );
OAI22xp5_ASAP7_75t_SL g617 ( .A1(n_571), .A2(n_618), .B1(n_619), .B2(n_621), .Y(n_617) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x4_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
INVx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OAI221xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_583), .B1(n_584), .B2(n_586), .C(n_587), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx8_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_583), .A2(n_621), .B1(n_653), .B2(n_655), .Y(n_652) );
BUFx3_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_586), .A2(n_657), .B1(n_661), .B2(n_662), .Y(n_656) );
BUFx6f_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AOI21xp33_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_597), .B(n_598), .Y(n_592) );
AND2x4_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x4_ASAP7_75t_L g598 ( .A(n_596), .B(n_599), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_597), .A2(n_627), .B1(n_628), .B2(n_633), .Y(n_626) );
INVx4_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x4_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx3_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
BUFx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OR2x6_ASAP7_75t_L g639 ( .A(n_614), .B(n_640), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g615 ( .A(n_616), .B(n_651), .C(n_682), .Y(n_615) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
BUFx12f_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_623), .Y(n_650) );
NAND2x1p5_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx3_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
BUFx3_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_632), .Y(n_660) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g647 ( .A(n_635), .Y(n_647) );
BUFx2_ASAP7_75t_L g663 ( .A(n_635), .Y(n_663) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_637), .Y(n_674) );
BUFx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OR2x6_ASAP7_75t_L g642 ( .A(n_643), .B(n_647), .Y(n_642) );
OR2x6_ASAP7_75t_L g686 ( .A(n_643), .B(n_687), .Y(n_686) );
OR2x6_ASAP7_75t_L g688 ( .A(n_643), .B(n_650), .Y(n_688) );
INVx4_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g668 ( .A(n_646), .Y(n_668) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx3_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVxp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
BUFx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
BUFx12f_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
INVx3_ASAP7_75t_L g687 ( .A(n_660), .Y(n_687) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
BUFx6f_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx3_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx4_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx5_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AND2x4_ASAP7_75t_L g676 ( .A(n_677), .B(n_681), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVxp67_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
BUFx6f_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_694), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
BUFx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g721 ( .A(n_693), .Y(n_721) );
AND2x2_ASAP7_75t_L g744 ( .A(n_694), .B(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_695), .B(n_721), .Y(n_720) );
XOR2xp5_ASAP7_75t_L g697 ( .A(n_698), .B(n_709), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_703), .B1(n_704), .B2(n_708), .Y(n_698) );
INVx1_ASAP7_75t_L g708 ( .A(n_699), .Y(n_708) );
INVx1_ASAP7_75t_L g702 ( .A(n_701), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
BUFx3_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx5_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx3_ASAP7_75t_L g739 ( .A(n_718), .Y(n_739) );
AND2x6_ASAP7_75t_L g718 ( .A(n_719), .B(n_726), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_722), .Y(n_719) );
INVxp67_ASAP7_75t_L g735 ( .A(n_720), .Y(n_735) );
INVx1_ASAP7_75t_L g745 ( .A(n_721), .Y(n_745) );
INVxp67_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_723), .B(n_730), .Y(n_736) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
CKINVDCx11_ASAP7_75t_R g728 ( .A(n_725), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_729), .Y(n_726) );
CKINVDCx5p33_ASAP7_75t_R g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
BUFx6f_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
BUFx4f_ASAP7_75t_SL g740 ( .A(n_733), .Y(n_740) );
INVx4_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_743), .Y(n_742) );
endmodule