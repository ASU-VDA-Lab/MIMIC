module real_jpeg_16572_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_508),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_0),
.B(n_509),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_1),
.Y(n_116)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_1),
.Y(n_128)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_1),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_2),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_2),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g358 ( 
.A(n_2),
.Y(n_358)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_3),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_3),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g386 ( 
.A(n_3),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_4),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_23)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g130 ( 
.A1(n_4),
.A2(n_26),
.B1(n_131),
.B2(n_133),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_4),
.A2(n_26),
.B1(n_148),
.B2(n_151),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_4),
.B(n_256),
.Y(n_257)
);

OAI22x1_ASAP7_75t_SL g238 ( 
.A1(n_5),
.A2(n_239),
.B1(n_244),
.B2(n_245),
.Y(n_238)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_5),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_5),
.A2(n_244),
.B1(n_288),
.B2(n_290),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_5),
.A2(n_244),
.B1(n_330),
.B2(n_333),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g367 ( 
.A1(n_5),
.A2(n_244),
.B1(n_368),
.B2(n_371),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_6),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_6),
.Y(n_89)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_6),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_6),
.Y(n_124)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_6),
.Y(n_150)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_6),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_6),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_7),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_8),
.A2(n_97),
.B1(n_102),
.B2(n_107),
.Y(n_96)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_8),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_8),
.A2(n_107),
.B1(n_185),
.B2(n_190),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_8),
.A2(n_107),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_8),
.A2(n_107),
.B1(n_315),
.B2(n_319),
.Y(n_314)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_9),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_10),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_11),
.Y(n_172)
);

BUFx4f_ASAP7_75t_L g318 ( 
.A(n_11),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_12),
.Y(n_52)
);

OAI22x1_ASAP7_75t_L g87 ( 
.A1(n_12),
.A2(n_52),
.B1(n_88),
.B2(n_90),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_12),
.A2(n_52),
.B1(n_175),
.B2(n_178),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_12),
.B(n_211),
.Y(n_210)
);

OAI32xp33_ASAP7_75t_L g343 ( 
.A1(n_12),
.A2(n_344),
.A3(n_345),
.B1(n_348),
.B2(n_352),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_12),
.B(n_121),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_12),
.B(n_384),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_12),
.B(n_61),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g220 ( 
.A(n_13),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g332 ( 
.A(n_13),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_229),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_227),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_200),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_18),
.B(n_200),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_137),
.C(n_154),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_19),
.A2(n_137),
.B1(n_138),
.B2(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_19),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_57),
.B2(n_58),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_20),
.B(n_60),
.C(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_20),
.A2(n_21),
.B1(n_204),
.B2(n_226),
.Y(n_203)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_41),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_22),
.B(n_433),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_32),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_23),
.B(n_42),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_26),
.B(n_255),
.Y(n_254)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_29),
.A2(n_44),
.B1(n_47),
.B2(n_50),
.Y(n_43)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_29),
.Y(n_333)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_32),
.B(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_43),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_33),
.A2(n_198),
.B(n_199),
.Y(n_197)
);

OAI21xp33_ASAP7_75t_SL g217 ( 
.A1(n_33),
.A2(n_218),
.B(n_223),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_33),
.B(n_52),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_L g476 ( 
.A1(n_33),
.A2(n_198),
.B1(n_199),
.B2(n_477),
.Y(n_476)
);

OA22x2_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_36),
.Y(n_120)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_41),
.B(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_51),
.Y(n_41)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_42),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_42),
.B(n_329),
.Y(n_433)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_46),
.Y(n_309)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_51),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B(n_55),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_52),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_52),
.B(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_52),
.B(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_52),
.B(n_349),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_54),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_55),
.A2(n_302),
.B1(n_306),
.B2(n_312),
.Y(n_301)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_95),
.B2(n_136),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_59),
.A2(n_206),
.B1(n_207),
.B2(n_215),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_59),
.A2(n_215),
.B1(n_335),
.B2(n_336),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_59),
.B(n_327),
.C(n_336),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

OA21x2_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_77),
.B(n_87),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_61),
.B(n_147),
.Y(n_195)
);

OA21x2_ASAP7_75t_L g215 ( 
.A1(n_61),
.A2(n_77),
.B(n_87),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_61),
.B(n_287),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_61),
.B(n_184),
.Y(n_439)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_62),
.B(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_62),
.B(n_145),
.Y(n_144)
);

AOI22x1_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_67),
.B1(n_70),
.B2(n_73),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_69),
.Y(n_181)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_72),
.Y(n_177)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_72),
.Y(n_256)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_72),
.Y(n_321)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_72),
.Y(n_347)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_72),
.Y(n_370)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_77),
.B(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_77),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_77),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_77),
.B(n_87),
.Y(n_361)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_81),
.B1(n_84),
.B2(n_86),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_86),
.Y(n_354)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_94),
.Y(n_189)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_94),
.Y(n_193)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_95),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_108),
.B(n_129),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_100),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_101),
.Y(n_243)
);

BUFx5_ASAP7_75t_L g269 ( 
.A(n_101),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2x1_ASAP7_75t_L g411 ( 
.A(n_108),
.B(n_412),
.Y(n_411)
);

AOI21x1_ASAP7_75t_L g449 ( 
.A1(n_108),
.A2(n_412),
.B(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_130),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_109),
.B(n_238),
.Y(n_237)
);

NOR2x1p5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_121),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_114),
.B1(n_117),
.B2(n_118),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_113),
.Y(n_214)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_114),
.Y(n_117)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_121),
.B(n_130),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_121),
.A2(n_140),
.B(n_141),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_121),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_121),
.B(n_238),
.Y(n_337)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_121),
.Y(n_450)
);

AO22x2_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_121)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_129),
.B(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_129),
.Y(n_475)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OA21x2_ASAP7_75t_L g489 ( 
.A1(n_138),
.A2(n_139),
.B(n_143),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g207 ( 
.A(n_142),
.B(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_142),
.B(n_337),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_144),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_146),
.B(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_146),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_153),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_154),
.B(n_503),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_196),
.B(n_197),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_156),
.B(n_491),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_182),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_157),
.B(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_157),
.B(n_265),
.Y(n_413)
);

XNOR2x2_ASAP7_75t_SL g470 ( 
.A(n_157),
.B(n_182),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_157),
.B(n_197),
.Y(n_491)
);

OA21x2_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_164),
.B(n_173),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx4_ASAP7_75t_SL g391 ( 
.A(n_161),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_163),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_165),
.B(n_174),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_165),
.B(n_257),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_165),
.B(n_367),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_165),
.A2(n_314),
.B(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

AO21x1_ASAP7_75t_L g363 ( 
.A1(n_173),
.A2(n_364),
.B(n_366),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_173),
.A2(n_325),
.B(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_177),
.Y(n_373)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_194),
.B(n_195),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_192),
.Y(n_289)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_195),
.B(n_286),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_195),
.B(n_361),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_203),
.Y(n_200)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_216),
.B1(n_217),
.B2(n_225),
.Y(n_204)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AND2x2_ASAP7_75t_SL g430 ( 
.A(n_208),
.B(n_237),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_209),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI32xp33_ASAP7_75t_L g265 ( 
.A1(n_213),
.A2(n_266),
.A3(n_270),
.B1(n_273),
.B2(n_279),
.Y(n_265)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_224),
.B(n_328),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_501),
.B(n_507),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

AO221x1_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_424),
.B1(n_494),
.B2(n_499),
.C(n_500),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_338),
.B(n_423),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_295),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_234),
.B(n_295),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_264),
.C(n_283),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_235),
.B(n_419),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_249),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_236),
.B(n_250),
.C(n_263),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_243),
.Y(n_248)
);

BUFx2_ASAP7_75t_SL g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_247),
.Y(n_312)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx8_ASAP7_75t_L g305 ( 
.A(n_248),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_262),
.B2(n_263),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_252),
.B(n_388),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_253),
.B(n_366),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_253),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_257),
.B(n_258),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_258),
.Y(n_365)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_264),
.A2(n_283),
.B1(n_284),
.B2(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_264),
.Y(n_420)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_269),
.Y(n_268)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_272),
.Y(n_282)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx6_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_326),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_297),
.B(n_300),
.C(n_326),
.Y(n_460)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_313),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_301),
.B(n_313),
.Y(n_429)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_310),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_314),
.A2(n_322),
.B(n_324),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_318),
.Y(n_351)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx6_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_323),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_324),
.B(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_334),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_329),
.Y(n_477)
);

INVx5_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx8_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_337),
.B(n_410),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_417),
.B(n_422),
.Y(n_338)
);

OAI21x1_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_402),
.B(n_416),
.Y(n_339)
);

AOI21x1_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_379),
.B(n_401),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_362),
.Y(n_341)
);

NOR2xp67_ASAP7_75t_SL g401 ( 
.A(n_342),
.B(n_362),
.Y(n_401)
);

NAND2xp33_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_359),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_343),
.B(n_359),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_345),
.B(n_383),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_355),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_360),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_374),
.Y(n_362)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_363),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_367),
.B(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_375),
.A2(n_376),
.B1(n_377),
.B2(n_378),
.Y(n_374)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_375),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_376),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_376),
.B(n_377),
.C(n_415),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_380),
.A2(n_396),
.B(n_400),
.Y(n_379)
);

AOI21x1_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_392),
.B(n_395),
.Y(n_380)
);

NOR2x1_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_387),
.Y(n_381)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_388),
.Y(n_398)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_393),
.B(n_394),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_393),
.B(n_394),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_399),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_397),
.B(n_399),
.Y(n_400)
);

NOR2xp67_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_414),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_403),
.B(n_414),
.Y(n_416)
);

XOR2x2_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_413),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_405),
.A2(n_406),
.B1(n_408),
.B2(n_409),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_405),
.B(n_409),
.C(n_413),
.Y(n_421)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

NOR2x1_ASAP7_75t_L g474 ( 
.A(n_411),
.B(n_475),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_418),
.B(n_421),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_418),
.B(n_421),
.Y(n_422)
);

NOR3xp33_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_463),
.C(n_480),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_426),
.B(n_459),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_426),
.B(n_497),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_427),
.B(n_452),
.Y(n_426)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_427),
.B(n_452),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_434),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_428),
.B(n_435),
.C(n_441),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.C(n_431),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_429),
.B(n_455),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_430),
.A2(n_431),
.B1(n_432),
.B2(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_430),
.Y(n_456)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_441),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_438),
.Y(n_435)
);

AOI21x1_ASAP7_75t_SL g472 ( 
.A1(n_436),
.A2(n_439),
.B(n_440),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_446),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_442),
.B(n_467),
.C(n_468),
.Y(n_466)
);

NAND2x1_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_445),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_443),
.B(n_445),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_447),
.A2(n_448),
.B1(n_449),
.B2(n_451),
.Y(n_446)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_447),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_448),
.Y(n_467)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_451),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_457),
.C(n_458),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_454),
.B(n_462),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_457),
.B(n_458),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_461),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_460),
.B(n_461),
.Y(n_497)
);

A2O1A1Ixp33_ASAP7_75t_L g494 ( 
.A1(n_463),
.A2(n_495),
.B(n_496),
.C(n_498),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_465),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_464),
.B(n_465),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_469),
.Y(n_465)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_466),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_470),
.A2(n_471),
.B1(n_478),
.B2(n_479),
.Y(n_469)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_470),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_470),
.B(n_478),
.C(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_471),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_472),
.B(n_485),
.C(n_487),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_476),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_474),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_476),
.Y(n_487)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_480),
.Y(n_499)
);

NOR2x1_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_483),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_481),
.B(n_483),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_488),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_484),
.B(n_489),
.C(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_489),
.A2(n_490),
.B1(n_492),
.B2(n_493),
.Y(n_488)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_489),
.Y(n_493)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_490),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_492),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_502),
.B(n_505),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_502),
.B(n_505),
.Y(n_507)
);


endmodule