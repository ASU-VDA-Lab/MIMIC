module fake_jpeg_12543_n_450 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_450);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_450;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_15),
.B(n_7),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_46),
.B(n_50),
.Y(n_98)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_15),
.B(n_7),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_48),
.B(n_80),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_25),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_49),
.B(n_55),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_25),
.B(n_6),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_52),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

BUFx4f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_56),
.Y(n_147)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_58),
.B(n_60),
.Y(n_106)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_37),
.B(n_6),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_64),
.B(n_69),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_67),
.Y(n_127)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_8),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_34),
.B(n_35),
.Y(n_70)
);

AOI21xp33_ASAP7_75t_SL g125 ( 
.A1(n_70),
.A2(n_30),
.B(n_28),
.Y(n_125)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_72),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_31),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_78),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_35),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_31),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_81),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_35),
.B(n_8),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_31),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_82),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_83),
.Y(n_133)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_85),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_38),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_90),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_33),
.Y(n_89)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_38),
.B(n_8),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_91),
.B(n_93),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_33),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_92),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_44),
.B(n_26),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_42),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_80),
.B(n_33),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_99),
.B(n_132),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_94),
.A2(n_78),
.B1(n_48),
.B2(n_68),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_100),
.A2(n_110),
.B1(n_93),
.B2(n_65),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_92),
.A2(n_44),
.B1(n_39),
.B2(n_17),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_101),
.A2(n_114),
.B1(n_118),
.B2(n_134),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_70),
.A2(n_23),
.B(n_24),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_104),
.A2(n_1),
.B(n_2),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_71),
.A2(n_39),
.B1(n_17),
.B2(n_27),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_89),
.A2(n_44),
.B1(n_39),
.B2(n_17),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_57),
.A2(n_27),
.B1(n_22),
.B2(n_17),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_116),
.A2(n_123),
.B1(n_124),
.B2(n_145),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_89),
.A2(n_27),
.B1(n_22),
.B2(n_23),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_61),
.A2(n_27),
.B1(n_22),
.B2(n_42),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_63),
.A2(n_22),
.B1(n_28),
.B2(n_30),
.Y(n_124)
);

NAND2x1_ASAP7_75t_L g178 ( 
.A(n_125),
.B(n_72),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_47),
.A2(n_24),
.B1(n_23),
.B2(n_16),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_70),
.B(n_16),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_59),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_74),
.A2(n_24),
.B1(n_41),
.B2(n_40),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_142),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_52),
.A2(n_40),
.B1(n_41),
.B2(n_9),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_56),
.A2(n_41),
.B1(n_9),
.B2(n_10),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_146),
.A2(n_87),
.B1(n_53),
.B2(n_91),
.Y(n_173)
);

O2A1O1Ixp33_ASAP7_75t_SL g149 ( 
.A1(n_100),
.A2(n_85),
.B(n_86),
.C(n_83),
.Y(n_149)
);

AO21x2_ASAP7_75t_SL g196 ( 
.A1(n_149),
.A2(n_174),
.B(n_123),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_154),
.Y(n_194)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_151),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_153),
.A2(n_155),
.B1(n_111),
.B2(n_108),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_110),
.A2(n_76),
.B1(n_51),
.B2(n_73),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_157),
.Y(n_223)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_158),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_132),
.A2(n_82),
.B1(n_66),
.B2(n_67),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_159),
.A2(n_180),
.B1(n_143),
.B2(n_138),
.Y(n_206)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_126),
.A2(n_62),
.B(n_54),
.C(n_83),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_161),
.A2(n_130),
.B(n_122),
.C(n_127),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_0),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_162),
.B(n_175),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_168),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_165),
.Y(n_212)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

BUFx12_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

BUFx24_ASAP7_75t_L g211 ( 
.A(n_167),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_135),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_170),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_99),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_171),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_129),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_172),
.B(n_176),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_173),
.A2(n_192),
.B1(n_145),
.B2(n_148),
.Y(n_205)
);

AO22x2_ASAP7_75t_L g174 ( 
.A1(n_99),
.A2(n_75),
.B1(n_72),
.B2(n_54),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_119),
.B(n_0),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_135),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_95),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_177),
.B(n_181),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_187),
.B(n_115),
.Y(n_204)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_105),
.Y(n_179)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_104),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_180)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_103),
.B(n_131),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_120),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_185),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_184),
.A2(n_107),
.B(n_113),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_98),
.B(n_9),
.Y(n_185)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_140),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_186),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_188),
.A2(n_148),
.B1(n_121),
.B2(n_109),
.Y(n_217)
);

OR2x4_ASAP7_75t_L g189 ( 
.A(n_117),
.B(n_10),
.Y(n_189)
);

NOR2x1_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_102),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_108),
.B(n_1),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_190),
.B(n_191),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_124),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_106),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_196),
.A2(n_205),
.B1(n_206),
.B2(n_174),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_198),
.A2(n_201),
.B1(n_203),
.B2(n_152),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_111),
.C(n_112),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_178),
.C(n_171),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_191),
.A2(n_144),
.B1(n_137),
.B2(n_117),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_179),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_163),
.A2(n_137),
.B1(n_116),
.B2(n_112),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_204),
.A2(n_208),
.B(n_220),
.Y(n_230)
);

AOI32xp33_ASAP7_75t_L g207 ( 
.A1(n_178),
.A2(n_130),
.A3(n_121),
.B1(n_122),
.B2(n_113),
.Y(n_207)
);

MAJx2_ASAP7_75t_L g247 ( 
.A(n_207),
.B(n_174),
.C(n_161),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_217),
.A2(n_222),
.B1(n_165),
.B2(n_211),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_154),
.A2(n_164),
.B1(n_149),
.B2(n_170),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_225),
.B(n_174),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_228),
.A2(n_220),
.B(n_208),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_203),
.A2(n_176),
.B1(n_169),
.B2(n_168),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_229),
.A2(n_249),
.B(n_251),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_231),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_211),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_232),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_162),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_233),
.B(n_235),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_234),
.B(n_255),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_196),
.A2(n_215),
.B1(n_206),
.B2(n_218),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_237),
.Y(n_283)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_238),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_194),
.B(n_160),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_239),
.B(n_246),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_245),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_196),
.A2(n_150),
.B1(n_149),
.B2(n_187),
.Y(n_241)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_241),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_198),
.A2(n_159),
.B1(n_160),
.B2(n_171),
.Y(n_242)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_242),
.Y(n_281)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_195),
.Y(n_243)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_243),
.Y(n_271)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_244),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_197),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_194),
.B(n_190),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_247),
.B(n_241),
.Y(n_282)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_214),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_248),
.B(n_250),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_225),
.A2(n_174),
.B(n_189),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_180),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_183),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_214),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_252),
.Y(n_267)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_195),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_253),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_218),
.B(n_175),
.C(n_97),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_204),
.C(n_197),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_221),
.B(n_200),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_223),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_256),
.Y(n_275)
);

NAND3xp33_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_177),
.C(n_158),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_257),
.A2(n_211),
.B(n_225),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_259),
.B(n_263),
.C(n_268),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_261),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_216),
.C(n_207),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_265),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_230),
.A2(n_208),
.B(n_196),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_266),
.A2(n_274),
.B(n_278),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_239),
.C(n_254),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_233),
.B(n_216),
.C(n_97),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_236),
.C(n_238),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_230),
.A2(n_210),
.B(n_201),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_237),
.A2(n_196),
.B(n_219),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_282),
.B(n_226),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_235),
.B(n_210),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_286),
.A2(n_227),
.B(n_213),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_251),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_287),
.B(n_289),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_260),
.A2(n_231),
.B1(n_242),
.B2(n_245),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_288),
.A2(n_290),
.B1(n_309),
.B2(n_314),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_193),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_285),
.A2(n_244),
.B1(n_250),
.B2(n_247),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_246),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_294),
.B(n_296),
.C(n_307),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_285),
.A2(n_249),
.B1(n_205),
.B2(n_247),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_295),
.A2(n_301),
.B1(n_302),
.B2(n_313),
.Y(n_319)
);

FAx1_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_249),
.CI(n_211),
.CON(n_297),
.SN(n_297)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_297),
.A2(n_303),
.B(n_266),
.Y(n_323)
);

A2O1A1Ixp33_ASAP7_75t_R g298 ( 
.A1(n_283),
.A2(n_240),
.B(n_252),
.C(n_248),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_298),
.B(n_299),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_269),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_262),
.Y(n_300)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_300),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_260),
.A2(n_232),
.B1(n_199),
.B2(n_219),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_281),
.A2(n_199),
.B1(n_232),
.B2(n_256),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_262),
.Y(n_304)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_304),
.Y(n_331)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_273),
.Y(n_305)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_305),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_270),
.B(n_227),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_306),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_268),
.B(n_213),
.C(n_253),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_273),
.Y(n_308)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_308),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_281),
.A2(n_212),
.B1(n_199),
.B2(n_165),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_311),
.B(n_277),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_277),
.B(n_226),
.C(n_156),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_277),
.C(n_259),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_279),
.A2(n_151),
.B1(n_188),
.B2(n_243),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_271),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_290),
.A2(n_279),
.B1(n_280),
.B2(n_278),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_318),
.A2(n_329),
.B1(n_293),
.B2(n_301),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_298),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_321),
.B(n_310),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_322),
.B(n_326),
.Y(n_344)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_323),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_325),
.B(n_327),
.C(n_332),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_291),
.B(n_259),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_291),
.B(n_263),
.C(n_282),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_295),
.A2(n_258),
.B1(n_280),
.B2(n_283),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_328),
.A2(n_330),
.B1(n_335),
.B2(n_342),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_293),
.A2(n_286),
.B1(n_258),
.B2(n_261),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_303),
.A2(n_274),
.B1(n_263),
.B2(n_284),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_294),
.B(n_270),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_307),
.B(n_269),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_334),
.B(n_314),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_292),
.A2(n_284),
.B1(n_286),
.B2(n_265),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_296),
.B(n_226),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_338),
.B(n_339),
.C(n_340),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_311),
.B(n_267),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_312),
.B(n_267),
.C(n_275),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_310),
.B(n_264),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_309),
.C(n_297),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_292),
.A2(n_275),
.B1(n_272),
.B2(n_264),
.Y(n_342)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_343),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_345),
.A2(n_349),
.B1(n_352),
.B2(n_353),
.Y(n_373)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_337),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_346),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_336),
.B(n_302),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_347),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_316),
.B(n_300),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_348),
.B(n_350),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_320),
.A2(n_318),
.B1(n_329),
.B2(n_323),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_324),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_331),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_351),
.A2(n_363),
.B1(n_165),
.B2(n_181),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_339),
.A2(n_313),
.B1(n_297),
.B2(n_304),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_341),
.A2(n_297),
.B1(n_308),
.B2(n_305),
.Y(n_353)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_333),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_361),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_359),
.B(n_360),
.C(n_364),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_315),
.A2(n_272),
.B1(n_271),
.B2(n_212),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_342),
.B(n_271),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_362),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_317),
.B(n_223),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_317),
.B(n_157),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_319),
.A2(n_212),
.B1(n_147),
.B2(n_138),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_365),
.A2(n_357),
.B1(n_340),
.B2(n_355),
.Y(n_371)
);

OAI321xp33_ASAP7_75t_L g370 ( 
.A1(n_354),
.A2(n_328),
.A3(n_335),
.B1(n_330),
.B2(n_319),
.C(n_322),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_370),
.B(n_376),
.Y(n_395)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_371),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_356),
.B(n_326),
.C(n_364),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_372),
.B(n_375),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_347),
.B(n_338),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_374),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_356),
.B(n_358),
.C(n_325),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_362),
.B(n_332),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_354),
.B(n_334),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_377),
.B(n_378),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_352),
.B(n_327),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_353),
.B(n_358),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_382),
.B(n_384),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_344),
.B(n_107),
.C(n_143),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_383),
.B(n_359),
.C(n_360),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_349),
.B(n_186),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_385),
.B(n_109),
.Y(n_401)
);

INVx11_ASAP7_75t_L g386 ( 
.A(n_368),
.Y(n_386)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_386),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_367),
.B(n_355),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_388),
.B(n_389),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_384),
.A2(n_345),
.B(n_344),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_390),
.A2(n_371),
.B(n_366),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_379),
.A2(n_365),
.B(n_167),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_391),
.A2(n_369),
.B(n_379),
.Y(n_406)
);

INVxp33_ASAP7_75t_L g392 ( 
.A(n_381),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_392),
.B(n_402),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_375),
.B(n_109),
.C(n_143),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_393),
.B(n_373),
.Y(n_416)
);

OAI221xp5_ASAP7_75t_L g394 ( 
.A1(n_382),
.A2(n_167),
.B1(n_14),
.B2(n_147),
.C(n_102),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_394),
.A2(n_380),
.B1(n_138),
.B2(n_369),
.Y(n_403)
);

NOR2xp67_ASAP7_75t_L g396 ( 
.A(n_372),
.B(n_167),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_396),
.B(n_366),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_367),
.B(n_102),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_399),
.B(n_401),
.Y(n_410)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_403),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_402),
.Y(n_404)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_404),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_406),
.B(n_413),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_386),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_407),
.B(n_408),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_397),
.B(n_378),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_395),
.B(n_377),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_411),
.B(n_412),
.Y(n_417)
);

INVx6_ASAP7_75t_L g412 ( 
.A(n_395),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_414),
.B(n_416),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_415),
.A2(n_400),
.B1(n_387),
.B2(n_376),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_405),
.B(n_388),
.C(n_400),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_420),
.B(n_421),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_412),
.A2(n_390),
.B(n_387),
.Y(n_424)
);

AOI21x1_ASAP7_75t_SL g429 ( 
.A1(n_424),
.A2(n_428),
.B(n_422),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_406),
.A2(n_374),
.B1(n_391),
.B2(n_370),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_425),
.B(n_426),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_405),
.B(n_399),
.C(n_398),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_413),
.A2(n_373),
.B(n_389),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_429),
.A2(n_383),
.B(n_410),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_419),
.B(n_414),
.Y(n_431)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_431),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_427),
.A2(n_404),
.B(n_409),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_432),
.A2(n_433),
.B(n_435),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_426),
.B(n_398),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_417),
.B(n_393),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_423),
.B(n_410),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_436),
.A2(n_437),
.B(n_3),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_420),
.B(n_428),
.C(n_422),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_437),
.A2(n_418),
.B1(n_424),
.B2(n_401),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_438),
.B(n_439),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_441),
.B(n_4),
.C(n_5),
.Y(n_444)
);

A2O1A1Ixp33_ASAP7_75t_L g443 ( 
.A1(n_442),
.A2(n_430),
.B(n_429),
.C(n_434),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_443),
.A2(n_444),
.B(n_440),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_446),
.A2(n_447),
.B(n_4),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_445),
.A2(n_4),
.B(n_5),
.Y(n_447)
);

BUFx24_ASAP7_75t_SL g449 ( 
.A(n_448),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_449),
.B(n_5),
.Y(n_450)
);


endmodule