module fake_jpeg_30621_n_324 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_324);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_7),
.A2(n_10),
.B(n_16),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_8),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_46),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_8),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_27),
.B(n_7),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_53),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_52),
.B(n_38),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_27),
.B(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_21),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_62),
.Y(n_71)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_21),
.B(n_1),
.Y(n_62)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_32),
.Y(n_88)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_28),
.B1(n_34),
.B2(n_40),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_75),
.A2(n_91),
.B1(n_112),
.B2(n_19),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_34),
.B1(n_37),
.B2(n_40),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_76),
.A2(n_85),
.B1(n_96),
.B2(n_110),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_42),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_80),
.B(n_105),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_28),
.B1(n_38),
.B2(n_42),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_84),
.A2(n_92),
.B1(n_1),
.B2(n_2),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_65),
.A2(n_40),
.B1(n_32),
.B2(n_26),
.Y(n_85)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_66),
.A2(n_32),
.B1(n_30),
.B2(n_36),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_52),
.A2(n_41),
.B1(n_39),
.B2(n_23),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_33),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_93),
.B(n_94),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_33),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_47),
.B(n_36),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_95),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_58),
.A2(n_70),
.B1(n_56),
.B2(n_49),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_51),
.Y(n_100)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_41),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_101),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_61),
.B(n_39),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_102),
.Y(n_131)
);

OR2x2_ASAP7_75t_SL g119 ( 
.A(n_103),
.B(n_104),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_51),
.B(n_35),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_57),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_69),
.A2(n_35),
.B1(n_31),
.B2(n_29),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_64),
.A2(n_31),
.B1(n_29),
.B2(n_23),
.Y(n_112)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_114),
.Y(n_181)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_68),
.B1(n_67),
.B2(n_54),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_116),
.A2(n_97),
.B1(n_113),
.B2(n_79),
.Y(n_156)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_71),
.A2(n_69),
.B1(n_45),
.B2(n_51),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_122),
.A2(n_136),
.B1(n_139),
.B2(n_150),
.Y(n_173)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_124),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_140),
.B1(n_142),
.B2(n_100),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_82),
.A2(n_19),
.B1(n_69),
.B2(n_3),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_75),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_127),
.A2(n_145),
.B1(n_97),
.B2(n_113),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_73),
.Y(n_153)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_80),
.A2(n_11),
.B1(n_3),
.B2(n_4),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_71),
.B(n_1),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_81),
.Y(n_162)
);

AO22x2_ASAP7_75t_L g138 ( 
.A1(n_98),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_138)
);

OAI32xp33_ASAP7_75t_L g177 ( 
.A1(n_138),
.A2(n_139),
.A3(n_122),
.B1(n_120),
.B2(n_124),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_82),
.A2(n_5),
.B1(n_7),
.B2(n_11),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_82),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_81),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_143),
.B(n_144),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_77),
.A2(n_17),
.B(n_18),
.C(n_74),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_112),
.A2(n_17),
.B1(n_99),
.B2(n_111),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_104),
.A2(n_17),
.B(n_92),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_147),
.A2(n_148),
.B(n_132),
.Y(n_176)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_99),
.Y(n_149)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_111),
.A2(n_109),
.B1(n_86),
.B2(n_83),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_86),
.A2(n_105),
.B1(n_89),
.B2(n_106),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_151),
.A2(n_150),
.B1(n_121),
.B2(n_115),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_152),
.A2(n_153),
.B1(n_156),
.B2(n_157),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_79),
.B1(n_87),
.B2(n_108),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_158),
.A2(n_175),
.B1(n_118),
.B2(n_138),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_108),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_159),
.B(n_162),
.Y(n_190)
);

BUFx24_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

INVxp67_ASAP7_75t_SL g193 ( 
.A(n_160),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_87),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_119),
.C(n_117),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_73),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_167),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_129),
.B(n_73),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_123),
.B(n_107),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_172),
.B(n_174),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_123),
.B(n_107),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_125),
.A2(n_127),
.B1(n_147),
.B2(n_145),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_176),
.A2(n_144),
.B(n_119),
.Y(n_195)
);

AOI21x1_ASAP7_75t_SL g189 ( 
.A1(n_177),
.A2(n_138),
.B(n_129),
.Y(n_189)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_121),
.Y(n_178)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_178),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_141),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_182),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_131),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_151),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_118),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_178),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_187),
.B(n_214),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_189),
.A2(n_196),
.B1(n_206),
.B2(n_190),
.Y(n_234)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_194),
.A2(n_209),
.B1(n_181),
.B2(n_170),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

OAI22x1_ASAP7_75t_L g196 ( 
.A1(n_154),
.A2(n_177),
.B1(n_182),
.B2(n_153),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_196),
.A2(n_205),
.B(n_211),
.Y(n_217)
);

INVx13_ASAP7_75t_L g198 ( 
.A(n_181),
.Y(n_198)
);

INVxp33_ASAP7_75t_L g235 ( 
.A(n_198),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_208),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_204),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_179),
.A2(n_114),
.B(n_149),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_201),
.A2(n_186),
.B(n_187),
.Y(n_236)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_184),
.Y(n_203)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_203),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_161),
.B(n_133),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_176),
.A2(n_134),
.B(n_135),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_155),
.Y(n_207)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_162),
.B(n_153),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_157),
.A2(n_173),
.B1(n_156),
.B2(n_154),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_165),
.B(n_173),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_188),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_160),
.A2(n_164),
.B(n_180),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_155),
.Y(n_212)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_160),
.B(n_164),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_204),
.C(n_200),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_168),
.B(n_163),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_169),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_215),
.B(n_185),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_219),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_202),
.B(n_160),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_168),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_222),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_189),
.A2(n_170),
.B1(n_171),
.B2(n_169),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_224),
.A2(n_228),
.B1(n_234),
.B2(n_191),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_225),
.B(n_191),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_197),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_227),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_194),
.A2(n_171),
.B1(n_185),
.B2(n_163),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_213),
.C(n_208),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_205),
.C(n_211),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_206),
.B(n_210),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_233),
.B(n_240),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_236),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_207),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_237),
.Y(n_255)
);

NOR2x1_ASAP7_75t_L g239 ( 
.A(n_188),
.B(n_209),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_239),
.Y(n_242)
);

NAND3xp33_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_195),
.C(n_186),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_230),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_250),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_192),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_224),
.Y(n_274)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_216),
.Y(n_247)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_247),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_240),
.A2(n_191),
.B1(n_234),
.B2(n_221),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_248),
.A2(n_251),
.B1(n_259),
.B2(n_228),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_225),
.C(n_229),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_252),
.B(n_260),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_193),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_253),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_218),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_256),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_233),
.B(n_203),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_258),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_239),
.A2(n_212),
.B1(n_215),
.B2(n_198),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_230),
.B(n_226),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_263),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_221),
.B1(n_239),
.B2(n_222),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_265),
.B1(n_270),
.B2(n_271),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_275),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_254),
.A2(n_257),
.B1(n_260),
.B2(n_242),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_245),
.A2(n_219),
.B1(n_236),
.B2(n_217),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_R g272 ( 
.A(n_258),
.B(n_217),
.Y(n_272)
);

AOI321xp33_ASAP7_75t_L g277 ( 
.A1(n_272),
.A2(n_248),
.A3(n_249),
.B1(n_254),
.B2(n_243),
.C(n_256),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_273),
.Y(n_278)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_278),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_272),
.A2(n_249),
.B(n_244),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_271),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_252),
.C(n_250),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_286),
.C(n_287),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_268),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_283),
.B(n_255),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_226),
.Y(n_284)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_284),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_246),
.C(n_251),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_259),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_255),
.Y(n_288)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_288),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_290),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_286),
.C(n_278),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_296),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_281),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_263),
.C(n_265),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_268),
.C(n_262),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_298),
.B(n_216),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_261),
.C(n_275),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_279),
.Y(n_300)
);

OAI221xp5_ASAP7_75t_L g305 ( 
.A1(n_300),
.A2(n_285),
.B1(n_279),
.B2(n_261),
.C(n_237),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_302),
.C(n_291),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_264),
.Y(n_302)
);

AOI21x1_ASAP7_75t_L g304 ( 
.A1(n_295),
.A2(n_277),
.B(n_285),
.Y(n_304)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_304),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_307),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_299),
.A2(n_223),
.B(n_232),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_308),
.A2(n_302),
.B(n_306),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_299),
.C(n_223),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_294),
.Y(n_312)
);

BUFx24_ASAP7_75t_SL g318 ( 
.A(n_312),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_292),
.Y(n_313)
);

AOI21x1_ASAP7_75t_L g317 ( 
.A1(n_313),
.A2(n_220),
.B(n_310),
.Y(n_317)
);

AOI21x1_ASAP7_75t_SL g316 ( 
.A1(n_314),
.A2(n_235),
.B(n_232),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_315),
.Y(n_319)
);

AO22x2_ASAP7_75t_L g321 ( 
.A1(n_316),
.A2(n_317),
.B1(n_311),
.B2(n_220),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_313),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_320),
.B(n_321),
.Y(n_322)
);

BUFx24_ASAP7_75t_SL g323 ( 
.A(n_322),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_319),
.Y(n_324)
);


endmodule