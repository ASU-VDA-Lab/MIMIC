module fake_jpeg_22180_n_178 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_178);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_SL g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_27),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_14),
.B(n_1),
.Y(n_28)
);

OAI21xp33_ASAP7_75t_L g46 ( 
.A1(n_28),
.A2(n_1),
.B(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_30),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_24),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_36),
.B(n_20),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_26),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_41),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_25),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_51),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_49),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_16),
.B(n_18),
.C(n_25),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_21),
.B1(n_15),
.B2(n_26),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_15),
.B1(n_16),
.B2(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_29),
.B(n_13),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_52),
.Y(n_60)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_22),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_56),
.Y(n_68)
);

OAI21xp33_ASAP7_75t_SL g79 ( 
.A1(n_54),
.A2(n_20),
.B(n_43),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_66),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_58),
.A2(n_42),
.B1(n_40),
.B2(n_39),
.Y(n_83)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_64),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_13),
.Y(n_63)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_44),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_16),
.Y(n_66)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_55),
.B(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_71),
.B(n_76),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_67),
.A2(n_47),
.B1(n_33),
.B2(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_67),
.A2(n_45),
.B1(n_44),
.B2(n_35),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_75),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_52),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_78),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NAND2xp33_ASAP7_75t_SL g90 ( 
.A(n_79),
.B(n_40),
.Y(n_90)
);

NOR2x1_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_49),
.Y(n_80)
);

NOR2x1_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_59),
.Y(n_91)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_82),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_83),
.B(n_66),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_57),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_71),
.B(n_68),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_85),
.B(n_69),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_32),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_23),
.B(n_14),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_73),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_64),
.B(n_60),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_95),
.B(n_96),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_60),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_70),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_94),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_30),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_37),
.B(n_65),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_51),
.Y(n_97)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_98),
.A2(n_53),
.B1(n_82),
.B2(n_39),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_101),
.A2(n_103),
.B(n_86),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_69),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_102),
.B(n_110),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_77),
.B(n_80),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_104),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_89),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_108),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_97),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_83),
.B1(n_37),
.B2(n_22),
.Y(n_111)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_114),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_19),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_115),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_84),
.C(n_87),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_122),
.C(n_106),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_93),
.Y(n_121)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_92),
.C(n_91),
.Y(n_122)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_125),
.A2(n_23),
.B(n_19),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_95),
.Y(n_126)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_30),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_95),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_107),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_134),
.C(n_122),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_124),
.B(n_107),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_133),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_103),
.C(n_100),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_114),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_139),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_116),
.A2(n_108),
.B1(n_110),
.B2(n_100),
.Y(n_138)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_111),
.Y(n_139)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_141),
.A2(n_125),
.B(n_129),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_143),
.C(n_151),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_135),
.B(n_117),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_146),
.B(n_149),
.Y(n_157)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_121),
.C(n_119),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_17),
.C(n_32),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_120),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_137),
.B1(n_132),
.B2(n_133),
.Y(n_152)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_142),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_159),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_9),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_158),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_150),
.A2(n_17),
.B1(n_31),
.B2(n_12),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_2),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_10),
.Y(n_158)
);

AOI211xp5_ASAP7_75t_L g162 ( 
.A1(n_154),
.A2(n_148),
.B(n_3),
.C(n_4),
.Y(n_162)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

NOR2xp67_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_32),
.Y(n_164)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

AO21x2_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_159),
.B(n_3),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_165),
.A2(n_4),
.B(n_5),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_166),
.B(n_3),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_2),
.Y(n_167)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_167),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_170),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_168),
.A2(n_160),
.B1(n_165),
.B2(n_163),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_5),
.C(n_7),
.Y(n_176)
);

AOI21xp33_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_171),
.B(n_6),
.Y(n_175)
);

AOI222xp33_ASAP7_75t_SL g177 ( 
.A1(n_175),
.A2(n_176),
.B1(n_172),
.B2(n_7),
.C1(n_5),
.C2(n_31),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_31),
.Y(n_178)
);


endmodule