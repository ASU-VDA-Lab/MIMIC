module real_jpeg_1230_n_16 (n_5, n_4, n_8, n_0, n_12, n_398, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_397, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_398;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_397;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_0),
.B(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_0),
.B(n_38),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_0),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_0),
.B(n_104),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_0),
.B(n_86),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_0),
.B(n_25),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_0),
.B(n_27),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_0),
.B(n_47),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_1),
.Y(n_87)
);

BUFx4f_ASAP7_75t_L g104 ( 
.A(n_2),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_3),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_3),
.B(n_104),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_3),
.B(n_86),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_3),
.B(n_27),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_3),
.B(n_47),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_3),
.B(n_43),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_3),
.B(n_38),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_4),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_4),
.B(n_43),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_4),
.B(n_38),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_6),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_6),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_6),
.B(n_47),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_6),
.B(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_6),
.B(n_32),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_6),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_6),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_6),
.B(n_38),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_9),
.B(n_104),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_9),
.B(n_25),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_9),
.B(n_86),
.Y(n_154)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_9),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_9),
.B(n_43),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_9),
.B(n_38),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_9),
.B(n_32),
.Y(n_308)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_13),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_13),
.B(n_32),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_13),
.B(n_27),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_13),
.B(n_47),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_13),
.B(n_104),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_13),
.B(n_25),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_14),
.B(n_86),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_14),
.B(n_25),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_14),
.B(n_27),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_14),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_14),
.B(n_47),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_15),
.B(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_15),
.B(n_43),
.Y(n_56)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_15),
.B(n_38),
.Y(n_66)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_15),
.B(n_27),
.Y(n_95)
);

AND2x2_ASAP7_75t_SL g218 ( 
.A(n_15),
.B(n_86),
.Y(n_218)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_125),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_123),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_74),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_20),
.B(n_74),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_57),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_41),
.C(n_49),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_22),
.B(n_122),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_34),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_23),
.B(n_35),
.C(n_40),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_26),
.C(n_29),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_24),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_24),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_24),
.A2(n_29),
.B1(n_78),
.B2(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_24),
.B(n_81),
.C(n_83),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_24),
.A2(n_78),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_24),
.B(n_212),
.C(n_213),
.Y(n_249)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_25),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_26),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_26),
.B(n_53),
.C(n_56),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_26),
.A2(n_52),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_26),
.A2(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_26),
.B(n_255),
.Y(n_256)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_27),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_29),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_30),
.B(n_109),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_30),
.B(n_170),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_31),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_31),
.B(n_141),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_31),
.B(n_169),
.Y(n_275)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_40),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_36),
.B(n_85),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_37),
.B(n_169),
.Y(n_241)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_41),
.B(n_49),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_45),
.C(n_48),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_42),
.A2(n_45),
.B1(n_46),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_42),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_43),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_45),
.A2(n_46),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_46),
.B(n_103),
.C(n_218),
.Y(n_341)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_47),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_55),
.B2(n_56),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_54),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_53),
.A2(n_54),
.B1(n_274),
.B2(n_277),
.Y(n_273)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_54),
.B(n_201),
.C(n_275),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_83),
.C(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_55),
.A2(n_56),
.B1(n_90),
.B2(n_347),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_67),
.B1(n_72),
.B2(n_73),
.Y(n_59)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_63),
.A2(n_64),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_64),
.B(n_309),
.C(n_310),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_65),
.A2(n_66),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_66),
.B(n_95),
.C(n_97),
.Y(n_119)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_68),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_69),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_114),
.C(n_121),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_75),
.B(n_393),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_98),
.C(n_101),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_76),
.B(n_389),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_89),
.C(n_91),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_77),
.B(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_88),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_81),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_82),
.A2(n_83),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_82),
.B(n_200),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_82),
.A2(n_83),
.B1(n_346),
.B2(n_348),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_85),
.B(n_141),
.Y(n_171)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_89),
.B(n_91),
.Y(n_359)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_90),
.Y(n_347)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_94),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_95),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_95),
.A2(n_96),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_95),
.B(n_294),
.C(n_295),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_98),
.B(n_101),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_110),
.C(n_113),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_102),
.B(n_366),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.C(n_107),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_103),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_103),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_103),
.B(n_159),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_103),
.A2(n_158),
.B1(n_218),
.B2(n_220),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_103),
.A2(n_105),
.B1(n_158),
.B2(n_354),
.Y(n_353)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_105),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_106),
.B(n_109),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_107),
.A2(n_108),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_107),
.B(n_263),
.C(n_264),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_107),
.A2(n_108),
.B1(n_352),
.B2(n_353),
.Y(n_351)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_109),
.B(n_141),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_110),
.A2(n_113),
.B1(n_338),
.B2(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_110),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_112),
.B(n_169),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_113),
.A2(n_338),
.B1(n_339),
.B2(n_340),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_113),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_113),
.B(n_339),
.C(n_341),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_114),
.B(n_121),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_119),
.C(n_120),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_115),
.B(n_387),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_119),
.B(n_120),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI321xp33_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_383),
.A3(n_391),
.B1(n_394),
.B2(n_395),
.C(n_397),
.Y(n_125)
);

AOI321xp33_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_328),
.A3(n_372),
.B1(n_377),
.B2(n_382),
.C(n_398),
.Y(n_126)
);

NOR3xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_266),
.C(n_324),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_234),
.B(n_265),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_204),
.B(n_233),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_183),
.B(n_203),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_162),
.B(n_182),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_143),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_133),
.B(n_143),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_138),
.C(n_142),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_134),
.A2(n_135),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_135),
.A2(n_136),
.B(n_137),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_138),
.A2(n_139),
.B1(n_142),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_140),
.B(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_151),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_142),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_152),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_153),
.C(n_157),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_150),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_146),
.B(n_149),
.C(n_150),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_151),
.B(n_194),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_156),
.B1(n_157),
.B2(n_161),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_161),
.A2(n_175),
.B(n_176),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_173),
.B(n_181),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_167),
.B(n_172),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_165),
.B(n_166),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_174),
.B(n_177),
.Y(n_181)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_184),
.B(n_185),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_196),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_195),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_195),
.C(n_196),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_193),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_189),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_192),
.C(n_193),
.Y(n_221)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_190),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_202),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_199),
.C(n_202),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_200),
.A2(n_201),
.B1(n_275),
.B2(n_276),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_205),
.B(n_206),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_222),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_223),
.C(n_224),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_214),
.B2(n_215),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_216),
.C(n_221),
.Y(n_238)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_221),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_217),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_218),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_219),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_227),
.B2(n_232),
.Y(n_224)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_225),
.Y(n_232)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_231),
.C(n_232),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_230),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_235),
.B(n_236),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_252),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_250),
.B2(n_251),
.Y(n_237)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_238),
.Y(n_251)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_239),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_239),
.B(n_251),
.C(n_252),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_247),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_248),
.C(n_249),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_241),
.B(n_244),
.C(n_246),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_242)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_243),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_260),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_253)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_254),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_280),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_256),
.B(n_281),
.C(n_284),
.Y(n_315)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_257),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_258),
.C(n_260),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_264),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

AOI21xp33_ASAP7_75t_L g378 ( 
.A1(n_267),
.A2(n_379),
.B(n_380),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_297),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_268),
.B(n_297),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_285),
.C(n_286),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_269),
.B(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_270),
.B(n_272),
.C(n_279),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_278),
.B2(n_279),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_274),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_275),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_283),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_285),
.B(n_286),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_296),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_291),
.C(n_296),
.Y(n_313)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_295),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_293),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_323),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_312),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_299),
.B(n_312),
.C(n_323),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_303),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_300),
.B(n_304),
.C(n_305),
.Y(n_332)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_308),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_309),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_313),
.B(n_315),
.C(n_316),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_322),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_319),
.B1(n_320),
.B2(n_321),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_318),
.B(n_321),
.C(n_322),
.Y(n_335)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_320),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_325),
.B(n_326),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_356),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_329),
.B(n_356),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_342),
.C(n_355),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_330),
.B(n_342),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_332),
.B1(n_333),
.B2(n_334),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_331),
.B(n_335),
.C(n_336),
.Y(n_369)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_341),
.Y(n_336)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_339),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_351),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_344),
.A2(n_345),
.B1(n_349),
.B2(n_350),
.Y(n_343)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_344),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_344),
.B(n_350),
.C(n_351),
.Y(n_362)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_345),
.Y(n_350)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_346),
.Y(n_348)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_355),
.B(n_376),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_357),
.A2(n_369),
.B1(n_370),
.B2(n_371),
.Y(n_356)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_357),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_360),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_358),
.B(n_360),
.C(n_371),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_362),
.B1(n_363),
.B2(n_368),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_361),
.B(n_364),
.C(n_365),
.Y(n_390)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_363),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_369),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_373),
.A2(n_378),
.B(n_381),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_374),
.B(n_375),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_385),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_384),
.B(n_385),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_385),
.B(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_385),
.B(n_392),
.Y(n_395)
);

FAx1_ASAP7_75t_SL g385 ( 
.A(n_386),
.B(n_388),
.CI(n_390),
.CON(n_385),
.SN(n_385)
);


endmodule