module fake_jpeg_9663_n_276 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_276);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_276;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_1),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_21),
.B(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_41),
.Y(n_46)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_45),
.B(n_32),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_29),
.Y(n_48)
);

OAI21xp33_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_2),
.B(n_3),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_31),
.B1(n_29),
.B2(n_17),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_50),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_69)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

AO21x1_ASAP7_75t_L g83 ( 
.A1(n_51),
.A2(n_53),
.B(n_56),
.Y(n_83)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_31),
.B1(n_18),
.B2(n_25),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_21),
.B1(n_22),
.B2(n_27),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_26),
.B1(n_20),
.B2(n_24),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_43),
.C(n_22),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_27),
.C(n_24),
.Y(n_94)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_18),
.B1(n_23),
.B2(n_32),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_65),
.A2(n_96),
.B1(n_9),
.B2(n_10),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_66),
.B(n_75),
.Y(n_110)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_33),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_68),
.B(n_74),
.Y(n_103)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_94),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_72),
.Y(n_123)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_73),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_33),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_33),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_76),
.B(n_82),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_2),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_77),
.A2(n_92),
.B(n_4),
.Y(n_112)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_48),
.B(n_16),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_2),
.Y(n_84)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_85),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_52),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_87),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_45),
.B(n_15),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_27),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_5),
.C(n_6),
.Y(n_115)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_3),
.Y(n_90)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_4),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_47),
.B(n_4),
.Y(n_93)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_52),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_98),
.B1(n_99),
.B2(n_43),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_47),
.A2(n_28),
.B1(n_26),
.B2(n_24),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_51),
.Y(n_98)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_61),
.A2(n_28),
.B1(n_26),
.B2(n_20),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_28),
.B1(n_34),
.B2(n_30),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_104),
.A2(n_80),
.B1(n_70),
.B2(n_78),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_108),
.B(n_85),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_112),
.B(n_114),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_66),
.A2(n_34),
.B1(n_30),
.B2(n_8),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_114),
.A2(n_88),
.B1(n_99),
.B2(n_73),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_117),
.C(n_112),
.Y(n_148)
);

MAJx2_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_5),
.C(n_6),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_67),
.A2(n_16),
.B1(n_6),
.B2(n_8),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_121),
.B1(n_128),
.B2(n_87),
.Y(n_137)
);

OAI32xp33_ASAP7_75t_L g121 ( 
.A1(n_82),
.A2(n_5),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_122),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_94),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_106),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_133),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_132),
.Y(n_179)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_134),
.A2(n_138),
.B(n_148),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_77),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_139),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_136),
.A2(n_150),
.B1(n_151),
.B2(n_131),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_137),
.B(n_140),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_95),
.B(n_86),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_92),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_81),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_141),
.Y(n_170)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_144),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_143),
.Y(n_182)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_102),
.A2(n_69),
.B1(n_100),
.B2(n_83),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_145),
.A2(n_156),
.B1(n_129),
.B2(n_126),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_92),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_146),
.A2(n_154),
.B(n_119),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_111),
.B(n_83),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_152),
.Y(n_160)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_109),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_104),
.A2(n_69),
.B1(n_101),
.B2(n_91),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_102),
.B(n_81),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_101),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_157),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_120),
.A2(n_79),
.B(n_89),
.Y(n_154)
);

AO21x1_ASAP7_75t_L g167 ( 
.A1(n_155),
.A2(n_126),
.B(n_105),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_79),
.B1(n_97),
.B2(n_72),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_113),
.B(n_97),
.Y(n_157)
);

NAND2xp33_ASAP7_75t_SL g158 ( 
.A(n_107),
.B(n_85),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_158),
.A2(n_123),
.B(n_127),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_169),
.B1(n_183),
.B2(n_151),
.Y(n_189)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_162),
.B(n_165),
.Y(n_186)
);

NAND2x1_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_121),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_163),
.A2(n_173),
.B(n_184),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_115),
.C(n_120),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_146),
.C(n_136),
.Y(n_201)
);

AO21x1_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_133),
.B(n_158),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_145),
.A2(n_105),
.B1(n_113),
.B2(n_119),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_157),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_172),
.B(n_174),
.Y(n_202)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_176),
.A2(n_182),
.B1(n_164),
.B2(n_181),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_130),
.B(n_125),
.Y(n_178)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_180),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_127),
.Y(n_181)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_185),
.Y(n_200)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_182),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_204),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_189),
.A2(n_176),
.B1(n_171),
.B2(n_182),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_148),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_195),
.C(n_201),
.Y(n_216)
);

AOI22x1_ASAP7_75t_L g217 ( 
.A1(n_194),
.A2(n_167),
.B1(n_184),
.B2(n_179),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_135),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_185),
.A2(n_134),
.B(n_147),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_196),
.A2(n_197),
.B(n_205),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_171),
.A2(n_146),
.B(n_137),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_142),
.Y(n_198)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_198),
.Y(n_210)
);

INVx13_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_177),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_178),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_164),
.Y(n_206)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_207),
.A2(n_161),
.B1(n_168),
.B2(n_162),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_195),
.B(n_173),
.Y(n_208)
);

NAND3xp33_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_159),
.C(n_193),
.Y(n_230)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_207),
.A2(n_168),
.B1(n_169),
.B2(n_163),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_211),
.A2(n_215),
.B1(n_223),
.B2(n_205),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_217),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_199),
.A2(n_179),
.B1(n_172),
.B2(n_167),
.Y(n_220)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_220),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_166),
.Y(n_221)
);

BUFx12_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_192),
.A2(n_174),
.B1(n_170),
.B2(n_160),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_224),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_159),
.C(n_160),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_225),
.B(n_206),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_190),
.C(n_225),
.Y(n_247)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_230),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_231),
.A2(n_211),
.B1(n_200),
.B2(n_220),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_188),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_188),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_234),
.A2(n_238),
.B(n_239),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_209),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_236),
.B(n_237),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_210),
.B(n_170),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_192),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_216),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_248),
.Y(n_254)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_243),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_216),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_212),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_247),
.B(n_190),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_221),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_208),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_228),
.C(n_235),
.Y(n_253)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_229),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_232),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_252),
.A2(n_246),
.B(n_200),
.Y(n_261)
);

MAJx2_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_256),
.C(n_197),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_255),
.B(n_257),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_242),
.B(n_229),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_240),
.C(n_238),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_258),
.A2(n_246),
.B(n_228),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_251),
.A2(n_244),
.B(n_239),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_261),
.Y(n_267)
);

NOR2xp67_ASAP7_75t_L g260 ( 
.A(n_258),
.B(n_217),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_189),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_262),
.A2(n_213),
.B1(n_253),
.B2(n_254),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_196),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_193),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_268),
.Y(n_271)
);

AOI322xp5_ASAP7_75t_L g269 ( 
.A1(n_267),
.A2(n_264),
.A3(n_186),
.B1(n_254),
.B2(n_249),
.C1(n_233),
.C2(n_194),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_269),
.A2(n_149),
.B(n_153),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_270),
.B(n_233),
.C(n_144),
.Y(n_272)
);

OA21x2_ASAP7_75t_L g274 ( 
.A1(n_272),
.A2(n_273),
.B(n_271),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_274),
.A2(n_85),
.B(n_12),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_275),
.B(n_14),
.Y(n_276)
);


endmodule