module real_aes_8922_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_393;
wire n_294;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g275 ( .A(n_0), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g151 ( .A1(n_1), .A2(n_50), .B1(n_152), .B2(n_158), .Y(n_151) );
AOI21xp33_ASAP7_75t_L g217 ( .A1(n_2), .A2(n_218), .B(n_224), .Y(n_217) );
INVx1_ASAP7_75t_L g198 ( .A(n_3), .Y(n_198) );
AND2x6_ASAP7_75t_L g223 ( .A(n_3), .B(n_196), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_3), .B(n_531), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_4), .A2(n_316), .B(n_317), .Y(n_315) );
INVx1_ASAP7_75t_L g234 ( .A(n_5), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_6), .B(n_308), .Y(n_307) );
AO22x2_ASAP7_75t_L g91 ( .A1(n_7), .A2(n_22), .B1(n_92), .B2(n_93), .Y(n_91) );
INVx1_ASAP7_75t_L g216 ( .A(n_8), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_9), .A2(n_178), .B1(n_184), .B2(n_185), .Y(n_177) );
INVx1_ASAP7_75t_L g184 ( .A(n_9), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_10), .B(n_263), .Y(n_336) );
AO22x2_ASAP7_75t_L g95 ( .A1(n_11), .A2(n_24), .B1(n_92), .B2(n_96), .Y(n_95) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_12), .B(n_218), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_13), .B(n_209), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g319 ( .A1(n_14), .A2(n_320), .B(n_321), .C(n_322), .Y(n_319) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_15), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_16), .A2(n_80), .B1(n_81), .B2(n_176), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_16), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_17), .B(n_232), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g116 ( .A1(n_18), .A2(n_20), .B1(n_117), .B2(n_124), .Y(n_116) );
INVx1_ASAP7_75t_L g253 ( .A(n_19), .Y(n_253) );
INVx2_ASAP7_75t_L g221 ( .A(n_21), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_23), .Y(n_133) );
OAI221xp5_ASAP7_75t_L g189 ( .A1(n_24), .A2(n_34), .B1(n_43), .B2(n_190), .C(n_191), .Y(n_189) );
INVxp67_ASAP7_75t_L g192 ( .A(n_24), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_L g288 ( .A1(n_25), .A2(n_223), .B(n_227), .C(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g251 ( .A(n_26), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g335 ( .A(n_27), .B(n_232), .Y(n_335) );
OAI22xp5_ASAP7_75t_SL g181 ( .A1(n_28), .A2(n_76), .B1(n_182), .B2(n_183), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_28), .Y(n_182) );
CKINVDCx16_ASAP7_75t_R g254 ( .A(n_29), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_30), .B(n_218), .Y(n_310) );
AOI22xp5_ASAP7_75t_L g246 ( .A1(n_31), .A2(n_227), .B1(n_247), .B2(n_249), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g297 ( .A(n_32), .Y(n_297) );
CKINVDCx16_ASAP7_75t_R g272 ( .A(n_33), .Y(n_272) );
AO22x2_ASAP7_75t_L g101 ( .A1(n_34), .A2(n_54), .B1(n_92), .B2(n_96), .Y(n_101) );
INVxp67_ASAP7_75t_L g193 ( .A(n_34), .Y(n_193) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_35), .A2(n_231), .B(n_233), .C(n_236), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g162 ( .A1(n_36), .A2(n_45), .B1(n_163), .B2(n_167), .Y(n_162) );
INVx1_ASAP7_75t_L g225 ( .A(n_37), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g339 ( .A(n_38), .Y(n_339) );
INVx1_ASAP7_75t_L g196 ( .A(n_39), .Y(n_196) );
INVx1_ASAP7_75t_L g215 ( .A(n_40), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_41), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g85 ( .A(n_42), .Y(n_85) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_43), .A2(n_59), .B1(n_92), .B2(n_93), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_44), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_SL g262 ( .A1(n_46), .A2(n_236), .B(n_263), .C(n_264), .Y(n_262) );
INVxp67_ASAP7_75t_L g265 ( .A(n_47), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_48), .Y(n_257) );
INVx1_ASAP7_75t_L g332 ( .A(n_49), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g143 ( .A1(n_51), .A2(n_63), .B1(n_144), .B2(n_147), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g333 ( .A1(n_52), .A2(n_223), .B(n_227), .C(n_334), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_53), .A2(n_179), .B1(n_180), .B2(n_181), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_53), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_55), .B(n_276), .Y(n_290) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_55), .A2(n_80), .B1(n_81), .B2(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_55), .Y(n_527) );
INVx2_ASAP7_75t_L g213 ( .A(n_56), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_57), .B(n_263), .Y(n_291) );
INVx1_ASAP7_75t_L g536 ( .A(n_57), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_L g273 ( .A1(n_58), .A2(n_223), .B(n_227), .C(n_274), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g171 ( .A1(n_60), .A2(n_70), .B1(n_172), .B2(n_174), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_61), .B(n_240), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g280 ( .A(n_62), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_L g304 ( .A1(n_64), .A2(n_223), .B(n_227), .C(n_305), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g312 ( .A(n_65), .Y(n_312) );
INVx1_ASAP7_75t_L g261 ( .A(n_66), .Y(n_261) );
CKINVDCx16_ASAP7_75t_R g318 ( .A(n_67), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_68), .B(n_276), .Y(n_306) );
INVx1_ASAP7_75t_L g92 ( .A(n_69), .Y(n_92) );
INVx1_ASAP7_75t_L g94 ( .A(n_69), .Y(n_94) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_71), .B(n_211), .Y(n_323) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_72), .Y(n_102) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_73), .A2(n_218), .B(n_260), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_74), .Y(n_109) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_75), .A2(n_80), .B1(n_81), .B2(n_538), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_75), .Y(n_538) );
INVx1_ASAP7_75t_L g183 ( .A(n_76), .Y(n_183) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_186), .B1(n_199), .B2(n_517), .C(n_525), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_177), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NAND2xp5_ASAP7_75t_L g82 ( .A(n_83), .B(n_141), .Y(n_82) );
NOR3xp33_ASAP7_75t_L g83 ( .A(n_84), .B(n_108), .C(n_127), .Y(n_83) );
OAI22xp5_ASAP7_75t_L g84 ( .A1(n_85), .A2(n_86), .B1(n_102), .B2(n_103), .Y(n_84) );
INVx1_ASAP7_75t_SL g86 ( .A(n_87), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
OR2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_97), .Y(n_88) );
INVx2_ASAP7_75t_L g166 ( .A(n_89), .Y(n_166) );
OR2x2_ASAP7_75t_L g89 ( .A(n_90), .B(n_95), .Y(n_89) );
AND2x2_ASAP7_75t_L g107 ( .A(n_90), .B(n_95), .Y(n_107) );
AND2x2_ASAP7_75t_L g146 ( .A(n_90), .B(n_122), .Y(n_146) );
INVx2_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
AND2x2_ASAP7_75t_L g113 ( .A(n_91), .B(n_95), .Y(n_113) );
AND2x2_ASAP7_75t_L g123 ( .A(n_91), .B(n_101), .Y(n_123) );
INVx1_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx1_ASAP7_75t_L g96 ( .A(n_94), .Y(n_96) );
INVx2_ASAP7_75t_L g122 ( .A(n_95), .Y(n_122) );
INVx1_ASAP7_75t_L g160 ( .A(n_95), .Y(n_160) );
INVx1_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
NAND2x1p5_ASAP7_75t_L g106 ( .A(n_98), .B(n_107), .Y(n_106) );
AND2x4_ASAP7_75t_L g170 ( .A(n_98), .B(n_146), .Y(n_170) );
AND2x2_ASAP7_75t_L g98 ( .A(n_99), .B(n_100), .Y(n_98) );
INVx1_ASAP7_75t_L g115 ( .A(n_99), .Y(n_115) );
INVx1_ASAP7_75t_L g121 ( .A(n_99), .Y(n_121) );
INVx1_ASAP7_75t_L g140 ( .A(n_99), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_99), .B(n_101), .Y(n_150) );
AND2x2_ASAP7_75t_L g114 ( .A(n_100), .B(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
AND2x2_ASAP7_75t_L g157 ( .A(n_101), .B(n_140), .Y(n_157) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
BUFx3_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g156 ( .A(n_107), .B(n_157), .Y(n_156) );
AND2x4_ASAP7_75t_L g173 ( .A(n_107), .B(n_114), .Y(n_173) );
OAI21xp33_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_110), .B(n_116), .Y(n_108) );
BUFx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx4_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x6_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
INVx1_ASAP7_75t_L g137 ( .A(n_113), .Y(n_137) );
AND2x2_ASAP7_75t_L g145 ( .A(n_114), .B(n_146), .Y(n_145) );
AND2x6_ASAP7_75t_L g165 ( .A(n_114), .B(n_166), .Y(n_165) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x4_ASAP7_75t_L g119 ( .A(n_120), .B(n_123), .Y(n_119) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
INVx1_ASAP7_75t_L g126 ( .A(n_121), .Y(n_126) );
INVx1_ASAP7_75t_L g132 ( .A(n_122), .Y(n_132) );
AND2x4_ASAP7_75t_L g125 ( .A(n_123), .B(n_126), .Y(n_125) );
NAND2x1p5_ASAP7_75t_L g131 ( .A(n_123), .B(n_132), .Y(n_131) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI22xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_129), .B1(n_133), .B2(n_134), .Y(n_127) );
INVx3_ASAP7_75t_SL g129 ( .A(n_130), .Y(n_129) );
INVx4_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
CKINVDCx16_ASAP7_75t_R g135 ( .A(n_136), .Y(n_135) );
OR2x6_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_142), .B(n_161), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_151), .Y(n_142) );
BUFx2_ASAP7_75t_SL g144 ( .A(n_145), .Y(n_144) );
AND2x4_ASAP7_75t_L g148 ( .A(n_146), .B(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g175 ( .A(n_146), .B(n_157), .Y(n_175) );
BUFx2_ASAP7_75t_SL g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
OR2x6_ASAP7_75t_L g159 ( .A(n_150), .B(n_160), .Y(n_159) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx4_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx8_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_162), .B(n_171), .Y(n_161) );
INVx2_ASAP7_75t_SL g163 ( .A(n_164), .Y(n_163) );
INVx11_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx4_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx4_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
BUFx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
BUFx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_178), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_181), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_184), .B(n_320), .Y(n_321) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_187), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_188), .Y(n_187) );
AND3x1_ASAP7_75t_SL g188 ( .A(n_189), .B(n_194), .C(n_197), .Y(n_188) );
INVxp67_ASAP7_75t_L g531 ( .A(n_189), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_192), .B(n_193), .Y(n_191) );
INVx1_ASAP7_75t_SL g532 ( .A(n_194), .Y(n_532) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_194), .A2(n_520), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g542 ( .A(n_194), .Y(n_542) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_195), .B(n_198), .Y(n_535) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
OR2x2_ASAP7_75t_SL g541 ( .A(n_197), .B(n_542), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_198), .Y(n_197) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND3x1_ASAP7_75t_L g203 ( .A(n_204), .B(n_439), .C(n_484), .Y(n_203) );
NOR4xp25_ASAP7_75t_L g204 ( .A(n_205), .B(n_362), .C(n_403), .D(n_420), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_267), .B(n_283), .C(n_324), .Y(n_205) );
OR2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_241), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_207), .B(n_268), .Y(n_267) );
NOR4xp25_ASAP7_75t_L g386 ( .A(n_207), .B(n_380), .C(n_387), .D(n_393), .Y(n_386) );
AND2x2_ASAP7_75t_L g459 ( .A(n_207), .B(n_348), .Y(n_459) );
AND2x2_ASAP7_75t_L g478 ( .A(n_207), .B(n_424), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_207), .B(n_473), .Y(n_487) );
AND2x2_ASAP7_75t_L g500 ( .A(n_207), .B(n_282), .Y(n_500) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx1_ASAP7_75t_SL g345 ( .A(n_208), .Y(n_345) );
AND2x2_ASAP7_75t_L g352 ( .A(n_208), .B(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g402 ( .A(n_208), .B(n_242), .Y(n_402) );
AND2x2_ASAP7_75t_SL g413 ( .A(n_208), .B(n_348), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_208), .B(n_242), .Y(n_417) );
AND2x2_ASAP7_75t_L g426 ( .A(n_208), .B(n_351), .Y(n_426) );
BUFx2_ASAP7_75t_L g449 ( .A(n_208), .Y(n_449) );
AND2x2_ASAP7_75t_L g453 ( .A(n_208), .B(n_258), .Y(n_453) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_217), .B(n_239), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_SL g296 ( .A(n_210), .B(n_297), .Y(n_296) );
INVx4_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
OA21x2_ASAP7_75t_L g258 ( .A1(n_211), .A2(n_259), .B(n_266), .Y(n_258) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g244 ( .A(n_212), .Y(n_244) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
AND2x2_ASAP7_75t_SL g240 ( .A(n_213), .B(n_214), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
BUFx2_ASAP7_75t_L g316 ( .A(n_218), .Y(n_316) );
AND2x4_ASAP7_75t_L g218 ( .A(n_219), .B(n_223), .Y(n_218) );
NAND2x1p5_ASAP7_75t_L g255 ( .A(n_219), .B(n_223), .Y(n_255) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_222), .Y(n_219) );
INVx1_ASAP7_75t_L g522 ( .A(n_220), .Y(n_522) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g228 ( .A(n_221), .Y(n_228) );
INVx1_ASAP7_75t_L g248 ( .A(n_221), .Y(n_248) );
INVx1_ASAP7_75t_L g229 ( .A(n_222), .Y(n_229) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_222), .Y(n_232) );
INVx3_ASAP7_75t_L g235 ( .A(n_222), .Y(n_235) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_222), .Y(n_250) );
INVx1_ASAP7_75t_L g263 ( .A(n_222), .Y(n_263) );
INVx4_ASAP7_75t_SL g238 ( .A(n_223), .Y(n_238) );
BUFx3_ASAP7_75t_L g519 ( .A(n_223), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_230), .C(n_238), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g260 ( .A1(n_226), .A2(n_238), .B(n_261), .C(n_262), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_L g317 ( .A1(n_226), .A2(n_238), .B(n_318), .C(n_319), .Y(n_317) );
INVx5_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x6_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_228), .Y(n_237) );
BUFx3_ASAP7_75t_L g294 ( .A(n_228), .Y(n_294) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx4_ASAP7_75t_L g308 ( .A(n_232), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_235), .B(n_265), .Y(n_264) );
INVx5_ASAP7_75t_L g276 ( .A(n_235), .Y(n_276) );
INVx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_237), .Y(n_309) );
OAI22xp33_ASAP7_75t_L g245 ( .A1(n_238), .A2(n_246), .B1(n_254), .B2(n_255), .Y(n_245) );
INVx1_ASAP7_75t_L g281 ( .A(n_240), .Y(n_281) );
INVx2_ASAP7_75t_L g302 ( .A(n_240), .Y(n_302) );
OA21x2_ASAP7_75t_L g314 ( .A1(n_240), .A2(n_315), .B(n_323), .Y(n_314) );
OR2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_258), .Y(n_241) );
AND2x2_ASAP7_75t_L g282 ( .A(n_242), .B(n_258), .Y(n_282) );
BUFx2_ASAP7_75t_L g355 ( .A(n_242), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_242), .A2(n_388), .B1(n_390), .B2(n_391), .Y(n_387) );
OR2x2_ASAP7_75t_L g409 ( .A(n_242), .B(n_270), .Y(n_409) );
AND2x2_ASAP7_75t_L g473 ( .A(n_242), .B(n_351), .Y(n_473) );
INVx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g341 ( .A(n_243), .B(n_270), .Y(n_341) );
AND2x2_ASAP7_75t_L g348 ( .A(n_243), .B(n_258), .Y(n_348) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_243), .Y(n_390) );
OR2x2_ASAP7_75t_L g425 ( .A(n_243), .B(n_269), .Y(n_425) );
AO21x2_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_256), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_244), .B(n_257), .Y(n_256) );
AO21x2_ASAP7_75t_L g270 ( .A1(n_244), .A2(n_271), .B(n_279), .Y(n_270) );
INVx2_ASAP7_75t_L g295 ( .A(n_244), .Y(n_295) );
INVx2_ASAP7_75t_L g278 ( .A(n_247), .Y(n_278) );
INVx3_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
OAI22xp5_ASAP7_75t_SL g249 ( .A1(n_250), .A2(n_251), .B1(n_252), .B2(n_253), .Y(n_249) );
INVx2_ASAP7_75t_L g252 ( .A(n_250), .Y(n_252) );
INVx4_ASAP7_75t_L g320 ( .A(n_250), .Y(n_320) );
INVx2_ASAP7_75t_L g524 ( .A(n_252), .Y(n_524) );
OAI21xp5_ASAP7_75t_L g271 ( .A1(n_255), .A2(n_272), .B(n_273), .Y(n_271) );
OAI21xp5_ASAP7_75t_L g331 ( .A1(n_255), .A2(n_332), .B(n_333), .Y(n_331) );
INVx1_ASAP7_75t_L g344 ( .A(n_258), .Y(n_344) );
INVx3_ASAP7_75t_L g353 ( .A(n_258), .Y(n_353) );
BUFx2_ASAP7_75t_L g377 ( .A(n_258), .Y(n_377) );
AND2x2_ASAP7_75t_L g410 ( .A(n_258), .B(n_345), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_267), .A2(n_496), .B1(n_497), .B2(n_498), .Y(n_495) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_282), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_269), .B(n_353), .Y(n_357) );
INVx1_ASAP7_75t_L g385 ( .A(n_269), .Y(n_385) );
INVx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx3_ASAP7_75t_L g351 ( .A(n_270), .Y(n_351) );
O2A1O1Ixp33_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_276), .B(n_277), .C(n_278), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_281), .B(n_312), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_281), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g363 ( .A(n_282), .Y(n_363) );
NAND2x1_ASAP7_75t_SL g283 ( .A(n_284), .B(n_298), .Y(n_283) );
AND2x2_ASAP7_75t_L g361 ( .A(n_284), .B(n_313), .Y(n_361) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_284), .Y(n_435) );
AND2x2_ASAP7_75t_L g462 ( .A(n_284), .B(n_382), .Y(n_462) );
AND2x2_ASAP7_75t_L g470 ( .A(n_284), .B(n_432), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_284), .B(n_327), .Y(n_497) );
INVx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g328 ( .A(n_285), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g346 ( .A(n_285), .B(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g367 ( .A(n_285), .Y(n_367) );
INVx1_ASAP7_75t_L g373 ( .A(n_285), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_285), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g406 ( .A(n_285), .B(n_330), .Y(n_406) );
OR2x2_ASAP7_75t_L g444 ( .A(n_285), .B(n_399), .Y(n_444) );
AOI32xp33_ASAP7_75t_L g456 ( .A1(n_285), .A2(n_457), .A3(n_460), .B1(n_461), .B2(n_462), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_285), .B(n_432), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_285), .B(n_392), .Y(n_507) );
OR2x6_ASAP7_75t_L g285 ( .A(n_286), .B(n_296), .Y(n_285) );
AOI21xp5_ASAP7_75t_SL g286 ( .A1(n_287), .A2(n_288), .B(n_295), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_291), .B(n_292), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_292), .A2(n_335), .B(n_336), .Y(n_334) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g322 ( .A(n_294), .Y(n_322) );
INVx1_ASAP7_75t_L g337 ( .A(n_295), .Y(n_337) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g418 ( .A(n_299), .B(n_419), .Y(n_418) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_313), .Y(n_299) );
INVx1_ASAP7_75t_L g380 ( .A(n_300), .Y(n_380) );
AND2x2_ASAP7_75t_L g382 ( .A(n_300), .B(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_300), .B(n_329), .Y(n_399) );
AND2x2_ASAP7_75t_L g432 ( .A(n_300), .B(n_408), .Y(n_432) );
AND2x2_ASAP7_75t_L g469 ( .A(n_300), .B(n_330), .Y(n_469) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g327 ( .A(n_301), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_301), .B(n_329), .Y(n_359) );
AND2x2_ASAP7_75t_L g366 ( .A(n_301), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g407 ( .A(n_301), .B(n_408), .Y(n_407) );
AO21x2_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_303), .B(n_311), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_310), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_307), .B(n_309), .Y(n_305) );
INVx2_ASAP7_75t_L g383 ( .A(n_313), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_313), .B(n_329), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_313), .B(n_374), .Y(n_455) );
INVx1_ASAP7_75t_L g477 ( .A(n_313), .Y(n_477) );
INVx1_ASAP7_75t_L g494 ( .A(n_313), .Y(n_494) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g347 ( .A(n_314), .B(n_329), .Y(n_347) );
AND2x2_ASAP7_75t_L g369 ( .A(n_314), .B(n_330), .Y(n_369) );
INVx1_ASAP7_75t_L g408 ( .A(n_314), .Y(n_408) );
AOI221x1_ASAP7_75t_SL g324 ( .A1(n_325), .A2(n_340), .B1(n_346), .B2(n_348), .C(n_349), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_325), .A2(n_413), .B1(n_480), .B2(n_481), .Y(n_479) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
AND2x2_ASAP7_75t_L g371 ( .A(n_326), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g466 ( .A(n_326), .B(n_346), .Y(n_466) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g422 ( .A(n_327), .B(n_347), .Y(n_422) );
INVx1_ASAP7_75t_L g434 ( .A(n_328), .Y(n_434) );
AND2x2_ASAP7_75t_L g445 ( .A(n_328), .B(n_432), .Y(n_445) );
AND2x2_ASAP7_75t_L g512 ( .A(n_328), .B(n_407), .Y(n_512) );
INVx2_ASAP7_75t_L g374 ( .A(n_329), .Y(n_374) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AO21x2_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_337), .B(n_338), .Y(n_330) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_341), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g464 ( .A(n_341), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_342), .B(n_425), .Y(n_428) );
INVx3_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_343), .A2(n_464), .B(n_509), .Y(n_508) );
AND2x4_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
NOR2xp33_ASAP7_75t_SL g486 ( .A(n_346), .B(n_372), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_347), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g438 ( .A(n_347), .B(n_366), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_347), .B(n_373), .Y(n_515) );
AND2x2_ASAP7_75t_L g384 ( .A(n_348), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g451 ( .A(n_348), .Y(n_451) );
AOI21xp33_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_354), .B(n_358), .Y(n_349) );
NAND2x1_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_351), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g400 ( .A(n_351), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g412 ( .A(n_351), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_351), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g436 ( .A(n_352), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_352), .B(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_352), .B(n_355), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
AOI211xp5_ASAP7_75t_L g423 ( .A1(n_355), .A2(n_394), .B(n_424), .C(n_426), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g441 ( .A1(n_355), .A2(n_442), .B1(n_445), .B2(n_446), .C(n_450), .Y(n_441) );
AND2x2_ASAP7_75t_L g437 ( .A(n_356), .B(n_390), .Y(n_437) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g397 ( .A(n_361), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g468 ( .A(n_361), .B(n_469), .Y(n_468) );
OAI211xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B(n_370), .C(n_395), .Y(n_362) );
NAND3xp33_ASAP7_75t_SL g481 ( .A(n_363), .B(n_482), .C(n_483), .Y(n_481) );
OR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_368), .Y(n_364) );
OR2x2_ASAP7_75t_L g454 ( .A(n_365), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AOI221xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_375), .B1(n_378), .B2(n_384), .C(n_386), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_372), .B(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_372), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g394 ( .A(n_377), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_377), .A2(n_434), .B1(n_435), .B2(n_436), .Y(n_433) );
OR2x2_ASAP7_75t_L g514 ( .A(n_377), .B(n_425), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g378 ( .A(n_379), .B(n_381), .Y(n_378) );
INVxp67_ASAP7_75t_L g488 ( .A(n_380), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_382), .B(n_503), .Y(n_502) );
INVxp67_ASAP7_75t_L g389 ( .A(n_383), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_385), .B(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_385), .B(n_432), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_385), .B(n_452), .Y(n_491) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_389), .Y(n_415) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g505 ( .A(n_394), .B(n_425), .Y(n_505) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_400), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_SL g483 ( .A(n_400), .Y(n_483) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OAI322xp33_ASAP7_75t_SL g403 ( .A1(n_404), .A2(n_409), .A3(n_410), .B1(n_411), .B2(n_414), .C1(n_416), .C2(n_418), .Y(n_403) );
OAI322xp33_ASAP7_75t_L g485 ( .A1(n_404), .A2(n_486), .A3(n_487), .B1(n_488), .B2(n_489), .C1(n_490), .C2(n_492), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g404 ( .A(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
INVx4_ASAP7_75t_L g419 ( .A(n_406), .Y(n_419) );
AND2x2_ASAP7_75t_L g480 ( .A(n_406), .B(n_432), .Y(n_480) );
AND2x2_ASAP7_75t_L g493 ( .A(n_406), .B(n_494), .Y(n_493) );
CKINVDCx16_ASAP7_75t_R g504 ( .A(n_409), .Y(n_504) );
INVx1_ASAP7_75t_L g482 ( .A(n_410), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
OR2x2_ASAP7_75t_L g416 ( .A(n_412), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g499 ( .A(n_412), .B(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_412), .B(n_453), .Y(n_510) );
OR2x2_ASAP7_75t_L g443 ( .A(n_415), .B(n_444), .Y(n_443) );
INVxp33_ASAP7_75t_L g460 ( .A(n_415), .Y(n_460) );
OAI221xp5_ASAP7_75t_SL g420 ( .A1(n_419), .A2(n_421), .B1(n_423), .B2(n_427), .C(n_429), .Y(n_420) );
NOR2xp67_ASAP7_75t_L g476 ( .A(n_419), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g503 ( .A(n_419), .Y(n_503) );
INVx1_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
INVx3_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
AOI322xp5_ASAP7_75t_L g467 ( .A1(n_426), .A2(n_451), .A3(n_468), .B1(n_470), .B2(n_471), .C1(n_474), .C2(n_478), .Y(n_467) );
INVxp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_433), .B1(n_437), .B2(n_438), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_440), .B(n_463), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_441), .B(n_456), .Y(n_440) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_444), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
NAND2xp33_ASAP7_75t_SL g461 ( .A(n_447), .B(n_458), .Y(n_461) );
INVx1_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
OAI322xp33_ASAP7_75t_L g501 ( .A1(n_449), .A2(n_502), .A3(n_504), .B1(n_505), .B2(n_506), .C1(n_508), .C2(n_511), .Y(n_501) );
AOI21xp33_ASAP7_75t_SL g450 ( .A1(n_451), .A2(n_452), .B(n_454), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_459), .B(n_507), .Y(n_516) );
OAI211xp5_ASAP7_75t_SL g463 ( .A1(n_464), .A2(n_465), .B(n_467), .C(n_479), .Y(n_463) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NOR4xp25_ASAP7_75t_L g484 ( .A(n_485), .B(n_495), .C(n_501), .D(n_513), .Y(n_484) );
INVxp67_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
INVxp67_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
CKINVDCx14_ASAP7_75t_R g511 ( .A(n_512), .Y(n_511) );
OAI21xp5_ASAP7_75t_SL g513 ( .A1(n_514), .A2(n_515), .B(n_516), .Y(n_513) );
CKINVDCx16_ASAP7_75t_R g517 ( .A(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_523), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
OAI322xp33_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_528), .A3(n_532), .B1(n_533), .B2(n_536), .C1(n_537), .C2(n_539), .Y(n_525) );
INVx1_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_530), .Y(n_529) );
CKINVDCx16_ASAP7_75t_R g533 ( .A(n_534), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_540), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_541), .Y(n_540) );
endmodule