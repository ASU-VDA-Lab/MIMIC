module fake_netlist_1_6577_n_35 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_35);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_35;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
NOR2xp33_ASAP7_75t_R g11 ( .A(n_4), .B(n_3), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_9), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_9), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_4), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_10), .Y(n_15) );
NAND2xp5_ASAP7_75t_SL g16 ( .A(n_6), .B(n_0), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_13), .B(n_0), .Y(n_17) );
OAI21xp5_ASAP7_75t_L g18 ( .A1(n_12), .A2(n_0), .B(n_1), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_13), .B(n_10), .Y(n_19) );
BUFx3_ASAP7_75t_L g20 ( .A(n_12), .Y(n_20) );
NOR2xp33_ASAP7_75t_L g21 ( .A(n_15), .B(n_1), .Y(n_21) );
HB1xp67_ASAP7_75t_L g22 ( .A(n_17), .Y(n_22) );
INVx2_ASAP7_75t_SL g23 ( .A(n_20), .Y(n_23) );
NOR2xp33_ASAP7_75t_L g24 ( .A(n_20), .B(n_14), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_22), .B(n_19), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_23), .B(n_18), .Y(n_26) );
INVx5_ASAP7_75t_SL g27 ( .A(n_23), .Y(n_27) );
OR2x2_ASAP7_75t_L g28 ( .A(n_25), .B(n_21), .Y(n_28) );
AOI22xp5_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_18), .B1(n_24), .B2(n_16), .Y(n_29) );
OAI221xp5_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_29), .B1(n_26), .B2(n_14), .C(n_11), .Y(n_30) );
AO22x2_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_27), .B1(n_5), .B2(n_7), .Y(n_31) );
BUFx2_ASAP7_75t_L g32 ( .A(n_31), .Y(n_32) );
AO22x2_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_2), .B1(n_7), .B2(n_8), .Y(n_33) );
HB1xp67_ASAP7_75t_L g34 ( .A(n_31), .Y(n_34) );
AOI22xp33_ASAP7_75t_L g35 ( .A1(n_32), .A2(n_27), .B1(n_34), .B2(n_33), .Y(n_35) );
endmodule