module fake_jpeg_12611_n_298 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_298);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_182;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_274;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_23),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_48),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_22),
.B(n_0),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_19),
.Y(n_50)
);

INVxp33_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_29),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_51),
.B(n_54),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

BUFx4f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_29),
.B(n_0),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_26),
.B(n_1),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_56),
.B(n_63),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_25),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_61),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_20),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_20),
.B(n_1),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_25),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_34),
.Y(n_95)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_67),
.B(n_68),
.Y(n_125)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_28),
.B1(n_39),
.B2(n_40),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_69),
.A2(n_83),
.B1(n_90),
.B2(n_91),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_39),
.B1(n_52),
.B2(n_35),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_75),
.A2(n_81),
.B1(n_87),
.B2(n_92),
.Y(n_115)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_52),
.A2(n_35),
.B1(n_40),
.B2(n_42),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_89),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_54),
.A2(n_28),
.B1(n_42),
.B2(n_36),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_48),
.A2(n_56),
.B(n_63),
.C(n_61),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_86),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_62),
.A2(n_42),
.B1(n_28),
.B2(n_33),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_48),
.A2(n_36),
.B1(n_24),
.B2(n_30),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_24),
.B1(n_64),
.B2(n_49),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_62),
.A2(n_55),
.B1(n_47),
.B2(n_44),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_100),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_50),
.B(n_34),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_97),
.B(n_18),
.Y(n_118)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_55),
.A2(n_33),
.B1(n_30),
.B2(n_22),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_99),
.A2(n_110),
.B1(n_71),
.B2(n_85),
.Y(n_144)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_55),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_104),
.Y(n_129)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_46),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_6),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_60),
.A2(n_41),
.B1(n_27),
.B2(n_21),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_108),
.A2(n_16),
.B1(n_87),
.B2(n_81),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_51),
.A2(n_41),
.B1(n_27),
.B2(n_21),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_109),
.A2(n_96),
.B(n_92),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_112),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

AOI32xp33_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_38),
.A3(n_12),
.B1(n_13),
.B2(n_18),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_113),
.B(n_130),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_38),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_114),
.B(n_119),
.Y(n_160)
);

OR2x2_ASAP7_75t_SL g147 ( 
.A(n_117),
.B(n_71),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_118),
.B(n_138),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_3),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_73),
.B(n_3),
.C(n_4),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_123),
.Y(n_159)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_78),
.B(n_5),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_74),
.B(n_6),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_135),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_7),
.B1(n_8),
.B2(n_14),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_133),
.A2(n_80),
.B1(n_84),
.B2(n_110),
.Y(n_146)
);

CKINVDCx12_ASAP7_75t_R g134 ( 
.A(n_77),
.Y(n_134)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

NOR2x1_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_8),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

NAND2xp33_ASAP7_75t_SL g137 ( 
.A(n_94),
.B(n_8),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_137),
.A2(n_85),
.B(n_72),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_79),
.B(n_15),
.Y(n_138)
);

CKINVDCx12_ASAP7_75t_R g140 ( 
.A(n_77),
.Y(n_140)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_141),
.A2(n_144),
.B1(n_70),
.B2(n_106),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_115),
.Y(n_168)
);

AND2x6_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_72),
.Y(n_145)
);

A2O1A1O1Ixp25_ASAP7_75t_L g203 ( 
.A1(n_145),
.A2(n_155),
.B(n_176),
.C(n_143),
.D(n_147),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_146),
.A2(n_158),
.B1(n_144),
.B2(n_143),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_172),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_149),
.Y(n_178)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

INVx11_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

AND2x6_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_93),
.Y(n_155)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_168),
.A2(n_135),
.B(n_137),
.Y(n_184)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_169),
.Y(n_204)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_170),
.B(n_173),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_93),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_171),
.B(n_174),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_112),
.A2(n_70),
.B1(n_76),
.B2(n_141),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_121),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_76),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_111),
.Y(n_177)
);

AND2x6_ASAP7_75t_L g176 ( 
.A(n_117),
.B(n_142),
.Y(n_176)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_123),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_179),
.B(n_181),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_125),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_184),
.A2(n_203),
.B(n_145),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_114),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_191),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_152),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_189),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_153),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_124),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_199),
.C(n_175),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_148),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_120),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_195),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_160),
.A2(n_124),
.B1(n_114),
.B2(n_135),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_198),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_146),
.A2(n_158),
.B1(n_155),
.B2(n_176),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_154),
.B(n_139),
.C(n_131),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_150),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_201),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_154),
.B(n_127),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_202),
.B(n_148),
.Y(n_225)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_178),
.A2(n_149),
.B(n_169),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_211),
.Y(n_243)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_200),
.Y(n_212)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_217),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_214),
.B(n_216),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_178),
.A2(n_165),
.B(n_153),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_177),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_163),
.B1(n_161),
.B2(n_173),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_220),
.A2(n_226),
.B1(n_192),
.B2(n_180),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_170),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_221),
.B(n_224),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_193),
.A2(n_161),
.B(n_163),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_193),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_221),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_186),
.A2(n_167),
.B1(n_143),
.B2(n_165),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_227),
.A2(n_233),
.B1(n_212),
.B2(n_209),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_187),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_235),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_238),
.C(n_241),
.Y(n_250)
);

OAI22x1_ASAP7_75t_L g230 ( 
.A1(n_211),
.A2(n_198),
.B1(n_196),
.B2(n_203),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_230),
.A2(n_226),
.B1(n_206),
.B2(n_191),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_223),
.B(n_185),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_225),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_185),
.Y(n_240)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_240),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_199),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_205),
.B(n_183),
.Y(n_242)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_242),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_184),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_216),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_233),
.A2(n_218),
.B1(n_219),
.B2(n_215),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_247),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_243),
.A2(n_218),
.B1(n_219),
.B2(n_215),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_243),
.A2(n_214),
.B1(n_222),
.B2(n_220),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_248),
.Y(n_261)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_251),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_238),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_234),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_254),
.B(n_183),
.Y(n_258)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_255),
.Y(n_264)
);

XNOR2x1_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_257),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_262),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_247),
.Y(n_260)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_260),
.Y(n_276)
);

CKINVDCx11_ASAP7_75t_R g262 ( 
.A(n_253),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_232),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_230),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_251),
.B(n_244),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_267),
.B(n_249),
.Y(n_269)
);

MAJx2_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_250),
.C(n_252),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_269),
.A2(n_263),
.B(n_239),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_261),
.A2(n_231),
.B(n_248),
.Y(n_270)
);

AOI21x1_ASAP7_75t_L g284 ( 
.A1(n_270),
.A2(n_273),
.B(n_227),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_275),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_261),
.A2(n_245),
.B(n_256),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_232),
.C(n_241),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_277),
.C(n_259),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_229),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_272),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_281),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_284),
.Y(n_288)
);

XNOR2x1_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_271),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_276),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_274),
.A2(n_265),
.B(n_260),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_282),
.B(n_275),
.Y(n_287)
);

BUFx24_ASAP7_75t_SL g285 ( 
.A(n_278),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_264),
.Y(n_291)
);

OAI21x1_ASAP7_75t_SL g292 ( 
.A1(n_287),
.A2(n_286),
.B(n_288),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_289),
.B(n_283),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_290),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_291),
.A2(n_292),
.B1(n_208),
.B2(n_213),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_246),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_293),
.C(n_197),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_204),
.B(n_180),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_204),
.C(n_182),
.Y(n_298)
);


endmodule