module fake_aes_9637_n_39 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
HB1xp67_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
HB1xp67_ASAP7_75t_L g13 ( .A(n_10), .Y(n_13) );
NOR2xp33_ASAP7_75t_L g14 ( .A(n_6), .B(n_9), .Y(n_14) );
AND2x4_ASAP7_75t_L g15 ( .A(n_11), .B(n_6), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_7), .B(n_4), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_8), .Y(n_17) );
AOI22xp5_ASAP7_75t_L g18 ( .A1(n_12), .A2(n_16), .B1(n_15), .B2(n_14), .Y(n_18) );
AND2x6_ASAP7_75t_L g19 ( .A(n_15), .B(n_0), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_17), .Y(n_20) );
BUFx3_ASAP7_75t_L g21 ( .A(n_13), .Y(n_21) );
AOI22xp5_ASAP7_75t_L g22 ( .A1(n_19), .A2(n_12), .B1(n_13), .B2(n_2), .Y(n_22) );
AND2x4_ASAP7_75t_L g23 ( .A(n_21), .B(n_0), .Y(n_23) );
AND2x4_ASAP7_75t_L g24 ( .A(n_23), .B(n_18), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_22), .Y(n_25) );
BUFx2_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
OR2x2_ASAP7_75t_L g27 ( .A(n_24), .B(n_18), .Y(n_27) );
AOI21xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_25), .B(n_20), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
NAND5xp2_ASAP7_75t_L g31 ( .A(n_29), .B(n_25), .C(n_19), .D(n_3), .E(n_5), .Y(n_31) );
OAI22xp5_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_19), .B1(n_2), .B2(n_3), .Y(n_32) );
NAND4xp75_ASAP7_75t_L g33 ( .A(n_31), .B(n_19), .C(n_5), .D(n_7), .Y(n_33) );
NAND3xp33_ASAP7_75t_L g34 ( .A(n_32), .B(n_1), .C(n_8), .Y(n_34) );
NAND4xp25_ASAP7_75t_L g35 ( .A(n_30), .B(n_1), .C(n_9), .D(n_31), .Y(n_35) );
NOR2x1p5_ASAP7_75t_L g36 ( .A(n_33), .B(n_30), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_35), .Y(n_37) );
INVx1_ASAP7_75t_L g38 ( .A(n_36), .Y(n_38) );
OAI21xp5_ASAP7_75t_SL g39 ( .A1(n_38), .A2(n_37), .B(n_34), .Y(n_39) );
endmodule