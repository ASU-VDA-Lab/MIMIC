module fake_jpeg_15457_n_156 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_156);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_156;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_62),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_0),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_70),
.B(n_60),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_45),
.C(n_60),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_78),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_48),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_56),
.B(n_61),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_79),
.A2(n_83),
.B(n_85),
.Y(n_104)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_84),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_66),
.Y(n_82)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_71),
.A2(n_63),
.B1(n_51),
.B2(n_53),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_50),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_66),
.A2(n_51),
.B1(n_55),
.B2(n_45),
.Y(n_85)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

FAx1_ASAP7_75t_SL g90 ( 
.A(n_75),
.B(n_0),
.CI(n_1),
.CON(n_90),
.SN(n_90)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_107),
.Y(n_115)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_86),
.A2(n_54),
.B1(n_57),
.B2(n_58),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_99),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_58),
.B1(n_54),
.B2(n_52),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_100),
.A2(n_85),
.B1(n_5),
.B2(n_6),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_2),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_102),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_74),
.B(n_2),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_73),
.B(n_3),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_4),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_106),
.Y(n_111)
);

OAI32xp33_ASAP7_75t_L g107 ( 
.A1(n_83),
.A2(n_22),
.A3(n_43),
.B1(n_40),
.B2(n_39),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_108),
.A2(n_116),
.B1(n_92),
.B2(n_9),
.Y(n_122)
);

MAJx2_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_104),
.C(n_90),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_96),
.C(n_89),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_7),
.Y(n_123)
);

FAx1_ASAP7_75t_SL g120 ( 
.A(n_114),
.B(n_92),
.CI(n_102),
.CON(n_120),
.SN(n_120)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_120),
.B(n_122),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_117),
.A2(n_93),
.B1(n_91),
.B2(n_105),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_121),
.A2(n_110),
.B1(n_111),
.B2(n_10),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_124),
.Y(n_126)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_125),
.A2(n_113),
.B1(n_109),
.B2(n_118),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_127),
.A2(n_129),
.B1(n_130),
.B2(n_121),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_124),
.A2(n_117),
.B1(n_115),
.B2(n_113),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_120),
.B(n_24),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_135),
.C(n_136),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_126),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_131),
.B(n_25),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_120),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_139),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_144),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_143),
.C(n_145),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_138),
.B(n_23),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_21),
.Y(n_150)
);

AO21x1_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_26),
.B(n_33),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_151),
.A2(n_20),
.B(n_32),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_18),
.B(n_31),
.Y(n_153)
);

A2O1A1O1Ixp25_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_17),
.B(n_30),
.C(n_13),
.D(n_14),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_16),
.C(n_28),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_29),
.Y(n_156)
);


endmodule