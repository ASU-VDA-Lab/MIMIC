module real_aes_8894_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_119;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_417;
wire n_182;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_679;
wire n_633;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g486 ( .A1(n_0), .A2(n_131), .B(n_487), .C(n_490), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_1), .B(n_481), .Y(n_492) );
INVx1_ASAP7_75t_L g424 ( .A(n_2), .Y(n_424) );
INVx1_ASAP7_75t_L g169 ( .A(n_3), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_4), .B(n_132), .Y(n_564) );
OAI22xp5_ASAP7_75t_SL g108 ( .A1(n_5), .A2(n_96), .B1(n_109), .B2(n_110), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_5), .Y(n_110) );
OAI22xp5_ASAP7_75t_SL g451 ( .A1(n_5), .A2(n_110), .B1(n_111), .B2(n_452), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_6), .A2(n_466), .B(n_513), .Y(n_512) );
AO21x2_ASAP7_75t_L g543 ( .A1(n_7), .A2(n_138), .B(n_544), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_8), .A2(n_39), .B1(n_135), .B2(n_187), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_9), .B(n_138), .Y(n_155) );
AND2x6_ASAP7_75t_L g140 ( .A(n_10), .B(n_141), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g536 ( .A1(n_11), .A2(n_140), .B(n_469), .C(n_537), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_12), .B(n_40), .Y(n_425) );
INVx1_ASAP7_75t_L g122 ( .A(n_13), .Y(n_122) );
INVx1_ASAP7_75t_L g161 ( .A(n_14), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_15), .B(n_128), .Y(n_181) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_16), .A2(n_104), .B1(n_431), .B2(n_439), .C1(n_442), .C2(n_748), .Y(n_103) );
AOI321xp33_ASAP7_75t_L g105 ( .A1(n_16), .A2(n_106), .A3(n_419), .B1(n_426), .B2(n_427), .C(n_429), .Y(n_105) );
INVx1_ASAP7_75t_L g426 ( .A(n_16), .Y(n_426) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_17), .B(n_132), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_18), .B(n_118), .Y(n_117) );
AO32x2_ASAP7_75t_L g198 ( .A1(n_19), .A2(n_138), .A3(n_139), .B1(n_158), .B2(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_20), .B(n_135), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_21), .B(n_118), .Y(n_171) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_22), .A2(n_55), .B1(n_135), .B2(n_187), .Y(n_201) );
AOI22xp33_ASAP7_75t_SL g195 ( .A1(n_23), .A2(n_80), .B1(n_128), .B2(n_135), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_24), .B(n_135), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_25), .A2(n_139), .B(n_469), .C(n_471), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_26), .A2(n_139), .B(n_469), .C(n_547), .Y(n_546) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_27), .Y(n_126) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_28), .A2(n_97), .B1(n_446), .B2(n_447), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_28), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_29), .B(n_177), .Y(n_235) );
AOI222xp33_ASAP7_75t_SL g443 ( .A1(n_30), .A2(n_444), .B1(n_450), .B2(n_742), .C1(n_743), .C2(n_745), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_31), .A2(n_466), .B(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_32), .B(n_177), .Y(n_214) );
INVx2_ASAP7_75t_L g130 ( .A(n_33), .Y(n_130) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_34), .A2(n_501), .B(n_502), .C(n_506), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_35), .B(n_135), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_36), .B(n_177), .Y(n_189) );
OAI22xp5_ASAP7_75t_SL g444 ( .A1(n_37), .A2(n_445), .B1(n_448), .B2(n_449), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_37), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_38), .B(n_183), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_41), .B(n_465), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_42), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_43), .B(n_132), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_44), .B(n_466), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_45), .A2(n_501), .B(n_506), .C(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_46), .B(n_135), .Y(n_148) );
INVx1_ASAP7_75t_L g488 ( .A(n_47), .Y(n_488) );
OAI22xp5_ASAP7_75t_SL g106 ( .A1(n_48), .A2(n_107), .B1(n_417), .B2(n_418), .Y(n_106) );
INVx1_ASAP7_75t_L g418 ( .A(n_48), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_49), .A2(n_88), .B1(n_187), .B2(n_194), .Y(n_193) );
INVx1_ASAP7_75t_L g527 ( .A(n_50), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_51), .B(n_135), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_52), .B(n_135), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_53), .B(n_466), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_54), .B(n_153), .Y(n_152) );
AOI22xp33_ASAP7_75t_SL g134 ( .A1(n_56), .A2(n_60), .B1(n_128), .B2(n_135), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_57), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_58), .B(n_135), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_59), .B(n_135), .Y(n_234) );
INVx1_ASAP7_75t_L g141 ( .A(n_61), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_62), .B(n_466), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_63), .B(n_481), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_64), .A2(n_153), .B(n_164), .C(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_65), .B(n_135), .Y(n_170) );
INVx1_ASAP7_75t_L g121 ( .A(n_66), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_67), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_68), .B(n_132), .Y(n_504) );
AO32x2_ASAP7_75t_L g191 ( .A1(n_69), .A2(n_138), .A3(n_139), .B1(n_192), .B2(n_196), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_70), .B(n_133), .Y(n_538) );
INVx1_ASAP7_75t_L g233 ( .A(n_71), .Y(n_233) );
INVx1_ASAP7_75t_L g209 ( .A(n_72), .Y(n_209) );
CKINVDCx16_ASAP7_75t_R g484 ( .A(n_73), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_74), .B(n_473), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g561 ( .A1(n_75), .A2(n_469), .B(n_506), .C(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_76), .B(n_128), .Y(n_210) );
CKINVDCx16_ASAP7_75t_R g514 ( .A(n_77), .Y(n_514) );
INVx1_ASAP7_75t_L g438 ( .A(n_78), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_79), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_81), .B(n_187), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_82), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_83), .B(n_128), .Y(n_213) );
INVx2_ASAP7_75t_L g119 ( .A(n_84), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_85), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_86), .B(n_125), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_87), .B(n_128), .Y(n_149) );
OR2x2_ASAP7_75t_L g421 ( .A(n_89), .B(n_422), .Y(n_421) );
OR2x2_ASAP7_75t_L g455 ( .A(n_89), .B(n_423), .Y(n_455) );
INVx2_ASAP7_75t_L g741 ( .A(n_89), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g127 ( .A1(n_90), .A2(n_102), .B1(n_128), .B2(n_129), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_91), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_92), .B(n_466), .Y(n_499) );
INVx1_ASAP7_75t_L g503 ( .A(n_93), .Y(n_503) );
INVxp67_ASAP7_75t_L g517 ( .A(n_94), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_95), .B(n_128), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_96), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_97), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_98), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g534 ( .A(n_99), .Y(n_534) );
INVx1_ASAP7_75t_L g563 ( .A(n_100), .Y(n_563) );
AND2x2_ASAP7_75t_L g529 ( .A(n_101), .B(n_177), .Y(n_529) );
INVxp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_106), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g417 ( .A(n_107), .Y(n_417) );
XNOR2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx2_ASAP7_75t_L g452 ( .A(n_111), .Y(n_452) );
AND2x2_ASAP7_75t_SL g111 ( .A(n_112), .B(n_351), .Y(n_111) );
NOR5xp2_ASAP7_75t_L g112 ( .A(n_113), .B(n_264), .C(n_310), .D(n_323), .E(n_335), .Y(n_112) );
OAI211xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_172), .B(n_218), .C(n_245), .Y(n_113) );
INVx1_ASAP7_75t_SL g346 ( .A(n_114), .Y(n_346) );
OR2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_142), .Y(n_114) );
AND2x2_ASAP7_75t_L g270 ( .A(n_115), .B(n_143), .Y(n_270) );
AND2x2_ASAP7_75t_L g298 ( .A(n_115), .B(n_244), .Y(n_298) );
AND2x2_ASAP7_75t_L g306 ( .A(n_115), .B(n_249), .Y(n_306) );
INVx3_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g236 ( .A(n_116), .B(n_144), .Y(n_236) );
INVx2_ASAP7_75t_L g248 ( .A(n_116), .Y(n_248) );
AND2x2_ASAP7_75t_L g373 ( .A(n_116), .B(n_315), .Y(n_373) );
OR2x2_ASAP7_75t_L g375 ( .A(n_116), .B(n_376), .Y(n_375) );
AND2x4_ASAP7_75t_L g116 ( .A(n_117), .B(n_123), .Y(n_116) );
INVx1_ASAP7_75t_L g242 ( .A(n_117), .Y(n_242) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_118), .Y(n_138) );
INVx1_ASAP7_75t_L g158 ( .A(n_118), .Y(n_158) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
AND2x2_ASAP7_75t_SL g177 ( .A(n_119), .B(n_120), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
NAND3xp33_ASAP7_75t_L g123 ( .A(n_124), .B(n_137), .C(n_139), .Y(n_123) );
AO21x1_ASAP7_75t_L g241 ( .A1(n_124), .A2(n_137), .B(n_242), .Y(n_241) );
OAI22xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_127), .B1(n_131), .B2(n_134), .Y(n_124) );
INVx2_ASAP7_75t_L g188 ( .A(n_125), .Y(n_188) );
OAI22xp5_ASAP7_75t_SL g192 ( .A1(n_125), .A2(n_133), .B1(n_193), .B2(n_195), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_125), .A2(n_131), .B1(n_200), .B2(n_201), .Y(n_199) );
INVx4_ASAP7_75t_L g489 ( .A(n_125), .Y(n_489) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx3_ASAP7_75t_L g133 ( .A(n_126), .Y(n_133) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_126), .Y(n_166) );
INVx1_ASAP7_75t_L g183 ( .A(n_126), .Y(n_183) );
AND2x2_ASAP7_75t_L g467 ( .A(n_126), .B(n_154), .Y(n_467) );
INVx1_ASAP7_75t_L g470 ( .A(n_126), .Y(n_470) );
INVx2_ASAP7_75t_L g162 ( .A(n_128), .Y(n_162) );
INVx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g136 ( .A(n_130), .Y(n_136) );
INVx1_ASAP7_75t_L g154 ( .A(n_130), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_131), .A2(n_151), .B(n_152), .Y(n_150) );
O2A1O1Ixp33_ASAP7_75t_L g167 ( .A1(n_131), .A2(n_168), .B(n_169), .C(n_170), .Y(n_167) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_132), .A2(n_148), .B(n_149), .Y(n_147) );
O2A1O1Ixp5_ASAP7_75t_SL g207 ( .A1(n_132), .A2(n_208), .B(n_209), .C(n_210), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_132), .A2(n_230), .B(n_231), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_132), .B(n_517), .Y(n_516) );
INVx5_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx3_ASAP7_75t_L g208 ( .A(n_135), .Y(n_208) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_135), .Y(n_565) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g187 ( .A(n_136), .Y(n_187) );
BUFx3_ASAP7_75t_L g194 ( .A(n_136), .Y(n_194) );
AND2x6_ASAP7_75t_L g469 ( .A(n_136), .B(n_470), .Y(n_469) );
INVx3_ASAP7_75t_L g481 ( .A(n_137), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_137), .B(n_508), .Y(n_507) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_137), .A2(n_533), .B(n_540), .Y(n_532) );
AO21x2_ASAP7_75t_L g559 ( .A1(n_137), .A2(n_560), .B(n_567), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_137), .B(n_568), .Y(n_567) );
INVx4_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OA21x2_ASAP7_75t_L g145 ( .A1(n_138), .A2(n_146), .B(n_155), .Y(n_145) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_138), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_138), .A2(n_545), .B(n_546), .Y(n_544) );
OAI21xp5_ASAP7_75t_L g228 ( .A1(n_139), .A2(n_229), .B(n_232), .Y(n_228) );
BUFx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OAI21xp5_ASAP7_75t_L g146 ( .A1(n_140), .A2(n_147), .B(n_150), .Y(n_146) );
OAI21xp5_ASAP7_75t_L g159 ( .A1(n_140), .A2(n_160), .B(n_167), .Y(n_159) );
OAI21xp5_ASAP7_75t_L g178 ( .A1(n_140), .A2(n_179), .B(n_184), .Y(n_178) );
OAI21xp5_ASAP7_75t_L g206 ( .A1(n_140), .A2(n_207), .B(n_211), .Y(n_206) );
AND2x4_ASAP7_75t_L g466 ( .A(n_140), .B(n_467), .Y(n_466) );
INVx4_ASAP7_75t_SL g491 ( .A(n_140), .Y(n_491) );
NAND2x1p5_ASAP7_75t_L g535 ( .A(n_140), .B(n_467), .Y(n_535) );
INVx2_ASAP7_75t_SL g142 ( .A(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g286 ( .A(n_143), .B(n_258), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_143), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g400 ( .A(n_143), .B(n_240), .Y(n_400) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_156), .Y(n_143) );
AND2x2_ASAP7_75t_L g243 ( .A(n_144), .B(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g290 ( .A(n_144), .Y(n_290) );
AND2x2_ASAP7_75t_L g315 ( .A(n_144), .B(n_227), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_144), .B(n_348), .Y(n_385) );
INVx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g249 ( .A(n_145), .B(n_227), .Y(n_249) );
AND2x2_ASAP7_75t_L g263 ( .A(n_145), .B(n_226), .Y(n_263) );
AND2x2_ASAP7_75t_L g280 ( .A(n_145), .B(n_156), .Y(n_280) );
AND2x2_ASAP7_75t_L g337 ( .A(n_145), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_145), .B(n_244), .Y(n_350) );
AND2x2_ASAP7_75t_L g402 ( .A(n_145), .B(n_327), .Y(n_402) );
INVx2_ASAP7_75t_L g168 ( .A(n_153), .Y(n_168) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_L g225 ( .A(n_156), .B(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g244 ( .A(n_156), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_156), .B(n_227), .Y(n_321) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_159), .B(n_171), .Y(n_156) );
OA21x2_ASAP7_75t_L g227 ( .A1(n_157), .A2(n_228), .B(n_235), .Y(n_227) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_158), .B(n_541), .Y(n_540) );
O2A1O1Ixp33_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .B(n_163), .C(n_164), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_162), .A2(n_538), .B(n_539), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_162), .A2(n_548), .B(n_549), .Y(n_547) );
O2A1O1Ixp33_ASAP7_75t_L g562 ( .A1(n_164), .A2(n_563), .B(n_564), .C(n_565), .Y(n_562) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_165), .A2(n_212), .B(n_213), .Y(n_211) );
INVx4_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g473 ( .A(n_166), .Y(n_473) );
O2A1O1Ixp5_ASAP7_75t_L g232 ( .A1(n_168), .A2(n_188), .B(n_233), .C(n_234), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_168), .A2(n_472), .B(n_474), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_202), .B(n_215), .Y(n_172) );
INVx1_ASAP7_75t_SL g334 ( .A(n_173), .Y(n_334) );
AND2x4_ASAP7_75t_L g173 ( .A(n_174), .B(n_190), .Y(n_173) );
BUFx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_SL g222 ( .A(n_175), .B(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g217 ( .A(n_176), .Y(n_217) );
INVx1_ASAP7_75t_L g254 ( .A(n_176), .Y(n_254) );
AND2x2_ASAP7_75t_L g275 ( .A(n_176), .B(n_197), .Y(n_275) );
AND2x2_ASAP7_75t_L g309 ( .A(n_176), .B(n_198), .Y(n_309) );
OR2x2_ASAP7_75t_L g328 ( .A(n_176), .B(n_204), .Y(n_328) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_176), .Y(n_342) );
AND2x2_ASAP7_75t_L g355 ( .A(n_176), .B(n_356), .Y(n_355) );
OA21x2_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_189), .Y(n_176) );
INVx2_ASAP7_75t_L g196 ( .A(n_177), .Y(n_196) );
OA21x2_ASAP7_75t_L g205 ( .A1(n_177), .A2(n_206), .B(n_214), .Y(n_205) );
INVx1_ASAP7_75t_L g479 ( .A(n_177), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_177), .A2(n_499), .B(n_500), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_177), .A2(n_524), .B(n_525), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_182), .Y(n_179) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_188), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_190), .A2(n_277), .B1(n_278), .B2(n_287), .Y(n_276) );
AND2x2_ASAP7_75t_L g360 ( .A(n_190), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_197), .Y(n_190) );
INVx1_ASAP7_75t_L g221 ( .A(n_191), .Y(n_221) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_191), .Y(n_258) );
INVx1_ASAP7_75t_L g269 ( .A(n_191), .Y(n_269) );
AND2x2_ASAP7_75t_L g284 ( .A(n_191), .B(n_198), .Y(n_284) );
INVx2_ASAP7_75t_L g490 ( .A(n_194), .Y(n_490) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_194), .Y(n_505) );
INVx1_ASAP7_75t_L g476 ( .A(n_196), .Y(n_476) );
OR2x2_ASAP7_75t_L g238 ( .A(n_197), .B(n_223), .Y(n_238) );
AND2x2_ASAP7_75t_L g268 ( .A(n_197), .B(n_269), .Y(n_268) );
NOR2xp67_ASAP7_75t_L g356 ( .A(n_197), .B(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g216 ( .A(n_198), .B(n_217), .Y(n_216) );
BUFx2_ASAP7_75t_L g325 ( .A(n_198), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_202), .B(n_341), .Y(n_340) );
BUFx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g303 ( .A(n_203), .B(n_269), .Y(n_303) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g215 ( .A(n_204), .B(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g274 ( .A(n_204), .Y(n_274) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g223 ( .A(n_205), .Y(n_223) );
OR2x2_ASAP7_75t_L g253 ( .A(n_205), .B(n_254), .Y(n_253) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_205), .Y(n_308) );
AOI32xp33_ASAP7_75t_L g345 ( .A1(n_215), .A2(n_275), .A3(n_346), .B1(n_347), .B2(n_349), .Y(n_345) );
AND2x2_ASAP7_75t_L g271 ( .A(n_216), .B(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_216), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_216), .B(n_303), .Y(n_389) );
INVx1_ASAP7_75t_L g394 ( .A(n_216), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_224), .B1(n_237), .B2(n_239), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_222), .Y(n_219) );
AND2x2_ASAP7_75t_L g324 ( .A(n_220), .B(n_325), .Y(n_324) );
HB1xp67_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_221), .B(n_223), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_222), .A2(n_246), .B1(n_250), .B2(n_260), .Y(n_245) );
AND2x2_ASAP7_75t_L g267 ( .A(n_222), .B(n_268), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g318 ( .A1(n_222), .A2(n_236), .B(n_284), .C(n_319), .Y(n_318) );
OAI332xp33_ASAP7_75t_L g323 ( .A1(n_222), .A2(n_324), .A3(n_326), .B1(n_328), .B2(n_329), .B3(n_331), .C1(n_332), .C2(n_334), .Y(n_323) );
INVx2_ASAP7_75t_L g364 ( .A(n_222), .Y(n_364) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_223), .Y(n_282) );
INVx1_ASAP7_75t_L g357 ( .A(n_223), .Y(n_357) );
AND2x2_ASAP7_75t_L g411 ( .A(n_223), .B(n_275), .Y(n_411) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_236), .Y(n_224) );
AND2x2_ASAP7_75t_L g291 ( .A(n_226), .B(n_241), .Y(n_291) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g240 ( .A(n_227), .B(n_241), .Y(n_240) );
OR2x2_ASAP7_75t_L g339 ( .A(n_227), .B(n_241), .Y(n_339) );
INVx1_ASAP7_75t_L g348 ( .A(n_227), .Y(n_348) );
INVx1_ASAP7_75t_L g322 ( .A(n_236), .Y(n_322) );
INVxp67_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
OR2x2_ASAP7_75t_L g406 ( .A(n_238), .B(n_258), .Y(n_406) );
INVx1_ASAP7_75t_SL g317 ( .A(n_239), .Y(n_317) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_243), .Y(n_239) );
AND2x2_ASAP7_75t_L g344 ( .A(n_240), .B(n_302), .Y(n_344) );
INVx1_ASAP7_75t_L g363 ( .A(n_240), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g365 ( .A(n_240), .B(n_330), .Y(n_365) );
INVx1_ASAP7_75t_L g262 ( .A(n_241), .Y(n_262) );
AND2x2_ASAP7_75t_L g266 ( .A(n_243), .B(n_247), .Y(n_266) );
AND2x2_ASAP7_75t_L g333 ( .A(n_243), .B(n_291), .Y(n_333) );
INVx2_ASAP7_75t_L g376 ( .A(n_243), .Y(n_376) );
INVx2_ASAP7_75t_L g259 ( .A(n_244), .Y(n_259) );
AND2x2_ASAP7_75t_L g261 ( .A(n_244), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_249), .Y(n_246) );
INVx1_ASAP7_75t_L g277 ( .A(n_247), .Y(n_277) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_248), .B(n_321), .Y(n_327) );
OR2x2_ASAP7_75t_L g391 ( .A(n_248), .B(n_350), .Y(n_391) );
INVx1_ASAP7_75t_L g415 ( .A(n_248), .Y(n_415) );
INVx1_ASAP7_75t_L g371 ( .A(n_249), .Y(n_371) );
AND2x2_ASAP7_75t_L g416 ( .A(n_249), .B(n_259), .Y(n_416) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_255), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_253), .A2(n_279), .B1(n_281), .B2(n_285), .Y(n_278) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OAI322xp33_ASAP7_75t_SL g362 ( .A1(n_256), .A2(n_363), .A3(n_364), .B1(n_365), .B2(n_366), .C1(n_369), .C2(n_371), .Y(n_362) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_259), .Y(n_256) );
AND2x2_ASAP7_75t_L g359 ( .A(n_257), .B(n_275), .Y(n_359) );
OR2x2_ASAP7_75t_L g393 ( .A(n_257), .B(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g396 ( .A(n_257), .B(n_328), .Y(n_396) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g341 ( .A(n_258), .B(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g397 ( .A(n_258), .B(n_328), .Y(n_397) );
INVx3_ASAP7_75t_L g330 ( .A(n_259), .Y(n_330) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
INVx1_ASAP7_75t_L g386 ( .A(n_261), .Y(n_386) );
AOI222xp33_ASAP7_75t_L g265 ( .A1(n_263), .A2(n_266), .B1(n_267), .B2(n_270), .C1(n_271), .C2(n_273), .Y(n_265) );
INVx1_ASAP7_75t_L g296 ( .A(n_263), .Y(n_296) );
NAND3xp33_ASAP7_75t_SL g264 ( .A(n_265), .B(n_276), .C(n_293), .Y(n_264) );
AND2x2_ASAP7_75t_L g381 ( .A(n_268), .B(n_282), .Y(n_381) );
BUFx2_ASAP7_75t_L g272 ( .A(n_269), .Y(n_272) );
INVx1_ASAP7_75t_L g313 ( .A(n_269), .Y(n_313) );
AOI221xp5_ASAP7_75t_L g358 ( .A1(n_270), .A2(n_306), .B1(n_359), .B2(n_360), .C(n_362), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_272), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_275), .Y(n_299) );
AND2x2_ASAP7_75t_L g312 ( .A(n_275), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_280), .B(n_291), .Y(n_292) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
OAI21xp33_ASAP7_75t_L g287 ( .A1(n_282), .A2(n_288), .B(n_292), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_282), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g379 ( .A(n_284), .B(n_361), .Y(n_379) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx1_ASAP7_75t_L g302 ( .A(n_290), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_291), .B(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g408 ( .A(n_291), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_299), .B1(n_300), .B2(n_303), .C(n_304), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_SL g383 ( .A(n_295), .B(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g404 ( .A(n_303), .B(n_309), .Y(n_404) );
INVxp67_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
OAI31xp33_ASAP7_75t_SL g372 ( .A1(n_307), .A2(n_346), .A3(n_373), .B(n_374), .Y(n_372) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx1_ASAP7_75t_L g361 ( .A(n_308), .Y(n_361) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_309), .B(n_313), .Y(n_412) );
OAI221xp5_ASAP7_75t_SL g310 ( .A1(n_311), .A2(n_314), .B1(n_316), .B2(n_317), .C(n_318), .Y(n_310) );
INVx1_ASAP7_75t_L g316 ( .A(n_312), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_315), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g331 ( .A(n_324), .Y(n_331) );
INVx2_ASAP7_75t_L g367 ( .A(n_325), .Y(n_367) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g353 ( .A(n_330), .B(n_339), .Y(n_353) );
A2O1A1Ixp33_ASAP7_75t_L g403 ( .A1(n_330), .A2(n_347), .B(n_404), .C(n_405), .Y(n_403) );
OAI221xp5_ASAP7_75t_SL g335 ( .A1(n_331), .A2(n_336), .B1(n_340), .B2(n_343), .C(n_345), .Y(n_335) );
INVx1_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
A2O1A1Ixp33_ASAP7_75t_L g398 ( .A1(n_334), .A2(n_399), .B(n_401), .C(n_403), .Y(n_398) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_337), .A2(n_388), .B1(n_390), .B2(n_392), .C(n_395), .Y(n_387) );
INVx1_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
NOR4xp25_ASAP7_75t_L g351 ( .A(n_352), .B(n_377), .C(n_398), .D(n_409), .Y(n_351) );
OAI211xp5_ASAP7_75t_SL g352 ( .A1(n_353), .A2(n_354), .B(n_358), .C(n_372), .Y(n_352) );
INVx1_ASAP7_75t_SL g407 ( .A(n_359), .Y(n_407) );
OR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
INVx1_ASAP7_75t_SL g370 ( .A(n_368), .Y(n_370) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_375), .A2(n_384), .B1(n_396), .B2(n_397), .Y(n_395) );
A2O1A1Ixp33_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_380), .B(n_382), .C(n_387), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AOI31xp33_ASAP7_75t_L g409 ( .A1(n_380), .A2(n_410), .A3(n_412), .B(n_413), .Y(n_409) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVxp67_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_407), .B(n_408), .Y(n_405) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_414), .B(n_416), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NAND2xp33_ASAP7_75t_L g749 ( .A(n_419), .B(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_SL g428 ( .A(n_421), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_421), .B(n_430), .Y(n_429) );
BUFx2_ASAP7_75t_L g441 ( .A(n_421), .Y(n_441) );
NOR2x2_ASAP7_75t_L g747 ( .A(n_422), .B(n_741), .Y(n_747) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OR2x2_ASAP7_75t_L g740 ( .A(n_423), .B(n_741), .Y(n_740) );
AND2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_436), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OA21x2_ASAP7_75t_L g440 ( .A1(n_435), .A2(n_436), .B(n_441), .Y(n_440) );
NOR2xp33_ASAP7_75t_SL g750 ( .A(n_435), .B(n_437), .Y(n_750) );
INVx1_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
INVxp67_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g742 ( .A(n_444), .Y(n_742) );
INVx1_ASAP7_75t_L g448 ( .A(n_445), .Y(n_448) );
OAI22xp5_ASAP7_75t_SL g450 ( .A1(n_451), .A2(n_453), .B1(n_456), .B2(n_738), .Y(n_450) );
INVx1_ASAP7_75t_L g744 ( .A(n_451), .Y(n_744) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_455), .A2(n_457), .B1(n_740), .B2(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_SL g457 ( .A(n_458), .B(n_674), .Y(n_457) );
NOR5xp2_ASAP7_75t_L g458 ( .A(n_459), .B(n_605), .C(n_634), .D(n_654), .E(n_661), .Y(n_458) );
OAI211xp5_ASAP7_75t_SL g459 ( .A1(n_460), .A2(n_493), .B(n_550), .C(n_592), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_461), .A2(n_677), .B1(n_679), .B2(n_680), .Y(n_676) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_480), .Y(n_461) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_462), .Y(n_553) );
AND2x4_ASAP7_75t_L g585 ( .A(n_462), .B(n_586), .Y(n_585) );
INVx5_ASAP7_75t_L g603 ( .A(n_462), .Y(n_603) );
AND2x2_ASAP7_75t_L g612 ( .A(n_462), .B(n_604), .Y(n_612) );
AND2x2_ASAP7_75t_L g624 ( .A(n_462), .B(n_497), .Y(n_624) );
AND2x2_ASAP7_75t_L g720 ( .A(n_462), .B(n_588), .Y(n_720) );
OR2x6_ASAP7_75t_L g462 ( .A(n_463), .B(n_477), .Y(n_462) );
AOI21xp5_ASAP7_75t_SL g463 ( .A1(n_464), .A2(n_468), .B(n_476), .Y(n_463) );
BUFx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx5_ASAP7_75t_L g485 ( .A(n_469), .Y(n_485) );
INVx2_ASAP7_75t_L g475 ( .A(n_473), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g502 ( .A1(n_475), .A2(n_503), .B(n_504), .C(n_505), .Y(n_502) );
O2A1O1Ixp33_ASAP7_75t_L g526 ( .A1(n_475), .A2(n_505), .B(n_527), .C(n_528), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
INVx2_ASAP7_75t_L g586 ( .A(n_480), .Y(n_586) );
AND2x2_ASAP7_75t_L g604 ( .A(n_480), .B(n_559), .Y(n_604) );
AND2x2_ASAP7_75t_L g623 ( .A(n_480), .B(n_558), .Y(n_623) );
AND2x2_ASAP7_75t_L g663 ( .A(n_480), .B(n_603), .Y(n_663) );
OA21x2_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_482), .B(n_492), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_SL g483 ( .A1(n_484), .A2(n_485), .B(n_486), .C(n_491), .Y(n_483) );
INVx2_ASAP7_75t_L g501 ( .A(n_485), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_L g513 ( .A1(n_485), .A2(n_491), .B(n_514), .C(n_515), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
INVx1_ASAP7_75t_L g506 ( .A(n_491), .Y(n_506) );
INVxp67_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_495), .B(n_519), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AOI322xp5_ASAP7_75t_L g722 ( .A1(n_496), .A2(n_530), .A3(n_577), .B1(n_585), .B2(n_639), .C1(n_723), .C2(n_726), .Y(n_722) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_509), .Y(n_496) );
INVx5_ASAP7_75t_L g555 ( .A(n_497), .Y(n_555) );
AND2x2_ASAP7_75t_L g571 ( .A(n_497), .B(n_557), .Y(n_571) );
BUFx2_ASAP7_75t_L g649 ( .A(n_497), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_497), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g726 ( .A(n_497), .B(n_633), .Y(n_726) );
OR2x6_ASAP7_75t_L g497 ( .A(n_498), .B(n_507), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_509), .B(n_521), .Y(n_580) );
INVx1_ASAP7_75t_L g607 ( .A(n_509), .Y(n_607) );
AND2x2_ASAP7_75t_L g620 ( .A(n_509), .B(n_542), .Y(n_620) );
AND2x2_ASAP7_75t_L g721 ( .A(n_509), .B(n_639), .Y(n_721) );
INVx3_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OR2x2_ASAP7_75t_L g575 ( .A(n_510), .B(n_521), .Y(n_575) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_510), .Y(n_583) );
OR2x2_ASAP7_75t_L g590 ( .A(n_510), .B(n_542), .Y(n_590) );
AND2x2_ASAP7_75t_L g600 ( .A(n_510), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_510), .B(n_532), .Y(n_629) );
INVxp67_ASAP7_75t_L g653 ( .A(n_510), .Y(n_653) );
AND2x2_ASAP7_75t_L g660 ( .A(n_510), .B(n_530), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_510), .B(n_542), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_510), .B(n_531), .Y(n_686) );
OA21x2_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B(n_518), .Y(n_510) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_530), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_521), .B(n_543), .Y(n_630) );
OR2x2_ASAP7_75t_L g652 ( .A(n_521), .B(n_531), .Y(n_652) );
AND2x2_ASAP7_75t_L g665 ( .A(n_521), .B(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_521), .B(n_620), .Y(n_671) );
OAI211xp5_ASAP7_75t_SL g675 ( .A1(n_521), .A2(n_676), .B(n_681), .C(n_690), .Y(n_675) );
AND2x2_ASAP7_75t_L g736 ( .A(n_521), .B(n_542), .Y(n_736) );
INVx5_ASAP7_75t_SL g521 ( .A(n_522), .Y(n_521) );
OR2x2_ASAP7_75t_L g589 ( .A(n_522), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_522), .B(n_595), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_522), .B(n_584), .Y(n_596) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_522), .Y(n_598) );
OR2x2_ASAP7_75t_L g609 ( .A(n_522), .B(n_531), .Y(n_609) );
AND2x2_ASAP7_75t_SL g614 ( .A(n_522), .B(n_600), .Y(n_614) );
AND2x2_ASAP7_75t_L g639 ( .A(n_522), .B(n_531), .Y(n_639) );
AND2x2_ASAP7_75t_L g659 ( .A(n_522), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g697 ( .A(n_522), .B(n_530), .Y(n_697) );
OR2x2_ASAP7_75t_L g700 ( .A(n_522), .B(n_686), .Y(n_700) );
OR2x6_ASAP7_75t_L g522 ( .A(n_523), .B(n_529), .Y(n_522) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_542), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g643 ( .A1(n_531), .A2(n_644), .B(n_647), .C(n_653), .Y(n_643) );
INVx5_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g574 ( .A(n_532), .B(n_542), .Y(n_574) );
AND2x2_ASAP7_75t_L g578 ( .A(n_532), .B(n_543), .Y(n_578) );
OR2x2_ASAP7_75t_L g584 ( .A(n_532), .B(n_542), .Y(n_584) );
OAI21xp5_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_535), .B(n_536), .Y(n_533) );
INVx1_ASAP7_75t_SL g601 ( .A(n_542), .Y(n_601) );
OR2x2_ASAP7_75t_L g729 ( .A(n_542), .B(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
O2A1O1Ixp33_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_569), .B(n_572), .C(n_581), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AOI31xp33_ASAP7_75t_L g654 ( .A1(n_552), .A2(n_655), .A3(n_657), .B(n_658), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_553), .B(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_554), .B(n_585), .Y(n_591) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_555), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g611 ( .A(n_555), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g616 ( .A(n_555), .B(n_586), .Y(n_616) );
AND2x2_ASAP7_75t_L g626 ( .A(n_555), .B(n_585), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_555), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g646 ( .A(n_555), .B(n_603), .Y(n_646) );
AND2x2_ASAP7_75t_L g651 ( .A(n_555), .B(n_623), .Y(n_651) );
OR2x2_ASAP7_75t_L g670 ( .A(n_555), .B(n_557), .Y(n_670) );
OR2x2_ASAP7_75t_L g672 ( .A(n_555), .B(n_673), .Y(n_672) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_555), .Y(n_719) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g619 ( .A(n_557), .B(n_586), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_557), .B(n_603), .Y(n_642) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
BUFx2_ASAP7_75t_L g588 ( .A(n_559), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_566), .Y(n_560) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g679 ( .A(n_571), .B(n_603), .Y(n_679) );
AOI322xp5_ASAP7_75t_L g681 ( .A1(n_571), .A2(n_585), .A3(n_623), .B1(n_682), .B2(n_683), .C1(n_684), .C2(n_687), .Y(n_681) );
INVx1_ASAP7_75t_L g689 ( .A(n_571), .Y(n_689) );
NAND2xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_576), .Y(n_572) );
INVx1_ASAP7_75t_SL g683 ( .A(n_573), .Y(n_683) );
OR2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
OR2x2_ASAP7_75t_L g635 ( .A(n_574), .B(n_580), .Y(n_635) );
INVx1_ASAP7_75t_L g666 ( .A(n_574), .Y(n_666) );
INVx2_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
AND2x4_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OAI32xp33_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_585), .A3(n_587), .B1(n_589), .B2(n_591), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
AOI21xp33_ASAP7_75t_SL g621 ( .A1(n_584), .A2(n_599), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_SL g636 ( .A(n_585), .Y(n_636) );
AND2x4_ASAP7_75t_L g633 ( .A(n_586), .B(n_603), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_586), .B(n_669), .Y(n_668) );
AOI322xp5_ASAP7_75t_L g698 ( .A1(n_587), .A2(n_614), .A3(n_633), .B1(n_666), .B2(n_699), .C1(n_701), .C2(n_702), .Y(n_698) );
OAI221xp5_ASAP7_75t_L g727 ( .A1(n_587), .A2(n_664), .B1(n_728), .B2(n_729), .C(n_731), .Y(n_727) );
AND2x2_ASAP7_75t_L g615 ( .A(n_588), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_SL g595 ( .A(n_590), .Y(n_595) );
OR2x2_ASAP7_75t_L g667 ( .A(n_590), .B(n_652), .Y(n_667) );
OAI31xp33_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_596), .A3(n_597), .B(n_602), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_593), .A2(n_626), .B1(n_627), .B2(n_631), .Y(n_625) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g638 ( .A(n_595), .B(n_639), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_597), .A2(n_638), .B1(n_691), .B2(n_694), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g680 ( .A(n_600), .B(n_649), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_600), .B(n_639), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_601), .B(n_707), .Y(n_706) );
OR2x2_ASAP7_75t_L g714 ( .A(n_601), .B(n_652), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_602), .A2(n_697), .B1(n_710), .B2(n_713), .Y(n_709) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
INVx2_ASAP7_75t_L g618 ( .A(n_603), .Y(n_618) );
AND2x2_ASAP7_75t_L g701 ( .A(n_603), .B(n_623), .Y(n_701) );
OR2x2_ASAP7_75t_L g703 ( .A(n_603), .B(n_670), .Y(n_703) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_603), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_604), .B(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_604), .B(n_649), .Y(n_657) );
OAI211xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_610), .B(n_613), .C(n_625), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_615), .B1(n_617), .B2(n_620), .C(n_621), .Y(n_613) );
INVxp67_ASAP7_75t_L g725 ( .A(n_616), .Y(n_725) );
INVx1_ASAP7_75t_L g692 ( .A(n_617), .Y(n_692) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
AND2x2_ASAP7_75t_L g656 ( .A(n_618), .B(n_623), .Y(n_656) );
INVx1_ASAP7_75t_L g673 ( .A(n_619), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_619), .B(n_646), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx1_ASAP7_75t_L g688 ( .A(n_623), .Y(n_688) );
AND2x2_ASAP7_75t_L g694 ( .A(n_623), .B(n_649), .Y(n_694) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx1_ASAP7_75t_SL g682 ( .A(n_630), .Y(n_682) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_633), .B(n_669), .Y(n_693) );
OAI221xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_636), .B1(n_637), .B2(n_640), .C(n_643), .Y(n_634) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g730 ( .A(n_639), .Y(n_730) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g648 ( .A(n_642), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_646), .B(n_705), .Y(n_704) );
AOI21xp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_650), .B(n_652), .Y(n_647) );
OAI211xp5_ASAP7_75t_SL g695 ( .A1(n_650), .A2(n_696), .B(n_698), .C(n_704), .Y(n_695) );
INVx1_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g707 ( .A(n_652), .Y(n_707) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OAI222xp33_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_664), .B1(n_667), .B2(n_668), .C1(n_671), .C2(n_672), .Y(n_661) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g737 ( .A(n_668), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_669), .B(n_712), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_669), .A2(n_716), .B1(n_718), .B2(n_721), .Y(n_715) );
INVx2_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
NOR4xp25_ASAP7_75t_L g674 ( .A(n_675), .B(n_695), .C(n_708), .D(n_727), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_677), .B(n_707), .Y(n_717) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g684 ( .A(n_682), .B(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_685), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVx1_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND3xp33_ASAP7_75t_L g708 ( .A(n_709), .B(n_715), .C(n_722), .Y(n_708) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
INVx2_ASAP7_75t_L g724 ( .A(n_720), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
OAI21xp5_ASAP7_75t_SL g731 ( .A1(n_732), .A2(n_734), .B(n_737), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
endmodule