module fake_ariane_326_n_1770 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1770);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1770;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_150;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx2_ASAP7_75t_L g150 ( 
.A(n_18),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_14),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_108),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_64),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_73),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_91),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_128),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_131),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_72),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_40),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_16),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_14),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_38),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_65),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_99),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_85),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_116),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_124),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_83),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_3),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_9),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_61),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_134),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_109),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_27),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_69),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_62),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_47),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_5),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_80),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_118),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_82),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_37),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_66),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_71),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_122),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_95),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_27),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_18),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_87),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_115),
.Y(n_197)
);

BUFx10_ASAP7_75t_L g198 ( 
.A(n_34),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_52),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_143),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_52),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_16),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_11),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_70),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_48),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_77),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_105),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_129),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_3),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_29),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_23),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_135),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_25),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_8),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_33),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_51),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_55),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_97),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_75),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_5),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_9),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_51),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_63),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_148),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_86),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_19),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_121),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_101),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_141),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_19),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_111),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_40),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_28),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_42),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_139),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_104),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_127),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_92),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_100),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_102),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_84),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_7),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_13),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_147),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_145),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_11),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_37),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_7),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_24),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_8),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_20),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_17),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_2),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_132),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_2),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_55),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_76),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_126),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_1),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_24),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_136),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_45),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_43),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_113),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_42),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_106),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_57),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_13),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_56),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_0),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_45),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_21),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_133),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_22),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_26),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_67),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_26),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_50),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_39),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_50),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_144),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_60),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_49),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_46),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_138),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_96),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_44),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_29),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_23),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_15),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_59),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_1),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_130),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_38),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_6),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_10),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_12),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_153),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_153),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_151),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_159),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_280),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_159),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_227),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_164),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_0),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_235),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_258),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_164),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_166),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_266),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_162),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_163),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_166),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_175),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_175),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_174),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_179),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_185),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_173),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_189),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_195),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_203),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_218),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_179),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_L g327 ( 
.A(n_191),
.B(n_4),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_199),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_198),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_201),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_180),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_180),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_178),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_182),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_182),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_205),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_215),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g338 ( 
.A(n_151),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_183),
.B(n_4),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_183),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_194),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_184),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_170),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_184),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_165),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_190),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_190),
.B(n_6),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_209),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_204),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_204),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_150),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_150),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_210),
.Y(n_353)
);

NOR2xp67_ASAP7_75t_L g354 ( 
.A(n_191),
.B(n_10),
.Y(n_354)
);

NOR2xp67_ASAP7_75t_L g355 ( 
.A(n_191),
.B(n_12),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_211),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_249),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_206),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_214),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_222),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_165),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_206),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_218),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_232),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_207),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_253),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_207),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_233),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_208),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_234),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_198),
.B(n_15),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_181),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_208),
.B(n_17),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_298),
.B(n_212),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_298),
.B(n_178),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_343),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_321),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_325),
.B(n_212),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_343),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_343),
.Y(n_380)
);

OA21x2_ASAP7_75t_L g381 ( 
.A1(n_321),
.A2(n_224),
.B(n_219),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_321),
.Y(n_382)
);

INVx4_ASAP7_75t_L g383 ( 
.A(n_343),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_343),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_343),
.Y(n_385)
);

OA21x2_ASAP7_75t_L g386 ( 
.A1(n_299),
.A2(n_224),
.B(n_219),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_341),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_299),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_301),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_301),
.B(n_241),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g391 ( 
.A(n_306),
.B(n_161),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_303),
.Y(n_392)
);

OA21x2_ASAP7_75t_L g393 ( 
.A1(n_303),
.A2(n_245),
.B(n_241),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_371),
.B(n_160),
.Y(n_394)
);

OA21x2_ASAP7_75t_L g395 ( 
.A1(n_305),
.A2(n_254),
.B(n_245),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_305),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_310),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_310),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_311),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_311),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_341),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_315),
.Y(n_402)
);

NAND2x1_ASAP7_75t_L g403 ( 
.A(n_327),
.B(n_170),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_315),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_316),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_325),
.B(n_254),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_316),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_317),
.B(n_261),
.Y(n_408)
);

OA21x2_ASAP7_75t_L g409 ( 
.A1(n_317),
.A2(n_326),
.B(n_319),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_319),
.Y(n_410)
);

NAND2xp33_ASAP7_75t_L g411 ( 
.A(n_371),
.B(n_173),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_326),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_331),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_331),
.B(n_226),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_332),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_332),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_334),
.B(n_226),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_334),
.B(n_230),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_335),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_335),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_302),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_340),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_340),
.B(n_261),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_342),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_333),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_342),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_344),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_344),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_325),
.B(n_267),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_346),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_346),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_349),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_349),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_350),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_350),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_358),
.B(n_267),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_327),
.B(n_173),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_358),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_362),
.B(n_230),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_306),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_362),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_363),
.B(n_286),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_401),
.B(n_313),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_389),
.B(n_363),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_392),
.Y(n_445)
);

AO22x2_ASAP7_75t_L g446 ( 
.A1(n_401),
.A2(n_307),
.B1(n_300),
.B2(n_338),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_392),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_389),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_392),
.Y(n_449)
);

INVx5_ASAP7_75t_L g450 ( 
.A(n_392),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_392),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_392),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_392),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_392),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_375),
.B(n_307),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_392),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_401),
.B(n_314),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_425),
.B(n_329),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_392),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_389),
.B(n_363),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_399),
.Y(n_461)
);

NAND3xp33_ASAP7_75t_L g462 ( 
.A(n_394),
.B(n_320),
.C(n_318),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_389),
.Y(n_463)
);

AND2x6_ASAP7_75t_L g464 ( 
.A(n_388),
.B(n_286),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_399),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_399),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_394),
.A2(n_373),
.B1(n_339),
.B2(n_347),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_399),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_394),
.A2(n_329),
.B1(n_370),
.B2(n_328),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_411),
.A2(n_369),
.B1(n_367),
.B2(n_365),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_425),
.B(n_322),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_389),
.B(n_365),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_389),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_399),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_399),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_399),
.Y(n_476)
);

INVxp33_ASAP7_75t_L g477 ( 
.A(n_387),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_L g478 ( 
.A1(n_411),
.A2(n_386),
.B1(n_395),
.B2(n_393),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_399),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_399),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_399),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_407),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_407),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_388),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_407),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_388),
.B(n_323),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_396),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_396),
.B(n_330),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_386),
.A2(n_369),
.B1(n_367),
.B2(n_355),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_433),
.B(n_336),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_407),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_387),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_421),
.B(n_308),
.Y(n_493)
);

OR2x6_ASAP7_75t_L g494 ( 
.A(n_421),
.B(n_345),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_407),
.Y(n_495)
);

AND2x6_ASAP7_75t_L g496 ( 
.A(n_396),
.B(n_291),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_421),
.A2(n_337),
.B1(n_324),
.B2(n_366),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_433),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_407),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_407),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_433),
.B(n_348),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_409),
.Y(n_502)
);

OR2x6_ASAP7_75t_L g503 ( 
.A(n_374),
.B(n_345),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_391),
.B(n_353),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_407),
.Y(n_505)
);

INVx6_ASAP7_75t_L g506 ( 
.A(n_375),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_433),
.B(n_356),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_407),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_398),
.B(n_359),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_375),
.B(n_300),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_407),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_433),
.B(n_441),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_398),
.B(n_360),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_391),
.A2(n_354),
.B1(n_355),
.B2(n_216),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_386),
.A2(n_354),
.B1(n_338),
.B2(n_161),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_440),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_375),
.B(n_361),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_420),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_433),
.Y(n_519)
);

INVxp67_ASAP7_75t_SL g520 ( 
.A(n_441),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_420),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_420),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_441),
.B(n_364),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_414),
.B(n_351),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_420),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_420),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_441),
.B(n_368),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_441),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_420),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_403),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_441),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_420),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_375),
.B(n_361),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_420),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_L g535 ( 
.A1(n_386),
.A2(n_288),
.B1(n_217),
.B2(n_213),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_398),
.B(n_304),
.Y(n_536)
);

AND2x6_ASAP7_75t_L g537 ( 
.A(n_400),
.B(n_291),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_403),
.Y(n_538)
);

INVx1_ASAP7_75t_SL g539 ( 
.A(n_440),
.Y(n_539)
);

A2O1A1Ixp33_ASAP7_75t_L g540 ( 
.A1(n_400),
.A2(n_269),
.B(n_181),
.C(n_202),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_400),
.B(n_351),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_420),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_391),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_420),
.Y(n_544)
);

INVx4_ASAP7_75t_L g545 ( 
.A(n_409),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_432),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_432),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_404),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_404),
.Y(n_549)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_409),
.Y(n_550)
);

NAND2xp33_ASAP7_75t_L g551 ( 
.A(n_432),
.B(n_404),
.Y(n_551)
);

INVxp33_ASAP7_75t_L g552 ( 
.A(n_391),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_432),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_405),
.B(n_309),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_432),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_432),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g557 ( 
.A(n_414),
.Y(n_557)
);

OAI22xp33_ASAP7_75t_SL g558 ( 
.A1(n_374),
.A2(n_277),
.B1(n_352),
.B2(n_372),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_409),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_SL g560 ( 
.A(n_414),
.B(n_312),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_405),
.B(n_415),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_437),
.A2(n_263),
.B1(n_296),
.B2(n_295),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_432),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_432),
.Y(n_564)
);

INVxp67_ASAP7_75t_SL g565 ( 
.A(n_409),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_405),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_432),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_432),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_415),
.Y(n_569)
);

NOR2x1p5_ASAP7_75t_L g570 ( 
.A(n_374),
.B(n_202),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_414),
.B(n_352),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_415),
.B(n_372),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_409),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_409),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_416),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_416),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_386),
.A2(n_395),
.B1(n_393),
.B2(n_375),
.Y(n_577)
);

NAND3xp33_ASAP7_75t_SL g578 ( 
.A(n_390),
.B(n_246),
.C(n_243),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_390),
.B(n_213),
.Y(n_579)
);

BUFx8_ASAP7_75t_SL g580 ( 
.A(n_375),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_416),
.Y(n_581)
);

OR2x6_ASAP7_75t_L g582 ( 
.A(n_390),
.B(n_217),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_422),
.B(n_231),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_403),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_422),
.B(n_264),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_422),
.B(n_293),
.Y(n_586)
);

OR2x6_ASAP7_75t_L g587 ( 
.A(n_408),
.B(n_288),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_402),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_424),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_424),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_424),
.B(n_293),
.Y(n_591)
);

OR2x6_ASAP7_75t_L g592 ( 
.A(n_408),
.B(n_220),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_486),
.A2(n_442),
.B1(n_406),
.B2(n_378),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_488),
.B(n_378),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_490),
.B(n_437),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_509),
.B(n_406),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_501),
.B(n_427),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_469),
.B(n_427),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_SL g599 ( 
.A(n_539),
.B(n_357),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_462),
.B(n_536),
.Y(n_600)
);

INVxp33_ASAP7_75t_L g601 ( 
.A(n_493),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_573),
.B(n_427),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_513),
.A2(n_467),
.B1(n_554),
.B2(n_503),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_572),
.B(n_429),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_510),
.B(n_429),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_573),
.B(n_428),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_510),
.B(n_442),
.Y(n_607)
);

OR2x2_ASAP7_75t_L g608 ( 
.A(n_492),
.B(n_494),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_510),
.B(n_428),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_446),
.A2(n_395),
.B1(n_386),
.B2(n_393),
.Y(n_610)
);

BUFx5_ASAP7_75t_L g611 ( 
.A(n_574),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_557),
.B(n_428),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_471),
.B(n_438),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_592),
.B(n_438),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_507),
.B(n_523),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_548),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_573),
.B(n_438),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_573),
.B(n_402),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_588),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_592),
.B(n_583),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_458),
.B(n_408),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_548),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_592),
.B(n_417),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_592),
.B(n_417),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_492),
.B(n_417),
.Y(n_625)
);

INVxp67_ASAP7_75t_L g626 ( 
.A(n_494),
.Y(n_626)
);

INVx1_ASAP7_75t_SL g627 ( 
.A(n_477),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_585),
.B(n_417),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_494),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_573),
.B(n_402),
.Y(n_630)
);

INVxp67_ASAP7_75t_SL g631 ( 
.A(n_559),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_520),
.A2(n_436),
.B(n_423),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_503),
.A2(n_439),
.B1(n_418),
.B2(n_436),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_575),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_503),
.A2(n_439),
.B1(n_418),
.B2(n_436),
.Y(n_635)
);

INVxp67_ASAP7_75t_L g636 ( 
.A(n_494),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_549),
.B(n_418),
.Y(n_637)
);

O2A1O1Ixp33_ASAP7_75t_L g638 ( 
.A1(n_565),
.A2(n_423),
.B(n_435),
.C(n_434),
.Y(n_638)
);

OAI21xp5_ASAP7_75t_L g639 ( 
.A1(n_574),
.A2(n_381),
.B(n_402),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_549),
.B(n_418),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_527),
.B(n_423),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_566),
.B(n_439),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_543),
.B(n_439),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_443),
.B(n_397),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_566),
.B(n_397),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_569),
.B(n_397),
.Y(n_646)
);

NOR3xp33_ASAP7_75t_L g647 ( 
.A(n_504),
.B(n_516),
.C(n_578),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_575),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_581),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_503),
.A2(n_435),
.B1(n_434),
.B2(n_431),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_569),
.B(n_397),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_590),
.Y(n_652)
);

NAND2xp33_ASAP7_75t_L g653 ( 
.A(n_464),
.B(n_402),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_590),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_455),
.B(n_410),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g656 ( 
.A(n_493),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_543),
.B(n_410),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_455),
.B(n_410),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_448),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_455),
.B(n_579),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_581),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_589),
.Y(n_662)
);

INVxp33_ASAP7_75t_L g663 ( 
.A(n_497),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_502),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_579),
.B(n_413),
.Y(n_665)
);

AND2x6_ASAP7_75t_SL g666 ( 
.A(n_517),
.B(n_220),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_502),
.B(n_545),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_589),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_484),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_487),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_506),
.B(n_413),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_502),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_576),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_579),
.B(n_413),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_524),
.Y(n_675)
);

INVx4_ASAP7_75t_L g676 ( 
.A(n_506),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_579),
.B(n_413),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_545),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_552),
.B(n_524),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_545),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_550),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_582),
.B(n_419),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_550),
.B(n_412),
.Y(n_683)
);

NAND2xp33_ASAP7_75t_L g684 ( 
.A(n_464),
.B(n_412),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_582),
.B(n_419),
.Y(n_685)
);

INVx4_ASAP7_75t_L g686 ( 
.A(n_506),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_457),
.B(n_419),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_550),
.B(n_448),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_463),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_582),
.B(n_419),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_577),
.B(n_463),
.Y(n_691)
);

OR2x6_ASAP7_75t_L g692 ( 
.A(n_446),
.B(n_426),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_582),
.A2(n_435),
.B1(n_434),
.B2(n_431),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_587),
.B(n_426),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_446),
.A2(n_515),
.B1(n_535),
.B2(n_496),
.Y(n_695)
);

BUFx10_ASAP7_75t_L g696 ( 
.A(n_517),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_473),
.Y(n_697)
);

INVxp67_ASAP7_75t_SL g698 ( 
.A(n_473),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_571),
.B(n_426),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_498),
.B(n_412),
.Y(n_700)
);

INVxp67_ASAP7_75t_L g701 ( 
.A(n_560),
.Y(n_701)
);

O2A1O1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_472),
.A2(n_435),
.B(n_434),
.C(n_431),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_498),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_519),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_519),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_528),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_528),
.B(n_531),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_531),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_587),
.A2(n_431),
.B1(n_430),
.B2(n_426),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_456),
.B(n_412),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_587),
.B(n_430),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_449),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_456),
.B(n_412),
.Y(n_713)
);

NAND2x1p5_ASAP7_75t_L g714 ( 
.A(n_530),
.B(n_386),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_512),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_561),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_449),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_451),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_446),
.A2(n_395),
.B1(n_393),
.B2(n_381),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_530),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_587),
.B(n_430),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_444),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_571),
.B(n_430),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_517),
.B(n_198),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_452),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_460),
.Y(n_726)
);

BUFx6f_ASAP7_75t_SL g727 ( 
.A(n_533),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_538),
.B(n_393),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_538),
.B(n_393),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_533),
.B(n_247),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_586),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_456),
.B(n_383),
.Y(n_732)
);

O2A1O1Ixp5_ASAP7_75t_L g733 ( 
.A1(n_459),
.A2(n_383),
.B(n_384),
.C(n_380),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_591),
.Y(n_734)
);

AO22x2_ASAP7_75t_L g735 ( 
.A1(n_514),
.A2(n_533),
.B1(n_584),
.B2(n_558),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_584),
.B(n_393),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_541),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_570),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_562),
.B(n_221),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_470),
.B(n_395),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_456),
.B(n_542),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_489),
.A2(n_268),
.B1(n_248),
.B2(n_255),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_551),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_540),
.B(n_221),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_452),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_551),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_474),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_456),
.B(n_383),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_464),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_542),
.B(n_383),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_464),
.B(n_395),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_464),
.B(n_395),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_542),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_474),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_464),
.B(n_381),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_542),
.B(n_383),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_496),
.B(n_250),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_496),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_496),
.B(n_198),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_496),
.B(n_381),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_496),
.B(n_381),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_580),
.B(n_256),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_662),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_594),
.B(n_537),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_596),
.B(n_537),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_604),
.B(n_537),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_696),
.B(n_542),
.Y(n_767)
);

INVx5_ASAP7_75t_L g768 ( 
.A(n_664),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_676),
.Y(n_769)
);

OAI21xp33_ASAP7_75t_L g770 ( 
.A1(n_603),
.A2(n_265),
.B(n_262),
.Y(n_770)
);

NOR3xp33_ASAP7_75t_L g771 ( 
.A(n_762),
.B(n_251),
.C(n_250),
.Y(n_771)
);

O2A1O1Ixp33_ASAP7_75t_SL g772 ( 
.A1(n_683),
.A2(n_479),
.B(n_568),
.C(n_454),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_676),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_696),
.B(n_478),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_618),
.A2(n_447),
.B(n_445),
.Y(n_775)
);

OR2x2_ASAP7_75t_L g776 ( 
.A(n_627),
.B(n_251),
.Y(n_776)
);

INVxp67_ASAP7_75t_L g777 ( 
.A(n_599),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_618),
.A2(n_447),
.B(n_445),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_641),
.B(n_537),
.Y(n_779)
);

INVx11_ASAP7_75t_L g780 ( 
.A(n_727),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_686),
.B(n_608),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_727),
.A2(n_537),
.B1(n_568),
.B2(n_508),
.Y(n_782)
);

O2A1O1Ixp33_ASAP7_75t_SL g783 ( 
.A1(n_683),
.A2(n_606),
.B(n_617),
.C(n_602),
.Y(n_783)
);

OAI21xp5_ASAP7_75t_L g784 ( 
.A1(n_639),
.A2(n_454),
.B(n_453),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_641),
.B(n_716),
.Y(n_785)
);

AOI21x1_ASAP7_75t_L g786 ( 
.A1(n_630),
.A2(n_465),
.B(n_453),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_620),
.A2(n_537),
.B1(n_465),
.B2(n_564),
.Y(n_787)
);

OAI21xp5_ASAP7_75t_L g788 ( 
.A1(n_630),
.A2(n_468),
.B(n_466),
.Y(n_788)
);

NAND2x1p5_ASAP7_75t_L g789 ( 
.A(n_686),
.B(n_450),
.Y(n_789)
);

OAI21xp5_ASAP7_75t_L g790 ( 
.A1(n_733),
.A2(n_468),
.B(n_466),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_667),
.A2(n_479),
.B(n_475),
.Y(n_791)
);

O2A1O1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_621),
.A2(n_723),
.B(n_640),
.C(n_642),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_629),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_657),
.B(n_459),
.Y(n_794)
);

O2A1O1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_637),
.A2(n_675),
.B(n_607),
.C(n_605),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_634),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_737),
.B(n_459),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_593),
.B(n_461),
.Y(n_798)
);

OR2x6_ASAP7_75t_L g799 ( 
.A(n_692),
.B(n_580),
.Y(n_799)
);

NAND2xp33_ASAP7_75t_L g800 ( 
.A(n_611),
.B(n_476),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_628),
.B(n_461),
.Y(n_801)
);

AOI21xp33_ASAP7_75t_L g802 ( 
.A1(n_692),
.A2(n_481),
.B(n_476),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_602),
.A2(n_483),
.B(n_475),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_606),
.A2(n_499),
.B(n_483),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_699),
.B(n_461),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_626),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_638),
.A2(n_500),
.B(n_499),
.Y(n_807)
);

INVxp67_ASAP7_75t_L g808 ( 
.A(n_643),
.Y(n_808)
);

A2O1A1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_615),
.A2(n_529),
.B(n_480),
.C(n_547),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_731),
.B(n_734),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_697),
.Y(n_811)
);

AO21x1_ASAP7_75t_L g812 ( 
.A1(n_615),
.A2(n_505),
.B(n_500),
.Y(n_812)
);

O2A1O1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_613),
.A2(n_283),
.B(n_279),
.C(n_275),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_634),
.Y(n_814)
);

AO21x1_ASAP7_75t_L g815 ( 
.A1(n_600),
.A2(n_508),
.B(n_505),
.Y(n_815)
);

A2O1A1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_595),
.A2(n_597),
.B(n_687),
.C(n_671),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_625),
.B(n_480),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_654),
.B(n_633),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_619),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_636),
.B(n_480),
.Y(n_820)
);

O2A1O1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_655),
.A2(n_283),
.B(n_259),
.C(n_260),
.Y(n_821)
);

INVxp67_ASAP7_75t_L g822 ( 
.A(n_730),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_617),
.A2(n_532),
.B(n_518),
.Y(n_823)
);

BUFx3_ASAP7_75t_L g824 ( 
.A(n_656),
.Y(n_824)
);

AO21x1_ASAP7_75t_L g825 ( 
.A1(n_597),
.A2(n_532),
.B(n_518),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_710),
.A2(n_553),
.B(n_534),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_632),
.A2(n_553),
.B(n_534),
.Y(n_827)
);

NAND3xp33_ASAP7_75t_L g828 ( 
.A(n_730),
.B(n_272),
.C(n_271),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_L g829 ( 
.A1(n_595),
.A2(n_563),
.B(n_555),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_648),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_609),
.A2(n_529),
.B1(n_547),
.B2(n_563),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_715),
.A2(n_564),
.B(n_555),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_710),
.A2(n_482),
.B(n_481),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_635),
.B(n_529),
.Y(n_834)
);

O2A1O1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_658),
.A2(n_297),
.B(n_252),
.C(n_259),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_648),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_649),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_654),
.B(n_547),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_679),
.B(n_482),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_649),
.Y(n_840)
);

AO21x1_ASAP7_75t_L g841 ( 
.A1(n_691),
.A2(n_172),
.B(n_168),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_661),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_738),
.B(n_252),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_713),
.A2(n_741),
.B(n_646),
.Y(n_844)
);

INVx1_ASAP7_75t_SL g845 ( 
.A(n_601),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_713),
.A2(n_741),
.B(n_651),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_661),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_645),
.A2(n_567),
.B(n_556),
.Y(n_848)
);

OAI21xp5_ASAP7_75t_L g849 ( 
.A1(n_751),
.A2(n_567),
.B(n_556),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_701),
.B(n_485),
.Y(n_850)
);

O2A1O1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_612),
.A2(n_292),
.B(n_279),
.C(n_297),
.Y(n_851)
);

BUFx4f_ASAP7_75t_L g852 ( 
.A(n_757),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_668),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_623),
.B(n_624),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_647),
.A2(n_546),
.B1(n_544),
.B2(n_526),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_667),
.A2(n_546),
.B(n_544),
.Y(n_856)
);

NAND2xp33_ASAP7_75t_L g857 ( 
.A(n_611),
.B(n_485),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_688),
.A2(n_748),
.B(n_732),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_688),
.A2(n_526),
.B(n_525),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_697),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_700),
.A2(n_525),
.B(n_522),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_697),
.Y(n_862)
);

O2A1O1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_614),
.A2(n_260),
.B(n_275),
.C(n_274),
.Y(n_863)
);

INVxp67_ASAP7_75t_L g864 ( 
.A(n_687),
.Y(n_864)
);

AOI33xp33_ASAP7_75t_L g865 ( 
.A1(n_739),
.A2(n_292),
.A3(n_269),
.B1(n_270),
.B2(n_274),
.B3(n_278),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_732),
.A2(n_522),
.B(n_521),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_748),
.A2(n_521),
.B(n_511),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_697),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_720),
.B(n_511),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_750),
.A2(n_495),
.B(n_491),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_750),
.A2(n_495),
.B(n_491),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_724),
.B(n_284),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_720),
.B(n_381),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_757),
.Y(n_874)
);

OAI21xp5_ASAP7_75t_L g875 ( 
.A1(n_752),
.A2(n_450),
.B(n_381),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_762),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_668),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_660),
.B(n_287),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_700),
.A2(n_450),
.B(n_383),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_712),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_669),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_659),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_691),
.A2(n_450),
.B(n_380),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_739),
.B(n_290),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_653),
.A2(n_450),
.B(n_380),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_684),
.A2(n_756),
.B(n_631),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_728),
.A2(n_384),
.B(n_380),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_671),
.A2(n_678),
.B1(n_680),
.B2(n_681),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_756),
.A2(n_384),
.B(n_377),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_729),
.A2(n_736),
.B(n_726),
.Y(n_890)
);

NOR2x2_ASAP7_75t_L g891 ( 
.A(n_692),
.B(n_294),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_722),
.A2(n_384),
.B(n_377),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_659),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_L g894 ( 
.A1(n_678),
.A2(n_173),
.B1(n_242),
.B2(n_384),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_680),
.A2(n_384),
.B(n_377),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_673),
.B(n_382),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_598),
.B(n_152),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_749),
.B(n_382),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_681),
.A2(n_156),
.B(n_285),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_735),
.B(n_382),
.Y(n_900)
);

OAI22xp5_ASAP7_75t_L g901 ( 
.A1(n_695),
.A2(n_173),
.B1(n_242),
.B2(n_281),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_SL g902 ( 
.A(n_663),
.B(n_154),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_664),
.B(n_155),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_664),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_747),
.A2(n_385),
.B(n_379),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_702),
.A2(n_223),
.B(n_158),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_743),
.A2(n_242),
.B(n_167),
.C(n_169),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_753),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_759),
.B(n_242),
.Y(n_909)
);

NOR2xp67_ASAP7_75t_L g910 ( 
.A(n_742),
.B(n_157),
.Y(n_910)
);

NOR2xp67_ASAP7_75t_L g911 ( 
.A(n_650),
.B(n_171),
.Y(n_911)
);

A2O1A1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_746),
.A2(n_242),
.B(n_176),
.C(n_177),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_717),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_735),
.A2(n_236),
.B1(n_186),
.B2(n_187),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_754),
.A2(n_385),
.B(n_379),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_664),
.B(n_188),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_753),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_669),
.A2(n_238),
.B(n_192),
.C(n_193),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_707),
.A2(n_239),
.B(n_196),
.Y(n_919)
);

INVx4_ASAP7_75t_L g920 ( 
.A(n_672),
.Y(n_920)
);

O2A1O1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_670),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_SL g922 ( 
.A1(n_707),
.A2(n_25),
.B(n_28),
.C(n_30),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_717),
.A2(n_385),
.B(n_379),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_718),
.A2(n_240),
.B(n_197),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_718),
.A2(n_244),
.B(n_200),
.Y(n_925)
);

OR2x2_ASAP7_75t_L g926 ( 
.A(n_744),
.B(n_30),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_670),
.Y(n_927)
);

BUFx2_ASAP7_75t_L g928 ( 
.A(n_666),
.Y(n_928)
);

AO21x1_ASAP7_75t_L g929 ( 
.A1(n_714),
.A2(n_170),
.B(n_225),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_672),
.B(n_257),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_644),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_689),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_672),
.B(n_273),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_725),
.A2(n_237),
.B(n_228),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_745),
.A2(n_385),
.B(n_379),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_616),
.B(n_229),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_622),
.B(n_276),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_745),
.A2(n_385),
.B(n_379),
.Y(n_938)
);

NAND3xp33_ASAP7_75t_L g939 ( 
.A(n_652),
.B(n_282),
.C(n_379),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_755),
.A2(n_385),
.B(n_379),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_665),
.A2(n_225),
.B(n_170),
.C(n_376),
.Y(n_941)
);

O2A1O1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_703),
.A2(n_31),
.B(n_32),
.C(n_33),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_672),
.Y(n_943)
);

A2O1A1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_674),
.A2(n_225),
.B(n_170),
.C(n_376),
.Y(n_944)
);

BUFx12f_ASAP7_75t_L g945 ( 
.A(n_928),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_822),
.B(n_611),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_852),
.B(n_785),
.Y(n_947)
);

BUFx8_ASAP7_75t_L g948 ( 
.A(n_884),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_763),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_793),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_816),
.B(n_611),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_908),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_908),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_808),
.B(n_876),
.Y(n_954)
);

INVx1_ASAP7_75t_SL g955 ( 
.A(n_845),
.Y(n_955)
);

OAI22xp5_ASAP7_75t_L g956 ( 
.A1(n_779),
.A2(n_695),
.B1(n_698),
.B2(n_689),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_800),
.A2(n_761),
.B(n_760),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_810),
.B(n_611),
.Y(n_958)
);

AOI22xp33_ASAP7_75t_L g959 ( 
.A1(n_771),
.A2(n_735),
.B1(n_758),
.B2(n_611),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_881),
.Y(n_960)
);

AOI221xp5_ASAP7_75t_L g961 ( 
.A1(n_770),
.A2(n_610),
.B1(n_682),
.B2(n_721),
.C(n_677),
.Y(n_961)
);

INVx4_ASAP7_75t_L g962 ( 
.A(n_780),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_830),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_857),
.A2(n_753),
.B(n_714),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_836),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_852),
.B(n_705),
.Y(n_966)
);

CKINVDCx6p67_ASAP7_75t_R g967 ( 
.A(n_824),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_864),
.B(n_705),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_927),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_764),
.A2(n_753),
.B(n_708),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_932),
.B(n_708),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_777),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_854),
.B(n_610),
.Y(n_973)
);

NOR2x1_ASAP7_75t_L g974 ( 
.A(n_811),
.B(n_706),
.Y(n_974)
);

NOR3xp33_ASAP7_75t_SL g975 ( 
.A(n_828),
.B(n_872),
.C(n_918),
.Y(n_975)
);

BUFx4f_ASAP7_75t_L g976 ( 
.A(n_799),
.Y(n_976)
);

OAI21x1_ASAP7_75t_SL g977 ( 
.A1(n_795),
.A2(n_685),
.B(n_711),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_R g978 ( 
.A(n_902),
.B(n_704),
.Y(n_978)
);

O2A1O1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_766),
.A2(n_694),
.B(n_690),
.C(n_740),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_806),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_847),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_796),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_765),
.A2(n_709),
.B(n_693),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_874),
.B(n_719),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_829),
.A2(n_719),
.B(n_385),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_798),
.A2(n_385),
.B(n_379),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_942),
.A2(n_31),
.B(n_32),
.C(n_34),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_843),
.A2(n_225),
.B1(n_379),
.B2(n_376),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_814),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_827),
.A2(n_385),
.B(n_379),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_860),
.Y(n_991)
);

BUFx2_ASAP7_75t_L g992 ( 
.A(n_799),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_768),
.B(n_385),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_837),
.B(n_35),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_840),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_768),
.B(n_376),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_859),
.A2(n_376),
.B(n_225),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_842),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_813),
.A2(n_35),
.B(n_36),
.C(n_39),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_897),
.A2(n_376),
.B(n_41),
.C(n_43),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_853),
.Y(n_1001)
);

OAI21xp33_ASAP7_75t_L g1002 ( 
.A1(n_878),
.A2(n_36),
.B(n_41),
.Y(n_1002)
);

NAND2x1p5_ASAP7_75t_L g1003 ( 
.A(n_768),
.B(n_376),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_799),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_877),
.Y(n_1005)
);

INVxp67_ASAP7_75t_L g1006 ( 
.A(n_776),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_768),
.B(n_44),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_896),
.Y(n_1008)
);

NOR3xp33_ASAP7_75t_L g1009 ( 
.A(n_921),
.B(n_46),
.C(n_47),
.Y(n_1009)
);

A2O1A1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_792),
.A2(n_376),
.B(n_49),
.C(n_53),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_794),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_819),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_926),
.A2(n_376),
.B(n_56),
.C(n_54),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_940),
.A2(n_376),
.B(n_68),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_844),
.A2(n_58),
.B(n_74),
.Y(n_1015)
);

INVxp67_ASAP7_75t_L g1016 ( 
.A(n_843),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_781),
.B(n_78),
.Y(n_1017)
);

NAND3xp33_ASAP7_75t_SL g1018 ( 
.A(n_914),
.B(n_851),
.C(n_863),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_839),
.B(n_890),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_880),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_900),
.A2(n_79),
.B1(n_81),
.B2(n_89),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_787),
.A2(n_90),
.B1(n_93),
.B2(n_94),
.Y(n_1022)
);

INVx4_ASAP7_75t_L g1023 ( 
.A(n_860),
.Y(n_1023)
);

AO32x1_ASAP7_75t_L g1024 ( 
.A1(n_901),
.A2(n_98),
.A3(n_103),
.B1(n_107),
.B2(n_112),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_769),
.B(n_773),
.Y(n_1025)
);

OR2x6_ASAP7_75t_L g1026 ( 
.A(n_920),
.B(n_114),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_891),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_882),
.B(n_117),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_913),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_818),
.B(n_119),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_R g1031 ( 
.A(n_811),
.B(n_123),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_844),
.A2(n_846),
.B(n_856),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_860),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_911),
.A2(n_137),
.B1(n_146),
.B2(n_936),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_805),
.B(n_801),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_908),
.Y(n_1036)
);

CKINVDCx16_ASAP7_75t_R g1037 ( 
.A(n_868),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_SL g1038 ( 
.A1(n_906),
.A2(n_807),
.B(n_790),
.C(n_893),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_797),
.B(n_817),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_937),
.B(n_931),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_865),
.B(n_850),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_SL g1042 ( 
.A1(n_782),
.A2(n_820),
.B1(n_934),
.B2(n_868),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_846),
.A2(n_809),
.B(n_784),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_821),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_862),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_917),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_917),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_769),
.B(n_773),
.Y(n_1048)
);

BUFx2_ASAP7_75t_L g1049 ( 
.A(n_868),
.Y(n_1049)
);

OAI21xp33_ASAP7_75t_L g1050 ( 
.A1(n_834),
.A2(n_832),
.B(n_907),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_917),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_862),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_882),
.Y(n_1053)
);

AND2x2_ASAP7_75t_SL g1054 ( 
.A(n_920),
.B(n_904),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_SL g1055 ( 
.A1(n_893),
.A2(n_788),
.B(n_858),
.C(n_803),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_835),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_904),
.Y(n_1057)
);

NOR3xp33_ASAP7_75t_L g1058 ( 
.A(n_903),
.B(n_933),
.C(n_930),
.Y(n_1058)
);

INVx1_ASAP7_75t_SL g1059 ( 
.A(n_774),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_943),
.Y(n_1060)
);

NOR2x1_ASAP7_75t_R g1061 ( 
.A(n_916),
.B(n_767),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_888),
.B(n_943),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_898),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_910),
.B(n_898),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_SL g1065 ( 
.A1(n_838),
.A2(n_912),
.B(n_831),
.C(n_886),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_886),
.A2(n_855),
.B1(n_873),
.B2(n_789),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_783),
.A2(n_848),
.B(n_791),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_786),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_848),
.A2(n_772),
.B(n_775),
.Y(n_1069)
);

AO21x2_ASAP7_75t_L g1070 ( 
.A1(n_812),
.A2(n_825),
.B(n_929),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_775),
.A2(n_778),
.B(n_871),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_922),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_778),
.A2(n_867),
.B(n_866),
.Y(n_1073)
);

INVx4_ASAP7_75t_L g1074 ( 
.A(n_789),
.Y(n_1074)
);

O2A1O1Ixp5_ASAP7_75t_L g1075 ( 
.A1(n_815),
.A2(n_915),
.B(n_905),
.C(n_883),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_892),
.B(n_802),
.Y(n_1076)
);

INVx4_ASAP7_75t_L g1077 ( 
.A(n_885),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_892),
.B(n_909),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_869),
.B(n_919),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_895),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_889),
.Y(n_1081)
);

O2A1O1Ixp5_ASAP7_75t_L g1082 ( 
.A1(n_905),
.A2(n_915),
.B(n_883),
.C(n_885),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_875),
.B(n_849),
.Y(n_1083)
);

INVx1_ASAP7_75t_SL g1084 ( 
.A(n_924),
.Y(n_1084)
);

INVxp33_ASAP7_75t_SL g1085 ( 
.A(n_894),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_870),
.A2(n_803),
.B(n_804),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_804),
.B(n_823),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_823),
.A2(n_861),
.B(n_826),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_887),
.Y(n_1089)
);

OAI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_983),
.A2(n_861),
.B(n_833),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_1008),
.A2(n_1085),
.B1(n_951),
.B2(n_958),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_1067),
.A2(n_938),
.B(n_935),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_976),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_951),
.A2(n_833),
.B(n_938),
.Y(n_1094)
);

OR2x2_ASAP7_75t_L g1095 ( 
.A(n_1006),
.B(n_899),
.Y(n_1095)
);

INVxp67_ASAP7_75t_SL g1096 ( 
.A(n_958),
.Y(n_1096)
);

NOR2xp67_ASAP7_75t_L g1097 ( 
.A(n_962),
.B(n_939),
.Y(n_1097)
);

AOI21x1_ASAP7_75t_L g1098 ( 
.A1(n_986),
.A2(n_841),
.B(n_923),
.Y(n_1098)
);

AO32x2_ASAP7_75t_L g1099 ( 
.A1(n_1077),
.A2(n_941),
.A3(n_944),
.B1(n_923),
.B2(n_935),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_975),
.A2(n_1002),
.B(n_1034),
.C(n_1050),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_1067),
.A2(n_826),
.B(n_879),
.Y(n_1101)
);

CKINVDCx20_ASAP7_75t_R g1102 ( 
.A(n_967),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1019),
.B(n_879),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_1016),
.B(n_925),
.Y(n_1104)
);

INVx4_ASAP7_75t_L g1105 ( 
.A(n_962),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_964),
.A2(n_1078),
.B(n_1038),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1019),
.B(n_973),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_1035),
.A2(n_959),
.B1(n_947),
.B2(n_1039),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_SL g1109 ( 
.A(n_976),
.B(n_1007),
.Y(n_1109)
);

AND2x4_ASAP7_75t_L g1110 ( 
.A(n_1063),
.B(n_992),
.Y(n_1110)
);

O2A1O1Ixp33_ASAP7_75t_SL g1111 ( 
.A1(n_946),
.A2(n_1055),
.B(n_1000),
.C(n_1010),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_SL g1112 ( 
.A(n_1007),
.B(n_1026),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1018),
.A2(n_1059),
.B1(n_948),
.B2(n_984),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_973),
.B(n_1035),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_964),
.A2(n_1078),
.B(n_957),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_957),
.A2(n_1043),
.B(n_1032),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1043),
.A2(n_1032),
.B(n_1014),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_949),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_954),
.B(n_980),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_960),
.Y(n_1120)
);

NAND2x1_ASAP7_75t_L g1121 ( 
.A(n_1074),
.B(n_1023),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_1027),
.B(n_950),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1073),
.A2(n_1066),
.B(n_1087),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1039),
.B(n_982),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_963),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_986),
.A2(n_1069),
.B(n_1086),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_969),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_955),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_1037),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_999),
.A2(n_987),
.B(n_1041),
.C(n_1013),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1089),
.A2(n_985),
.B(n_1076),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_972),
.B(n_1004),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_989),
.Y(n_1133)
);

AO21x2_ASAP7_75t_L g1134 ( 
.A1(n_1070),
.A2(n_1069),
.B(n_985),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_995),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_998),
.B(n_1044),
.Y(n_1136)
);

OR2x2_ASAP7_75t_L g1137 ( 
.A(n_1040),
.B(n_971),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_948),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1086),
.A2(n_1071),
.B(n_1073),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_1071),
.A2(n_1088),
.B(n_1082),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1087),
.A2(n_1077),
.B(n_1083),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1056),
.A2(n_994),
.B1(n_1062),
.B2(n_1011),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1030),
.A2(n_1079),
.B(n_1064),
.C(n_1017),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_994),
.A2(n_1062),
.B1(n_1042),
.B2(n_1083),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_990),
.A2(n_1065),
.B(n_970),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1075),
.A2(n_1076),
.B(n_997),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_991),
.Y(n_1147)
);

O2A1O1Ixp5_ASAP7_75t_L g1148 ( 
.A1(n_1022),
.A2(n_1072),
.B(n_1015),
.C(n_968),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1009),
.A2(n_977),
.B(n_1058),
.C(n_1030),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1081),
.A2(n_1080),
.B(n_956),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1080),
.A2(n_1068),
.B(n_979),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1052),
.B(n_1053),
.Y(n_1152)
);

A2O1A1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_1028),
.A2(n_1084),
.B(n_961),
.C(n_1021),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_965),
.B(n_1001),
.Y(n_1154)
);

INVx3_ASAP7_75t_SL g1155 ( 
.A(n_1054),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1024),
.A2(n_1070),
.B(n_1025),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_961),
.A2(n_966),
.B(n_1045),
.C(n_974),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_981),
.B(n_1005),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1012),
.B(n_1029),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1024),
.A2(n_1048),
.B(n_996),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1026),
.A2(n_988),
.B1(n_1057),
.B2(n_1003),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1020),
.B(n_1057),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1060),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1024),
.A2(n_993),
.B(n_1003),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1026),
.A2(n_1061),
.B(n_1074),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1023),
.A2(n_1049),
.B(n_1033),
.Y(n_1166)
);

OAI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1031),
.A2(n_1060),
.B(n_978),
.Y(n_1167)
);

BUFx2_ASAP7_75t_L g1168 ( 
.A(n_952),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1060),
.A2(n_952),
.B(n_953),
.C(n_1036),
.Y(n_1169)
);

BUFx5_ASAP7_75t_L g1170 ( 
.A(n_952),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_953),
.A2(n_1036),
.B(n_1046),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_953),
.A2(n_1036),
.B(n_1046),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_945),
.B(n_1047),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1047),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1047),
.A2(n_816),
.B(n_983),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1051),
.A2(n_857),
.B(n_800),
.Y(n_1176)
);

AOI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1051),
.A2(n_876),
.B1(n_603),
.B2(n_599),
.Y(n_1177)
);

AO31x2_ASAP7_75t_L g1178 ( 
.A1(n_1051),
.A2(n_812),
.A3(n_825),
.B(n_841),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_958),
.A2(n_857),
.B(n_800),
.Y(n_1179)
);

NAND2x1p5_ASAP7_75t_L g1180 ( 
.A(n_1054),
.B(n_768),
.Y(n_1180)
);

AO31x2_ASAP7_75t_L g1181 ( 
.A1(n_1068),
.A2(n_812),
.A3(n_825),
.B(n_841),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1067),
.A2(n_986),
.B(n_1032),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1008),
.B(n_785),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1016),
.B(n_492),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_963),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_967),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1016),
.B(n_492),
.Y(n_1187)
);

INVx2_ASAP7_75t_SL g1188 ( 
.A(n_976),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_958),
.A2(n_857),
.B(n_800),
.Y(n_1189)
);

AO31x2_ASAP7_75t_L g1190 ( 
.A1(n_1068),
.A2(n_812),
.A3(n_825),
.B(n_841),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1008),
.A2(n_603),
.B1(n_785),
.B2(n_816),
.Y(n_1191)
);

AO32x2_ASAP7_75t_L g1192 ( 
.A1(n_1077),
.A2(n_1066),
.A3(n_901),
.B1(n_1011),
.B2(n_1042),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1067),
.A2(n_986),
.B(n_1032),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_958),
.A2(n_857),
.B(n_800),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_958),
.A2(n_857),
.B(n_800),
.Y(n_1195)
);

OA21x2_ASAP7_75t_L g1196 ( 
.A1(n_1032),
.A2(n_986),
.B(n_1069),
.Y(n_1196)
);

INVxp67_ASAP7_75t_SL g1197 ( 
.A(n_958),
.Y(n_1197)
);

AO21x2_ASAP7_75t_L g1198 ( 
.A1(n_986),
.A2(n_929),
.B(n_1070),
.Y(n_1198)
);

BUFx3_ASAP7_75t_L g1199 ( 
.A(n_967),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_983),
.A2(n_816),
.B(n_779),
.Y(n_1200)
);

INVx2_ASAP7_75t_SL g1201 ( 
.A(n_976),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1067),
.A2(n_986),
.B(n_1032),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1067),
.A2(n_986),
.B(n_1032),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1016),
.B(n_492),
.Y(n_1204)
);

BUFx2_ASAP7_75t_R g1205 ( 
.A(n_980),
.Y(n_1205)
);

O2A1O1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_947),
.A2(n_822),
.B(n_596),
.C(n_594),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_958),
.A2(n_857),
.B(n_800),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1054),
.B(n_852),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1067),
.A2(n_986),
.B(n_1032),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_958),
.A2(n_857),
.B(n_800),
.Y(n_1210)
);

INVx4_ASAP7_75t_L g1211 ( 
.A(n_962),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_975),
.A2(n_603),
.B(n_897),
.C(n_1002),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_958),
.A2(n_857),
.B(n_800),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1008),
.B(n_785),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_1074),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1008),
.B(n_785),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_980),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1016),
.B(n_492),
.Y(n_1218)
);

AO31x2_ASAP7_75t_L g1219 ( 
.A1(n_1068),
.A2(n_812),
.A3(n_825),
.B(n_841),
.Y(n_1219)
);

NAND3xp33_ASAP7_75t_L g1220 ( 
.A(n_1002),
.B(n_603),
.C(n_467),
.Y(n_1220)
);

AOI21xp33_ASAP7_75t_L g1221 ( 
.A1(n_1002),
.A2(n_603),
.B(n_692),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_949),
.Y(n_1222)
);

AO21x2_ASAP7_75t_L g1223 ( 
.A1(n_986),
.A2(n_929),
.B(n_1070),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_967),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_958),
.A2(n_857),
.B(n_800),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_949),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1067),
.A2(n_986),
.B(n_1032),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_980),
.Y(n_1228)
);

AOI21x1_ASAP7_75t_L g1229 ( 
.A1(n_986),
.A2(n_1067),
.B(n_1069),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_949),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1016),
.B(n_492),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1067),
.A2(n_986),
.B(n_1032),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_949),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_958),
.A2(n_857),
.B(n_800),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_975),
.A2(n_603),
.B(n_897),
.C(n_1002),
.Y(n_1235)
);

CKINVDCx11_ASAP7_75t_R g1236 ( 
.A(n_945),
.Y(n_1236)
);

AOI221x1_ASAP7_75t_L g1237 ( 
.A1(n_1002),
.A2(n_1009),
.B1(n_1000),
.B2(n_1010),
.C(n_1018),
.Y(n_1237)
);

OAI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1112),
.A2(n_1220),
.B1(n_1109),
.B2(n_1144),
.Y(n_1238)
);

AOI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1112),
.A2(n_1177),
.B1(n_1109),
.B2(n_1144),
.Y(n_1239)
);

OAI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1191),
.A2(n_1183),
.B1(n_1216),
.B2(n_1214),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_1129),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_1186),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_1093),
.B(n_1188),
.Y(n_1243)
);

OAI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1191),
.A2(n_1183),
.B1(n_1216),
.B2(n_1214),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1212),
.A2(n_1235),
.B1(n_1130),
.B2(n_1100),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1221),
.A2(n_1113),
.B1(n_1108),
.B2(n_1142),
.Y(n_1246)
);

INVx1_ASAP7_75t_SL g1247 ( 
.A(n_1217),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1118),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_SL g1249 ( 
.A1(n_1091),
.A2(n_1108),
.B1(n_1142),
.B2(n_1161),
.Y(n_1249)
);

BUFx10_ASAP7_75t_L g1250 ( 
.A(n_1119),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1125),
.Y(n_1251)
);

CKINVDCx8_ASAP7_75t_R g1252 ( 
.A(n_1138),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1185),
.Y(n_1253)
);

CKINVDCx11_ASAP7_75t_R g1254 ( 
.A(n_1236),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1091),
.A2(n_1206),
.B1(n_1153),
.B2(n_1143),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_1152),
.Y(n_1256)
);

INVx6_ASAP7_75t_L g1257 ( 
.A(n_1105),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1149),
.A2(n_1095),
.B1(n_1200),
.B2(n_1155),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1140),
.Y(n_1259)
);

OR2x2_ASAP7_75t_L g1260 ( 
.A(n_1114),
.B(n_1107),
.Y(n_1260)
);

BUFx4_ASAP7_75t_R g1261 ( 
.A(n_1170),
.Y(n_1261)
);

INVx6_ASAP7_75t_L g1262 ( 
.A(n_1105),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1199),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1221),
.A2(n_1114),
.B1(n_1200),
.B2(n_1107),
.Y(n_1264)
);

BUFx12f_ASAP7_75t_L g1265 ( 
.A(n_1211),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1222),
.Y(n_1266)
);

CKINVDCx20_ASAP7_75t_R g1267 ( 
.A(n_1102),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1151),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_1205),
.Y(n_1269)
);

BUFx2_ASAP7_75t_SL g1270 ( 
.A(n_1224),
.Y(n_1270)
);

BUFx4f_ASAP7_75t_SL g1271 ( 
.A(n_1211),
.Y(n_1271)
);

OAI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1237),
.A2(n_1124),
.B1(n_1136),
.B2(n_1137),
.Y(n_1272)
);

INVx6_ASAP7_75t_L g1273 ( 
.A(n_1110),
.Y(n_1273)
);

BUFx10_ASAP7_75t_L g1274 ( 
.A(n_1173),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_1228),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1226),
.Y(n_1276)
);

NAND2x1p5_ASAP7_75t_L g1277 ( 
.A(n_1208),
.B(n_1201),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1104),
.A2(n_1218),
.B1(n_1204),
.B2(n_1187),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1120),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_SL g1280 ( 
.A1(n_1161),
.A2(n_1167),
.B1(n_1165),
.B2(n_1175),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1184),
.A2(n_1231),
.B1(n_1132),
.B2(n_1110),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1230),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1124),
.A2(n_1233),
.B1(n_1135),
.B2(n_1127),
.Y(n_1283)
);

BUFx10_ASAP7_75t_L g1284 ( 
.A(n_1174),
.Y(n_1284)
);

INVx6_ASAP7_75t_L g1285 ( 
.A(n_1170),
.Y(n_1285)
);

OAI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1136),
.A2(n_1175),
.B1(n_1197),
.B2(n_1096),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1133),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1159),
.A2(n_1128),
.B1(n_1167),
.B2(n_1131),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1147),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1159),
.A2(n_1131),
.B1(n_1154),
.B2(n_1158),
.Y(n_1290)
);

CKINVDCx11_ASAP7_75t_R g1291 ( 
.A(n_1168),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_SL g1292 ( 
.A1(n_1192),
.A2(n_1122),
.B1(n_1154),
.B2(n_1158),
.Y(n_1292)
);

OAI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1103),
.A2(n_1162),
.B1(n_1141),
.B2(n_1192),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1097),
.A2(n_1234),
.B1(n_1225),
.B2(n_1179),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1162),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1103),
.A2(n_1134),
.B1(n_1156),
.B2(n_1192),
.Y(n_1296)
);

INVx4_ASAP7_75t_L g1297 ( 
.A(n_1170),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1166),
.Y(n_1298)
);

INVx4_ASAP7_75t_L g1299 ( 
.A(n_1170),
.Y(n_1299)
);

INVx6_ASAP7_75t_L g1300 ( 
.A(n_1170),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1163),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1166),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1157),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1215),
.B(n_1169),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1134),
.A2(n_1123),
.B1(n_1090),
.B2(n_1160),
.Y(n_1305)
);

INVx3_ASAP7_75t_L g1306 ( 
.A(n_1121),
.Y(n_1306)
);

BUFx10_ASAP7_75t_L g1307 ( 
.A(n_1170),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1189),
.A2(n_1194),
.B1(n_1213),
.B2(n_1210),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1195),
.A2(n_1207),
.B1(n_1106),
.B2(n_1176),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1178),
.Y(n_1310)
);

BUFx3_ASAP7_75t_L g1311 ( 
.A(n_1215),
.Y(n_1311)
);

CKINVDCx20_ASAP7_75t_R g1312 ( 
.A(n_1171),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1090),
.A2(n_1094),
.B1(n_1150),
.B2(n_1223),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1094),
.A2(n_1223),
.B1(n_1198),
.B2(n_1146),
.Y(n_1314)
);

CKINVDCx11_ASAP7_75t_R g1315 ( 
.A(n_1172),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1181),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1190),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1190),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1190),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_1139),
.Y(n_1320)
);

CKINVDCx11_ASAP7_75t_R g1321 ( 
.A(n_1111),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1198),
.A2(n_1115),
.B1(n_1116),
.B2(n_1164),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_SL g1323 ( 
.A1(n_1196),
.A2(n_1148),
.B1(n_1099),
.B2(n_1117),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1145),
.A2(n_1196),
.B1(n_1229),
.B2(n_1098),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1219),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1101),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1092),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1099),
.Y(n_1328)
);

BUFx6f_ASAP7_75t_SL g1329 ( 
.A(n_1099),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1126),
.A2(n_1182),
.B1(n_1193),
.B2(n_1202),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1203),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1209),
.A2(n_692),
.B1(n_446),
.B2(n_603),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_SL g1333 ( 
.A1(n_1227),
.A2(n_603),
.B(n_1212),
.Y(n_1333)
);

INVxp67_ASAP7_75t_SL g1334 ( 
.A(n_1232),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1183),
.B(n_1214),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_SL g1336 ( 
.A1(n_1112),
.A2(n_497),
.B1(n_308),
.B2(n_312),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1118),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1118),
.Y(n_1338)
);

BUFx10_ASAP7_75t_L g1339 ( 
.A(n_1119),
.Y(n_1339)
);

CKINVDCx11_ASAP7_75t_R g1340 ( 
.A(n_1236),
.Y(n_1340)
);

BUFx6f_ASAP7_75t_SL g1341 ( 
.A(n_1186),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1217),
.Y(n_1342)
);

CKINVDCx11_ASAP7_75t_R g1343 ( 
.A(n_1236),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1118),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1220),
.A2(n_692),
.B1(n_446),
.B2(n_603),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1212),
.A2(n_603),
.B1(n_1235),
.B2(n_822),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1212),
.A2(n_603),
.B1(n_1235),
.B2(n_822),
.Y(n_1347)
);

INVxp33_ASAP7_75t_L g1348 ( 
.A(n_1119),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1147),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1118),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1220),
.A2(n_692),
.B1(n_446),
.B2(n_603),
.Y(n_1351)
);

INVx1_ASAP7_75t_SL g1352 ( 
.A(n_1217),
.Y(n_1352)
);

BUFx2_ASAP7_75t_SL g1353 ( 
.A(n_1102),
.Y(n_1353)
);

CKINVDCx20_ASAP7_75t_R g1354 ( 
.A(n_1236),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_1236),
.Y(n_1355)
);

CKINVDCx6p67_ASAP7_75t_R g1356 ( 
.A(n_1236),
.Y(n_1356)
);

INVxp67_ASAP7_75t_SL g1357 ( 
.A(n_1112),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1129),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1236),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1220),
.A2(n_692),
.B1(n_446),
.B2(n_603),
.Y(n_1360)
);

BUFx6f_ASAP7_75t_L g1361 ( 
.A(n_1180),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1220),
.A2(n_692),
.B1(n_446),
.B2(n_603),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1129),
.Y(n_1363)
);

CKINVDCx6p67_ASAP7_75t_R g1364 ( 
.A(n_1236),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1212),
.A2(n_603),
.B1(n_1235),
.B2(n_822),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1316),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1317),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1318),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1295),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1325),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1310),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1297),
.B(n_1299),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1324),
.A2(n_1309),
.B(n_1308),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1249),
.B(n_1296),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1294),
.A2(n_1322),
.B(n_1314),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1322),
.A2(n_1314),
.B(n_1331),
.Y(n_1376)
);

CKINVDCx6p67_ASAP7_75t_R g1377 ( 
.A(n_1254),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1296),
.B(n_1248),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1302),
.Y(n_1379)
);

AOI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1327),
.A2(n_1259),
.B(n_1255),
.Y(n_1380)
);

OA21x2_ASAP7_75t_L g1381 ( 
.A1(n_1305),
.A2(n_1313),
.B(n_1333),
.Y(n_1381)
);

BUFx3_ASAP7_75t_L g1382 ( 
.A(n_1298),
.Y(n_1382)
);

NAND3x1_ASAP7_75t_L g1383 ( 
.A(n_1239),
.B(n_1281),
.C(n_1335),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1266),
.B(n_1276),
.Y(n_1384)
);

INVx1_ASAP7_75t_SL g1385 ( 
.A(n_1291),
.Y(n_1385)
);

INVx3_ASAP7_75t_L g1386 ( 
.A(n_1320),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1305),
.A2(n_1313),
.B(n_1268),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1312),
.Y(n_1388)
);

AO21x2_ASAP7_75t_L g1389 ( 
.A1(n_1293),
.A2(n_1286),
.B(n_1319),
.Y(n_1389)
);

BUFx3_ASAP7_75t_L g1390 ( 
.A(n_1349),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1245),
.A2(n_1246),
.B1(n_1347),
.B2(n_1346),
.Y(n_1391)
);

NOR2x1_ASAP7_75t_SL g1392 ( 
.A(n_1258),
.B(n_1261),
.Y(n_1392)
);

OA21x2_ASAP7_75t_L g1393 ( 
.A1(n_1328),
.A2(n_1334),
.B(n_1268),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1320),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1348),
.B(n_1250),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1282),
.Y(n_1396)
);

BUFx2_ASAP7_75t_L g1397 ( 
.A(n_1326),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1326),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1337),
.B(n_1338),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1240),
.A2(n_1244),
.B(n_1286),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1344),
.Y(n_1401)
);

AO21x2_ASAP7_75t_L g1402 ( 
.A1(n_1293),
.A2(n_1272),
.B(n_1238),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1329),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1329),
.Y(n_1404)
);

AOI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1259),
.A2(n_1304),
.B(n_1303),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1350),
.Y(n_1406)
);

INVxp67_ASAP7_75t_L g1407 ( 
.A(n_1241),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1279),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1287),
.Y(n_1409)
);

CKINVDCx14_ASAP7_75t_R g1410 ( 
.A(n_1340),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1240),
.Y(n_1411)
);

OAI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1365),
.A2(n_1244),
.B(n_1246),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1260),
.B(n_1272),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1283),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1278),
.B(n_1283),
.Y(n_1415)
);

AO31x2_ASAP7_75t_L g1416 ( 
.A1(n_1251),
.A2(n_1253),
.A3(n_1301),
.B(n_1323),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1285),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1290),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1264),
.A2(n_1290),
.B(n_1306),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1357),
.B(n_1311),
.Y(n_1420)
);

BUFx2_ASAP7_75t_L g1421 ( 
.A(n_1311),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1278),
.B(n_1264),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1292),
.B(n_1332),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1288),
.B(n_1358),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1261),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1363),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1306),
.A2(n_1332),
.B(n_1277),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1330),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1285),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1238),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1300),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1300),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1280),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1307),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1284),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1284),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1277),
.A2(n_1362),
.B(n_1360),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_SL g1438 ( 
.A(n_1355),
.B(n_1359),
.Y(n_1438)
);

AOI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1243),
.A2(n_1289),
.B(n_1256),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1345),
.A2(n_1360),
.B(n_1351),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_1361),
.B(n_1349),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1315),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1321),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1247),
.B(n_1342),
.Y(n_1444)
);

CKINVDCx11_ASAP7_75t_R g1445 ( 
.A(n_1354),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1345),
.A2(n_1351),
.B(n_1362),
.Y(n_1446)
);

AO32x1_ASAP7_75t_L g1447 ( 
.A1(n_1391),
.A2(n_1242),
.A3(n_1263),
.B1(n_1348),
.B2(n_1352),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1390),
.B(n_1339),
.Y(n_1448)
);

O2A1O1Ixp33_ASAP7_75t_SL g1449 ( 
.A1(n_1412),
.A2(n_1267),
.B(n_1271),
.C(n_1364),
.Y(n_1449)
);

OR2x6_ASAP7_75t_L g1450 ( 
.A(n_1400),
.B(n_1425),
.Y(n_1450)
);

AO32x1_ASAP7_75t_L g1451 ( 
.A1(n_1374),
.A2(n_1250),
.A3(n_1339),
.B1(n_1273),
.B2(n_1336),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1390),
.B(n_1274),
.Y(n_1452)
);

AND2x4_ASAP7_75t_L g1453 ( 
.A(n_1390),
.B(n_1275),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1382),
.B(n_1274),
.Y(n_1454)
);

NOR2x1_ASAP7_75t_SL g1455 ( 
.A(n_1439),
.B(n_1265),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1382),
.B(n_1269),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1426),
.B(n_1273),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1396),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1388),
.B(n_1353),
.Y(n_1459)
);

A2O1A1Ixp33_ASAP7_75t_L g1460 ( 
.A1(n_1374),
.A2(n_1270),
.B(n_1341),
.C(n_1271),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1379),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1439),
.B(n_1424),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1388),
.B(n_1252),
.Y(n_1463)
);

INVx4_ASAP7_75t_L g1464 ( 
.A(n_1372),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1411),
.B(n_1257),
.Y(n_1465)
);

BUFx2_ASAP7_75t_L g1466 ( 
.A(n_1441),
.Y(n_1466)
);

OA21x2_ASAP7_75t_L g1467 ( 
.A1(n_1373),
.A2(n_1262),
.B(n_1341),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1396),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1393),
.Y(n_1469)
);

OAI211xp5_ASAP7_75t_L g1470 ( 
.A1(n_1428),
.A2(n_1343),
.B(n_1356),
.C(n_1262),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1420),
.B(n_1429),
.Y(n_1471)
);

OAI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1433),
.A2(n_1422),
.B1(n_1430),
.B2(n_1411),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1384),
.B(n_1399),
.Y(n_1473)
);

AO21x2_ASAP7_75t_L g1474 ( 
.A1(n_1405),
.A2(n_1402),
.B(n_1428),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1429),
.B(n_1392),
.Y(n_1475)
);

OA21x2_ASAP7_75t_L g1476 ( 
.A1(n_1375),
.A2(n_1376),
.B(n_1387),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1401),
.Y(n_1477)
);

AOI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1433),
.A2(n_1383),
.B1(n_1402),
.B2(n_1430),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1421),
.Y(n_1479)
);

AOI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1383),
.A2(n_1402),
.B1(n_1415),
.B2(n_1423),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1401),
.B(n_1406),
.Y(n_1481)
);

OAI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1419),
.A2(n_1413),
.B(n_1375),
.Y(n_1482)
);

AO32x2_ASAP7_75t_L g1483 ( 
.A1(n_1378),
.A2(n_1415),
.A3(n_1422),
.B1(n_1414),
.B2(n_1418),
.Y(n_1483)
);

AO21x2_ASAP7_75t_L g1484 ( 
.A1(n_1380),
.A2(n_1389),
.B(n_1376),
.Y(n_1484)
);

OAI21xp33_ASAP7_75t_L g1485 ( 
.A1(n_1419),
.A2(n_1423),
.B(n_1369),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_SL g1486 ( 
.A1(n_1392),
.A2(n_1440),
.B1(n_1446),
.B2(n_1381),
.Y(n_1486)
);

A2O1A1Ixp33_ASAP7_75t_L g1487 ( 
.A1(n_1446),
.A2(n_1437),
.B(n_1427),
.C(n_1387),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1397),
.B(n_1398),
.Y(n_1488)
);

O2A1O1Ixp33_ASAP7_75t_SL g1489 ( 
.A1(n_1385),
.A2(n_1443),
.B(n_1436),
.C(n_1435),
.Y(n_1489)
);

O2A1O1Ixp33_ASAP7_75t_SL g1490 ( 
.A1(n_1443),
.A2(n_1435),
.B(n_1436),
.C(n_1395),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1407),
.B(n_1444),
.Y(n_1491)
);

AOI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1434),
.A2(n_1442),
.B(n_1397),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1408),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1398),
.B(n_1417),
.Y(n_1494)
);

OAI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1381),
.A2(n_1427),
.B(n_1434),
.Y(n_1495)
);

OAI21xp33_ASAP7_75t_SL g1496 ( 
.A1(n_1369),
.A2(n_1442),
.B(n_1432),
.Y(n_1496)
);

OA21x2_ASAP7_75t_L g1497 ( 
.A1(n_1437),
.A2(n_1370),
.B(n_1366),
.Y(n_1497)
);

AOI221xp5_ASAP7_75t_L g1498 ( 
.A1(n_1370),
.A2(n_1366),
.B1(n_1367),
.B2(n_1368),
.C(n_1371),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1408),
.B(n_1409),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_1459),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1473),
.B(n_1381),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1461),
.B(n_1381),
.Y(n_1502)
);

BUFx4f_ASAP7_75t_L g1503 ( 
.A(n_1467),
.Y(n_1503)
);

NOR3xp33_ASAP7_75t_L g1504 ( 
.A(n_1470),
.B(n_1410),
.C(n_1445),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1461),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1469),
.Y(n_1506)
);

NAND3xp33_ASAP7_75t_L g1507 ( 
.A(n_1478),
.B(n_1431),
.C(n_1432),
.Y(n_1507)
);

BUFx2_ASAP7_75t_SL g1508 ( 
.A(n_1456),
.Y(n_1508)
);

BUFx2_ASAP7_75t_L g1509 ( 
.A(n_1488),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1458),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1475),
.B(n_1394),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1468),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1477),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1479),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1488),
.B(n_1386),
.Y(n_1515)
);

INVx1_ASAP7_75t_SL g1516 ( 
.A(n_1479),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_1467),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1481),
.B(n_1389),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1462),
.B(n_1416),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1493),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1471),
.B(n_1386),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_SL g1522 ( 
.A(n_1460),
.B(n_1377),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1497),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1497),
.Y(n_1524)
);

NOR2xp67_ASAP7_75t_L g1525 ( 
.A(n_1469),
.B(n_1496),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1497),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1462),
.B(n_1416),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1499),
.Y(n_1528)
);

OAI221xp5_ASAP7_75t_L g1529 ( 
.A1(n_1480),
.A2(n_1440),
.B1(n_1403),
.B2(n_1404),
.C(n_1438),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1471),
.B(n_1393),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1472),
.A2(n_1440),
.B1(n_1403),
.B2(n_1404),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1492),
.Y(n_1532)
);

AOI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1472),
.A2(n_1440),
.B1(n_1404),
.B2(n_1403),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1482),
.B(n_1416),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_SL g1535 ( 
.A1(n_1508),
.A2(n_1456),
.B1(n_1529),
.B2(n_1450),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1502),
.B(n_1491),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1525),
.B(n_1475),
.Y(n_1537)
);

NAND4xp25_ASAP7_75t_SL g1538 ( 
.A(n_1504),
.B(n_1463),
.C(n_1486),
.D(n_1377),
.Y(n_1538)
);

AOI331xp33_ASAP7_75t_L g1539 ( 
.A1(n_1510),
.A2(n_1449),
.A3(n_1483),
.B1(n_1489),
.B2(n_1447),
.B3(n_1453),
.C1(n_1451),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1505),
.Y(n_1540)
);

INVx3_ASAP7_75t_L g1541 ( 
.A(n_1511),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1509),
.B(n_1454),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1509),
.B(n_1454),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1501),
.B(n_1498),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1501),
.B(n_1456),
.Y(n_1545)
);

AOI221xp5_ASAP7_75t_SL g1546 ( 
.A1(n_1502),
.A2(n_1485),
.B1(n_1495),
.B2(n_1457),
.C(n_1487),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1525),
.B(n_1464),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1505),
.B(n_1474),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1518),
.B(n_1466),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1510),
.Y(n_1550)
);

AOI221xp5_ASAP7_75t_L g1551 ( 
.A1(n_1519),
.A2(n_1527),
.B1(n_1534),
.B2(n_1529),
.C(n_1507),
.Y(n_1551)
);

NOR3xp33_ASAP7_75t_L g1552 ( 
.A(n_1507),
.B(n_1490),
.C(n_1489),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1512),
.Y(n_1553)
);

BUFx6f_ASAP7_75t_L g1554 ( 
.A(n_1517),
.Y(n_1554)
);

INVx1_ASAP7_75t_SL g1555 ( 
.A(n_1516),
.Y(n_1555)
);

OR2x6_ASAP7_75t_L g1556 ( 
.A(n_1508),
.B(n_1450),
.Y(n_1556)
);

INVxp67_ASAP7_75t_SL g1557 ( 
.A(n_1519),
.Y(n_1557)
);

AOI211xp5_ASAP7_75t_L g1558 ( 
.A1(n_1522),
.A2(n_1449),
.B(n_1490),
.C(n_1487),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1531),
.A2(n_1474),
.B1(n_1450),
.B2(n_1451),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1531),
.A2(n_1450),
.B1(n_1451),
.B2(n_1484),
.Y(n_1560)
);

OAI211xp5_ASAP7_75t_L g1561 ( 
.A1(n_1527),
.A2(n_1448),
.B(n_1465),
.C(n_1452),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1515),
.B(n_1471),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1533),
.A2(n_1451),
.B1(n_1484),
.B2(n_1476),
.Y(n_1563)
);

AOI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1522),
.A2(n_1447),
.B(n_1455),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1513),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1530),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1528),
.B(n_1494),
.Y(n_1567)
);

NAND4xp25_ASAP7_75t_SL g1568 ( 
.A(n_1504),
.B(n_1447),
.C(n_1483),
.D(n_1453),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1550),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1566),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_SL g1571 ( 
.A(n_1539),
.B(n_1500),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1544),
.B(n_1506),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1544),
.B(n_1506),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1537),
.B(n_1511),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1550),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1536),
.B(n_1528),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1536),
.B(n_1534),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1540),
.B(n_1516),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1553),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1557),
.B(n_1520),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1547),
.B(n_1530),
.Y(n_1581)
);

NOR2x1_ASAP7_75t_L g1582 ( 
.A(n_1538),
.B(n_1453),
.Y(n_1582)
);

AOI221xp5_ASAP7_75t_L g1583 ( 
.A1(n_1568),
.A2(n_1526),
.B1(n_1524),
.B2(n_1523),
.C(n_1532),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1547),
.B(n_1530),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1547),
.B(n_1514),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1547),
.B(n_1514),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_SL g1587 ( 
.A(n_1558),
.B(n_1537),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1553),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1540),
.B(n_1520),
.Y(n_1589)
);

INVx1_ASAP7_75t_SL g1590 ( 
.A(n_1555),
.Y(n_1590)
);

INVx5_ASAP7_75t_L g1591 ( 
.A(n_1554),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1537),
.B(n_1511),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1548),
.Y(n_1593)
);

INVx3_ASAP7_75t_L g1594 ( 
.A(n_1554),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1541),
.B(n_1514),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1541),
.B(n_1521),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1565),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1570),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1571),
.B(n_1561),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1574),
.B(n_1545),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1574),
.B(n_1545),
.Y(n_1601)
);

NAND2x1_ASAP7_75t_L g1602 ( 
.A(n_1574),
.B(n_1537),
.Y(n_1602)
);

NAND2x1p5_ASAP7_75t_L g1603 ( 
.A(n_1591),
.B(n_1503),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1572),
.B(n_1565),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1569),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1572),
.B(n_1548),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1569),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1590),
.B(n_1555),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1573),
.B(n_1551),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1575),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1592),
.B(n_1542),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1573),
.B(n_1567),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1575),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1579),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1590),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1579),
.B(n_1588),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1570),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1592),
.B(n_1542),
.Y(n_1618)
);

INVxp67_ASAP7_75t_L g1619 ( 
.A(n_1587),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1570),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1592),
.B(n_1552),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1591),
.B(n_1556),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1585),
.B(n_1543),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1588),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1597),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1578),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1585),
.B(n_1543),
.Y(n_1627)
);

BUFx2_ASAP7_75t_L g1628 ( 
.A(n_1582),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1585),
.B(n_1562),
.Y(n_1629)
);

AOI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1583),
.A2(n_1533),
.B1(n_1559),
.B2(n_1546),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1576),
.B(n_1567),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1591),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1576),
.B(n_1549),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1586),
.B(n_1562),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1591),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1597),
.B(n_1546),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1583),
.A2(n_1560),
.B1(n_1558),
.B2(n_1563),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1605),
.Y(n_1638)
);

OAI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1637),
.A2(n_1630),
.B1(n_1609),
.B2(n_1619),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1609),
.B(n_1593),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1615),
.B(n_1582),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1636),
.B(n_1593),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1628),
.B(n_1586),
.Y(n_1643)
);

NOR2xp67_ASAP7_75t_L g1644 ( 
.A(n_1630),
.B(n_1591),
.Y(n_1644)
);

INVx1_ASAP7_75t_SL g1645 ( 
.A(n_1628),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1636),
.B(n_1580),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1637),
.B(n_1626),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1605),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1611),
.B(n_1591),
.Y(n_1649)
);

NAND2xp33_ASAP7_75t_R g1650 ( 
.A(n_1621),
.B(n_1586),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_SL g1651 ( 
.A(n_1621),
.B(n_1591),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1604),
.B(n_1577),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1611),
.B(n_1581),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1618),
.B(n_1581),
.Y(n_1654)
);

INVx2_ASAP7_75t_SL g1655 ( 
.A(n_1602),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1618),
.B(n_1581),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1600),
.B(n_1584),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1600),
.B(n_1584),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1604),
.B(n_1577),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1601),
.B(n_1584),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1607),
.B(n_1580),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1598),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1601),
.B(n_1629),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1612),
.B(n_1589),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1629),
.B(n_1595),
.Y(n_1665)
);

NAND2xp33_ASAP7_75t_SL g1666 ( 
.A(n_1602),
.B(n_1595),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1634),
.B(n_1595),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1634),
.B(n_1596),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1612),
.B(n_1589),
.Y(n_1669)
);

INVx1_ASAP7_75t_SL g1670 ( 
.A(n_1621),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1621),
.B(n_1594),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1607),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1662),
.Y(n_1673)
);

O2A1O1Ixp33_ASAP7_75t_SL g1674 ( 
.A1(n_1639),
.A2(n_1599),
.B(n_1608),
.C(n_1635),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1638),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1639),
.B(n_1631),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1663),
.B(n_1623),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1638),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1640),
.B(n_1631),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1648),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1662),
.Y(n_1681)
);

OAI322xp33_ASAP7_75t_L g1682 ( 
.A1(n_1647),
.A2(n_1606),
.A3(n_1633),
.B1(n_1616),
.B2(n_1613),
.C1(n_1614),
.C2(n_1625),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_SL g1683 ( 
.A(n_1644),
.B(n_1622),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1640),
.B(n_1623),
.Y(n_1684)
);

OAI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1644),
.A2(n_1641),
.B1(n_1647),
.B2(n_1670),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1648),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1646),
.B(n_1627),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1672),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1672),
.Y(n_1689)
);

INVxp67_ASAP7_75t_SL g1690 ( 
.A(n_1642),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1664),
.Y(n_1691)
);

OAI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1646),
.A2(n_1564),
.B1(n_1554),
.B2(n_1603),
.Y(n_1692)
);

OAI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1642),
.A2(n_1554),
.B1(n_1603),
.B2(n_1633),
.Y(n_1693)
);

AOI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1645),
.A2(n_1447),
.B(n_1535),
.Y(n_1694)
);

OAI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1645),
.A2(n_1606),
.B(n_1603),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1670),
.B(n_1627),
.Y(n_1696)
);

OAI21xp33_ASAP7_75t_L g1697 ( 
.A1(n_1643),
.A2(n_1616),
.B(n_1614),
.Y(n_1697)
);

INVxp67_ASAP7_75t_L g1698 ( 
.A(n_1676),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1674),
.B(n_1655),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1690),
.B(n_1663),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1673),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1673),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1676),
.A2(n_1650),
.B1(n_1662),
.B2(n_1535),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1677),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1696),
.A2(n_1655),
.B1(n_1658),
.B2(n_1657),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1681),
.Y(n_1706)
);

OA21x2_ASAP7_75t_L g1707 ( 
.A1(n_1681),
.A2(n_1651),
.B(n_1635),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1675),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1677),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1691),
.Y(n_1710)
);

INVx2_ASAP7_75t_SL g1711 ( 
.A(n_1683),
.Y(n_1711)
);

OAI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1685),
.A2(n_1660),
.B1(n_1657),
.B2(n_1658),
.Y(n_1712)
);

AOI322xp5_ASAP7_75t_L g1713 ( 
.A1(n_1679),
.A2(n_1661),
.A3(n_1643),
.B1(n_1617),
.B2(n_1620),
.C1(n_1598),
.C2(n_1666),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1684),
.B(n_1660),
.Y(n_1714)
);

OAI22xp33_ASAP7_75t_SL g1715 ( 
.A1(n_1683),
.A2(n_1669),
.B1(n_1664),
.B2(n_1661),
.Y(n_1715)
);

AOI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1674),
.A2(n_1598),
.B1(n_1620),
.B2(n_1617),
.Y(n_1716)
);

NAND2xp33_ASAP7_75t_SL g1717 ( 
.A(n_1711),
.B(n_1687),
.Y(n_1717)
);

AOI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1698),
.A2(n_1694),
.B1(n_1692),
.B2(n_1695),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1704),
.B(n_1669),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1714),
.B(n_1653),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1707),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1702),
.Y(n_1722)
);

AOI22xp33_ASAP7_75t_L g1723 ( 
.A1(n_1698),
.A2(n_1682),
.B1(n_1678),
.B2(n_1680),
.Y(n_1723)
);

INVx1_ASAP7_75t_SL g1724 ( 
.A(n_1700),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1708),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1702),
.Y(n_1726)
);

XOR2xp5_ASAP7_75t_L g1727 ( 
.A(n_1712),
.B(n_1671),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1707),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1720),
.B(n_1709),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1719),
.Y(n_1730)
);

OAI32xp33_ASAP7_75t_L g1731 ( 
.A1(n_1721),
.A2(n_1699),
.A3(n_1728),
.B1(n_1723),
.B2(n_1717),
.Y(n_1731)
);

NOR3x1_ASAP7_75t_SL g1732 ( 
.A(n_1725),
.B(n_1708),
.C(n_1715),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1721),
.Y(n_1733)
);

NOR2x1_ASAP7_75t_L g1734 ( 
.A(n_1728),
.B(n_1699),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1724),
.B(n_1710),
.Y(n_1735)
);

AOI21xp33_ASAP7_75t_L g1736 ( 
.A1(n_1723),
.A2(n_1710),
.B(n_1706),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1725),
.B(n_1701),
.Y(n_1737)
);

AOI211xp5_ASAP7_75t_L g1738 ( 
.A1(n_1718),
.A2(n_1693),
.B(n_1705),
.C(n_1703),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1731),
.A2(n_1727),
.B(n_1707),
.Y(n_1739)
);

AOI221xp5_ASAP7_75t_L g1740 ( 
.A1(n_1736),
.A2(n_1732),
.B1(n_1733),
.B2(n_1735),
.C(n_1722),
.Y(n_1740)
);

OAI211xp5_ASAP7_75t_L g1741 ( 
.A1(n_1734),
.A2(n_1713),
.B(n_1697),
.C(n_1726),
.Y(n_1741)
);

AOI322xp5_ASAP7_75t_L g1742 ( 
.A1(n_1730),
.A2(n_1716),
.A3(n_1689),
.B1(n_1686),
.B2(n_1688),
.C1(n_1617),
.C2(n_1620),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1729),
.Y(n_1743)
);

OAI211xp5_ASAP7_75t_SL g1744 ( 
.A1(n_1740),
.A2(n_1738),
.B(n_1737),
.C(n_1632),
.Y(n_1744)
);

AOI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1739),
.A2(n_1671),
.B(n_1649),
.Y(n_1745)
);

AOI221xp5_ASAP7_75t_L g1746 ( 
.A1(n_1741),
.A2(n_1671),
.B1(n_1652),
.B2(n_1659),
.C(n_1632),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1743),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1742),
.B(n_1665),
.Y(n_1748)
);

AOI221xp5_ASAP7_75t_L g1749 ( 
.A1(n_1740),
.A2(n_1671),
.B1(n_1652),
.B2(n_1659),
.C(n_1632),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1747),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1748),
.Y(n_1751)
);

OAI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1745),
.A2(n_1635),
.B(n_1649),
.Y(n_1752)
);

INVxp67_ASAP7_75t_SL g1753 ( 
.A(n_1749),
.Y(n_1753)
);

NAND2x1_ASAP7_75t_L g1754 ( 
.A(n_1744),
.B(n_1649),
.Y(n_1754)
);

NOR3xp33_ASAP7_75t_L g1755 ( 
.A(n_1750),
.B(n_1746),
.C(n_1649),
.Y(n_1755)
);

NOR3xp33_ASAP7_75t_SL g1756 ( 
.A(n_1753),
.B(n_1613),
.C(n_1624),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1752),
.B(n_1653),
.Y(n_1757)
);

INVxp67_ASAP7_75t_L g1758 ( 
.A(n_1755),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1758),
.Y(n_1759)
);

INVx3_ASAP7_75t_L g1760 ( 
.A(n_1759),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1759),
.Y(n_1761)
);

OAI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1760),
.A2(n_1751),
.B1(n_1754),
.B2(n_1756),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1760),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1763),
.B(n_1761),
.Y(n_1764)
);

OAI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1762),
.A2(n_1757),
.B1(n_1654),
.B2(n_1656),
.Y(n_1765)
);

OAI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1764),
.A2(n_1610),
.B1(n_1625),
.B2(n_1624),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_SL g1767 ( 
.A(n_1766),
.B(n_1765),
.Y(n_1767)
);

HB1xp67_ASAP7_75t_L g1768 ( 
.A(n_1767),
.Y(n_1768)
);

AOI221xp5_ASAP7_75t_L g1769 ( 
.A1(n_1768),
.A2(n_1610),
.B1(n_1654),
.B2(n_1656),
.C(n_1665),
.Y(n_1769)
);

AOI211xp5_ASAP7_75t_L g1770 ( 
.A1(n_1769),
.A2(n_1667),
.B(n_1668),
.C(n_1622),
.Y(n_1770)
);


endmodule