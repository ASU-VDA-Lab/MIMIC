module fake_jpeg_8849_n_295 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_19),
.Y(n_55)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_41),
.Y(n_46)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_29),
.Y(n_56)
);

OAI21xp33_ASAP7_75t_L g84 ( 
.A1(n_56),
.A2(n_67),
.B(n_68),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_29),
.B1(n_31),
.B2(n_28),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_57),
.A2(n_62),
.B1(n_32),
.B2(n_22),
.Y(n_92)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_29),
.B1(n_27),
.B2(n_20),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_31),
.B1(n_18),
.B2(n_27),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_17),
.B1(n_28),
.B2(n_31),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_51),
.B1(n_17),
.B2(n_56),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_20),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_34),
.B(n_26),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_34),
.B(n_33),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_SL g87 ( 
.A(n_69),
.B(n_28),
.Y(n_87)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_45),
.A2(n_55),
.B1(n_28),
.B2(n_63),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_76),
.A2(n_81),
.B1(n_90),
.B2(n_92),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_44),
.Y(n_79)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_69),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_46),
.A2(n_22),
.B1(n_32),
.B2(n_19),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_83),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_94),
.B(n_30),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_70),
.A2(n_47),
.B1(n_65),
.B2(n_67),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_95),
.A2(n_112),
.B1(n_22),
.B2(n_32),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_17),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_98),
.A2(n_107),
.B(n_115),
.Y(n_127)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_103),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_84),
.C(n_89),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_110),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_86),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_117),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_105),
.B(n_108),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_17),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_88),
.B(n_65),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_88),
.A2(n_47),
.B1(n_73),
.B2(n_78),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_65),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_73),
.B(n_26),
.Y(n_116)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_77),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_102),
.A2(n_91),
.B1(n_89),
.B2(n_75),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_118),
.A2(n_130),
.B1(n_135),
.B2(n_136),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_71),
.B1(n_52),
.B2(n_53),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_138),
.B1(n_104),
.B2(n_99),
.Y(n_151)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_124),
.Y(n_165)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_37),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_137),
.Y(n_159)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_128),
.B(n_129),
.Y(n_166)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_111),
.A2(n_91),
.B1(n_78),
.B2(n_79),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_132),
.B(n_93),
.Y(n_147)
);

AO22x1_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_43),
.B1(n_42),
.B2(n_59),
.Y(n_133)
);

AO22x1_ASAP7_75t_L g152 ( 
.A1(n_133),
.A2(n_61),
.B1(n_49),
.B2(n_64),
.Y(n_152)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_115),
.A2(n_42),
.B1(n_43),
.B2(n_58),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_107),
.A2(n_43),
.B1(n_60),
.B2(n_19),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_16),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_141),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_30),
.B(n_24),
.C(n_25),
.Y(n_140)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_23),
.Y(n_141)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_93),
.B(n_105),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_144),
.A2(n_154),
.B(n_0),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_108),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_145),
.A2(n_24),
.B(n_1),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_12),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_146),
.B(n_150),
.Y(n_176)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_139),
.A2(n_109),
.B1(n_101),
.B2(n_106),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_148),
.A2(n_160),
.B1(n_163),
.B2(n_169),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_137),
.B(n_9),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_151),
.Y(n_184)
);

OA22x2_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_161),
.B1(n_0),
.B2(n_1),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_127),
.A2(n_23),
.B(n_21),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_156),
.Y(n_177)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_130),
.A2(n_61),
.B1(n_64),
.B2(n_100),
.Y(n_160)
);

OA22x2_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_133),
.A2(n_61),
.B1(n_64),
.B2(n_74),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_127),
.A2(n_25),
.B1(n_24),
.B2(n_23),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_164),
.A2(n_142),
.B1(n_143),
.B2(n_122),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_23),
.Y(n_173)
);

AO22x1_ASAP7_75t_L g168 ( 
.A1(n_135),
.A2(n_140),
.B1(n_136),
.B2(n_118),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_169),
.Y(n_182)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_170),
.B(n_179),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_120),
.C(n_126),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_172),
.C(n_175),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_120),
.C(n_141),
.Y(n_172)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_113),
.C(n_114),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_114),
.C(n_74),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_181),
.C(n_188),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_23),
.Y(n_179)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_23),
.C(n_25),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_153),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_183),
.B(n_191),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_185),
.B(n_161),
.Y(n_209)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_194),
.Y(n_202)
);

NAND2xp33_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_161),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_7),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_144),
.A2(n_7),
.B1(n_13),
.B2(n_11),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_189),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_149),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_153),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_165),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_192),
.B(n_146),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_1),
.C(n_2),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_150),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_145),
.B(n_1),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_177),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_196),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_177),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_203),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_209),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_145),
.Y(n_205)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_155),
.Y(n_206)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_168),
.Y(n_207)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_168),
.Y(n_210)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_184),
.A2(n_160),
.B1(n_149),
.B2(n_163),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_211),
.A2(n_201),
.B1(n_210),
.B2(n_207),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_156),
.Y(n_212)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_213),
.A2(n_187),
.B1(n_148),
.B2(n_161),
.Y(n_219)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_214),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_158),
.Y(n_216)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_219),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_171),
.C(n_172),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_225),
.C(n_227),
.Y(n_244)
);

FAx1_ASAP7_75t_SL g224 ( 
.A(n_205),
.B(n_182),
.CI(n_190),
.CON(n_224),
.SN(n_224)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_229),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_182),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_175),
.C(n_178),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_199),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_201),
.A2(n_188),
.B1(n_180),
.B2(n_193),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_231),
.A2(n_195),
.B1(n_197),
.B2(n_202),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_185),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_233),
.B(n_212),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_235),
.A2(n_209),
.B1(n_197),
.B2(n_203),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_196),
.Y(n_236)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_225),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_238),
.B(n_245),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_239),
.Y(n_259)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_242),
.Y(n_257)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_235),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_246),
.B(n_247),
.Y(n_258)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_248),
.B(n_249),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_217),
.A2(n_203),
.B1(n_200),
.B2(n_211),
.Y(n_249)
);

AOI21xp33_ASAP7_75t_L g250 ( 
.A1(n_232),
.A2(n_202),
.B(n_198),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_218),
.C(n_230),
.Y(n_254)
);

NAND2xp33_ASAP7_75t_SL g252 ( 
.A(n_249),
.B(n_224),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_252),
.A2(n_256),
.B1(n_257),
.B2(n_236),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_181),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_254),
.A2(n_243),
.B(n_234),
.Y(n_263)
);

A2O1A1Ixp33_ASAP7_75t_SL g256 ( 
.A1(n_242),
.A2(n_226),
.B(n_224),
.C(n_219),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_222),
.C(n_227),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_238),
.C(n_239),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_233),
.C(n_226),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_176),
.C(n_187),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_263),
.B(n_268),
.Y(n_276)
);

NOR2xp67_ASAP7_75t_SL g264 ( 
.A(n_262),
.B(n_237),
.Y(n_264)
);

NOR2xp67_ASAP7_75t_SL g277 ( 
.A(n_264),
.B(n_9),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_266),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_240),
.C(n_231),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_260),
.B1(n_255),
.B2(n_258),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_267),
.B(n_256),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_270),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_200),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_271),
.A2(n_9),
.B(n_13),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_252),
.A2(n_187),
.B(n_152),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_272),
.A2(n_8),
.B(n_11),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_268),
.B1(n_280),
.B2(n_276),
.Y(n_283)
);

NAND4xp25_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_256),
.C(n_152),
.D(n_4),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_274),
.A2(n_277),
.B(n_278),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_279),
.B(n_10),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_282),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_275),
.B(n_269),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_283),
.A2(n_285),
.B(n_286),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_4),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_6),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_284),
.A2(n_6),
.B(n_8),
.Y(n_289)
);

NOR3xp33_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_290),
.C(n_2),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_284),
.A2(n_6),
.B1(n_11),
.B2(n_14),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_287),
.A2(n_2),
.B(n_3),
.Y(n_291)
);

BUFx24_ASAP7_75t_SL g293 ( 
.A(n_291),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_288),
.B(n_292),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_3),
.Y(n_295)
);


endmodule