module fake_jpeg_27329_n_329 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx8_ASAP7_75t_SL g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g66 ( 
.A(n_36),
.Y(n_66)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_8),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_45),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_29),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_50),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_29),
.B1(n_23),
.B2(n_24),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_51),
.A2(n_19),
.B1(n_20),
.B2(n_17),
.Y(n_91)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

NAND2xp33_ASAP7_75t_SL g58 ( 
.A(n_36),
.B(n_32),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_36),
.Y(n_78)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_63),
.Y(n_90)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_24),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_67),
.Y(n_76)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_24),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_68),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_23),
.B1(n_30),
.B2(n_32),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_72),
.A2(n_81),
.B1(n_91),
.B2(n_17),
.Y(n_100)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_73),
.B(n_83),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_57),
.A2(n_38),
.B1(n_23),
.B2(n_19),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_77),
.A2(n_95),
.B1(n_33),
.B2(n_63),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_40),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_19),
.B1(n_21),
.B2(n_17),
.Y(n_81)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_48),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_85),
.Y(n_98)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

BUFx12_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_57),
.A2(n_20),
.B1(n_25),
.B2(n_31),
.Y(n_95)
);

CKINVDCx6p67_ASAP7_75t_R g96 ( 
.A(n_66),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_89),
.A2(n_56),
.B1(n_20),
.B2(n_55),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_100),
.A2(n_101),
.B1(n_70),
.B2(n_85),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_90),
.A2(n_55),
.B1(n_58),
.B2(n_49),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_106),
.B(n_92),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_67),
.B1(n_64),
.B2(n_54),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_107),
.A2(n_114),
.B1(n_85),
.B2(n_74),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_66),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_43),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_87),
.B(n_33),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_111),
.B(n_123),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_36),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_43),
.C(n_41),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_113),
.A2(n_16),
.B(n_22),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_91),
.A2(n_64),
.B1(n_53),
.B2(n_60),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_79),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_74),
.Y(n_125)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_119),
.Y(n_137)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_71),
.A2(n_33),
.B1(n_28),
.B2(n_8),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_120),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_78),
.A2(n_26),
.B(n_28),
.C(n_8),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_71),
.A2(n_28),
.B1(n_15),
.B2(n_14),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_96),
.B1(n_94),
.B2(n_13),
.Y(n_141)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_78),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_121),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_128),
.A2(n_138),
.B1(n_108),
.B2(n_117),
.Y(n_178)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_143),
.Y(n_161)
);

NOR2xp67_ASAP7_75t_SL g131 ( 
.A(n_123),
.B(n_76),
.Y(n_131)
);

XOR2x2_ASAP7_75t_L g180 ( 
.A(n_131),
.B(n_149),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_114),
.A2(n_83),
.B1(n_70),
.B2(n_86),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_139),
.B1(n_141),
.B2(n_150),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_40),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_136),
.Y(n_162)
);

MAJx2_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_88),
.C(n_96),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_146),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_116),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_140),
.Y(n_166)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_145),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_103),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_84),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_106),
.B(n_94),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_151),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_96),
.C(n_41),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_110),
.C(n_115),
.Y(n_160)
);

XNOR2x1_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_26),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_93),
.B1(n_82),
.B2(n_43),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_102),
.B(n_41),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_102),
.B(n_16),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_118),
.Y(n_171)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_157),
.B(n_169),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_142),
.A2(n_126),
.B1(n_147),
.B2(n_128),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_159),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_156),
.C(n_135),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_110),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_163),
.B(n_160),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_140),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_168),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_151),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_137),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_173),
.Y(n_204)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_105),
.Y(n_172)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_150),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_105),
.Y(n_174)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_152),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_181),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_126),
.A2(n_136),
.B1(n_134),
.B2(n_133),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_133),
.A2(n_108),
.B1(n_115),
.B2(n_118),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_139),
.A2(n_99),
.B1(n_122),
.B2(n_104),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_179),
.A2(n_88),
.B1(n_21),
.B2(n_27),
.Y(n_200)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_131),
.A2(n_99),
.B1(n_122),
.B2(n_21),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_183),
.A2(n_129),
.B1(n_149),
.B2(n_141),
.Y(n_191)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_130),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_187),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_146),
.A2(n_82),
.B1(n_104),
.B2(n_21),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_185),
.A2(n_26),
.B1(n_22),
.B2(n_16),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_154),
.Y(n_186)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_130),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_191),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_161),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_194),
.Y(n_227)
);

OA22x2_ASAP7_75t_L g193 ( 
.A1(n_173),
.A2(n_135),
.B1(n_144),
.B2(n_153),
.Y(n_193)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_193),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_175),
.A2(n_165),
.B1(n_180),
.B2(n_166),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_158),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_195),
.A2(n_212),
.B(n_216),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_213),
.C(n_214),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_156),
.B(n_144),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_201),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_200),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_22),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_165),
.A2(n_31),
.B1(n_27),
.B2(n_25),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_203),
.A2(n_209),
.B1(n_215),
.B2(n_187),
.Y(n_222)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_184),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_158),
.A2(n_31),
.B1(n_27),
.B2(n_25),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_179),
.A2(n_31),
.B1(n_27),
.B2(n_25),
.Y(n_211)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_211),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_176),
.A2(n_26),
.B1(n_9),
.B2(n_10),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_22),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_26),
.C(n_22),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_159),
.A2(n_15),
.B1(n_12),
.B2(n_11),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_204),
.A2(n_162),
.B(n_164),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_221),
.Y(n_250)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_222),
.A2(n_235),
.B1(n_241),
.B2(n_198),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_189),
.A2(n_195),
.B1(n_199),
.B2(n_164),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_224),
.A2(n_229),
.B1(n_203),
.B2(n_200),
.Y(n_247)
);

NAND3xp33_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_199),
.C(n_216),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_230),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_189),
.A2(n_162),
.B1(n_167),
.B2(n_155),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_238),
.Y(n_258)
);

INVxp33_ASAP7_75t_SL g233 ( 
.A(n_206),
.Y(n_233)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_192),
.A2(n_168),
.B(n_166),
.Y(n_234)
);

INVxp33_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

XNOR2x1_ASAP7_75t_L g235 ( 
.A(n_196),
.B(n_208),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_182),
.C(n_185),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_237),
.C(n_239),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_182),
.C(n_157),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_202),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_197),
.B(n_155),
.C(n_177),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_214),
.Y(n_246)
);

NAND2x1_ASAP7_75t_L g241 ( 
.A(n_193),
.B(n_16),
.Y(n_241)
);

NOR3xp33_ASAP7_75t_SL g243 ( 
.A(n_241),
.B(n_212),
.C(n_193),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_243),
.B(n_260),
.Y(n_268)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_241),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_252),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_249),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_247),
.A2(n_227),
.B1(n_232),
.B2(n_248),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_259),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_190),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_242),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_227),
.A2(n_188),
.B1(n_193),
.B2(n_215),
.Y(n_254)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_254),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_15),
.Y(n_255)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_16),
.C(n_12),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_263),
.C(n_236),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_223),
.B(n_235),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_219),
.B(n_11),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_10),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_256),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_220),
.B(n_0),
.C(n_1),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_262),
.A2(n_228),
.B1(n_224),
.B2(n_231),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_265),
.A2(n_237),
.B1(n_220),
.B2(n_244),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_267),
.A2(n_243),
.B1(n_247),
.B2(n_253),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_258),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_269),
.B(n_274),
.Y(n_289)
);

O2A1O1Ixp33_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_231),
.B(n_217),
.C(n_218),
.Y(n_270)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_272),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_242),
.Y(n_275)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_257),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_276),
.B(n_278),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_222),
.Y(n_279)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_280),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_283),
.B(n_291),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_264),
.A2(n_263),
.B1(n_249),
.B2(n_261),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_265),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_267),
.A2(n_246),
.B1(n_244),
.B2(n_259),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_288),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_6),
.C(n_1),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_268),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_2),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_5),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_3),
.C(n_4),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_274),
.C(n_278),
.Y(n_294)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_294),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_275),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_296),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_273),
.C(n_266),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_287),
.B(n_273),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_297),
.B(n_305),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_300),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_270),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_3),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_303),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_3),
.C(n_5),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_298),
.A2(n_285),
.B1(n_286),
.B2(n_282),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_306),
.B(n_308),
.Y(n_318)
);

NOR2xp67_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_289),
.Y(n_307)
);

OAI21x1_ASAP7_75t_L g316 ( 
.A1(n_307),
.A2(n_285),
.B(n_302),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_280),
.C(n_286),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_299),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_5),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_314),
.B(n_305),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_317),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_319),
.Y(n_322)
);

INVx11_ASAP7_75t_L g317 ( 
.A(n_309),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_5),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_312),
.B(n_311),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_321),
.B(n_310),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_318),
.B(n_322),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_323),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_318),
.B(n_313),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_6),
.B(n_318),
.Y(n_328)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_328),
.Y(n_329)
);


endmodule