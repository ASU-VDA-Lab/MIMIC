module fake_jpeg_1096_n_137 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_137);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx11_ASAP7_75t_SL g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_20),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_49),
.Y(n_60)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_16),
.C(n_32),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_58),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_51),
.A2(n_42),
.B1(n_45),
.B2(n_50),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_69),
.B1(n_40),
.B2(n_48),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_40),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_46),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_43),
.C(n_39),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_46),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_57),
.A2(n_42),
.B1(n_45),
.B2(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_73),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_71),
.A2(n_74),
.B1(n_76),
.B2(n_79),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_48),
.B(n_43),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_77),
.Y(n_95)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_81),
.C(n_0),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_76),
.B(n_64),
.Y(n_85)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

NOR2x1_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_82),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_65),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_39),
.B(n_15),
.C(n_17),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_30),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_35),
.C(n_31),
.Y(n_81)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_85),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_68),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_86),
.B(n_88),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_80),
.A2(n_68),
.B1(n_64),
.B2(n_2),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_78),
.B1(n_77),
.B2(n_7),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_94),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_0),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_92),
.B(n_93),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_1),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_2),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_3),
.B(n_4),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_4),
.Y(n_101)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_101),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_120)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_104),
.Y(n_118)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_108),
.Y(n_116)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

A2O1A1O1Ixp25_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_18),
.B(n_28),
.C(n_27),
.D(n_26),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_109),
.B(n_21),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_95),
.Y(n_111)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_111),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_29),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_89),
.C(n_25),
.Y(n_119)
);

AND2x4_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_87),
.Y(n_117)
);

NOR3xp33_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_119),
.C(n_121),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_120),
.Y(n_127)
);

AO221x1_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.C(n_11),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_122),
.A2(n_123),
.B(n_109),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_23),
.A3(n_24),
.B1(n_13),
.B2(n_14),
.C1(n_11),
.C2(n_12),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_116),
.A2(n_113),
.B1(n_99),
.B2(n_102),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_124),
.B(n_126),
.Y(n_128)
);

AOI321xp33_ASAP7_75t_L g129 ( 
.A1(n_124),
.A2(n_116),
.A3(n_114),
.B1(n_110),
.B2(n_115),
.C(n_98),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_130),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_118),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_128),
.A2(n_101),
.B(n_125),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_130),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_131),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_112),
.B(n_122),
.Y(n_135)
);

OAI21x1_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_117),
.B(n_13),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_14),
.Y(n_137)
);


endmodule