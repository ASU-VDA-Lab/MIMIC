module fake_ariane_1069_n_197 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_30, n_31, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_197);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_30;
input n_31;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_197;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_190;
wire n_160;
wire n_64;
wire n_179;
wire n_180;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_195;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_187;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_189;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_82;
wire n_178;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_101;
wire n_94;
wire n_134;
wire n_188;
wire n_185;
wire n_32;
wire n_58;
wire n_37;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_121;
wire n_93;
wire n_118;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_196;
wire n_125;
wire n_168;
wire n_43;
wire n_87;
wire n_81;
wire n_41;
wire n_140;
wire n_55;
wire n_191;
wire n_151;
wire n_136;
wire n_192;
wire n_80;
wire n_146;
wire n_194;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_193;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

INVxp67_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVxp33_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVxp67_ASAP7_75t_SL g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVxp67_ASAP7_75t_SL g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

INVxp33_ASAP7_75t_SL g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_29),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

INVxp33_ASAP7_75t_SL g47 ( 
.A(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

INVxp67_ASAP7_75t_SL g52 ( 
.A(n_28),
.Y(n_52)
);

INVxp67_ASAP7_75t_SL g53 ( 
.A(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_R g55 ( 
.A(n_38),
.B(n_31),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_42),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_51),
.Y(n_60)
);

AOI21x1_ASAP7_75t_L g61 ( 
.A1(n_33),
.A2(n_0),
.B(n_1),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_33),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_R g68 ( 
.A(n_45),
.B(n_26),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_R g69 ( 
.A(n_45),
.B(n_27),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_47),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_47),
.Y(n_71)
);

NAND2xp33_ASAP7_75t_R g72 ( 
.A(n_46),
.B(n_2),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_R g73 ( 
.A(n_46),
.B(n_23),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_50),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

AND2x6_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_39),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_34),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NAND2xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_34),
.Y(n_84)
);

NAND2x1p5_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_39),
.Y(n_85)
);

NAND2x1p5_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_39),
.Y(n_86)
);

BUFx6f_ASAP7_75t_SL g87 ( 
.A(n_58),
.Y(n_87)
);

AO22x2_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_41),
.B1(n_37),
.B2(n_53),
.Y(n_88)
);

AO22x2_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_41),
.B1(n_37),
.B2(n_53),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_36),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_R g93 ( 
.A(n_87),
.B(n_71),
.Y(n_93)
);

NOR2xp67_ASAP7_75t_SL g94 ( 
.A(n_80),
.B(n_35),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_92),
.A2(n_32),
.B(n_49),
.C(n_40),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_32),
.B(n_49),
.C(n_40),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_35),
.B(n_44),
.C(n_52),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_79),
.B(n_62),
.Y(n_98)
);

AOI33xp33_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_44),
.A3(n_70),
.B1(n_59),
.B2(n_48),
.B3(n_36),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_52),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_72),
.B1(n_48),
.B2(n_75),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_89),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_103),
.A2(n_101),
.B(n_97),
.C(n_95),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_SL g107 ( 
.A1(n_98),
.A2(n_91),
.B(n_90),
.C(n_83),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_104),
.A2(n_89),
.B1(n_88),
.B2(n_60),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_82),
.Y(n_110)
);

OAI21x1_ASAP7_75t_L g111 ( 
.A1(n_102),
.A2(n_86),
.B(n_85),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_100),
.A2(n_85),
.B(n_86),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_R g113 ( 
.A(n_109),
.B(n_87),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_111),
.Y(n_114)
);

NOR3xp33_ASAP7_75t_SL g115 ( 
.A(n_106),
.B(n_72),
.C(n_96),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

NAND3xp33_ASAP7_75t_SL g117 ( 
.A(n_110),
.B(n_69),
.C(n_68),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_105),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_116),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_105),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_105),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_108),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_115),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_108),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_118),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_110),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_88),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_88),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

NOR2xp67_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_131),
.Y(n_143)
);

OAI211xp5_ASAP7_75t_L g144 ( 
.A1(n_142),
.A2(n_117),
.B(n_55),
.C(n_69),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_140),
.A2(n_116),
.B(n_112),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_130),
.Y(n_147)
);

NAND2x1_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_116),
.Y(n_148)
);

AOI321xp33_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_127),
.A3(n_125),
.B1(n_135),
.B2(n_126),
.C(n_88),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_135),
.Y(n_151)
);

AOI221xp5_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_89),
.B1(n_117),
.B2(n_55),
.C(n_107),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_144),
.A2(n_140),
.B(n_94),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_136),
.C(n_140),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_136),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_151),
.A2(n_89),
.B1(n_138),
.B2(n_87),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_138),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_89),
.B1(n_87),
.B2(n_126),
.Y(n_163)
);

OAI211xp5_ASAP7_75t_L g164 ( 
.A1(n_157),
.A2(n_148),
.B(n_149),
.C(n_73),
.Y(n_164)
);

OAI211xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_148),
.B(n_113),
.C(n_146),
.Y(n_165)
);

INVxp67_ASAP7_75t_SL g166 ( 
.A(n_159),
.Y(n_166)
);

AOI222xp33_ASAP7_75t_L g167 ( 
.A1(n_160),
.A2(n_77),
.B1(n_99),
.B2(n_91),
.C1(n_90),
.C2(n_94),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_2),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_161),
.A2(n_77),
.B1(n_81),
.B2(n_86),
.Y(n_169)
);

NAND3xp33_ASAP7_75t_SL g170 ( 
.A(n_154),
.B(n_85),
.C(n_5),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_R g171 ( 
.A(n_153),
.B(n_3),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_171),
.B(n_112),
.Y(n_172)
);

NAND2x1p5_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_76),
.Y(n_173)
);

AOI211x1_ASAP7_75t_SL g174 ( 
.A1(n_170),
.A2(n_162),
.B(n_6),
.C(n_7),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_166),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_5),
.Y(n_176)
);

O2A1O1Ixp5_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_8),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_173),
.Y(n_180)
);

NOR2x1_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_167),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_179),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_R g183 ( 
.A(n_178),
.B(n_9),
.Y(n_183)
);

AND2x4_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_11),
.Y(n_184)
);

O2A1O1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_182),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_174),
.Y(n_187)
);

AO21x1_ASAP7_75t_L g188 ( 
.A1(n_184),
.A2(n_174),
.B(n_16),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_180),
.A2(n_13),
.B1(n_17),
.B2(n_18),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_186),
.Y(n_190)
);

OAI22x1_ASAP7_75t_L g191 ( 
.A1(n_187),
.A2(n_183),
.B1(n_185),
.B2(n_17),
.Y(n_191)
);

OAI31xp67_ASAP7_75t_SL g192 ( 
.A1(n_188),
.A2(n_189),
.A3(n_18),
.B(n_77),
.Y(n_192)
);

AOI221xp5_ASAP7_75t_L g193 ( 
.A1(n_191),
.A2(n_76),
.B1(n_77),
.B2(n_102),
.C(n_190),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_191),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_77),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_R g196 ( 
.A1(n_194),
.A2(n_102),
.B1(n_77),
.B2(n_76),
.Y(n_196)
);

AOI221xp5_ASAP7_75t_L g197 ( 
.A1(n_196),
.A2(n_77),
.B1(n_193),
.B2(n_195),
.C(n_194),
.Y(n_197)
);


endmodule