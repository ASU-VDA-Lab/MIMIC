module fake_jpeg_6971_n_99 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_99);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_99;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx2_ASAP7_75t_SL g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_4),
.B(n_7),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_8),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_19),
.B(n_0),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_24),
.A2(n_31),
.B(n_5),
.Y(n_53)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_25),
.B(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_28),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_0),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_14),
.Y(n_35)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_12),
.Y(n_46)
);

AOI21xp33_ASAP7_75t_L g31 ( 
.A1(n_15),
.A2(n_0),
.B(n_1),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_21),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_32),
.A2(n_3),
.B(n_4),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_33),
.Y(n_37)
);

OAI22x1_ASAP7_75t_SL g34 ( 
.A1(n_29),
.A2(n_18),
.B1(n_12),
.B2(n_21),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_48),
.B(n_52),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_49),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_18),
.C(n_22),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_42),
.C(n_44),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_24),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_17),
.Y(n_60)
);

AND2x6_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_14),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_14),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_47),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_30),
.A2(n_20),
.B1(n_23),
.B2(n_17),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_25),
.B(n_1),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_27),
.B(n_12),
.C(n_20),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_6),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_45),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_59),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_60),
.B(n_35),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_48),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVxp33_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_66),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_42),
.B1(n_34),
.B2(n_53),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_74),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_38),
.C(n_52),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_73),
.Y(n_86)
);

XOR2x2_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_41),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_40),
.C(n_37),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_78),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_77),
.A2(n_57),
.B(n_61),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_41),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_82),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_80),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_77),
.C(n_78),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_81),
.Y(n_92)
);

MAJx2_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_86),
.C(n_85),
.Y(n_88)
);

AOI322xp5_ASAP7_75t_L g93 ( 
.A1(n_88),
.A2(n_56),
.A3(n_72),
.B1(n_60),
.B2(n_35),
.C1(n_66),
.C2(n_55),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_66),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_95),
.Y(n_96)
);

AOI322xp5_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_94),
.A3(n_91),
.B1(n_87),
.B2(n_66),
.C1(n_63),
.C2(n_36),
.Y(n_97)
);

AOI322xp5_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_67),
.A3(n_56),
.B1(n_55),
.B2(n_64),
.C1(n_84),
.C2(n_54),
.Y(n_94)
);

OAI21x1_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_90),
.B(n_23),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_96),
.C(n_9),
.Y(n_99)
);


endmodule